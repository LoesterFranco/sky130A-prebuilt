magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 257 1234 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 96 93 126 177
rect 195 93 225 177
rect 393 47 423 177
rect 503 47 533 177
rect 597 47 627 177
rect 681 47 711 177
rect 795 47 825 177
rect 889 47 919 177
rect 983 47 1013 177
rect 1087 47 1117 177
<< pmoshvt >>
rect 81 410 117 494
rect 188 297 224 381
rect 389 297 425 497
rect 495 297 531 497
rect 589 297 625 497
rect 683 297 719 497
rect 797 297 833 497
rect 891 297 927 497
rect 985 297 1021 497
rect 1079 297 1115 497
<< ndiff >>
rect 34 149 96 177
rect 34 115 42 149
rect 76 115 96 149
rect 34 93 96 115
rect 126 149 195 177
rect 126 115 141 149
rect 175 115 195 149
rect 126 93 195 115
rect 225 149 277 177
rect 225 115 235 149
rect 269 115 277 149
rect 225 93 277 115
rect 331 96 393 177
rect 331 62 339 96
rect 373 62 393 96
rect 331 47 393 62
rect 423 115 503 177
rect 423 81 449 115
rect 483 81 503 115
rect 423 47 503 81
rect 533 97 597 177
rect 533 63 543 97
rect 577 63 597 97
rect 533 47 597 63
rect 627 115 681 177
rect 627 81 637 115
rect 671 81 681 115
rect 627 47 681 81
rect 711 97 795 177
rect 711 63 749 97
rect 783 63 795 97
rect 711 47 795 63
rect 825 114 889 177
rect 825 80 845 114
rect 879 80 889 114
rect 825 47 889 80
rect 919 95 983 177
rect 919 61 939 95
rect 973 61 983 95
rect 919 47 983 61
rect 1013 163 1087 177
rect 1013 129 1033 163
rect 1067 129 1087 163
rect 1013 95 1087 129
rect 1013 61 1033 95
rect 1067 61 1087 95
rect 1013 47 1087 61
rect 1117 95 1169 177
rect 1117 61 1127 95
rect 1161 61 1169 95
rect 1117 47 1169 61
<< pdiff >>
rect 27 475 81 494
rect 27 441 35 475
rect 69 441 81 475
rect 27 410 81 441
rect 117 482 171 494
rect 117 448 129 482
rect 163 448 171 482
rect 117 410 171 448
rect 134 381 171 410
rect 335 425 389 497
rect 335 391 343 425
rect 377 391 389 425
rect 134 297 188 381
rect 224 346 278 381
rect 224 312 236 346
rect 270 312 278 346
rect 224 297 278 312
rect 335 297 389 391
rect 425 297 495 497
rect 531 297 589 497
rect 625 297 683 497
rect 719 477 797 497
rect 719 443 740 477
rect 774 443 797 477
rect 719 409 797 443
rect 719 375 740 409
rect 774 375 797 409
rect 719 297 797 375
rect 833 477 891 497
rect 833 443 845 477
rect 879 443 891 477
rect 833 409 891 443
rect 833 375 845 409
rect 879 375 891 409
rect 833 341 891 375
rect 833 307 845 341
rect 879 307 891 341
rect 833 297 891 307
rect 927 477 985 497
rect 927 443 939 477
rect 973 443 985 477
rect 927 409 985 443
rect 927 375 939 409
rect 973 375 985 409
rect 927 297 985 375
rect 1021 477 1079 497
rect 1021 443 1033 477
rect 1067 443 1079 477
rect 1021 409 1079 443
rect 1021 375 1033 409
rect 1067 375 1079 409
rect 1021 341 1079 375
rect 1021 307 1033 341
rect 1067 307 1079 341
rect 1021 297 1079 307
rect 1115 477 1169 497
rect 1115 443 1127 477
rect 1161 443 1169 477
rect 1115 409 1169 443
rect 1115 375 1127 409
rect 1161 375 1169 409
rect 1115 297 1169 375
<< ndiffc >>
rect 42 115 76 149
rect 141 115 175 149
rect 235 115 269 149
rect 339 62 373 96
rect 449 81 483 115
rect 543 63 577 97
rect 637 81 671 115
rect 749 63 783 97
rect 845 80 879 114
rect 939 61 973 95
rect 1033 129 1067 163
rect 1033 61 1067 95
rect 1127 61 1161 95
<< pdiffc >>
rect 35 441 69 475
rect 129 448 163 482
rect 343 391 377 425
rect 236 312 270 346
rect 740 443 774 477
rect 740 375 774 409
rect 845 443 879 477
rect 845 375 879 409
rect 845 307 879 341
rect 939 443 973 477
rect 939 375 973 409
rect 1033 443 1067 477
rect 1033 375 1067 409
rect 1033 307 1067 341
rect 1127 443 1161 477
rect 1127 375 1161 409
<< poly >>
rect 81 494 117 520
rect 389 497 425 523
rect 495 497 531 523
rect 589 497 625 523
rect 683 497 719 523
rect 797 497 833 523
rect 891 497 927 523
rect 985 497 1021 523
rect 1079 497 1115 523
rect 81 395 117 410
rect 79 265 119 395
rect 188 381 224 407
rect 188 282 224 297
rect 389 282 425 297
rect 495 282 531 297
rect 589 282 625 297
rect 683 282 719 297
rect 797 282 833 297
rect 891 282 927 297
rect 985 282 1021 297
rect 1079 282 1115 297
rect 186 265 226 282
rect 387 265 427 282
rect 493 265 533 282
rect 587 265 627 282
rect 681 265 721 282
rect 795 265 835 282
rect 889 265 929 282
rect 983 265 1023 282
rect 1077 265 1117 282
rect 75 249 139 265
rect 75 215 87 249
rect 121 215 139 249
rect 75 199 139 215
rect 186 249 259 265
rect 186 215 199 249
rect 233 215 259 249
rect 186 199 259 215
rect 315 249 427 265
rect 315 215 325 249
rect 359 215 427 249
rect 315 199 427 215
rect 469 249 533 265
rect 469 215 479 249
rect 513 215 533 249
rect 469 199 533 215
rect 575 249 639 265
rect 575 215 585 249
rect 619 215 639 249
rect 575 199 639 215
rect 681 249 745 265
rect 681 215 691 249
rect 725 215 745 249
rect 681 199 745 215
rect 795 249 1117 265
rect 795 215 805 249
rect 839 215 883 249
rect 917 215 961 249
rect 995 215 1039 249
rect 1073 215 1117 249
rect 795 199 1117 215
rect 96 177 126 199
rect 195 177 225 199
rect 393 177 423 199
rect 503 177 533 199
rect 597 177 627 199
rect 681 177 711 199
rect 795 177 825 199
rect 889 177 919 199
rect 983 177 1013 199
rect 1087 177 1117 199
rect 96 67 126 93
rect 195 67 225 93
rect 393 21 423 47
rect 503 21 533 47
rect 597 21 627 47
rect 681 21 711 47
rect 795 21 825 47
rect 889 21 919 47
rect 983 21 1013 47
rect 1087 21 1117 47
<< polycont >>
rect 87 215 121 249
rect 199 215 233 249
rect 325 215 359 249
rect 479 215 513 249
rect 585 215 619 249
rect 691 215 725 249
rect 805 215 839 249
rect 883 215 917 249
rect 961 215 995 249
rect 1039 215 1073 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 19 475 69 491
rect 19 441 35 475
rect 103 482 179 527
rect 103 448 129 482
rect 163 448 179 482
rect 245 459 513 493
rect 732 477 782 527
rect 19 414 69 441
rect 245 414 279 459
rect 19 380 279 414
rect 322 391 343 425
rect 377 391 445 425
rect 19 165 53 380
rect 87 249 165 339
rect 208 312 236 346
rect 270 312 339 346
rect 301 265 339 312
rect 121 215 165 249
rect 87 199 165 215
rect 199 249 267 265
rect 233 215 267 249
rect 199 199 267 215
rect 301 249 359 265
rect 301 215 325 249
rect 301 199 359 215
rect 301 165 339 199
rect 19 149 80 165
rect 19 115 42 149
rect 76 115 80 149
rect 19 90 80 115
rect 141 149 175 165
rect 141 17 175 115
rect 235 149 339 165
rect 269 131 339 149
rect 407 165 445 391
rect 479 249 513 459
rect 479 199 513 215
rect 569 249 629 475
rect 732 443 740 477
rect 774 443 782 477
rect 732 409 782 443
rect 732 375 740 409
rect 774 375 782 409
rect 732 359 782 375
rect 837 477 887 493
rect 837 443 845 477
rect 879 443 887 477
rect 837 409 887 443
rect 837 375 845 409
rect 879 375 887 409
rect 837 341 887 375
rect 931 477 981 527
rect 931 443 939 477
rect 973 443 981 477
rect 931 409 981 443
rect 931 375 939 409
rect 973 375 981 409
rect 931 359 981 375
rect 1025 477 1075 493
rect 1025 443 1033 477
rect 1067 443 1075 477
rect 1025 409 1075 443
rect 1025 375 1033 409
rect 1067 375 1075 409
rect 663 280 735 323
rect 837 307 845 341
rect 879 325 887 341
rect 1025 341 1075 375
rect 1119 477 1169 527
rect 1119 443 1127 477
rect 1161 443 1169 477
rect 1119 409 1169 443
rect 1119 375 1127 409
rect 1161 375 1169 409
rect 1119 359 1169 375
rect 1025 325 1033 341
rect 879 307 1033 325
rect 1067 325 1075 341
rect 1067 307 1171 325
rect 837 291 1171 307
rect 569 215 585 249
rect 619 215 629 249
rect 569 199 629 215
rect 691 249 735 280
rect 725 215 735 249
rect 691 199 735 215
rect 769 215 805 249
rect 839 215 883 249
rect 917 215 961 249
rect 995 215 1039 249
rect 1073 215 1089 249
rect 769 165 803 215
rect 1125 181 1171 291
rect 407 131 803 165
rect 845 163 1171 181
rect 845 145 1033 163
rect 235 90 269 115
rect 449 115 483 131
rect 323 62 339 96
rect 373 62 389 96
rect 323 17 389 62
rect 637 115 671 131
rect 449 61 483 81
rect 517 63 543 97
rect 577 63 593 97
rect 517 17 593 63
rect 845 114 895 145
rect 637 61 671 81
rect 723 63 749 97
rect 783 63 799 97
rect 723 17 799 63
rect 879 80 895 114
rect 1007 129 1033 145
rect 1067 145 1171 163
rect 1067 129 1083 145
rect 845 51 895 80
rect 939 95 973 111
rect 939 17 973 61
rect 1007 95 1083 129
rect 1007 61 1033 95
rect 1067 61 1083 95
rect 1007 51 1083 61
rect 1127 95 1161 111
rect 1127 17 1161 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
flabel corelocali s 213 221 247 255 0 FreeSans 400 0 0 0 D_N
port 4 nsew
flabel corelocali s 581 425 615 459 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel corelocali s 581 357 615 391 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel corelocali s 673 289 707 323 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 121 221 155 255 0 FreeSans 400 0 0 0 C_N
port 3 nsew
flabel corelocali s 1133 153 1167 187 0 FreeSans 400 0 0 0 X
port 9 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 1196 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 165908
string GDS_START 156888
<< end >>
