magic
tech sky130A
magscale 1 2
timestamp 1599588218
<< nwell >>
rect -38 335 2822 704
rect -38 332 800 335
rect 1129 332 2822 335
rect 1129 328 1903 332
rect 1601 311 1903 328
<< pwell >>
rect 0 0 2784 49
<< scpmos >>
rect 205 464 241 592
rect 305 464 341 592
rect 389 464 425 592
rect 479 464 515 592
rect 587 464 623 592
rect 701 464 737 592
rect 911 387 947 611
rect 1001 387 1037 611
rect 1205 463 1241 547
rect 1295 463 1331 547
rect 1373 463 1409 547
rect 1493 463 1529 547
rect 1691 347 1727 547
rect 1781 347 1817 547
rect 1936 489 1972 573
rect 2014 489 2050 573
rect 2141 489 2177 573
rect 2231 489 2267 573
rect 2367 368 2403 592
rect 2565 424 2601 592
rect 2669 368 2705 592
<< nmoslvt >>
rect 84 74 114 158
rect 282 90 312 174
rect 383 90 413 174
rect 515 97 545 181
rect 587 97 617 181
rect 682 88 712 172
rect 893 119 923 267
rect 1007 119 1037 267
rect 1205 119 1235 203
rect 1291 119 1321 203
rect 1369 119 1399 203
rect 1447 119 1477 203
rect 1631 74 1661 202
rect 1717 74 1747 202
rect 1936 74 1966 158
rect 2008 74 2038 158
rect 2094 74 2124 158
rect 2166 74 2196 158
rect 2378 74 2408 222
rect 2571 74 2601 184
rect 2669 74 2699 222
<< ndiff >>
rect 843 234 893 267
rect 458 174 515 181
rect 27 133 84 158
rect 27 99 39 133
rect 73 99 84 133
rect 27 74 84 99
rect 114 133 171 158
rect 114 99 125 133
rect 159 99 171 133
rect 114 74 171 99
rect 225 141 282 174
rect 225 107 237 141
rect 271 107 282 141
rect 225 90 282 107
rect 312 90 383 174
rect 413 169 515 174
rect 413 135 470 169
rect 504 135 515 169
rect 413 97 515 135
rect 545 97 587 181
rect 617 172 667 181
rect 819 186 893 234
rect 617 150 682 172
rect 617 116 628 150
rect 662 116 682 150
rect 617 97 682 116
rect 413 90 463 97
rect 632 88 682 97
rect 712 134 765 172
rect 712 100 723 134
rect 757 100 765 134
rect 819 152 845 186
rect 879 152 893 186
rect 819 119 893 152
rect 923 134 1007 267
rect 923 119 948 134
rect 712 88 765 100
rect 938 100 948 119
rect 982 119 1007 134
rect 1037 239 1091 267
rect 1037 205 1047 239
rect 1081 205 1091 239
rect 1037 165 1091 205
rect 1037 131 1047 165
rect 1081 131 1091 165
rect 1037 119 1091 131
rect 1152 176 1205 203
rect 1152 142 1160 176
rect 1194 142 1205 176
rect 1152 119 1205 142
rect 1235 169 1291 203
rect 1235 135 1246 169
rect 1280 135 1291 169
rect 1235 119 1291 135
rect 1321 119 1369 203
rect 1399 119 1447 203
rect 1477 202 1581 203
rect 1477 119 1631 202
rect 982 100 992 119
rect 938 84 992 100
rect 1492 85 1631 119
rect 1492 51 1504 85
rect 1538 74 1631 85
rect 1661 179 1717 202
rect 1661 145 1672 179
rect 1706 145 1717 179
rect 1661 74 1717 145
rect 1747 158 1797 202
rect 1747 131 1936 158
rect 1747 97 1857 131
rect 1891 97 1936 131
rect 1747 74 1936 97
rect 1966 74 2008 158
rect 2038 133 2094 158
rect 2038 99 2049 133
rect 2083 99 2094 133
rect 2038 74 2094 99
rect 2124 74 2166 158
rect 2196 127 2253 158
rect 2196 93 2207 127
rect 2241 93 2253 127
rect 2196 74 2253 93
rect 2307 82 2378 222
rect 1538 51 1550 74
rect 1492 39 1550 51
rect 2307 48 2318 82
rect 2352 74 2378 82
rect 2408 210 2464 222
rect 2408 176 2419 210
rect 2453 176 2464 210
rect 2616 210 2669 222
rect 2616 184 2624 210
rect 2408 120 2464 176
rect 2408 86 2419 120
rect 2453 86 2464 120
rect 2408 74 2464 86
rect 2518 146 2571 184
rect 2518 112 2526 146
rect 2560 112 2571 146
rect 2518 74 2571 112
rect 2601 176 2624 184
rect 2658 176 2669 210
rect 2601 120 2669 176
rect 2601 86 2624 120
rect 2658 86 2669 120
rect 2601 74 2669 86
rect 2699 210 2756 222
rect 2699 176 2710 210
rect 2744 176 2756 210
rect 2699 120 2756 176
rect 2699 86 2710 120
rect 2744 86 2756 120
rect 2699 74 2756 86
rect 2352 48 2363 74
rect 2307 36 2363 48
<< pdiff >>
rect 27 579 205 592
rect 27 545 39 579
rect 73 545 161 579
rect 195 545 205 579
rect 27 510 205 545
rect 27 476 39 510
rect 73 476 161 510
rect 195 476 205 510
rect 27 464 205 476
rect 241 584 305 592
rect 241 550 261 584
rect 295 550 305 584
rect 241 512 305 550
rect 241 478 261 512
rect 295 478 305 512
rect 241 464 305 478
rect 341 464 389 592
rect 425 584 479 592
rect 425 550 435 584
rect 469 550 479 584
rect 425 512 479 550
rect 425 478 435 512
rect 469 478 479 512
rect 425 464 479 478
rect 515 464 587 592
rect 623 580 701 592
rect 623 546 636 580
rect 670 546 701 580
rect 623 464 701 546
rect 737 584 793 592
rect 737 550 747 584
rect 781 550 793 584
rect 737 512 793 550
rect 737 478 747 512
rect 781 478 793 512
rect 737 464 793 478
rect 855 439 911 611
rect 855 405 867 439
rect 901 405 911 439
rect 855 387 911 405
rect 947 593 1001 611
rect 947 559 957 593
rect 991 559 1001 593
rect 947 387 1001 559
rect 1037 439 1091 611
rect 1037 405 1047 439
rect 1081 405 1091 439
rect 1037 387 1091 405
rect 1424 582 1478 594
rect 1424 548 1434 582
rect 1468 548 1478 582
rect 1424 547 1478 548
rect 2065 582 2126 594
rect 2065 573 2078 582
rect 1880 547 1936 573
rect 1151 522 1205 547
rect 1151 488 1161 522
rect 1195 488 1205 522
rect 1151 463 1205 488
rect 1241 534 1295 547
rect 1241 500 1251 534
rect 1285 500 1295 534
rect 1241 463 1295 500
rect 1331 463 1373 547
rect 1409 463 1493 547
rect 1529 524 1583 547
rect 1529 490 1539 524
rect 1573 490 1583 524
rect 1529 463 1583 490
rect 1637 535 1691 547
rect 1637 501 1647 535
rect 1681 501 1691 535
rect 1637 464 1691 501
rect 1637 430 1647 464
rect 1681 430 1691 464
rect 1637 393 1691 430
rect 1637 359 1647 393
rect 1681 359 1691 393
rect 1637 347 1691 359
rect 1727 535 1781 547
rect 1727 501 1737 535
rect 1771 501 1781 535
rect 1727 464 1781 501
rect 1727 430 1737 464
rect 1771 430 1781 464
rect 1727 393 1781 430
rect 1727 359 1737 393
rect 1771 359 1781 393
rect 1727 347 1781 359
rect 1817 535 1936 547
rect 1817 501 1892 535
rect 1926 501 1936 535
rect 1817 489 1936 501
rect 1972 489 2014 573
rect 2050 548 2078 573
rect 2112 573 2126 582
rect 2282 580 2367 592
rect 2282 573 2290 580
rect 2112 548 2141 573
rect 2050 489 2141 548
rect 2177 548 2231 573
rect 2177 514 2187 548
rect 2221 514 2231 548
rect 2177 489 2231 514
rect 2267 546 2290 573
rect 2324 546 2367 580
rect 2267 512 2367 546
rect 2267 489 2322 512
rect 1817 481 1869 489
rect 1817 447 1827 481
rect 1861 447 1869 481
rect 1817 401 1869 447
rect 1817 367 1827 401
rect 1861 367 1869 401
rect 2310 478 2322 489
rect 2356 478 2367 512
rect 1817 347 1869 367
rect 2310 444 2367 478
rect 2310 410 2322 444
rect 2356 410 2367 444
rect 2310 368 2367 410
rect 2403 580 2459 592
rect 2403 546 2413 580
rect 2447 546 2459 580
rect 2403 500 2459 546
rect 2403 466 2413 500
rect 2447 466 2459 500
rect 2403 428 2459 466
rect 2403 394 2413 428
rect 2447 394 2459 428
rect 2513 580 2565 592
rect 2513 546 2521 580
rect 2555 546 2565 580
rect 2513 470 2565 546
rect 2513 436 2521 470
rect 2555 436 2565 470
rect 2513 424 2565 436
rect 2601 580 2669 592
rect 2601 546 2618 580
rect 2652 546 2669 580
rect 2601 497 2669 546
rect 2601 463 2618 497
rect 2652 463 2669 497
rect 2601 424 2669 463
rect 2403 368 2459 394
rect 2617 414 2669 424
rect 2617 380 2625 414
rect 2659 380 2669 414
rect 2617 368 2669 380
rect 2705 580 2757 592
rect 2705 546 2715 580
rect 2749 546 2757 580
rect 2705 497 2757 546
rect 2705 463 2715 497
rect 2749 463 2757 497
rect 2705 414 2757 463
rect 2705 380 2715 414
rect 2749 380 2757 414
rect 2705 368 2757 380
<< ndiffc >>
rect 39 99 73 133
rect 125 99 159 133
rect 237 107 271 141
rect 470 135 504 169
rect 628 116 662 150
rect 723 100 757 134
rect 845 152 879 186
rect 948 100 982 134
rect 1047 205 1081 239
rect 1047 131 1081 165
rect 1160 142 1194 176
rect 1246 135 1280 169
rect 1504 51 1538 85
rect 1672 145 1706 179
rect 1857 97 1891 131
rect 2049 99 2083 133
rect 2207 93 2241 127
rect 2318 48 2352 82
rect 2419 176 2453 210
rect 2419 86 2453 120
rect 2526 112 2560 146
rect 2624 176 2658 210
rect 2624 86 2658 120
rect 2710 176 2744 210
rect 2710 86 2744 120
<< pdiffc >>
rect 39 545 73 579
rect 161 545 195 579
rect 39 476 73 510
rect 161 476 195 510
rect 261 550 295 584
rect 261 478 295 512
rect 435 550 469 584
rect 435 478 469 512
rect 636 546 670 580
rect 747 550 781 584
rect 747 478 781 512
rect 867 405 901 439
rect 957 559 991 593
rect 1047 405 1081 439
rect 1434 548 1468 582
rect 1161 488 1195 522
rect 1251 500 1285 534
rect 1539 490 1573 524
rect 1647 501 1681 535
rect 1647 430 1681 464
rect 1647 359 1681 393
rect 1737 501 1771 535
rect 1737 430 1771 464
rect 1737 359 1771 393
rect 1892 501 1926 535
rect 2078 548 2112 582
rect 2187 514 2221 548
rect 2290 546 2324 580
rect 1827 447 1861 481
rect 1827 367 1861 401
rect 2322 478 2356 512
rect 2322 410 2356 444
rect 2413 546 2447 580
rect 2413 466 2447 500
rect 2413 394 2447 428
rect 2521 546 2555 580
rect 2521 436 2555 470
rect 2618 546 2652 580
rect 2618 463 2652 497
rect 2625 380 2659 414
rect 2715 546 2749 580
rect 2715 463 2749 497
rect 2715 380 2749 414
<< poly >>
rect 205 592 241 618
rect 305 592 341 618
rect 389 592 425 618
rect 479 592 515 618
rect 587 592 623 618
rect 701 592 737 618
rect 911 611 947 637
rect 1001 611 1037 637
rect 1106 615 1817 645
rect 205 376 241 464
rect 305 376 341 464
rect 84 360 341 376
rect 84 326 137 360
rect 171 326 205 360
rect 239 326 273 360
rect 307 326 341 360
rect 84 310 341 326
rect 84 158 114 310
rect 389 262 425 464
rect 479 432 515 464
rect 587 449 623 464
rect 467 416 533 432
rect 467 382 483 416
rect 517 382 533 416
rect 467 366 533 382
rect 575 422 623 449
rect 701 430 737 464
rect 701 422 823 430
rect 575 406 641 422
rect 575 372 591 406
rect 625 372 641 406
rect 575 338 641 372
rect 213 246 279 262
rect 213 212 229 246
rect 263 226 279 246
rect 354 246 425 262
rect 467 302 533 318
rect 467 268 483 302
rect 517 268 533 302
rect 467 252 533 268
rect 263 212 312 226
rect 213 196 312 212
rect 354 212 370 246
rect 404 212 425 246
rect 354 196 425 212
rect 503 221 533 252
rect 575 304 591 338
rect 625 304 641 338
rect 575 288 641 304
rect 683 414 823 422
rect 683 380 773 414
rect 807 380 823 414
rect 683 364 823 380
rect 575 251 617 288
rect 503 196 545 221
rect 282 174 312 196
rect 383 174 413 196
rect 515 181 545 196
rect 587 181 617 251
rect 683 229 713 364
rect 911 355 947 387
rect 1001 372 1037 387
rect 879 339 947 355
rect 879 322 895 339
rect 755 306 895 322
rect 755 272 771 306
rect 805 305 895 306
rect 929 305 947 339
rect 805 282 947 305
rect 993 339 1059 372
rect 993 305 1009 339
rect 1043 312 1059 339
rect 1106 312 1136 615
rect 1205 547 1241 573
rect 1295 547 1331 615
rect 1373 547 1409 573
rect 1493 547 1529 573
rect 1691 547 1727 573
rect 1781 547 1817 615
rect 1936 573 1972 599
rect 2014 573 2050 599
rect 1205 381 1241 463
rect 1295 437 1331 463
rect 1178 365 1244 381
rect 1178 331 1194 365
rect 1228 345 1244 365
rect 1373 356 1409 463
rect 1493 430 1529 463
rect 1493 414 1605 430
rect 1493 400 1555 414
rect 1506 380 1555 400
rect 1589 380 1605 414
rect 1506 364 1605 380
rect 1228 331 1321 345
rect 1178 315 1321 331
rect 1043 305 1136 312
rect 993 282 1136 305
rect 805 272 821 282
rect 755 256 821 272
rect 893 267 923 282
rect 1007 267 1037 282
rect 682 187 713 229
rect 682 172 712 187
rect 84 48 114 74
rect 282 64 312 90
rect 383 64 413 90
rect 515 71 545 97
rect 587 71 617 97
rect 893 93 923 119
rect 1106 248 1136 282
rect 1106 218 1235 248
rect 1205 203 1235 218
rect 1291 203 1321 315
rect 1369 340 1458 356
rect 1369 306 1408 340
rect 1442 306 1458 340
rect 1369 290 1458 306
rect 1369 203 1399 290
rect 1506 248 1536 364
rect 2141 573 2177 599
rect 2231 573 2267 599
rect 2367 592 2403 618
rect 2565 592 2601 618
rect 2669 592 2705 618
rect 1936 446 1972 489
rect 1901 430 1972 446
rect 1901 396 1917 430
rect 1951 396 1972 430
rect 1901 380 1972 396
rect 2014 396 2050 489
rect 2141 474 2177 489
rect 2231 474 2267 489
rect 2141 444 2183 474
rect 2231 444 2285 474
rect 2153 402 2183 444
rect 2014 380 2105 396
rect 1691 319 1727 347
rect 1588 299 1727 319
rect 1781 332 1817 347
rect 2014 346 2055 380
rect 2089 346 2105 380
rect 1781 302 1966 332
rect 2014 330 2105 346
rect 2147 386 2213 402
rect 2147 352 2163 386
rect 2197 352 2213 386
rect 2147 336 2213 352
rect 2255 337 2285 444
rect 2367 337 2403 368
rect 2565 337 2601 424
rect 1588 265 1604 299
rect 1638 289 1727 299
rect 1638 265 1661 289
rect 1588 249 1661 265
rect 1447 218 1536 248
rect 1447 203 1477 218
rect 1631 202 1661 249
rect 1717 231 1887 247
rect 1717 217 1837 231
rect 1717 202 1747 217
rect 682 51 712 88
rect 1007 93 1037 119
rect 1205 93 1235 119
rect 1291 93 1321 119
rect 1369 93 1399 119
rect 1447 51 1477 119
rect 682 21 1477 51
rect 1821 197 1837 217
rect 1871 197 1887 231
rect 1821 181 1887 197
rect 1936 158 1966 302
rect 2008 300 2044 330
rect 2008 158 2038 300
rect 2147 282 2177 336
rect 2255 287 2601 337
rect 2669 326 2705 368
rect 2094 252 2177 282
rect 2219 271 2601 287
rect 2094 158 2124 252
rect 2219 237 2235 271
rect 2269 247 2408 271
rect 2269 237 2285 247
rect 2219 204 2285 237
rect 2378 222 2408 247
rect 2166 174 2285 204
rect 2166 158 2196 174
rect 1631 48 1661 74
rect 1717 48 1747 74
rect 1936 48 1966 74
rect 2008 48 2038 74
rect 2094 48 2124 74
rect 2166 48 2196 74
rect 2571 184 2601 271
rect 2643 310 2709 326
rect 2643 276 2659 310
rect 2693 276 2709 310
rect 2643 260 2709 276
rect 2669 222 2699 260
rect 2378 48 2408 74
rect 2571 48 2601 74
rect 2669 48 2699 74
<< polycont >>
rect 137 326 171 360
rect 205 326 239 360
rect 273 326 307 360
rect 483 382 517 416
rect 591 372 625 406
rect 229 212 263 246
rect 483 268 517 302
rect 370 212 404 246
rect 591 304 625 338
rect 773 380 807 414
rect 771 272 805 306
rect 895 305 929 339
rect 1009 305 1043 339
rect 1194 331 1228 365
rect 1555 380 1589 414
rect 1408 306 1442 340
rect 1917 396 1951 430
rect 2055 346 2089 380
rect 2163 352 2197 386
rect 1604 265 1638 299
rect 1837 197 1871 231
rect 2235 237 2269 271
rect 2659 276 2693 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 23 579 211 595
rect 23 545 39 579
rect 73 545 161 579
rect 195 545 211 579
rect 23 510 211 545
rect 23 476 39 510
rect 73 476 161 510
rect 195 476 211 510
rect 245 584 311 649
rect 245 550 261 584
rect 295 550 311 584
rect 245 512 311 550
rect 245 478 261 512
rect 295 478 311 512
rect 419 584 485 600
rect 419 550 435 584
rect 469 550 485 584
rect 419 512 485 550
rect 617 580 689 649
rect 617 546 636 580
rect 670 546 689 580
rect 723 584 797 600
rect 723 550 747 584
rect 781 550 797 584
rect 941 593 1007 649
rect 941 559 957 593
rect 991 559 1007 593
rect 1418 582 1484 649
rect 723 525 797 550
rect 1145 525 1195 551
rect 723 522 1195 525
rect 723 512 1161 522
rect 419 478 435 512
rect 469 478 747 512
rect 781 489 1161 512
rect 781 478 797 489
rect 23 444 211 476
rect 689 464 797 478
rect 1158 488 1161 489
rect 23 416 539 444
rect 23 410 483 416
rect 23 262 57 410
rect 473 382 483 410
rect 517 382 539 416
rect 121 360 359 376
rect 473 366 539 382
rect 587 406 653 430
rect 587 372 591 406
rect 625 372 653 406
rect 121 326 137 360
rect 171 326 205 360
rect 239 326 273 360
rect 307 332 359 360
rect 587 338 653 372
rect 307 326 545 332
rect 121 302 545 326
rect 121 298 483 302
rect 479 268 483 298
rect 517 268 545 302
rect 587 304 591 338
rect 625 304 653 338
rect 587 288 653 304
rect 23 246 279 262
rect 23 212 229 246
rect 263 212 279 246
rect 23 196 279 212
rect 313 246 420 262
rect 479 252 545 268
rect 313 212 370 246
rect 404 212 420 246
rect 689 218 723 464
rect 867 439 917 455
rect 757 424 833 430
rect 757 414 799 424
rect 757 380 773 414
rect 807 380 833 390
rect 901 423 917 439
rect 1031 439 1124 455
rect 901 405 997 423
rect 867 389 997 405
rect 1031 405 1047 439
rect 1081 405 1124 439
rect 1158 449 1195 488
rect 1235 534 1369 551
rect 1235 500 1251 534
rect 1285 500 1369 534
rect 1418 548 1434 582
rect 1468 548 1484 582
rect 1418 532 1484 548
rect 1235 498 1369 500
rect 1523 524 1589 551
rect 1523 498 1539 524
rect 1235 490 1539 498
rect 1573 490 1589 524
rect 1235 483 1589 490
rect 1335 464 1589 483
rect 1647 535 1697 649
rect 2061 582 2130 649
rect 1681 501 1697 535
rect 1647 464 1697 501
rect 1158 415 1301 449
rect 1031 389 1124 405
rect 757 364 833 380
rect 963 355 997 389
rect 1077 381 1124 389
rect 1077 365 1233 381
rect 879 339 929 355
rect 879 330 895 339
rect 757 306 895 330
rect 757 272 771 306
rect 805 305 895 306
rect 805 272 929 305
rect 757 236 929 272
rect 963 339 1043 355
rect 963 305 1009 339
rect 963 289 1043 305
rect 1077 331 1194 365
rect 1228 331 1233 365
rect 1077 315 1233 331
rect 23 133 73 196
rect 313 162 420 212
rect 454 184 723 218
rect 963 202 997 289
rect 1077 255 1124 315
rect 845 186 997 202
rect 454 169 520 184
rect 23 99 39 133
rect 23 70 73 99
rect 109 133 175 162
rect 109 99 125 133
rect 159 99 175 133
rect 109 17 175 99
rect 221 141 271 162
rect 221 107 237 141
rect 454 135 470 169
rect 504 135 520 169
rect 879 168 997 186
rect 1034 239 1124 255
rect 1267 253 1301 415
rect 1034 205 1047 239
rect 1081 221 1124 239
rect 1081 205 1084 221
rect 879 152 898 168
rect 454 119 520 135
rect 221 85 271 107
rect 612 116 628 150
rect 662 116 678 150
rect 612 85 678 116
rect 221 51 678 85
rect 712 134 773 150
rect 712 100 723 134
rect 757 100 773 134
rect 845 119 898 152
rect 1034 165 1084 205
rect 712 17 773 100
rect 932 100 948 134
rect 982 100 998 134
rect 932 17 998 100
rect 1034 131 1047 165
rect 1081 131 1084 165
rect 1034 85 1084 131
rect 1160 219 1301 253
rect 1160 176 1196 219
rect 1335 185 1369 464
rect 1403 340 1447 356
rect 1403 306 1408 340
rect 1442 306 1447 340
rect 1403 221 1447 306
rect 1481 309 1515 464
rect 1681 430 1697 464
rect 1549 424 1607 430
rect 1549 414 1567 424
rect 1549 380 1555 414
rect 1601 390 1607 424
rect 1589 380 1607 390
rect 1549 364 1607 380
rect 1647 393 1697 430
rect 1681 359 1697 393
rect 1647 343 1697 359
rect 1737 535 1787 551
rect 1771 501 1787 535
rect 1737 464 1787 501
rect 1771 430 1787 464
rect 1737 393 1787 430
rect 1771 359 1787 393
rect 1481 299 1654 309
rect 1481 265 1604 299
rect 1638 265 1654 299
rect 1737 283 1787 359
rect 1821 535 2019 551
rect 1821 501 1892 535
rect 1926 501 2019 535
rect 2061 548 2078 582
rect 2112 548 2130 582
rect 2274 580 2363 649
rect 2061 532 2130 548
rect 2171 548 2237 577
rect 1821 485 2019 501
rect 2171 514 2187 548
rect 2221 514 2237 548
rect 2274 546 2290 580
rect 2324 546 2363 580
rect 2274 539 2363 546
rect 2171 498 2237 514
rect 2317 512 2363 539
rect 1821 481 1865 485
rect 1821 447 1827 481
rect 1861 447 1865 481
rect 1821 401 1865 447
rect 1821 367 1827 401
rect 1861 367 1865 401
rect 1821 351 1865 367
rect 1901 430 1951 446
rect 1901 396 1917 430
rect 1901 315 1951 396
rect 1481 255 1654 265
rect 1688 249 1787 283
rect 1821 269 1951 315
rect 1985 287 2019 485
rect 2053 464 2281 498
rect 2053 380 2105 464
rect 2053 346 2055 380
rect 2089 346 2105 380
rect 2053 330 2105 346
rect 2139 424 2213 430
rect 2139 390 2143 424
rect 2177 390 2213 424
rect 2139 386 2213 390
rect 2139 352 2163 386
rect 2197 352 2213 386
rect 2139 337 2213 352
rect 2247 360 2281 464
rect 2317 478 2322 512
rect 2356 478 2363 512
rect 2317 444 2363 478
rect 2317 410 2322 444
rect 2356 410 2363 444
rect 2317 394 2363 410
rect 2403 580 2469 596
rect 2403 546 2413 580
rect 2447 546 2469 580
rect 2403 500 2469 546
rect 2403 466 2413 500
rect 2447 466 2469 500
rect 2403 428 2469 466
rect 2403 394 2413 428
rect 2447 394 2469 428
rect 2247 326 2369 360
rect 1985 271 2285 287
rect 1688 221 1722 249
rect 1403 187 1722 221
rect 1821 231 1887 269
rect 1985 237 2235 271
rect 2269 237 2285 271
rect 1985 235 2285 237
rect 1821 215 1837 231
rect 1194 142 1196 176
rect 1160 119 1196 142
rect 1230 169 1369 185
rect 1230 135 1246 169
rect 1280 135 1369 169
rect 1656 179 1722 187
rect 1230 119 1369 135
rect 1403 119 1622 153
rect 1656 145 1672 179
rect 1706 145 1722 179
rect 1656 119 1722 145
rect 1756 197 1837 215
rect 1871 197 1887 231
rect 1756 181 1887 197
rect 1921 201 2285 235
rect 1403 85 1437 119
rect 1588 85 1622 119
rect 1756 85 1790 181
rect 1921 147 1955 201
rect 1034 51 1437 85
rect 1488 51 1504 85
rect 1538 51 1554 85
rect 1588 51 1790 85
rect 1827 131 1955 147
rect 1827 97 1857 131
rect 1891 97 1955 131
rect 1827 81 1955 97
rect 2033 133 2099 152
rect 2335 150 2369 326
rect 2033 99 2049 133
rect 2083 99 2099 133
rect 1488 17 1554 51
rect 2033 17 2099 99
rect 2191 127 2369 150
rect 2191 93 2207 127
rect 2241 116 2369 127
rect 2403 210 2469 394
rect 2403 176 2419 210
rect 2453 176 2469 210
rect 2403 120 2469 176
rect 2241 93 2257 116
rect 2191 70 2257 93
rect 2403 86 2419 120
rect 2453 86 2469 120
rect 2514 580 2571 596
rect 2514 546 2521 580
rect 2555 546 2571 580
rect 2514 470 2571 546
rect 2514 436 2521 470
rect 2555 436 2571 470
rect 2514 326 2571 436
rect 2609 580 2665 649
rect 2609 546 2618 580
rect 2652 546 2665 580
rect 2609 497 2665 546
rect 2609 463 2618 497
rect 2652 463 2665 497
rect 2609 414 2665 463
rect 2609 380 2625 414
rect 2659 380 2665 414
rect 2609 364 2665 380
rect 2711 580 2767 596
rect 2711 546 2715 580
rect 2749 546 2767 580
rect 2711 497 2767 546
rect 2711 463 2715 497
rect 2749 463 2767 497
rect 2711 414 2767 463
rect 2711 380 2715 414
rect 2749 380 2767 414
rect 2711 364 2767 380
rect 2514 310 2697 326
rect 2514 276 2659 310
rect 2693 276 2697 310
rect 2514 260 2697 276
rect 2514 146 2571 260
rect 2733 226 2767 364
rect 2514 112 2526 146
rect 2560 112 2571 146
rect 2514 91 2571 112
rect 2624 210 2658 226
rect 2624 120 2658 176
rect 2302 48 2318 82
rect 2352 48 2368 82
rect 2403 70 2469 86
rect 2302 17 2368 48
rect 2624 17 2658 86
rect 2694 210 2767 226
rect 2694 176 2710 210
rect 2744 176 2767 210
rect 2694 120 2767 176
rect 2694 86 2710 120
rect 2744 86 2767 120
rect 2694 70 2767 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 799 414 833 424
rect 799 390 807 414
rect 807 390 833 414
rect 1567 414 1601 424
rect 1567 390 1589 414
rect 1589 390 1601 414
rect 2143 390 2177 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
<< metal1 >>
rect 0 683 2784 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 0 617 2784 649
rect 787 424 845 430
rect 787 390 799 424
rect 833 421 845 424
rect 1555 424 1613 430
rect 1555 421 1567 424
rect 833 393 1567 421
rect 833 390 845 393
rect 787 384 845 390
rect 1555 390 1567 393
rect 1601 421 1613 424
rect 2131 424 2189 430
rect 2131 421 2143 424
rect 1601 393 2143 421
rect 1601 390 1613 393
rect 1555 384 1613 390
rect 2131 390 2143 393
rect 2177 390 2189 424
rect 2131 384 2189 390
rect 0 17 2784 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
rect 0 -49 2784 -17
<< labels >>
flabel pwell s 0 0 2784 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nwell s 0 617 2784 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
rlabel comment s 0 0 0 0 4 sdfrbp_1
flabel comment s 1498 630 1498 630 0 FreeSans 300 0 0 0 no_jumper_check
flabel comment s 1102 36 1102 36 0 FreeSans 300 0 0 0 no_jumper_check
flabel metal1 s 2143 390 2177 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew
flabel metal1 s 0 617 2784 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 2784 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 2431 390 2465 424 0 FreeSans 340 0 0 0 Q_N
port 11 nsew
flabel corelocali s 2431 464 2465 498 0 FreeSans 340 0 0 0 Q_N
port 11 nsew
flabel corelocali s 2431 538 2465 572 0 FreeSans 340 0 0 0 Q_N
port 11 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 799 242 833 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 SCD
port 4 nsew
flabel corelocali s 607 390 641 424 0 FreeSans 340 0 0 0 SCD
port 4 nsew
flabel corelocali s 319 168 353 202 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 2719 168 2753 202 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2719 390 2753 424 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2719 464 2753 498 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2719 538 2753 572 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2719 94 2753 128 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2431 94 2465 128 0 FreeSans 340 0 0 0 Q_N
port 11 nsew
flabel corelocali s 2431 168 2465 202 0 FreeSans 340 0 0 0 Q_N
port 11 nsew
flabel corelocali s 2431 242 2465 276 0 FreeSans 340 0 0 0 Q_N
port 11 nsew
flabel corelocali s 2431 316 2465 350 0 FreeSans 340 0 0 0 Q_N
port 11 nsew
<< properties >>
string FIXED_BBOX 0 0 2784 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1011134
string GDS_START 989280
<< end >>
