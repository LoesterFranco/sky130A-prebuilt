magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 229 401 281 493
rect 421 401 473 493
rect 229 367 473 401
rect 85 151 165 265
rect 421 330 473 367
rect 421 283 582 330
rect 482 181 582 283
rect 210 147 582 181
rect 210 69 281 147
rect 421 69 473 147
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 17 333 79 493
rect 123 367 185 527
rect 325 435 376 527
rect 509 369 575 527
rect 17 299 243 333
rect 17 117 51 299
rect 199 249 243 299
rect 199 215 448 249
rect 17 51 77 117
rect 121 17 176 113
rect 325 17 376 113
rect 517 17 573 113
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 85 151 165 265 6 A
port 1 nsew signal input
rlabel locali s 482 181 582 283 6 X
port 2 nsew signal output
rlabel locali s 421 401 473 493 6 X
port 2 nsew signal output
rlabel locali s 421 330 473 367 6 X
port 2 nsew signal output
rlabel locali s 421 283 582 330 6 X
port 2 nsew signal output
rlabel locali s 421 69 473 147 6 X
port 2 nsew signal output
rlabel locali s 229 401 281 493 6 X
port 2 nsew signal output
rlabel locali s 229 367 473 401 6 X
port 2 nsew signal output
rlabel locali s 210 147 582 181 6 X
port 2 nsew signal output
rlabel locali s 210 69 281 147 6 X
port 2 nsew signal output
rlabel metal1 s 0 -48 644 48 8 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 4 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1770928
string GDS_START 1765484
<< end >>
