magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 1326 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 112 47 142 177
rect 206 47 236 177
rect 300 47 330 177
rect 394 47 424 177
rect 488 47 518 177
rect 582 47 612 177
rect 676 47 706 177
rect 770 47 800 177
rect 864 47 894 177
rect 958 47 988 177
rect 1052 47 1082 177
rect 1156 47 1186 177
<< pmoshvt >>
rect 114 297 150 497
rect 208 297 244 497
rect 302 297 338 497
rect 396 297 432 497
rect 490 297 526 497
rect 584 297 620 497
rect 678 297 714 497
rect 772 297 808 497
rect 866 297 902 497
rect 960 297 996 497
rect 1054 297 1090 497
rect 1148 297 1184 497
<< ndiff >>
rect 60 93 112 177
rect 60 59 68 93
rect 102 59 112 93
rect 60 47 112 59
rect 142 161 206 177
rect 142 127 162 161
rect 196 127 206 161
rect 142 93 206 127
rect 142 59 162 93
rect 196 59 206 93
rect 142 47 206 59
rect 236 93 300 177
rect 236 59 256 93
rect 290 59 300 93
rect 236 47 300 59
rect 330 161 394 177
rect 330 127 350 161
rect 384 127 394 161
rect 330 93 394 127
rect 330 59 350 93
rect 384 59 394 93
rect 330 47 394 59
rect 424 93 488 177
rect 424 59 444 93
rect 478 59 488 93
rect 424 47 488 59
rect 518 161 582 177
rect 518 127 538 161
rect 572 127 582 161
rect 518 93 582 127
rect 518 59 538 93
rect 572 59 582 93
rect 518 47 582 59
rect 612 93 676 177
rect 612 59 632 93
rect 666 59 676 93
rect 612 47 676 59
rect 706 161 770 177
rect 706 127 726 161
rect 760 127 770 161
rect 706 93 770 127
rect 706 59 726 93
rect 760 59 770 93
rect 706 47 770 59
rect 800 93 864 177
rect 800 59 820 93
rect 854 59 864 93
rect 800 47 864 59
rect 894 161 958 177
rect 894 127 914 161
rect 948 127 958 161
rect 894 93 958 127
rect 894 59 914 93
rect 948 59 958 93
rect 894 47 958 59
rect 988 93 1052 177
rect 988 59 1008 93
rect 1042 59 1052 93
rect 988 47 1052 59
rect 1082 161 1156 177
rect 1082 127 1102 161
rect 1136 127 1156 161
rect 1082 93 1156 127
rect 1082 59 1102 93
rect 1136 59 1156 93
rect 1082 47 1156 59
rect 1186 93 1240 177
rect 1186 59 1196 93
rect 1230 59 1240 93
rect 1186 47 1240 59
<< pdiff >>
rect 60 485 114 497
rect 60 451 68 485
rect 102 451 114 485
rect 60 417 114 451
rect 60 383 68 417
rect 102 383 114 417
rect 60 297 114 383
rect 150 485 208 497
rect 150 451 162 485
rect 196 451 208 485
rect 150 417 208 451
rect 150 383 162 417
rect 196 383 208 417
rect 150 349 208 383
rect 150 315 162 349
rect 196 315 208 349
rect 150 297 208 315
rect 244 485 302 497
rect 244 451 256 485
rect 290 451 302 485
rect 244 417 302 451
rect 244 383 256 417
rect 290 383 302 417
rect 244 297 302 383
rect 338 485 396 497
rect 338 451 350 485
rect 384 451 396 485
rect 338 417 396 451
rect 338 383 350 417
rect 384 383 396 417
rect 338 349 396 383
rect 338 315 350 349
rect 384 315 396 349
rect 338 297 396 315
rect 432 485 490 497
rect 432 451 444 485
rect 478 451 490 485
rect 432 417 490 451
rect 432 383 444 417
rect 478 383 490 417
rect 432 297 490 383
rect 526 485 584 497
rect 526 451 538 485
rect 572 451 584 485
rect 526 417 584 451
rect 526 383 538 417
rect 572 383 584 417
rect 526 349 584 383
rect 526 315 538 349
rect 572 315 584 349
rect 526 297 584 315
rect 620 485 678 497
rect 620 451 632 485
rect 666 451 678 485
rect 620 417 678 451
rect 620 383 632 417
rect 666 383 678 417
rect 620 297 678 383
rect 714 485 772 497
rect 714 451 726 485
rect 760 451 772 485
rect 714 417 772 451
rect 714 383 726 417
rect 760 383 772 417
rect 714 349 772 383
rect 714 315 726 349
rect 760 315 772 349
rect 714 297 772 315
rect 808 485 866 497
rect 808 451 820 485
rect 854 451 866 485
rect 808 417 866 451
rect 808 383 820 417
rect 854 383 866 417
rect 808 297 866 383
rect 902 485 960 497
rect 902 451 914 485
rect 948 451 960 485
rect 902 417 960 451
rect 902 383 914 417
rect 948 383 960 417
rect 902 349 960 383
rect 902 315 914 349
rect 948 315 960 349
rect 902 297 960 315
rect 996 485 1054 497
rect 996 451 1008 485
rect 1042 451 1054 485
rect 996 417 1054 451
rect 996 383 1008 417
rect 1042 383 1054 417
rect 996 297 1054 383
rect 1090 485 1148 497
rect 1090 451 1102 485
rect 1136 451 1148 485
rect 1090 417 1148 451
rect 1090 383 1102 417
rect 1136 383 1148 417
rect 1090 349 1148 383
rect 1090 315 1102 349
rect 1136 315 1148 349
rect 1090 297 1148 315
rect 1184 485 1240 497
rect 1184 451 1196 485
rect 1230 451 1240 485
rect 1184 417 1240 451
rect 1184 383 1196 417
rect 1230 383 1240 417
rect 1184 297 1240 383
<< ndiffc >>
rect 68 59 102 93
rect 162 127 196 161
rect 162 59 196 93
rect 256 59 290 93
rect 350 127 384 161
rect 350 59 384 93
rect 444 59 478 93
rect 538 127 572 161
rect 538 59 572 93
rect 632 59 666 93
rect 726 127 760 161
rect 726 59 760 93
rect 820 59 854 93
rect 914 127 948 161
rect 914 59 948 93
rect 1008 59 1042 93
rect 1102 127 1136 161
rect 1102 59 1136 93
rect 1196 59 1230 93
<< pdiffc >>
rect 68 451 102 485
rect 68 383 102 417
rect 162 451 196 485
rect 162 383 196 417
rect 162 315 196 349
rect 256 451 290 485
rect 256 383 290 417
rect 350 451 384 485
rect 350 383 384 417
rect 350 315 384 349
rect 444 451 478 485
rect 444 383 478 417
rect 538 451 572 485
rect 538 383 572 417
rect 538 315 572 349
rect 632 451 666 485
rect 632 383 666 417
rect 726 451 760 485
rect 726 383 760 417
rect 726 315 760 349
rect 820 451 854 485
rect 820 383 854 417
rect 914 451 948 485
rect 914 383 948 417
rect 914 315 948 349
rect 1008 451 1042 485
rect 1008 383 1042 417
rect 1102 451 1136 485
rect 1102 383 1136 417
rect 1102 315 1136 349
rect 1196 451 1230 485
rect 1196 383 1230 417
<< poly >>
rect 114 497 150 523
rect 208 497 244 523
rect 302 497 338 523
rect 396 497 432 523
rect 490 497 526 523
rect 584 497 620 523
rect 678 497 714 523
rect 772 497 808 523
rect 866 497 902 523
rect 960 497 996 523
rect 1054 497 1090 523
rect 1148 497 1184 523
rect 114 282 150 297
rect 208 282 244 297
rect 302 282 338 297
rect 396 282 432 297
rect 490 282 526 297
rect 584 282 620 297
rect 678 282 714 297
rect 772 282 808 297
rect 866 282 902 297
rect 960 282 996 297
rect 1054 282 1090 297
rect 1148 282 1184 297
rect 112 265 152 282
rect 206 265 246 282
rect 300 265 340 282
rect 394 265 434 282
rect 488 265 528 282
rect 582 265 622 282
rect 676 265 716 282
rect 770 265 810 282
rect 864 265 904 282
rect 958 265 998 282
rect 1052 265 1092 282
rect 1146 265 1186 282
rect 112 249 1186 265
rect 112 215 162 249
rect 196 215 256 249
rect 290 215 350 249
rect 384 215 444 249
rect 478 215 538 249
rect 572 215 632 249
rect 666 215 726 249
rect 760 215 820 249
rect 854 215 914 249
rect 948 215 1008 249
rect 1042 215 1102 249
rect 1136 215 1186 249
rect 112 199 1186 215
rect 112 177 142 199
rect 206 177 236 199
rect 300 177 330 199
rect 394 177 424 199
rect 488 177 518 199
rect 582 177 612 199
rect 676 177 706 199
rect 770 177 800 199
rect 864 177 894 199
rect 958 177 988 199
rect 1052 177 1082 199
rect 1156 177 1186 199
rect 112 21 142 47
rect 206 21 236 47
rect 300 21 330 47
rect 394 21 424 47
rect 488 21 518 47
rect 582 21 612 47
rect 676 21 706 47
rect 770 21 800 47
rect 864 21 894 47
rect 958 21 988 47
rect 1052 21 1082 47
rect 1156 21 1186 47
<< polycont >>
rect 162 215 196 249
rect 256 215 290 249
rect 350 215 384 249
rect 444 215 478 249
rect 538 215 572 249
rect 632 215 666 249
rect 726 215 760 249
rect 820 215 854 249
rect 914 215 948 249
rect 1008 215 1042 249
rect 1102 215 1136 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 51 485 102 527
rect 51 451 68 485
rect 51 417 102 451
rect 51 383 68 417
rect 51 367 102 383
rect 136 485 212 493
rect 136 451 162 485
rect 196 451 212 485
rect 136 417 212 451
rect 136 383 162 417
rect 196 383 212 417
rect 136 349 212 383
rect 256 485 290 527
rect 256 417 290 451
rect 256 367 290 383
rect 324 485 400 493
rect 324 451 350 485
rect 384 451 400 485
rect 324 417 400 451
rect 324 383 350 417
rect 384 383 400 417
rect 136 333 162 349
rect 17 315 162 333
rect 196 333 212 349
rect 324 349 400 383
rect 444 485 478 527
rect 444 417 478 451
rect 444 367 478 383
rect 512 485 588 493
rect 512 451 538 485
rect 572 451 588 485
rect 512 417 588 451
rect 512 383 538 417
rect 572 383 588 417
rect 324 333 350 349
rect 196 315 350 333
rect 384 333 400 349
rect 512 349 588 383
rect 632 485 666 527
rect 632 417 666 451
rect 632 367 666 383
rect 700 485 776 493
rect 700 451 726 485
rect 760 451 776 485
rect 700 417 776 451
rect 700 383 726 417
rect 760 383 776 417
rect 512 333 538 349
rect 384 315 538 333
rect 572 333 588 349
rect 700 349 776 383
rect 820 485 854 527
rect 820 417 854 451
rect 820 367 854 383
rect 888 485 964 493
rect 888 451 914 485
rect 948 451 964 485
rect 888 417 964 451
rect 888 383 914 417
rect 948 383 964 417
rect 700 333 726 349
rect 572 315 726 333
rect 760 333 776 349
rect 888 349 964 383
rect 1008 485 1042 527
rect 1008 417 1042 451
rect 1008 367 1042 383
rect 1076 485 1152 493
rect 1076 451 1102 485
rect 1136 451 1152 485
rect 1076 417 1152 451
rect 1076 383 1102 417
rect 1136 383 1152 417
rect 888 333 914 349
rect 760 315 914 333
rect 948 333 964 349
rect 1076 349 1152 383
rect 1195 485 1246 527
rect 1195 451 1196 485
rect 1230 451 1246 485
rect 1195 417 1246 451
rect 1195 383 1196 417
rect 1230 383 1246 417
rect 1195 367 1246 383
rect 1076 333 1102 349
rect 948 315 1102 333
rect 1136 333 1152 349
rect 1136 315 1264 333
rect 17 299 1264 315
rect 17 181 102 299
rect 136 249 1160 265
rect 136 215 162 249
rect 196 215 256 249
rect 290 215 350 249
rect 384 215 444 249
rect 478 215 538 249
rect 572 215 632 249
rect 666 215 726 249
rect 760 215 820 249
rect 854 215 914 249
rect 948 215 1008 249
rect 1042 215 1102 249
rect 1136 215 1160 249
rect 1194 181 1264 299
rect 17 161 1264 181
rect 17 143 162 161
rect 136 127 162 143
rect 196 143 350 161
rect 196 127 212 143
rect 51 93 102 109
rect 51 59 68 93
rect 51 17 102 59
rect 136 93 212 127
rect 324 127 350 143
rect 384 143 538 161
rect 384 127 400 143
rect 136 59 162 93
rect 196 59 212 93
rect 136 51 212 59
rect 256 93 290 109
rect 256 17 290 59
rect 324 93 400 127
rect 512 127 538 143
rect 572 143 726 161
rect 572 127 588 143
rect 324 59 350 93
rect 384 59 400 93
rect 324 51 400 59
rect 444 93 478 109
rect 444 17 478 59
rect 512 93 588 127
rect 700 127 726 143
rect 760 143 914 161
rect 760 127 776 143
rect 512 59 538 93
rect 572 59 588 93
rect 512 51 588 59
rect 632 93 666 109
rect 632 17 666 59
rect 700 93 776 127
rect 888 127 914 143
rect 948 143 1102 161
rect 948 127 964 143
rect 700 59 726 93
rect 760 59 776 93
rect 700 51 776 59
rect 820 93 854 109
rect 820 17 854 59
rect 888 93 964 127
rect 1076 127 1102 143
rect 1136 143 1264 161
rect 1136 127 1152 143
rect 888 59 914 93
rect 948 59 964 93
rect 888 51 964 59
rect 1008 93 1042 109
rect 1008 17 1042 59
rect 1076 93 1152 127
rect 1076 59 1102 93
rect 1136 59 1152 93
rect 1076 51 1152 59
rect 1192 93 1246 109
rect 1192 59 1196 93
rect 1230 59 1246 93
rect 1192 17 1246 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
flabel corelocali s 213 221 257 255 0 FreeSans 250 0 0 0 A
port 1 nsew
flabel corelocali s 305 221 349 255 0 FreeSans 250 0 0 0 A
port 1 nsew
flabel corelocali s 397 221 431 255 0 FreeSans 250 0 0 0 A
port 1 nsew
flabel corelocali s 490 221 524 255 0 FreeSans 250 0 0 0 A
port 1 nsew
flabel corelocali s 584 221 618 255 0 FreeSans 250 0 0 0 A
port 1 nsew
flabel corelocali s 676 221 710 255 0 FreeSans 250 0 0 0 A
port 1 nsew
flabel corelocali s 1218 221 1252 255 0 FreeSans 250 0 0 0 Y
port 6 nsew
flabel corelocali s 29 221 63 255 0 FreeSans 250 0 0 0 Y
port 6 nsew
flabel corelocali s 829 221 863 255 0 FreeSans 250 0 0 0 A
port 1 nsew
flabel corelocali s 931 221 965 255 0 FreeSans 250 0 0 0 A
port 1 nsew
flabel corelocali s 1017 221 1051 255 0 FreeSans 250 0 0 0 A
port 1 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 1288 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2085522
string GDS_START 2074868
<< end >>
