magic
tech sky130A
magscale 1 2
timestamp 1604502741
<< locali >>
rect 21 236 87 310
rect 215 270 281 430
rect 315 412 691 478
rect 315 226 349 412
rect 383 270 455 356
rect 793 290 869 356
rect 289 210 355 226
rect 289 176 647 210
rect 289 70 355 176
rect 572 70 647 176
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 130 580 269 649
rect 23 512 759 546
rect 23 364 155 512
rect 121 202 155 364
rect 725 378 759 512
rect 793 420 837 649
rect 871 420 937 596
rect 497 344 759 378
rect 497 270 563 344
rect 614 252 748 310
rect 903 252 937 420
rect 614 244 937 252
rect 23 136 155 202
rect 189 17 255 226
rect 714 218 937 244
rect 389 17 538 136
rect 681 17 835 184
rect 871 108 937 218
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
rlabel locali s 215 270 281 430 6 A
port 1 nsew signal input
rlabel locali s 383 270 455 356 6 B
port 2 nsew signal input
rlabel locali s 21 236 87 310 6 C_N
port 3 nsew signal input
rlabel locali s 793 290 869 356 6 D_N
port 4 nsew signal input
rlabel locali s 572 70 647 176 6 Y
port 5 nsew signal output
rlabel locali s 315 412 691 478 6 Y
port 5 nsew signal output
rlabel locali s 315 226 349 412 6 Y
port 5 nsew signal output
rlabel locali s 289 210 355 226 6 Y
port 5 nsew signal output
rlabel locali s 289 176 647 210 6 Y
port 5 nsew signal output
rlabel locali s 289 70 355 176 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -49 960 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 960 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1581160
string GDS_START 1573906
<< end >>
