magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< obsli1 >>
rect 21160 1071 45080 1105
rect 21214 966 21272 1071
rect 21314 923 21364 1032
rect 21398 966 21456 1071
rect 21557 1003 21963 1037
rect 21557 934 21607 1003
rect 21177 823 21296 889
rect 21330 875 21364 923
rect 21641 875 21707 969
rect 21741 934 21775 1003
rect 21809 911 21875 969
rect 21909 945 21963 1003
rect 21997 979 22047 1071
rect 22081 945 22147 1037
rect 22181 979 22235 1071
rect 22269 945 22335 1037
rect 21909 911 22335 945
rect 22369 911 22435 1071
rect 22469 945 22535 1037
rect 22569 979 22623 1071
rect 22657 945 22723 1037
rect 22757 979 22807 1071
rect 22841 1003 23247 1037
rect 22841 945 22895 1003
rect 22469 911 22895 945
rect 22929 911 22995 969
rect 23029 934 23063 1003
rect 21809 875 21855 911
rect 21330 809 21567 875
rect 21601 815 21855 875
rect 22091 823 22369 877
rect 22435 823 22713 877
rect 22949 875 22995 911
rect 23097 875 23163 969
rect 23197 934 23247 1003
rect 23348 966 23406 1071
rect 23440 923 23490 1032
rect 23532 966 23590 1071
rect 23698 966 23756 1071
rect 23798 923 23848 1032
rect 23882 966 23940 1071
rect 24041 1003 24447 1037
rect 24041 934 24091 1003
rect 23440 875 23474 923
rect 21330 767 21364 809
rect 21204 561 21264 767
rect 21298 595 21364 767
rect 21403 561 21458 767
rect 21507 595 21567 775
rect 0 527 21567 561
rect 18 299 85 493
rect 129 299 163 527
rect 214 459 683 493
rect 18 51 69 299
rect 214 265 254 459
rect 103 165 137 265
rect 199 199 254 265
rect 288 391 577 425
rect 288 165 322 391
rect 103 131 322 165
rect 356 323 615 357
rect 356 162 390 323
rect 287 124 322 131
rect 103 17 179 97
rect 287 51 391 124
rect 458 51 523 283
rect 557 51 615 323
rect 649 326 683 459
rect 717 367 763 527
rect 797 367 877 493
rect 649 288 799 326
rect 665 173 699 237
rect 761 211 799 288
rect 843 173 877 367
rect 947 299 996 527
rect 1031 299 1099 493
rect 1135 299 1185 527
rect 1226 459 1695 493
rect 665 139 877 173
rect 650 17 753 105
rect 807 51 856 139
rect 947 17 997 131
rect 1031 51 1081 299
rect 1226 265 1266 459
rect 1115 165 1149 265
rect 1211 199 1266 265
rect 1300 391 1589 425
rect 1300 165 1334 391
rect 1115 131 1334 165
rect 1368 323 1627 357
rect 1368 162 1402 323
rect 1299 124 1334 131
rect 1115 17 1191 97
rect 1299 51 1436 124
rect 1470 51 1535 283
rect 1569 51 1627 323
rect 1661 326 1695 459
rect 1729 367 1775 527
rect 1809 367 1889 493
rect 1661 288 1811 326
rect 1677 173 1711 237
rect 1773 211 1811 288
rect 1855 173 1889 367
rect 1959 299 2011 527
rect 2045 299 2111 493
rect 2145 299 2193 527
rect 2227 299 2299 493
rect 2333 299 2388 527
rect 2422 459 2891 493
rect 1677 139 1889 173
rect 2050 265 2102 299
rect 2227 265 2281 299
rect 2422 265 2462 459
rect 2050 213 2281 265
rect 1662 17 1765 105
rect 1819 51 1868 139
rect 1967 17 2016 131
rect 2050 51 2102 213
rect 2143 17 2193 131
rect 2227 51 2281 213
rect 2315 165 2349 265
rect 2407 199 2462 265
rect 2496 391 2785 425
rect 2496 165 2530 391
rect 2315 131 2530 165
rect 2564 323 2823 357
rect 2564 162 2598 323
rect 2495 124 2530 131
rect 2315 17 2387 97
rect 2495 51 2632 124
rect 2666 51 2731 283
rect 2765 51 2823 323
rect 2857 326 2891 459
rect 2925 367 2971 527
rect 3005 367 3085 493
rect 2857 288 3007 326
rect 2873 173 2907 237
rect 2969 211 3007 288
rect 3051 173 3085 367
rect 3147 299 3213 527
rect 3346 397 3412 493
rect 3308 361 3412 397
rect 3308 351 3387 361
rect 3195 211 3274 265
rect 2873 139 3085 173
rect 2858 17 2961 105
rect 3015 51 3064 139
rect 3154 17 3206 177
rect 3240 125 3274 211
rect 3308 201 3342 351
rect 3450 327 3516 493
rect 3420 301 3516 327
rect 3376 293 3516 301
rect 3561 293 3621 527
rect 3660 327 3726 493
rect 3764 397 3830 493
rect 3764 361 3868 397
rect 3789 351 3868 361
rect 3660 301 3756 327
rect 3660 293 3800 301
rect 3376 235 3454 293
rect 3308 167 3386 201
rect 3240 79 3295 125
rect 3337 66 3386 167
rect 3420 151 3454 235
rect 3489 189 3559 259
rect 3617 189 3687 259
rect 3722 235 3800 293
rect 3722 151 3756 235
rect 3834 201 3868 351
rect 3963 299 4041 527
rect 4174 397 4240 493
rect 4136 361 4240 397
rect 4136 351 4215 361
rect 3420 117 3508 151
rect 3458 66 3508 117
rect 3555 17 3621 132
rect 3668 117 3756 151
rect 3790 167 3868 201
rect 3902 211 3981 265
rect 4023 211 4102 265
rect 3668 66 3718 117
rect 3790 66 3839 167
rect 3902 125 3936 211
rect 3881 79 3936 125
rect 3970 17 4034 177
rect 4068 125 4102 211
rect 4136 201 4170 351
rect 4278 327 4344 493
rect 4248 301 4344 327
rect 4204 293 4344 301
rect 4383 293 4443 527
rect 4488 327 4554 493
rect 4592 397 4658 493
rect 4592 361 4696 397
rect 4617 351 4696 361
rect 4488 301 4584 327
rect 4488 293 4628 301
rect 4204 235 4282 293
rect 4136 167 4214 201
rect 4068 79 4123 125
rect 4165 66 4214 167
rect 4248 151 4282 235
rect 4317 189 4387 259
rect 4445 189 4515 259
rect 4550 235 4628 293
rect 4550 151 4584 235
rect 4662 201 4696 351
rect 4791 299 4857 527
rect 4895 442 4961 493
rect 4895 333 4955 442
rect 4995 421 5055 527
rect 4989 367 5055 421
rect 5099 459 5332 493
rect 5099 333 5133 459
rect 5169 351 5255 425
rect 4895 299 5133 333
rect 4248 117 4336 151
rect 4286 66 4336 117
rect 4383 17 4449 132
rect 4496 117 4584 151
rect 4618 167 4696 201
rect 4730 211 4809 265
rect 4895 211 5059 265
rect 4496 66 4546 117
rect 4618 66 4667 167
rect 4730 125 4764 211
rect 5082 177 5143 185
rect 5193 177 5227 351
rect 5298 329 5332 459
rect 5386 327 5452 493
rect 5366 295 5452 327
rect 5296 293 5452 295
rect 5487 293 5553 527
rect 5588 327 5654 493
rect 5708 459 5941 493
rect 5708 329 5742 459
rect 5785 351 5871 425
rect 5588 295 5674 327
rect 5588 293 5744 295
rect 5296 261 5400 293
rect 5640 261 5744 293
rect 5296 241 5379 261
rect 4709 79 4764 125
rect 4798 17 4850 177
rect 4905 143 5143 177
rect 4905 51 4971 143
rect 5005 17 5048 109
rect 5082 85 5143 143
rect 5177 119 5243 177
rect 5277 85 5311 154
rect 5345 151 5379 241
rect 5434 205 5501 259
rect 5539 205 5606 259
rect 5661 241 5744 261
rect 5661 151 5695 241
rect 5813 177 5847 351
rect 5907 333 5941 459
rect 5985 421 6045 527
rect 6079 442 6145 493
rect 5985 367 6051 421
rect 6085 333 6145 442
rect 5907 299 6145 333
rect 6183 442 6249 493
rect 6183 333 6243 442
rect 6283 421 6343 527
rect 6277 367 6343 421
rect 6387 459 6620 493
rect 6387 333 6421 459
rect 6457 351 6543 425
rect 6183 299 6421 333
rect 5981 211 6145 265
rect 6183 211 6347 265
rect 5897 177 5958 185
rect 6370 177 6431 185
rect 6481 177 6515 351
rect 6586 329 6620 459
rect 6674 327 6740 493
rect 6654 295 6740 327
rect 6584 293 6740 295
rect 6775 293 6841 527
rect 6876 327 6942 493
rect 6996 459 7229 493
rect 6996 329 7030 459
rect 7073 351 7159 425
rect 6876 295 6962 327
rect 6876 293 7032 295
rect 6584 261 6688 293
rect 6928 261 7032 293
rect 6584 241 6667 261
rect 5345 117 5461 151
rect 5082 51 5311 85
rect 5411 66 5461 117
rect 5495 17 5545 132
rect 5579 117 5695 151
rect 5579 66 5629 117
rect 5729 85 5763 154
rect 5797 119 5863 177
rect 5897 143 6135 177
rect 5897 85 5958 143
rect 5729 51 5958 85
rect 5992 17 6035 109
rect 6069 51 6135 143
rect 6193 143 6431 177
rect 6193 51 6259 143
rect 6293 17 6336 109
rect 6370 85 6431 143
rect 6465 119 6531 177
rect 6565 85 6599 154
rect 6633 151 6667 241
rect 6722 205 6789 259
rect 6827 205 6894 259
rect 6949 241 7032 261
rect 6949 151 6983 241
rect 7101 177 7135 351
rect 7195 333 7229 459
rect 7273 421 7333 527
rect 7367 442 7433 493
rect 7273 367 7339 421
rect 7373 333 7433 442
rect 7195 299 7433 333
rect 7477 299 7531 527
rect 7565 333 7631 493
rect 7665 367 7719 527
rect 7753 333 7819 493
rect 7853 367 7907 527
rect 7951 459 8393 493
rect 7951 333 8011 459
rect 7565 299 8011 333
rect 8045 273 8111 425
rect 8145 307 8199 459
rect 8233 273 8299 425
rect 8333 313 8393 459
rect 8442 321 8497 527
rect 8536 321 8602 493
rect 8636 321 8696 527
rect 8784 321 8844 527
rect 8878 321 8944 493
rect 8983 321 9038 527
rect 9087 459 9529 493
rect 8536 279 8570 321
rect 7269 211 7433 265
rect 7531 211 7809 265
rect 8045 213 8299 273
rect 8333 213 8570 279
rect 8910 279 8944 321
rect 9087 313 9147 459
rect 7185 177 7246 185
rect 8045 177 8091 213
rect 6633 117 6749 151
rect 6370 51 6599 85
rect 6699 66 6749 117
rect 6783 17 6833 132
rect 6867 117 6983 151
rect 6867 66 6917 117
rect 7017 85 7051 154
rect 7085 119 7151 177
rect 7185 143 7423 177
rect 7185 85 7246 143
rect 7017 51 7246 85
rect 7280 17 7323 109
rect 7357 51 7423 143
rect 7481 17 7531 177
rect 7565 143 7991 177
rect 7565 51 7631 143
rect 7665 17 7719 109
rect 7753 51 7819 143
rect 7853 17 7903 109
rect 7937 85 7991 143
rect 8025 119 8091 177
rect 8125 85 8159 154
rect 8193 119 8259 213
rect 8536 165 8570 213
rect 8604 199 8723 265
rect 8757 199 8876 265
rect 8910 213 9147 279
rect 9181 273 9247 425
rect 9281 307 9335 459
rect 9369 273 9435 425
rect 9469 333 9529 459
rect 9573 367 9627 527
rect 9661 333 9727 493
rect 9761 367 9815 527
rect 9849 333 9915 493
rect 9469 299 9915 333
rect 9949 299 10003 527
rect 10053 299 10107 527
rect 10141 333 10207 493
rect 10241 367 10295 527
rect 10329 333 10395 493
rect 10429 367 10483 527
rect 10527 459 10969 493
rect 10527 333 10587 459
rect 10141 299 10587 333
rect 9181 213 9435 273
rect 10621 273 10687 425
rect 10721 307 10775 459
rect 10809 273 10875 425
rect 10909 313 10969 459
rect 11018 321 11073 527
rect 11112 321 11178 493
rect 11212 321 11272 527
rect 11360 321 11420 527
rect 11454 321 11520 493
rect 11559 321 11614 527
rect 11663 459 12105 493
rect 11112 279 11146 321
rect 8910 165 8944 213
rect 8293 85 8343 154
rect 7937 51 8343 85
rect 8444 17 8502 122
rect 8536 56 8586 165
rect 8628 17 8686 122
rect 8794 17 8852 122
rect 8894 56 8944 165
rect 8978 17 9036 122
rect 9137 85 9187 154
rect 9221 119 9287 213
rect 9389 177 9435 213
rect 9671 211 9949 265
rect 10107 211 10385 265
rect 10621 213 10875 273
rect 10909 213 11146 279
rect 11486 279 11520 321
rect 11663 313 11723 459
rect 10621 177 10667 213
rect 9321 85 9355 154
rect 9389 119 9455 177
rect 9489 143 9915 177
rect 9489 85 9543 143
rect 9137 51 9543 85
rect 9577 17 9627 109
rect 9661 51 9727 143
rect 9761 17 9815 109
rect 9849 51 9915 143
rect 9949 17 9999 177
rect 10057 17 10107 177
rect 10141 143 10567 177
rect 10141 51 10207 143
rect 10241 17 10295 109
rect 10329 51 10395 143
rect 10429 17 10479 109
rect 10513 85 10567 143
rect 10601 119 10667 177
rect 10701 85 10735 154
rect 10769 119 10835 213
rect 11112 165 11146 213
rect 11180 199 11299 265
rect 11333 199 11452 265
rect 11486 213 11723 279
rect 11757 273 11823 425
rect 11857 307 11911 459
rect 11945 273 12011 425
rect 12045 333 12105 459
rect 12149 367 12203 527
rect 12237 333 12303 493
rect 12337 367 12391 527
rect 12425 333 12491 493
rect 12045 299 12491 333
rect 12525 299 12579 527
rect 12623 299 12689 527
rect 12822 397 12888 493
rect 12784 361 12888 397
rect 12784 351 12863 361
rect 11757 213 12011 273
rect 11486 165 11520 213
rect 10869 85 10919 154
rect 10513 51 10919 85
rect 11020 17 11078 122
rect 11112 56 11162 165
rect 11204 17 11262 122
rect 11370 17 11428 122
rect 11470 56 11520 165
rect 11554 17 11612 122
rect 11713 85 11763 154
rect 11797 119 11863 213
rect 11965 177 12011 213
rect 12247 211 12525 265
rect 12671 211 12750 265
rect 11897 85 11931 154
rect 11965 119 12031 177
rect 12065 143 12491 177
rect 12065 85 12119 143
rect 11713 51 12119 85
rect 12153 17 12203 109
rect 12237 51 12303 143
rect 12337 17 12391 109
rect 12425 51 12491 143
rect 12525 17 12575 177
rect 12630 17 12682 177
rect 12716 125 12750 211
rect 12784 201 12818 351
rect 12926 327 12992 493
rect 12896 301 12992 327
rect 12852 293 12992 301
rect 13031 293 13097 527
rect 13136 327 13202 493
rect 13240 397 13306 493
rect 13240 361 13344 397
rect 13265 351 13344 361
rect 13136 301 13232 327
rect 13136 293 13276 301
rect 12852 235 12930 293
rect 12784 167 12862 201
rect 12716 79 12771 125
rect 12813 66 12862 167
rect 12896 151 12930 235
rect 12965 189 13045 259
rect 13083 189 13163 259
rect 13198 235 13276 293
rect 13198 151 13232 235
rect 13310 201 13344 351
rect 13439 299 13517 527
rect 13650 397 13716 493
rect 13612 361 13716 397
rect 13612 351 13691 361
rect 12896 117 12984 151
rect 12934 66 12984 117
rect 13031 17 13097 132
rect 13144 117 13232 151
rect 13266 167 13344 201
rect 13378 211 13457 265
rect 13499 211 13578 265
rect 13144 66 13194 117
rect 13266 66 13315 167
rect 13378 125 13412 211
rect 13357 79 13412 125
rect 13446 17 13510 177
rect 13544 125 13578 211
rect 13612 201 13646 351
rect 13754 327 13820 493
rect 13724 301 13820 327
rect 13680 293 13820 301
rect 13859 293 13925 527
rect 13964 327 14030 493
rect 14068 397 14134 493
rect 14068 361 14172 397
rect 14093 351 14172 361
rect 13964 301 14060 327
rect 13964 293 14104 301
rect 13680 235 13758 293
rect 13612 167 13690 201
rect 13544 79 13599 125
rect 13641 66 13690 167
rect 13724 151 13758 235
rect 13793 189 13873 259
rect 13911 189 13991 259
rect 14026 235 14104 293
rect 14026 151 14060 235
rect 14138 201 14172 351
rect 14267 299 14345 527
rect 14478 397 14544 493
rect 14440 361 14544 397
rect 14440 351 14519 361
rect 13724 117 13812 151
rect 13762 66 13812 117
rect 13859 17 13925 132
rect 13972 117 14060 151
rect 14094 167 14172 201
rect 14206 211 14285 265
rect 14327 211 14406 265
rect 13972 66 14022 117
rect 14094 66 14143 167
rect 14206 125 14240 211
rect 14185 79 14240 125
rect 14274 17 14338 177
rect 14372 125 14406 211
rect 14440 201 14474 351
rect 14582 327 14648 493
rect 14552 301 14648 327
rect 14508 293 14648 301
rect 14687 293 14753 527
rect 14792 327 14858 493
rect 14896 397 14962 493
rect 14896 361 15000 397
rect 14921 351 15000 361
rect 14792 301 14888 327
rect 14792 293 14932 301
rect 14508 235 14586 293
rect 14440 167 14518 201
rect 14372 79 14427 125
rect 14469 66 14518 167
rect 14552 151 14586 235
rect 14621 189 14701 259
rect 14739 189 14819 259
rect 14854 235 14932 293
rect 14854 151 14888 235
rect 14966 201 15000 351
rect 15095 299 15173 527
rect 15306 397 15372 493
rect 15268 361 15372 397
rect 15268 351 15347 361
rect 14552 117 14640 151
rect 14590 66 14640 117
rect 14687 17 14753 132
rect 14800 117 14888 151
rect 14922 167 15000 201
rect 15034 211 15113 265
rect 15155 211 15234 265
rect 14800 66 14850 117
rect 14922 66 14971 167
rect 15034 125 15068 211
rect 15013 79 15068 125
rect 15102 17 15166 177
rect 15200 125 15234 211
rect 15268 201 15302 351
rect 15410 327 15476 493
rect 15380 301 15476 327
rect 15336 293 15476 301
rect 15515 293 15581 527
rect 15620 327 15686 493
rect 15724 397 15790 493
rect 15724 361 15828 397
rect 15749 351 15828 361
rect 15620 301 15716 327
rect 15620 293 15760 301
rect 15336 235 15414 293
rect 15268 167 15346 201
rect 15200 79 15255 125
rect 15297 66 15346 167
rect 15380 151 15414 235
rect 15449 189 15529 259
rect 15567 189 15647 259
rect 15682 235 15760 293
rect 15682 151 15716 235
rect 15794 201 15828 351
rect 15923 299 15989 527
rect 16027 442 16093 493
rect 16027 333 16087 442
rect 16127 421 16187 527
rect 16121 367 16187 421
rect 16231 459 16464 493
rect 16231 333 16265 459
rect 16301 351 16387 425
rect 16027 299 16265 333
rect 15380 117 15468 151
rect 15418 66 15468 117
rect 15515 17 15581 132
rect 15628 117 15716 151
rect 15750 167 15828 201
rect 15862 211 15941 265
rect 16027 211 16191 265
rect 15628 66 15678 117
rect 15750 66 15799 167
rect 15862 125 15896 211
rect 16214 177 16275 185
rect 16325 177 16359 351
rect 16430 329 16464 459
rect 16518 327 16584 493
rect 16498 295 16584 327
rect 16428 293 16584 295
rect 16619 293 16685 527
rect 16720 327 16786 493
rect 16840 459 17073 493
rect 16840 329 16874 459
rect 16917 351 17003 425
rect 16720 295 16806 327
rect 16720 293 16876 295
rect 16428 261 16532 293
rect 16772 261 16876 293
rect 16428 241 16511 261
rect 15841 79 15896 125
rect 15930 17 15982 177
rect 16037 143 16275 177
rect 16037 51 16103 143
rect 16137 17 16180 109
rect 16214 85 16275 143
rect 16309 119 16375 177
rect 16409 85 16443 154
rect 16477 151 16511 241
rect 16566 205 16633 259
rect 16671 205 16738 259
rect 16793 241 16876 261
rect 16793 151 16827 241
rect 16945 177 16979 351
rect 17039 333 17073 459
rect 17117 421 17177 527
rect 17211 442 17277 493
rect 17117 367 17183 421
rect 17217 333 17277 442
rect 17039 299 17277 333
rect 17315 442 17381 493
rect 17315 333 17375 442
rect 17415 421 17475 527
rect 17409 367 17475 421
rect 17519 459 17752 493
rect 17519 333 17553 459
rect 17589 351 17675 425
rect 17315 299 17553 333
rect 17113 211 17277 265
rect 17315 211 17479 265
rect 17029 177 17090 185
rect 17502 177 17563 185
rect 17613 177 17647 351
rect 17718 329 17752 459
rect 17806 327 17872 493
rect 17786 295 17872 327
rect 17716 293 17872 295
rect 17907 293 17973 527
rect 18008 327 18074 493
rect 18128 459 18361 493
rect 18128 329 18162 459
rect 18205 351 18291 425
rect 18008 295 18094 327
rect 18008 293 18164 295
rect 17716 261 17820 293
rect 18060 261 18164 293
rect 17716 241 17799 261
rect 16477 117 16593 151
rect 16214 51 16443 85
rect 16543 66 16593 117
rect 16627 17 16677 132
rect 16711 117 16827 151
rect 16711 66 16761 117
rect 16861 85 16895 154
rect 16929 119 16995 177
rect 17029 143 17267 177
rect 17029 85 17090 143
rect 16861 51 17090 85
rect 17124 17 17167 109
rect 17201 51 17267 143
rect 17325 143 17563 177
rect 17325 51 17391 143
rect 17425 17 17468 109
rect 17502 85 17563 143
rect 17597 119 17663 177
rect 17697 85 17731 154
rect 17765 151 17799 241
rect 17854 205 17921 259
rect 17959 205 18026 259
rect 18081 241 18164 261
rect 18081 151 18115 241
rect 18233 177 18267 351
rect 18327 333 18361 459
rect 18405 421 18465 527
rect 18499 442 18565 493
rect 18405 367 18471 421
rect 18505 333 18565 442
rect 18327 299 18565 333
rect 18603 442 18669 493
rect 18603 333 18663 442
rect 18703 421 18763 527
rect 18697 367 18763 421
rect 18807 459 19040 493
rect 18807 333 18841 459
rect 18877 351 18963 425
rect 18603 299 18841 333
rect 18401 211 18565 265
rect 18603 211 18767 265
rect 18317 177 18378 185
rect 18790 177 18851 185
rect 18901 177 18935 351
rect 19006 329 19040 459
rect 19094 327 19160 493
rect 19074 295 19160 327
rect 19004 293 19160 295
rect 19195 293 19261 527
rect 19296 327 19362 493
rect 19416 459 19649 493
rect 19416 329 19450 459
rect 19493 351 19579 425
rect 19296 295 19382 327
rect 19296 293 19452 295
rect 19004 261 19108 293
rect 19348 261 19452 293
rect 19004 241 19087 261
rect 17765 117 17881 151
rect 17502 51 17731 85
rect 17831 66 17881 117
rect 17915 17 17965 132
rect 17999 117 18115 151
rect 17999 66 18049 117
rect 18149 85 18183 154
rect 18217 119 18283 177
rect 18317 143 18555 177
rect 18317 85 18378 143
rect 18149 51 18378 85
rect 18412 17 18455 109
rect 18489 51 18555 143
rect 18613 143 18851 177
rect 18613 51 18679 143
rect 18713 17 18756 109
rect 18790 85 18851 143
rect 18885 119 18951 177
rect 18985 85 19019 154
rect 19053 151 19087 241
rect 19142 205 19209 259
rect 19247 205 19314 259
rect 19369 241 19452 261
rect 19369 151 19403 241
rect 19521 177 19555 351
rect 19615 333 19649 459
rect 19693 421 19753 527
rect 19787 442 19853 493
rect 19693 367 19759 421
rect 19793 333 19853 442
rect 19615 299 19853 333
rect 19891 442 19957 493
rect 19891 333 19951 442
rect 19991 421 20051 527
rect 19985 367 20051 421
rect 20095 459 20328 493
rect 20095 333 20129 459
rect 20165 351 20251 425
rect 19891 299 20129 333
rect 19689 211 19853 265
rect 19891 211 20055 265
rect 19605 177 19666 185
rect 20078 177 20139 185
rect 20189 177 20223 351
rect 20294 329 20328 459
rect 20382 327 20448 493
rect 20362 295 20448 327
rect 20292 293 20448 295
rect 20483 293 20549 527
rect 20584 327 20650 493
rect 20704 459 20937 493
rect 20704 329 20738 459
rect 20781 351 20867 425
rect 20584 295 20670 327
rect 20584 293 20740 295
rect 20292 261 20396 293
rect 20636 261 20740 293
rect 20292 241 20375 261
rect 19053 117 19169 151
rect 18790 51 19019 85
rect 19119 66 19169 117
rect 19203 17 19253 132
rect 19287 117 19403 151
rect 19287 66 19337 117
rect 19437 85 19471 154
rect 19505 119 19571 177
rect 19605 143 19843 177
rect 19605 85 19666 143
rect 19437 51 19666 85
rect 19700 17 19743 109
rect 19777 51 19843 143
rect 19901 143 20139 177
rect 19901 51 19967 143
rect 20001 17 20044 109
rect 20078 85 20139 143
rect 20173 119 20239 177
rect 20273 85 20307 154
rect 20341 151 20375 241
rect 20430 205 20497 259
rect 20535 205 20602 259
rect 20657 241 20740 261
rect 20657 151 20691 241
rect 20809 177 20843 351
rect 20903 333 20937 459
rect 20981 421 21041 527
rect 21075 442 21141 493
rect 20981 367 21047 421
rect 21081 333 21141 442
rect 20903 299 21141 333
rect 21204 321 21264 527
rect 21298 321 21364 493
rect 21403 321 21458 527
rect 21330 279 21364 321
rect 21507 313 21567 493
rect 20977 211 21141 265
rect 21177 199 21296 265
rect 21330 213 21567 279
rect 21601 273 21667 815
rect 21701 595 21755 781
rect 21701 307 21755 493
rect 21789 273 21855 815
rect 22949 815 23203 875
rect 21889 755 22335 789
rect 21889 595 21949 755
rect 21993 561 22047 721
rect 22081 595 22147 755
rect 22181 561 22235 721
rect 22269 595 22335 755
rect 22369 561 22435 789
rect 22469 755 22915 789
rect 22469 595 22535 755
rect 22569 561 22623 721
rect 22657 595 22723 755
rect 22757 561 22811 721
rect 22855 595 22915 755
rect 21889 527 22915 561
rect 21889 333 21949 493
rect 21993 367 22047 527
rect 22081 333 22147 493
rect 22181 367 22235 527
rect 22269 333 22335 493
rect 21889 299 22335 333
rect 22369 299 22435 527
rect 22469 333 22535 493
rect 22569 367 22623 527
rect 22657 333 22723 493
rect 22757 367 22811 527
rect 22855 333 22915 493
rect 22469 299 22915 333
rect 21601 213 21855 273
rect 22949 273 23015 815
rect 23049 595 23103 781
rect 23049 307 23103 493
rect 23137 273 23203 815
rect 23237 809 23474 875
rect 23508 823 23627 889
rect 23661 823 23780 889
rect 23814 875 23848 923
rect 24125 875 24191 969
rect 24225 934 24259 1003
rect 24293 911 24359 969
rect 24393 945 24447 1003
rect 24481 979 24531 1071
rect 24565 945 24631 1037
rect 24665 979 24719 1071
rect 24753 945 24819 1037
rect 24393 911 24819 945
rect 24853 911 24919 1071
rect 24953 945 25019 1037
rect 25053 979 25107 1071
rect 25141 945 25207 1037
rect 25241 979 25291 1071
rect 25325 1003 25731 1037
rect 25325 945 25379 1003
rect 24953 911 25379 945
rect 25413 911 25479 969
rect 25513 934 25547 1003
rect 24293 875 24339 911
rect 23237 595 23297 775
rect 23440 767 23474 809
rect 23814 809 24051 875
rect 24085 815 24339 875
rect 24575 823 24853 877
rect 24919 823 25197 877
rect 25433 875 25479 911
rect 25581 875 25647 969
rect 25681 934 25731 1003
rect 25832 966 25890 1071
rect 25924 923 25974 1032
rect 26016 966 26074 1071
rect 25924 875 25958 923
rect 26154 911 26206 1071
rect 26240 963 26295 1009
rect 23814 767 23848 809
rect 23346 561 23401 767
rect 23440 595 23506 767
rect 23540 561 23600 767
rect 23688 561 23748 767
rect 23782 595 23848 767
rect 23887 561 23942 767
rect 23991 595 24051 775
rect 23237 527 24051 561
rect 23237 313 23297 493
rect 23346 321 23401 527
rect 23440 321 23506 493
rect 23540 321 23600 527
rect 23688 321 23748 527
rect 23782 321 23848 493
rect 23887 321 23942 527
rect 23440 279 23474 321
rect 20893 177 20954 185
rect 20341 117 20457 151
rect 20078 51 20307 85
rect 20407 66 20457 117
rect 20491 17 20541 132
rect 20575 117 20691 151
rect 20575 66 20625 117
rect 20725 85 20759 154
rect 20793 119 20859 177
rect 20893 143 21131 177
rect 21330 165 21364 213
rect 20893 85 20954 143
rect 20725 51 20954 85
rect 20988 17 21031 109
rect 21065 51 21131 143
rect 21214 17 21272 122
rect 21314 56 21364 165
rect 21398 17 21456 122
rect 21557 85 21607 154
rect 21641 119 21707 213
rect 21809 177 21855 213
rect 22091 211 22369 265
rect 22435 211 22713 265
rect 22949 213 23203 273
rect 23237 213 23474 279
rect 23814 279 23848 321
rect 23991 313 24051 493
rect 22949 177 22995 213
rect 21741 85 21775 154
rect 21809 119 21875 177
rect 21909 143 22335 177
rect 21909 85 21963 143
rect 21557 51 21963 85
rect 21997 17 22047 109
rect 22081 51 22147 143
rect 22181 17 22235 109
rect 22269 51 22335 143
rect 22369 17 22435 177
rect 22469 143 22895 177
rect 22469 51 22535 143
rect 22569 17 22623 109
rect 22657 51 22723 143
rect 22757 17 22807 109
rect 22841 85 22895 143
rect 22929 119 22995 177
rect 23029 85 23063 154
rect 23097 119 23163 213
rect 23440 165 23474 213
rect 23508 199 23627 265
rect 23661 199 23780 265
rect 23814 213 24051 279
rect 24085 273 24151 815
rect 24185 595 24239 781
rect 24185 307 24239 493
rect 24273 273 24339 815
rect 25433 815 25687 875
rect 24373 755 24819 789
rect 24373 595 24433 755
rect 24477 561 24531 721
rect 24565 595 24631 755
rect 24665 561 24719 721
rect 24753 595 24819 755
rect 24853 561 24919 789
rect 24953 755 25399 789
rect 24953 595 25019 755
rect 25053 561 25107 721
rect 25141 595 25207 755
rect 25241 561 25295 721
rect 25339 595 25399 755
rect 24373 527 25399 561
rect 24373 333 24433 493
rect 24477 367 24531 527
rect 24565 333 24631 493
rect 24665 367 24719 527
rect 24753 333 24819 493
rect 24373 299 24819 333
rect 24853 299 24919 527
rect 24953 333 25019 493
rect 25053 367 25107 527
rect 25141 333 25207 493
rect 25241 367 25295 527
rect 25339 333 25399 493
rect 24953 299 25399 333
rect 24085 213 24339 273
rect 25433 273 25499 815
rect 25533 595 25587 781
rect 25533 307 25587 493
rect 25621 273 25687 815
rect 25721 809 25958 875
rect 25992 823 26111 889
rect 26240 877 26274 963
rect 26337 921 26386 1022
rect 26458 971 26508 1022
rect 26195 823 26274 877
rect 26308 887 26386 921
rect 26420 937 26508 971
rect 26555 956 26621 1071
rect 26668 971 26718 1022
rect 26668 937 26756 971
rect 25721 595 25781 775
rect 25924 767 25958 809
rect 25830 561 25885 767
rect 25924 595 25990 767
rect 26024 561 26084 767
rect 26147 561 26213 789
rect 26308 737 26342 887
rect 26420 853 26454 937
rect 26376 795 26454 853
rect 26489 829 26569 899
rect 26607 829 26687 899
rect 26722 853 26756 937
rect 26790 921 26839 1022
rect 26881 963 26936 1009
rect 26790 887 26868 921
rect 26722 795 26800 853
rect 26376 787 26516 795
rect 26420 761 26516 787
rect 26308 727 26387 737
rect 26308 691 26412 727
rect 26346 595 26412 691
rect 26450 595 26516 761
rect 25721 527 26312 561
rect 25721 313 25781 493
rect 25830 321 25885 527
rect 25924 321 25990 493
rect 26024 321 26084 527
rect 25924 279 25958 321
rect 26147 299 26213 527
rect 26346 493 26387 595
rect 26555 561 26621 795
rect 26660 787 26800 795
rect 26660 761 26756 787
rect 26660 595 26726 761
rect 26834 737 26868 887
rect 26902 877 26936 963
rect 26970 911 27034 1071
rect 27068 963 27123 1009
rect 27068 877 27102 963
rect 27165 921 27214 1022
rect 27286 971 27336 1022
rect 26902 823 26981 877
rect 27023 823 27102 877
rect 27136 887 27214 921
rect 27248 937 27336 971
rect 27383 956 27449 1071
rect 27496 971 27546 1022
rect 27496 937 27584 971
rect 26789 727 26868 737
rect 26764 691 26868 727
rect 26764 595 26830 691
rect 26421 527 26755 561
rect 26346 397 26412 493
rect 26308 361 26412 397
rect 26308 351 26387 361
rect 23814 165 23848 213
rect 23197 85 23247 154
rect 22841 51 23247 85
rect 23348 17 23406 122
rect 23440 56 23490 165
rect 23532 17 23590 122
rect 23698 17 23756 122
rect 23798 56 23848 165
rect 23882 17 23940 122
rect 24041 85 24091 154
rect 24125 119 24191 213
rect 24293 177 24339 213
rect 24575 211 24853 265
rect 24919 211 25197 265
rect 25433 213 25687 273
rect 25721 213 25958 279
rect 25433 177 25479 213
rect 24225 85 24259 154
rect 24293 119 24359 177
rect 24393 143 24819 177
rect 24393 85 24447 143
rect 24041 51 24447 85
rect 24481 17 24531 109
rect 24565 51 24631 143
rect 24665 17 24719 109
rect 24753 51 24819 143
rect 24853 17 24919 177
rect 24953 143 25379 177
rect 24953 51 25019 143
rect 25053 17 25107 109
rect 25141 51 25207 143
rect 25241 17 25291 109
rect 25325 85 25379 143
rect 25413 119 25479 177
rect 25513 85 25547 154
rect 25581 119 25647 213
rect 25924 165 25958 213
rect 25992 199 26111 265
rect 26195 211 26274 265
rect 25681 85 25731 154
rect 25325 51 25731 85
rect 25832 17 25890 122
rect 25924 56 25974 165
rect 26016 17 26074 122
rect 26154 17 26206 177
rect 26240 125 26274 211
rect 26308 201 26342 351
rect 26450 327 26516 493
rect 26420 301 26516 327
rect 26376 293 26516 301
rect 26555 293 26621 527
rect 26789 493 26830 595
rect 26963 561 27041 789
rect 27136 737 27170 887
rect 27248 853 27282 937
rect 27204 795 27282 853
rect 27317 829 27397 899
rect 27435 829 27515 899
rect 27550 853 27584 937
rect 27618 921 27667 1022
rect 27709 963 27764 1009
rect 27618 887 27696 921
rect 27550 795 27628 853
rect 27204 787 27344 795
rect 27248 761 27344 787
rect 27136 727 27215 737
rect 27136 691 27240 727
rect 27174 595 27240 691
rect 27278 595 27344 761
rect 26864 527 27140 561
rect 26660 327 26726 493
rect 26764 397 26830 493
rect 26764 361 26868 397
rect 26789 351 26868 361
rect 26660 301 26756 327
rect 26660 293 26800 301
rect 26376 235 26454 293
rect 26308 167 26386 201
rect 26240 79 26295 125
rect 26337 66 26386 167
rect 26420 151 26454 235
rect 26489 189 26569 259
rect 26607 189 26687 259
rect 26722 235 26800 293
rect 26722 151 26756 235
rect 26834 201 26868 351
rect 26963 299 27041 527
rect 27174 493 27215 595
rect 27383 561 27449 795
rect 27488 787 27628 795
rect 27488 761 27584 787
rect 27488 595 27554 761
rect 27662 737 27696 887
rect 27730 877 27764 963
rect 27798 911 27862 1071
rect 27896 963 27951 1009
rect 27896 877 27930 963
rect 27993 921 28042 1022
rect 28114 971 28164 1022
rect 27730 823 27809 877
rect 27851 823 27930 877
rect 27964 887 28042 921
rect 28076 937 28164 971
rect 28211 956 28277 1071
rect 28324 971 28374 1022
rect 28324 937 28412 971
rect 27617 727 27696 737
rect 27592 691 27696 727
rect 27592 595 27658 691
rect 27249 527 27583 561
rect 27174 397 27240 493
rect 27136 361 27240 397
rect 27136 351 27215 361
rect 26420 117 26508 151
rect 26458 66 26508 117
rect 26555 17 26621 132
rect 26668 117 26756 151
rect 26790 167 26868 201
rect 26902 211 26981 265
rect 27023 211 27102 265
rect 26668 66 26718 117
rect 26790 66 26839 167
rect 26902 125 26936 211
rect 26881 79 26936 125
rect 26970 17 27034 177
rect 27068 125 27102 211
rect 27136 201 27170 351
rect 27278 327 27344 493
rect 27248 301 27344 327
rect 27204 293 27344 301
rect 27383 293 27449 527
rect 27617 493 27658 595
rect 27791 561 27869 789
rect 27964 737 27998 887
rect 28076 853 28110 937
rect 28032 795 28110 853
rect 28145 829 28225 899
rect 28263 829 28343 899
rect 28378 853 28412 937
rect 28446 921 28495 1022
rect 28537 963 28592 1009
rect 28446 887 28524 921
rect 28378 795 28456 853
rect 28032 787 28172 795
rect 28076 761 28172 787
rect 27964 727 28043 737
rect 27964 691 28068 727
rect 28002 595 28068 691
rect 28106 595 28172 761
rect 27692 527 27968 561
rect 27488 327 27554 493
rect 27592 397 27658 493
rect 27592 361 27696 397
rect 27617 351 27696 361
rect 27488 301 27584 327
rect 27488 293 27628 301
rect 27204 235 27282 293
rect 27136 167 27214 201
rect 27068 79 27123 125
rect 27165 66 27214 167
rect 27248 151 27282 235
rect 27317 189 27397 259
rect 27435 189 27515 259
rect 27550 235 27628 293
rect 27550 151 27584 235
rect 27662 201 27696 351
rect 27791 299 27869 527
rect 28002 493 28043 595
rect 28211 561 28277 795
rect 28316 787 28456 795
rect 28316 761 28412 787
rect 28316 595 28382 761
rect 28490 737 28524 887
rect 28558 877 28592 963
rect 28626 911 28690 1071
rect 28724 963 28779 1009
rect 28724 877 28758 963
rect 28821 921 28870 1022
rect 28942 971 28992 1022
rect 28558 823 28637 877
rect 28679 823 28758 877
rect 28792 887 28870 921
rect 28904 937 28992 971
rect 29039 956 29105 1071
rect 29152 971 29202 1022
rect 29152 937 29240 971
rect 28445 727 28524 737
rect 28420 691 28524 727
rect 28420 595 28486 691
rect 28077 527 28411 561
rect 28002 397 28068 493
rect 27964 361 28068 397
rect 27964 351 28043 361
rect 27248 117 27336 151
rect 27286 66 27336 117
rect 27383 17 27449 132
rect 27496 117 27584 151
rect 27618 167 27696 201
rect 27730 211 27809 265
rect 27851 211 27930 265
rect 27496 66 27546 117
rect 27618 66 27667 167
rect 27730 125 27764 211
rect 27709 79 27764 125
rect 27798 17 27862 177
rect 27896 125 27930 211
rect 27964 201 27998 351
rect 28106 327 28172 493
rect 28076 301 28172 327
rect 28032 293 28172 301
rect 28211 293 28277 527
rect 28445 493 28486 595
rect 28619 561 28697 789
rect 28792 737 28826 887
rect 28904 853 28938 937
rect 28860 795 28938 853
rect 28973 829 29053 899
rect 29091 829 29171 899
rect 29206 853 29240 937
rect 29274 921 29323 1022
rect 29365 963 29420 1009
rect 29274 887 29352 921
rect 29206 795 29284 853
rect 28860 787 29000 795
rect 28904 761 29000 787
rect 28792 727 28871 737
rect 28792 691 28896 727
rect 28830 595 28896 691
rect 28934 595 29000 761
rect 28520 527 28796 561
rect 28316 327 28382 493
rect 28420 397 28486 493
rect 28420 361 28524 397
rect 28445 351 28524 361
rect 28316 301 28412 327
rect 28316 293 28456 301
rect 28032 235 28110 293
rect 27964 167 28042 201
rect 27896 79 27951 125
rect 27993 66 28042 167
rect 28076 151 28110 235
rect 28145 189 28225 259
rect 28263 189 28343 259
rect 28378 235 28456 293
rect 28378 151 28412 235
rect 28490 201 28524 351
rect 28619 299 28697 527
rect 28830 493 28871 595
rect 29039 561 29105 795
rect 29144 787 29284 795
rect 29144 761 29240 787
rect 29144 595 29210 761
rect 29318 737 29352 887
rect 29386 877 29420 963
rect 29454 911 29506 1071
rect 29561 945 29627 1037
rect 29661 979 29704 1071
rect 29738 1003 29967 1037
rect 29738 945 29799 1003
rect 29561 911 29799 945
rect 29833 911 29899 969
rect 29933 934 29967 1003
rect 30067 971 30117 1022
rect 30001 937 30117 971
rect 30151 956 30201 1071
rect 30235 971 30285 1022
rect 30385 1003 30614 1037
rect 30235 937 30351 971
rect 29738 903 29799 911
rect 29386 823 29465 877
rect 29551 823 29715 877
rect 29273 727 29352 737
rect 29248 691 29352 727
rect 29248 595 29314 691
rect 28905 527 29239 561
rect 28830 397 28896 493
rect 28792 361 28896 397
rect 28792 351 28871 361
rect 28076 117 28164 151
rect 28114 66 28164 117
rect 28211 17 28277 132
rect 28324 117 28412 151
rect 28446 167 28524 201
rect 28558 211 28637 265
rect 28679 211 28758 265
rect 28324 66 28374 117
rect 28446 66 28495 167
rect 28558 125 28592 211
rect 28537 79 28592 125
rect 28626 17 28690 177
rect 28724 125 28758 211
rect 28792 201 28826 351
rect 28934 327 29000 493
rect 28904 301 29000 327
rect 28860 293 29000 301
rect 29039 293 29105 527
rect 29273 493 29314 595
rect 29447 561 29513 789
rect 29551 755 29789 789
rect 29551 646 29611 755
rect 29645 667 29711 721
rect 29551 595 29617 646
rect 29651 561 29711 667
rect 29755 629 29789 755
rect 29849 737 29883 911
rect 30001 847 30035 937
rect 29952 827 30035 847
rect 30090 829 30157 883
rect 30195 829 30262 883
rect 30317 847 30351 937
rect 30385 934 30419 1003
rect 30453 911 30519 969
rect 30553 945 30614 1003
rect 30648 979 30691 1071
rect 30725 945 30791 1037
rect 30553 911 30791 945
rect 30849 945 30915 1037
rect 30949 979 30992 1071
rect 31026 1003 31255 1037
rect 31026 945 31087 1003
rect 30849 911 31087 945
rect 31121 911 31187 969
rect 31221 934 31255 1003
rect 31355 971 31405 1022
rect 31289 937 31405 971
rect 31439 956 31489 1071
rect 31523 971 31573 1022
rect 31673 1003 31902 1037
rect 31523 937 31639 971
rect 30317 827 30400 847
rect 29952 795 30056 827
rect 30296 795 30400 827
rect 29952 793 30108 795
rect 30022 761 30108 793
rect 29825 663 29911 737
rect 29755 595 29815 629
rect 29348 527 29815 561
rect 29144 327 29210 493
rect 29248 397 29314 493
rect 29248 361 29352 397
rect 29273 351 29352 361
rect 29144 301 29240 327
rect 29144 293 29284 301
rect 28860 235 28938 293
rect 28792 167 28870 201
rect 28724 79 28779 125
rect 28821 66 28870 167
rect 28904 151 28938 235
rect 28973 189 29053 259
rect 29091 189 29171 259
rect 29206 235 29284 293
rect 29206 151 29240 235
rect 29318 201 29352 351
rect 29447 299 29513 527
rect 29551 442 29617 493
rect 29551 333 29611 442
rect 29651 421 29711 527
rect 29645 367 29711 421
rect 29755 459 29815 493
rect 29755 333 29789 459
rect 29849 425 29883 663
rect 29954 629 29988 759
rect 29917 595 29988 629
rect 30042 595 30108 761
rect 30143 561 30209 795
rect 30244 793 30400 795
rect 30244 761 30330 793
rect 30244 595 30310 761
rect 30364 629 30398 759
rect 30469 737 30503 911
rect 30553 903 30614 911
rect 31026 903 31087 911
rect 30637 823 30801 877
rect 30839 823 31003 877
rect 30563 755 30801 789
rect 30441 663 30527 737
rect 30364 595 30435 629
rect 29917 527 30435 561
rect 29917 459 29988 493
rect 29825 351 29911 425
rect 29551 299 29789 333
rect 28904 117 28992 151
rect 28942 66 28992 117
rect 29039 17 29105 132
rect 29152 117 29240 151
rect 29274 167 29352 201
rect 29386 211 29465 265
rect 29551 211 29715 265
rect 29152 66 29202 117
rect 29274 66 29323 167
rect 29386 125 29420 211
rect 29738 177 29799 185
rect 29849 177 29883 351
rect 29954 329 29988 459
rect 30042 327 30108 493
rect 30022 295 30108 327
rect 29952 293 30108 295
rect 30143 293 30209 527
rect 30244 327 30310 493
rect 30364 459 30435 493
rect 30364 329 30398 459
rect 30469 425 30503 663
rect 30563 629 30597 755
rect 30537 595 30597 629
rect 30641 667 30707 721
rect 30641 561 30701 667
rect 30741 646 30801 755
rect 30735 595 30801 646
rect 30839 755 31077 789
rect 30839 646 30899 755
rect 30933 667 30999 721
rect 30839 595 30905 646
rect 30939 561 30999 667
rect 31043 629 31077 755
rect 31137 737 31171 911
rect 31289 847 31323 937
rect 31240 827 31323 847
rect 31378 829 31445 883
rect 31483 829 31550 883
rect 31605 847 31639 937
rect 31673 934 31707 1003
rect 31741 911 31807 969
rect 31841 945 31902 1003
rect 31936 979 31979 1071
rect 32013 945 32079 1037
rect 31841 911 32079 945
rect 32137 945 32203 1037
rect 32237 979 32280 1071
rect 32314 1003 32543 1037
rect 32314 945 32375 1003
rect 32137 911 32375 945
rect 32409 911 32475 969
rect 32509 934 32543 1003
rect 32643 971 32693 1022
rect 32577 937 32693 971
rect 32727 956 32777 1071
rect 32811 971 32861 1022
rect 32961 1003 33190 1037
rect 32811 937 32927 971
rect 31605 827 31688 847
rect 31240 795 31344 827
rect 31584 795 31688 827
rect 31240 793 31396 795
rect 31310 761 31396 793
rect 31113 663 31199 737
rect 31043 595 31103 629
rect 30537 527 31103 561
rect 30537 459 30597 493
rect 30441 351 30527 425
rect 30244 295 30330 327
rect 30244 293 30400 295
rect 29952 261 30056 293
rect 30296 261 30400 293
rect 29952 241 30035 261
rect 29365 79 29420 125
rect 29454 17 29506 177
rect 29561 143 29799 177
rect 29561 51 29627 143
rect 29661 17 29704 109
rect 29738 85 29799 143
rect 29833 119 29899 177
rect 29933 85 29967 154
rect 30001 151 30035 241
rect 30090 205 30157 259
rect 30195 205 30262 259
rect 30317 241 30400 261
rect 30317 151 30351 241
rect 30469 177 30503 351
rect 30563 333 30597 459
rect 30641 421 30701 527
rect 30735 442 30801 493
rect 30641 367 30707 421
rect 30741 333 30801 442
rect 30563 299 30801 333
rect 30839 442 30905 493
rect 30839 333 30899 442
rect 30939 421 30999 527
rect 30933 367 30999 421
rect 31043 459 31103 493
rect 31043 333 31077 459
rect 31137 425 31171 663
rect 31242 629 31276 759
rect 31205 595 31276 629
rect 31330 595 31396 761
rect 31431 561 31497 795
rect 31532 793 31688 795
rect 31532 761 31618 793
rect 31532 595 31598 761
rect 31652 629 31686 759
rect 31757 737 31791 911
rect 31841 903 31902 911
rect 32314 903 32375 911
rect 31925 823 32089 877
rect 32127 823 32291 877
rect 31851 755 32089 789
rect 31729 663 31815 737
rect 31652 595 31723 629
rect 31205 527 31723 561
rect 31205 459 31276 493
rect 31113 351 31199 425
rect 30839 299 31077 333
rect 30637 211 30801 265
rect 30839 211 31003 265
rect 30553 177 30614 185
rect 31026 177 31087 185
rect 31137 177 31171 351
rect 31242 329 31276 459
rect 31330 327 31396 493
rect 31310 295 31396 327
rect 31240 293 31396 295
rect 31431 293 31497 527
rect 31532 327 31598 493
rect 31652 459 31723 493
rect 31652 329 31686 459
rect 31757 425 31791 663
rect 31851 629 31885 755
rect 31825 595 31885 629
rect 31929 667 31995 721
rect 31929 561 31989 667
rect 32029 646 32089 755
rect 32023 595 32089 646
rect 32127 755 32365 789
rect 32127 646 32187 755
rect 32221 667 32287 721
rect 32127 595 32193 646
rect 32227 561 32287 667
rect 32331 629 32365 755
rect 32425 737 32459 911
rect 32577 847 32611 937
rect 32528 827 32611 847
rect 32666 829 32733 883
rect 32771 829 32838 883
rect 32893 847 32927 937
rect 32961 934 32995 1003
rect 33029 911 33095 969
rect 33129 945 33190 1003
rect 33224 979 33267 1071
rect 33301 945 33367 1037
rect 33129 911 33367 945
rect 33425 945 33491 1037
rect 33525 979 33568 1071
rect 33602 1003 33831 1037
rect 33602 945 33663 1003
rect 33425 911 33663 945
rect 33697 911 33763 969
rect 33797 934 33831 1003
rect 33931 971 33981 1022
rect 33865 937 33981 971
rect 34015 956 34065 1071
rect 34099 971 34149 1022
rect 34249 1003 34478 1037
rect 34099 937 34215 971
rect 32893 827 32976 847
rect 32528 795 32632 827
rect 32872 795 32976 827
rect 32528 793 32684 795
rect 32598 761 32684 793
rect 32401 663 32487 737
rect 32331 595 32391 629
rect 31825 527 32391 561
rect 31825 459 31885 493
rect 31729 351 31815 425
rect 31532 295 31618 327
rect 31532 293 31688 295
rect 31240 261 31344 293
rect 31584 261 31688 293
rect 31240 241 31323 261
rect 30001 117 30117 151
rect 29738 51 29967 85
rect 30067 66 30117 117
rect 30151 17 30201 132
rect 30235 117 30351 151
rect 30235 66 30285 117
rect 30385 85 30419 154
rect 30453 119 30519 177
rect 30553 143 30791 177
rect 30553 85 30614 143
rect 30385 51 30614 85
rect 30648 17 30691 109
rect 30725 51 30791 143
rect 30849 143 31087 177
rect 30849 51 30915 143
rect 30949 17 30992 109
rect 31026 85 31087 143
rect 31121 119 31187 177
rect 31221 85 31255 154
rect 31289 151 31323 241
rect 31378 205 31445 259
rect 31483 205 31550 259
rect 31605 241 31688 261
rect 31605 151 31639 241
rect 31757 177 31791 351
rect 31851 333 31885 459
rect 31929 421 31989 527
rect 32023 442 32089 493
rect 31929 367 31995 421
rect 32029 333 32089 442
rect 31851 299 32089 333
rect 32127 442 32193 493
rect 32127 333 32187 442
rect 32227 421 32287 527
rect 32221 367 32287 421
rect 32331 459 32391 493
rect 32331 333 32365 459
rect 32425 425 32459 663
rect 32530 629 32564 759
rect 32493 595 32564 629
rect 32618 595 32684 761
rect 32719 561 32785 795
rect 32820 793 32976 795
rect 32820 761 32906 793
rect 32820 595 32886 761
rect 32940 629 32974 759
rect 33045 737 33079 911
rect 33129 903 33190 911
rect 33602 903 33663 911
rect 33213 823 33377 877
rect 33415 823 33579 877
rect 33139 755 33377 789
rect 33017 663 33103 737
rect 32940 595 33011 629
rect 32493 527 33011 561
rect 32493 459 32564 493
rect 32401 351 32487 425
rect 32127 299 32365 333
rect 31925 211 32089 265
rect 32127 211 32291 265
rect 31841 177 31902 185
rect 32314 177 32375 185
rect 32425 177 32459 351
rect 32530 329 32564 459
rect 32618 327 32684 493
rect 32598 295 32684 327
rect 32528 293 32684 295
rect 32719 293 32785 527
rect 32820 327 32886 493
rect 32940 459 33011 493
rect 32940 329 32974 459
rect 33045 425 33079 663
rect 33139 629 33173 755
rect 33113 595 33173 629
rect 33217 667 33283 721
rect 33217 561 33277 667
rect 33317 646 33377 755
rect 33311 595 33377 646
rect 33415 755 33653 789
rect 33415 646 33475 755
rect 33509 667 33575 721
rect 33415 595 33481 646
rect 33515 561 33575 667
rect 33619 629 33653 755
rect 33713 737 33747 911
rect 33865 847 33899 937
rect 33816 827 33899 847
rect 33954 829 34021 883
rect 34059 829 34126 883
rect 34181 847 34215 937
rect 34249 934 34283 1003
rect 34317 911 34383 969
rect 34417 945 34478 1003
rect 34512 979 34555 1071
rect 34589 945 34655 1037
rect 34417 911 34655 945
rect 34713 911 34763 1071
rect 34797 945 34863 1037
rect 34897 979 34951 1071
rect 34985 945 35051 1037
rect 35085 979 35135 1071
rect 35169 1003 35575 1037
rect 35169 945 35223 1003
rect 34797 911 35223 945
rect 35257 911 35323 969
rect 35357 934 35391 1003
rect 34181 827 34264 847
rect 33816 795 33920 827
rect 34160 795 34264 827
rect 33816 793 33972 795
rect 33886 761 33972 793
rect 33689 663 33775 737
rect 33619 595 33679 629
rect 33113 527 33679 561
rect 33113 459 33173 493
rect 33017 351 33103 425
rect 32820 295 32906 327
rect 32820 293 32976 295
rect 32528 261 32632 293
rect 32872 261 32976 293
rect 32528 241 32611 261
rect 31289 117 31405 151
rect 31026 51 31255 85
rect 31355 66 31405 117
rect 31439 17 31489 132
rect 31523 117 31639 151
rect 31523 66 31573 117
rect 31673 85 31707 154
rect 31741 119 31807 177
rect 31841 143 32079 177
rect 31841 85 31902 143
rect 31673 51 31902 85
rect 31936 17 31979 109
rect 32013 51 32079 143
rect 32137 143 32375 177
rect 32137 51 32203 143
rect 32237 17 32280 109
rect 32314 85 32375 143
rect 32409 119 32475 177
rect 32509 85 32543 154
rect 32577 151 32611 241
rect 32666 205 32733 259
rect 32771 205 32838 259
rect 32893 241 32976 261
rect 32893 151 32927 241
rect 33045 177 33079 351
rect 33139 333 33173 459
rect 33217 421 33277 527
rect 33311 442 33377 493
rect 33217 367 33283 421
rect 33317 333 33377 442
rect 33139 299 33377 333
rect 33415 442 33481 493
rect 33415 333 33475 442
rect 33515 421 33575 527
rect 33509 367 33575 421
rect 33619 459 33679 493
rect 33619 333 33653 459
rect 33713 425 33747 663
rect 33818 629 33852 759
rect 33781 595 33852 629
rect 33906 595 33972 761
rect 34007 561 34073 795
rect 34108 793 34264 795
rect 34108 761 34194 793
rect 34108 595 34174 761
rect 34228 629 34262 759
rect 34333 737 34367 911
rect 34417 903 34478 911
rect 34501 823 34665 877
rect 34763 823 35041 877
rect 35277 875 35323 911
rect 35425 875 35491 969
rect 35525 934 35575 1003
rect 35676 966 35734 1071
rect 35768 923 35818 1032
rect 35860 966 35918 1071
rect 36026 966 36084 1071
rect 36126 923 36176 1032
rect 36210 966 36268 1071
rect 36369 1003 36775 1037
rect 36369 934 36419 1003
rect 35768 875 35802 923
rect 35277 815 35531 875
rect 34427 755 34665 789
rect 34305 663 34391 737
rect 34228 595 34299 629
rect 33781 527 34299 561
rect 33781 459 33852 493
rect 33689 351 33775 425
rect 33415 299 33653 333
rect 33213 211 33377 265
rect 33415 211 33579 265
rect 33129 177 33190 185
rect 33602 177 33663 185
rect 33713 177 33747 351
rect 33818 329 33852 459
rect 33906 327 33972 493
rect 33886 295 33972 327
rect 33816 293 33972 295
rect 34007 293 34073 527
rect 34108 327 34174 493
rect 34228 459 34299 493
rect 34228 329 34262 459
rect 34333 425 34367 663
rect 34427 629 34461 755
rect 34401 595 34461 629
rect 34505 667 34571 721
rect 34505 561 34565 667
rect 34605 646 34665 755
rect 34599 595 34665 646
rect 34709 561 34763 789
rect 34797 755 35243 789
rect 34797 595 34863 755
rect 34897 561 34951 721
rect 34985 595 35051 755
rect 35085 561 35139 721
rect 35183 595 35243 755
rect 34401 527 35243 561
rect 34401 459 34461 493
rect 34305 351 34391 425
rect 34108 295 34194 327
rect 34108 293 34264 295
rect 33816 261 33920 293
rect 34160 261 34264 293
rect 33816 241 33899 261
rect 32577 117 32693 151
rect 32314 51 32543 85
rect 32643 66 32693 117
rect 32727 17 32777 132
rect 32811 117 32927 151
rect 32811 66 32861 117
rect 32961 85 32995 154
rect 33029 119 33095 177
rect 33129 143 33367 177
rect 33129 85 33190 143
rect 32961 51 33190 85
rect 33224 17 33267 109
rect 33301 51 33367 143
rect 33425 143 33663 177
rect 33425 51 33491 143
rect 33525 17 33568 109
rect 33602 85 33663 143
rect 33697 119 33763 177
rect 33797 85 33831 154
rect 33865 151 33899 241
rect 33954 205 34021 259
rect 34059 205 34126 259
rect 34181 241 34264 261
rect 34181 151 34215 241
rect 34333 177 34367 351
rect 34427 333 34461 459
rect 34505 421 34565 527
rect 34599 442 34665 493
rect 34505 367 34571 421
rect 34605 333 34665 442
rect 34427 299 34665 333
rect 34709 299 34763 527
rect 34797 333 34863 493
rect 34897 367 34951 527
rect 34985 333 35051 493
rect 35085 367 35139 527
rect 35183 333 35243 493
rect 34797 299 35243 333
rect 35277 273 35343 815
rect 35377 595 35431 781
rect 35377 307 35431 493
rect 35465 273 35531 815
rect 35565 809 35802 875
rect 35836 823 35955 889
rect 35989 823 36108 889
rect 36142 875 36176 923
rect 36453 875 36519 969
rect 36553 934 36587 1003
rect 36621 911 36687 969
rect 36721 945 36775 1003
rect 36809 979 36859 1071
rect 36893 945 36959 1037
rect 36993 979 37047 1071
rect 37081 945 37147 1037
rect 36721 911 37147 945
rect 37181 911 37231 1071
rect 37289 911 37339 1071
rect 37373 945 37439 1037
rect 37473 979 37527 1071
rect 37561 945 37627 1037
rect 37661 979 37711 1071
rect 37745 1003 38151 1037
rect 37745 945 37799 1003
rect 37373 911 37799 945
rect 37833 911 37899 969
rect 37933 934 37967 1003
rect 36621 875 36667 911
rect 35565 595 35625 775
rect 35768 767 35802 809
rect 36142 809 36379 875
rect 36413 815 36667 875
rect 36903 823 37181 877
rect 37339 823 37617 877
rect 37853 875 37899 911
rect 38001 875 38067 969
rect 38101 934 38151 1003
rect 38252 966 38310 1071
rect 38344 923 38394 1032
rect 38436 966 38494 1071
rect 38602 966 38660 1071
rect 38702 923 38752 1032
rect 38786 966 38844 1071
rect 38945 1003 39351 1037
rect 38945 934 38995 1003
rect 38344 875 38378 923
rect 36142 767 36176 809
rect 35674 561 35729 767
rect 35768 595 35834 767
rect 35868 561 35928 767
rect 36016 561 36076 767
rect 36110 595 36176 767
rect 36215 561 36270 767
rect 36319 595 36379 775
rect 35565 527 36379 561
rect 35565 313 35625 493
rect 35674 321 35729 527
rect 35768 321 35834 493
rect 35868 321 35928 527
rect 36016 321 36076 527
rect 36110 321 36176 493
rect 36215 321 36270 527
rect 35768 279 35802 321
rect 34501 211 34665 265
rect 34763 211 35041 265
rect 35277 213 35531 273
rect 35565 213 35802 279
rect 36142 279 36176 321
rect 36319 313 36379 493
rect 34417 177 34478 185
rect 35277 177 35323 213
rect 33865 117 33981 151
rect 33602 51 33831 85
rect 33931 66 33981 117
rect 34015 17 34065 132
rect 34099 117 34215 151
rect 34099 66 34149 117
rect 34249 85 34283 154
rect 34317 119 34383 177
rect 34417 143 34655 177
rect 34417 85 34478 143
rect 34249 51 34478 85
rect 34512 17 34555 109
rect 34589 51 34655 143
rect 34713 17 34763 177
rect 34797 143 35223 177
rect 34797 51 34863 143
rect 34897 17 34951 109
rect 34985 51 35051 143
rect 35085 17 35135 109
rect 35169 85 35223 143
rect 35257 119 35323 177
rect 35357 85 35391 154
rect 35425 119 35491 213
rect 35768 165 35802 213
rect 35836 199 35955 265
rect 35989 199 36108 265
rect 36142 213 36379 279
rect 36413 273 36479 815
rect 36513 595 36567 781
rect 36513 307 36567 493
rect 36601 273 36667 815
rect 37853 815 38107 875
rect 36701 755 37147 789
rect 36701 595 36761 755
rect 36805 561 36859 721
rect 36893 595 36959 755
rect 36993 561 37047 721
rect 37081 595 37147 755
rect 37181 561 37235 789
rect 37285 561 37339 789
rect 37373 755 37819 789
rect 37373 595 37439 755
rect 37473 561 37527 721
rect 37561 595 37627 755
rect 37661 561 37715 721
rect 37759 595 37819 755
rect 36701 527 37819 561
rect 36701 333 36761 493
rect 36805 367 36859 527
rect 36893 333 36959 493
rect 36993 367 37047 527
rect 37081 333 37147 493
rect 36701 299 37147 333
rect 37181 299 37235 527
rect 37285 299 37339 527
rect 37373 333 37439 493
rect 37473 367 37527 527
rect 37561 333 37627 493
rect 37661 367 37715 527
rect 37759 333 37819 493
rect 37373 299 37819 333
rect 36413 213 36667 273
rect 37853 273 37919 815
rect 37953 595 38007 781
rect 37953 307 38007 493
rect 38041 273 38107 815
rect 38141 809 38378 875
rect 38412 823 38531 889
rect 38565 823 38684 889
rect 38718 875 38752 923
rect 39029 875 39095 969
rect 39129 934 39163 1003
rect 39197 911 39263 969
rect 39297 945 39351 1003
rect 39385 979 39435 1071
rect 39469 945 39535 1037
rect 39569 979 39623 1071
rect 39657 945 39723 1037
rect 39297 911 39723 945
rect 39757 911 39807 1071
rect 39853 926 39911 1035
rect 39957 911 40007 1071
rect 40041 945 40107 1037
rect 40141 979 40195 1071
rect 40229 945 40295 1037
rect 40329 979 40379 1071
rect 40413 1003 40819 1037
rect 40413 945 40467 1003
rect 40041 911 40467 945
rect 40501 911 40567 969
rect 40601 934 40635 1003
rect 39197 875 39243 911
rect 38141 595 38201 775
rect 38344 767 38378 809
rect 38718 809 38955 875
rect 38989 815 39243 875
rect 39479 823 39757 877
rect 40007 823 40285 877
rect 40521 875 40567 911
rect 40669 875 40735 969
rect 40769 934 40819 1003
rect 40920 966 40978 1071
rect 41012 923 41062 1032
rect 41104 966 41162 1071
rect 41270 966 41328 1071
rect 41370 923 41420 1032
rect 41454 966 41512 1071
rect 41613 1003 42019 1037
rect 41613 934 41663 1003
rect 41012 875 41046 923
rect 38718 767 38752 809
rect 38250 561 38305 767
rect 38344 595 38410 767
rect 38444 561 38504 767
rect 38592 561 38652 767
rect 38686 595 38752 767
rect 38791 561 38846 767
rect 38895 595 38955 775
rect 38141 527 38955 561
rect 38141 313 38201 493
rect 38250 321 38305 527
rect 38344 321 38410 493
rect 38444 321 38504 527
rect 38592 321 38652 527
rect 38686 321 38752 493
rect 38791 321 38846 527
rect 38344 279 38378 321
rect 36142 165 36176 213
rect 35525 85 35575 154
rect 35169 51 35575 85
rect 35676 17 35734 122
rect 35768 56 35818 165
rect 35860 17 35918 122
rect 36026 17 36084 122
rect 36126 56 36176 165
rect 36210 17 36268 122
rect 36369 85 36419 154
rect 36453 119 36519 213
rect 36621 177 36667 213
rect 36903 211 37181 265
rect 37339 211 37617 265
rect 37853 213 38107 273
rect 38141 213 38378 279
rect 38718 279 38752 321
rect 38895 313 38955 493
rect 37853 177 37899 213
rect 36553 85 36587 154
rect 36621 119 36687 177
rect 36721 143 37147 177
rect 36721 85 36775 143
rect 36369 51 36775 85
rect 36809 17 36859 109
rect 36893 51 36959 143
rect 36993 17 37047 109
rect 37081 51 37147 143
rect 37181 17 37231 177
rect 37289 17 37339 177
rect 37373 143 37799 177
rect 37373 51 37439 143
rect 37473 17 37527 109
rect 37561 51 37627 143
rect 37661 17 37711 109
rect 37745 85 37799 143
rect 37833 119 37899 177
rect 37933 85 37967 154
rect 38001 119 38067 213
rect 38344 165 38378 213
rect 38412 199 38531 265
rect 38565 199 38684 265
rect 38718 213 38955 279
rect 38989 273 39055 815
rect 39089 595 39143 781
rect 39089 307 39143 493
rect 39177 273 39243 815
rect 40521 815 40775 875
rect 39277 755 39723 789
rect 39277 595 39337 755
rect 39381 561 39435 721
rect 39469 595 39535 755
rect 39569 561 39623 721
rect 39657 595 39723 755
rect 39757 561 39811 789
rect 39853 597 39911 794
rect 39953 561 40007 789
rect 40041 755 40487 789
rect 40041 595 40107 755
rect 40141 561 40195 721
rect 40229 595 40295 755
rect 40329 561 40383 721
rect 40427 595 40487 755
rect 39277 527 40487 561
rect 39277 333 39337 493
rect 39381 367 39435 527
rect 39469 333 39535 493
rect 39569 367 39623 527
rect 39657 333 39723 493
rect 39277 299 39723 333
rect 39757 299 39811 527
rect 39853 294 39911 491
rect 39953 299 40007 527
rect 40041 333 40107 493
rect 40141 367 40195 527
rect 40229 333 40295 493
rect 40329 367 40383 527
rect 40427 333 40487 493
rect 40041 299 40487 333
rect 38989 213 39243 273
rect 40521 273 40587 815
rect 40621 595 40675 781
rect 40621 307 40675 493
rect 40709 273 40775 815
rect 40809 809 41046 875
rect 41080 823 41199 889
rect 41233 823 41352 889
rect 41386 875 41420 923
rect 41697 875 41763 969
rect 41797 934 41831 1003
rect 41865 911 41931 969
rect 41965 945 42019 1003
rect 42053 979 42103 1071
rect 42137 945 42203 1037
rect 42237 979 42291 1071
rect 42325 945 42391 1037
rect 41965 911 42391 945
rect 42425 911 42475 1071
rect 42533 911 42583 1071
rect 42617 945 42683 1037
rect 42717 979 42771 1071
rect 42805 945 42871 1037
rect 42905 979 42955 1071
rect 42989 1003 43395 1037
rect 42989 945 43043 1003
rect 42617 911 43043 945
rect 43077 911 43143 969
rect 43177 934 43211 1003
rect 41865 875 41911 911
rect 40809 595 40869 775
rect 41012 767 41046 809
rect 41386 809 41623 875
rect 41657 815 41911 875
rect 42147 823 42425 877
rect 42583 823 42861 877
rect 43097 875 43143 911
rect 43245 875 43311 969
rect 43345 934 43395 1003
rect 43496 966 43554 1071
rect 43588 923 43638 1032
rect 43680 966 43738 1071
rect 43846 966 43904 1071
rect 43946 923 43996 1032
rect 44030 966 44088 1071
rect 44189 1003 44595 1037
rect 44189 934 44239 1003
rect 43588 875 43622 923
rect 41386 767 41420 809
rect 40918 561 40973 767
rect 41012 595 41078 767
rect 41112 561 41172 767
rect 41260 561 41320 767
rect 41354 595 41420 767
rect 41459 561 41514 767
rect 41563 595 41623 775
rect 40809 527 41623 561
rect 40809 313 40869 493
rect 40918 321 40973 527
rect 41012 321 41078 493
rect 41112 321 41172 527
rect 41260 321 41320 527
rect 41354 321 41420 493
rect 41459 321 41514 527
rect 41012 279 41046 321
rect 38718 165 38752 213
rect 38101 85 38151 154
rect 37745 51 38151 85
rect 38252 17 38310 122
rect 38344 56 38394 165
rect 38436 17 38494 122
rect 38602 17 38660 122
rect 38702 56 38752 165
rect 38786 17 38844 122
rect 38945 85 38995 154
rect 39029 119 39095 213
rect 39197 177 39243 213
rect 39479 211 39757 265
rect 40007 211 40285 265
rect 40521 213 40775 273
rect 40809 213 41046 279
rect 41386 279 41420 321
rect 41563 313 41623 493
rect 40521 177 40567 213
rect 39129 85 39163 154
rect 39197 119 39263 177
rect 39297 143 39723 177
rect 39297 85 39351 143
rect 38945 51 39351 85
rect 39385 17 39435 109
rect 39469 51 39535 143
rect 39569 17 39623 109
rect 39657 51 39723 143
rect 39757 17 39807 177
rect 39853 53 39911 162
rect 39957 17 40007 177
rect 40041 143 40467 177
rect 40041 51 40107 143
rect 40141 17 40195 109
rect 40229 51 40295 143
rect 40329 17 40379 109
rect 40413 85 40467 143
rect 40501 119 40567 177
rect 40601 85 40635 154
rect 40669 119 40735 213
rect 41012 165 41046 213
rect 41080 199 41199 265
rect 41233 199 41352 265
rect 41386 213 41623 279
rect 41657 273 41723 815
rect 41757 595 41811 781
rect 41757 307 41811 493
rect 41845 273 41911 815
rect 43097 815 43351 875
rect 41945 755 42391 789
rect 41945 595 42005 755
rect 42049 561 42103 721
rect 42137 595 42203 755
rect 42237 561 42291 721
rect 42325 595 42391 755
rect 42425 561 42479 789
rect 42529 561 42583 789
rect 42617 755 43063 789
rect 42617 595 42683 755
rect 42717 561 42771 721
rect 42805 595 42871 755
rect 42905 561 42959 721
rect 43003 595 43063 755
rect 41945 527 43063 561
rect 41945 333 42005 493
rect 42049 367 42103 527
rect 42137 333 42203 493
rect 42237 367 42291 527
rect 42325 333 42391 493
rect 41945 299 42391 333
rect 42425 299 42479 527
rect 42529 299 42583 527
rect 42617 333 42683 493
rect 42717 367 42771 527
rect 42805 333 42871 493
rect 42905 367 42959 527
rect 43003 333 43063 493
rect 42617 299 43063 333
rect 41657 213 41911 273
rect 43097 273 43163 815
rect 43197 595 43251 781
rect 43197 307 43251 493
rect 43285 273 43351 815
rect 43385 809 43622 875
rect 43656 823 43775 889
rect 43809 823 43928 889
rect 43962 875 43996 923
rect 44273 875 44339 969
rect 44373 934 44407 1003
rect 44441 911 44507 969
rect 44541 945 44595 1003
rect 44629 979 44679 1071
rect 44713 945 44779 1037
rect 44813 979 44867 1071
rect 44901 945 44967 1037
rect 44541 911 44967 945
rect 45001 911 45051 1071
rect 44441 875 44487 911
rect 43385 595 43445 775
rect 43588 767 43622 809
rect 43962 809 44199 875
rect 44233 815 44487 875
rect 44723 823 45001 877
rect 43962 767 43996 809
rect 43494 561 43549 767
rect 43588 595 43654 767
rect 43688 561 43748 767
rect 43836 561 43896 767
rect 43930 595 43996 767
rect 44035 561 44090 767
rect 44139 595 44199 775
rect 43385 527 44199 561
rect 43385 313 43445 493
rect 43494 321 43549 527
rect 43588 321 43654 493
rect 43688 321 43748 527
rect 43836 321 43896 527
rect 43930 321 43996 493
rect 44035 321 44090 527
rect 43588 279 43622 321
rect 41386 165 41420 213
rect 40769 85 40819 154
rect 40413 51 40819 85
rect 40920 17 40978 122
rect 41012 56 41062 165
rect 41104 17 41162 122
rect 41270 17 41328 122
rect 41370 56 41420 165
rect 41454 17 41512 122
rect 41613 85 41663 154
rect 41697 119 41763 213
rect 41865 177 41911 213
rect 42147 211 42425 265
rect 42583 211 42861 265
rect 43097 213 43351 273
rect 43385 213 43622 279
rect 43962 279 43996 321
rect 44139 313 44199 493
rect 43097 177 43143 213
rect 41797 85 41831 154
rect 41865 119 41931 177
rect 41965 143 42391 177
rect 41965 85 42019 143
rect 41613 51 42019 85
rect 42053 17 42103 109
rect 42137 51 42203 143
rect 42237 17 42291 109
rect 42325 51 42391 143
rect 42425 17 42475 177
rect 42533 17 42583 177
rect 42617 143 43043 177
rect 42617 51 42683 143
rect 42717 17 42771 109
rect 42805 51 42871 143
rect 42905 17 42955 109
rect 42989 85 43043 143
rect 43077 119 43143 177
rect 43177 85 43211 154
rect 43245 119 43311 213
rect 43588 165 43622 213
rect 43656 199 43775 265
rect 43809 199 43928 265
rect 43962 213 44199 279
rect 44233 273 44299 815
rect 44333 595 44387 781
rect 44333 307 44387 493
rect 44421 273 44487 815
rect 44521 755 44967 789
rect 44521 595 44581 755
rect 44625 561 44679 721
rect 44713 595 44779 755
rect 44813 561 44867 721
rect 44901 595 44967 755
rect 45001 561 45055 789
rect 44521 527 45080 561
rect 44521 333 44581 493
rect 44625 367 44679 527
rect 44713 333 44779 493
rect 44813 367 44867 527
rect 44901 333 44967 493
rect 44521 299 44967 333
rect 45001 299 45055 527
rect 44233 213 44487 273
rect 43962 165 43996 213
rect 43345 85 43395 154
rect 42989 51 43395 85
rect 43496 17 43554 122
rect 43588 56 43638 165
rect 43680 17 43738 122
rect 43846 17 43904 122
rect 43946 56 43996 165
rect 44030 17 44088 122
rect 44189 85 44239 154
rect 44273 119 44339 213
rect 44441 177 44487 213
rect 44723 211 45001 265
rect 44373 85 44407 154
rect 44441 119 44507 177
rect 44541 143 44967 177
rect 44541 85 44595 143
rect 44189 51 44595 85
rect 44629 17 44679 109
rect 44713 51 44779 143
rect 44813 17 44867 109
rect 44901 51 44967 143
rect 45001 17 45051 177
rect 0 -17 45080 17
<< obsm1 >>
rect 21160 1040 45080 1136
rect 21605 728 21663 737
rect 21793 728 21851 737
rect 22953 728 23011 737
rect 23141 728 23199 737
rect 24089 728 24147 737
rect 24277 728 24335 737
rect 25437 728 25495 737
rect 25625 728 25683 737
rect 21605 700 25683 728
rect 21605 691 21663 700
rect 21793 691 21851 700
rect 22953 691 23011 700
rect 23141 691 23199 700
rect 24089 691 24147 700
rect 24277 691 24335 700
rect 25437 691 25495 700
rect 25625 691 25683 700
rect 26329 728 26387 737
rect 26789 728 26847 737
rect 27157 728 27215 737
rect 27617 728 27675 737
rect 27985 728 28043 737
rect 28445 728 28503 737
rect 28813 728 28871 737
rect 29273 728 29331 737
rect 26329 700 29331 728
rect 26329 691 26387 700
rect 26789 691 26847 700
rect 27157 691 27215 700
rect 27617 691 27675 700
rect 27985 691 28043 700
rect 28445 691 28503 700
rect 28813 691 28871 700
rect 29273 691 29331 700
rect 29825 728 29883 737
rect 30469 728 30527 737
rect 31113 728 31171 737
rect 31757 728 31815 737
rect 32401 728 32459 737
rect 33045 728 33103 737
rect 33689 728 33747 737
rect 34333 728 34391 737
rect 29825 700 34391 728
rect 29825 691 29883 700
rect 30469 691 30527 700
rect 31113 691 31171 700
rect 31757 691 31815 700
rect 32401 691 32459 700
rect 33045 691 33103 700
rect 33689 691 33747 700
rect 34333 691 34391 700
rect 35281 728 35339 737
rect 35469 728 35527 737
rect 36417 728 36475 737
rect 36605 728 36663 737
rect 37857 728 37915 737
rect 38045 728 38103 737
rect 38993 728 39051 737
rect 39181 728 39239 737
rect 40525 728 40583 737
rect 40713 728 40771 737
rect 41661 728 41719 737
rect 41849 728 41907 737
rect 43101 728 43159 737
rect 43289 728 43347 737
rect 44237 728 44295 737
rect 44425 728 44483 737
rect 35281 700 44483 728
rect 35281 691 35339 700
rect 35469 691 35527 700
rect 36417 691 36475 700
rect 36605 691 36663 700
rect 37857 691 37915 700
rect 38045 691 38103 700
rect 38993 691 39051 700
rect 39181 691 39239 700
rect 40525 691 40583 700
rect 40713 691 40771 700
rect 41661 691 41719 700
rect 41849 691 41907 700
rect 43101 691 43159 700
rect 43289 691 43347 700
rect 44237 691 44295 700
rect 44425 691 44483 700
rect 21509 657 21567 666
rect 21699 657 21757 666
rect 21889 657 21947 666
rect 22085 657 22143 666
rect 22273 657 22331 666
rect 21509 629 22331 657
rect 21509 620 21567 629
rect 21699 620 21757 629
rect 21889 620 21947 629
rect 22085 620 22143 629
rect 22273 620 22331 629
rect 22473 657 22531 666
rect 22661 657 22719 666
rect 22857 657 22915 666
rect 23047 657 23105 666
rect 23237 657 23295 666
rect 22473 629 23295 657
rect 22473 620 22531 629
rect 22661 620 22719 629
rect 22857 620 22915 629
rect 23047 620 23105 629
rect 23237 620 23295 629
rect 23993 657 24051 666
rect 24183 657 24241 666
rect 24373 657 24431 666
rect 24569 657 24627 666
rect 24757 657 24815 666
rect 23993 629 24815 657
rect 23993 620 24051 629
rect 24183 620 24241 629
rect 24373 620 24431 629
rect 24569 620 24627 629
rect 24757 620 24815 629
rect 24957 657 25015 666
rect 25145 657 25203 666
rect 25341 657 25399 666
rect 25531 657 25589 666
rect 25721 657 25779 666
rect 24957 629 25779 657
rect 24957 620 25015 629
rect 25145 620 25203 629
rect 25341 620 25399 629
rect 25531 620 25589 629
rect 25721 620 25779 629
rect 29555 657 29613 666
rect 29743 657 29801 666
rect 29942 657 30000 666
rect 29555 629 30000 657
rect 29555 620 29613 629
rect 29743 620 29801 629
rect 29942 620 30000 629
rect 30352 657 30410 666
rect 30551 657 30609 666
rect 30739 657 30797 666
rect 30352 629 30797 657
rect 30352 620 30410 629
rect 30551 620 30609 629
rect 30739 620 30797 629
rect 30843 657 30901 666
rect 31031 657 31089 666
rect 31230 657 31288 666
rect 30843 629 31288 657
rect 30843 620 30901 629
rect 31031 620 31089 629
rect 31230 620 31288 629
rect 31640 657 31698 666
rect 31839 657 31897 666
rect 32027 657 32085 666
rect 31640 629 32085 657
rect 31640 620 31698 629
rect 31839 620 31897 629
rect 32027 620 32085 629
rect 32131 657 32189 666
rect 32319 657 32377 666
rect 32518 657 32576 666
rect 32131 629 32576 657
rect 32131 620 32189 629
rect 32319 620 32377 629
rect 32518 620 32576 629
rect 32928 657 32986 666
rect 33127 657 33185 666
rect 33315 657 33373 666
rect 32928 629 33373 657
rect 32928 620 32986 629
rect 33127 620 33185 629
rect 33315 620 33373 629
rect 33419 657 33477 666
rect 33607 657 33665 666
rect 33806 657 33864 666
rect 33419 629 33864 657
rect 33419 620 33477 629
rect 33607 620 33665 629
rect 33806 620 33864 629
rect 34216 657 34274 666
rect 34415 657 34473 666
rect 34603 657 34661 666
rect 34216 629 34661 657
rect 34216 620 34274 629
rect 34415 620 34473 629
rect 34603 620 34661 629
rect 34801 657 34859 666
rect 34989 657 35047 666
rect 35185 657 35243 666
rect 35375 657 35433 666
rect 35565 657 35623 666
rect 34801 629 35623 657
rect 34801 620 34859 629
rect 34989 620 35047 629
rect 35185 620 35243 629
rect 35375 620 35433 629
rect 35565 620 35623 629
rect 36321 657 36379 666
rect 36511 657 36569 666
rect 36701 657 36759 666
rect 36897 657 36955 666
rect 37085 657 37143 666
rect 36321 629 37143 657
rect 36321 620 36379 629
rect 36511 620 36569 629
rect 36701 620 36759 629
rect 36897 620 36955 629
rect 37085 620 37143 629
rect 37377 657 37435 666
rect 37565 657 37623 666
rect 37761 657 37819 666
rect 37951 657 38009 666
rect 38141 657 38199 666
rect 37377 629 38199 657
rect 37377 620 37435 629
rect 37565 620 37623 629
rect 37761 620 37819 629
rect 37951 620 38009 629
rect 38141 620 38199 629
rect 38897 657 38955 666
rect 39087 657 39145 666
rect 39277 657 39335 666
rect 39473 657 39531 666
rect 39661 657 39719 666
rect 38897 629 39719 657
rect 38897 620 38955 629
rect 39087 620 39145 629
rect 39277 620 39335 629
rect 39473 620 39531 629
rect 39661 620 39719 629
rect 40045 657 40103 666
rect 40233 657 40291 666
rect 40429 657 40487 666
rect 40619 657 40677 666
rect 40809 657 40867 666
rect 40045 629 40867 657
rect 40045 620 40103 629
rect 40233 620 40291 629
rect 40429 620 40487 629
rect 40619 620 40677 629
rect 40809 620 40867 629
rect 41565 657 41623 666
rect 41755 657 41813 666
rect 41945 657 42003 666
rect 42141 657 42199 666
rect 42329 657 42387 666
rect 41565 629 42387 657
rect 41565 620 41623 629
rect 41755 620 41813 629
rect 41945 620 42003 629
rect 42141 620 42199 629
rect 42329 620 42387 629
rect 42621 657 42679 666
rect 42809 657 42867 666
rect 43005 657 43063 666
rect 43195 657 43253 666
rect 43385 657 43443 666
rect 42621 629 43443 657
rect 42621 620 42679 629
rect 42809 620 42867 629
rect 43005 620 43063 629
rect 43195 620 43253 629
rect 43385 620 43443 629
rect 44141 657 44199 666
rect 44331 657 44389 666
rect 44521 657 44579 666
rect 44717 657 44775 666
rect 44905 657 44963 666
rect 44141 629 44963 657
rect 44141 620 44199 629
rect 44331 620 44389 629
rect 44521 620 44579 629
rect 44717 620 44775 629
rect 44905 620 44963 629
rect 0 496 45080 592
rect 21509 459 21567 468
rect 21699 459 21757 468
rect 21889 459 21947 468
rect 22085 459 22143 468
rect 22273 459 22331 468
rect 21509 431 22331 459
rect 21509 422 21567 431
rect 21699 422 21757 431
rect 21889 422 21947 431
rect 22085 422 22143 431
rect 22273 422 22331 431
rect 22473 459 22531 468
rect 22661 459 22719 468
rect 22857 459 22915 468
rect 23047 459 23105 468
rect 23237 459 23295 468
rect 22473 431 23295 459
rect 22473 422 22531 431
rect 22661 422 22719 431
rect 22857 422 22915 431
rect 23047 422 23105 431
rect 23237 422 23295 431
rect 23993 459 24051 468
rect 24183 459 24241 468
rect 24373 459 24431 468
rect 24569 459 24627 468
rect 24757 459 24815 468
rect 23993 431 24815 459
rect 23993 422 24051 431
rect 24183 422 24241 431
rect 24373 422 24431 431
rect 24569 422 24627 431
rect 24757 422 24815 431
rect 24957 459 25015 468
rect 25145 459 25203 468
rect 25341 459 25399 468
rect 25531 459 25589 468
rect 25721 459 25779 468
rect 24957 431 25779 459
rect 24957 422 25015 431
rect 25145 422 25203 431
rect 25341 422 25399 431
rect 25531 422 25589 431
rect 25721 422 25779 431
rect 29555 459 29613 468
rect 29743 459 29801 468
rect 29942 459 30000 468
rect 29555 431 30000 459
rect 29555 422 29613 431
rect 29743 422 29801 431
rect 29942 422 30000 431
rect 30352 459 30410 468
rect 30551 459 30609 468
rect 30739 459 30797 468
rect 30352 431 30797 459
rect 30352 422 30410 431
rect 30551 422 30609 431
rect 30739 422 30797 431
rect 30843 459 30901 468
rect 31031 459 31089 468
rect 31230 459 31288 468
rect 30843 431 31288 459
rect 30843 422 30901 431
rect 31031 422 31089 431
rect 31230 422 31288 431
rect 31640 459 31698 468
rect 31839 459 31897 468
rect 32027 459 32085 468
rect 31640 431 32085 459
rect 31640 422 31698 431
rect 31839 422 31897 431
rect 32027 422 32085 431
rect 32131 459 32189 468
rect 32319 459 32377 468
rect 32518 459 32576 468
rect 32131 431 32576 459
rect 32131 422 32189 431
rect 32319 422 32377 431
rect 32518 422 32576 431
rect 32928 459 32986 468
rect 33127 459 33185 468
rect 33315 459 33373 468
rect 32928 431 33373 459
rect 32928 422 32986 431
rect 33127 422 33185 431
rect 33315 422 33373 431
rect 33419 459 33477 468
rect 33607 459 33665 468
rect 33806 459 33864 468
rect 33419 431 33864 459
rect 33419 422 33477 431
rect 33607 422 33665 431
rect 33806 422 33864 431
rect 34216 459 34274 468
rect 34415 459 34473 468
rect 34603 459 34661 468
rect 34216 431 34661 459
rect 34216 422 34274 431
rect 34415 422 34473 431
rect 34603 422 34661 431
rect 34801 459 34859 468
rect 34989 459 35047 468
rect 35185 459 35243 468
rect 35375 459 35433 468
rect 35565 459 35623 468
rect 34801 431 35623 459
rect 34801 422 34859 431
rect 34989 422 35047 431
rect 35185 422 35243 431
rect 35375 422 35433 431
rect 35565 422 35623 431
rect 36321 459 36379 468
rect 36511 459 36569 468
rect 36701 459 36759 468
rect 36897 459 36955 468
rect 37085 459 37143 468
rect 36321 431 37143 459
rect 36321 422 36379 431
rect 36511 422 36569 431
rect 36701 422 36759 431
rect 36897 422 36955 431
rect 37085 422 37143 431
rect 37377 459 37435 468
rect 37565 459 37623 468
rect 37761 459 37819 468
rect 37951 459 38009 468
rect 38141 459 38199 468
rect 37377 431 38199 459
rect 37377 422 37435 431
rect 37565 422 37623 431
rect 37761 422 37819 431
rect 37951 422 38009 431
rect 38141 422 38199 431
rect 38897 459 38955 468
rect 39087 459 39145 468
rect 39277 459 39335 468
rect 39473 459 39531 468
rect 39661 459 39719 468
rect 38897 431 39719 459
rect 38897 422 38955 431
rect 39087 422 39145 431
rect 39277 422 39335 431
rect 39473 422 39531 431
rect 39661 422 39719 431
rect 40045 459 40103 468
rect 40233 459 40291 468
rect 40429 459 40487 468
rect 40619 459 40677 468
rect 40809 459 40867 468
rect 40045 431 40867 459
rect 40045 422 40103 431
rect 40233 422 40291 431
rect 40429 422 40487 431
rect 40619 422 40677 431
rect 40809 422 40867 431
rect 41565 459 41623 468
rect 41755 459 41813 468
rect 41945 459 42003 468
rect 42141 459 42199 468
rect 42329 459 42387 468
rect 41565 431 42387 459
rect 41565 422 41623 431
rect 41755 422 41813 431
rect 41945 422 42003 431
rect 42141 422 42199 431
rect 42329 422 42387 431
rect 42621 459 42679 468
rect 42809 459 42867 468
rect 43005 459 43063 468
rect 43195 459 43253 468
rect 43385 459 43443 468
rect 42621 431 43443 459
rect 42621 422 42679 431
rect 42809 422 42867 431
rect 43005 422 43063 431
rect 43195 422 43253 431
rect 43385 422 43443 431
rect 44141 459 44199 468
rect 44331 459 44389 468
rect 44521 459 44579 468
rect 44717 459 44775 468
rect 44905 459 44963 468
rect 44141 431 44963 459
rect 44141 422 44199 431
rect 44331 422 44389 431
rect 44521 422 44579 431
rect 44717 422 44775 431
rect 44905 422 44963 431
rect 3329 388 3387 397
rect 3789 388 3847 397
rect 4157 388 4215 397
rect 4617 388 4675 397
rect 3329 360 4675 388
rect 3329 351 3387 360
rect 3789 351 3847 360
rect 4157 351 4215 360
rect 4617 351 4675 360
rect 5169 388 5227 397
rect 5813 388 5871 397
rect 6457 388 6515 397
rect 7101 388 7159 397
rect 5169 360 7159 388
rect 5169 351 5227 360
rect 5813 351 5871 360
rect 6457 351 6515 360
rect 7101 351 7159 360
rect 8049 388 8107 397
rect 8237 388 8295 397
rect 9185 388 9243 397
rect 9373 388 9431 397
rect 10625 388 10683 397
rect 10813 388 10871 397
rect 11761 388 11819 397
rect 11949 388 12007 397
rect 8049 360 12007 388
rect 8049 351 8107 360
rect 8237 351 8295 360
rect 9185 351 9243 360
rect 9373 351 9431 360
rect 10625 351 10683 360
rect 10813 351 10871 360
rect 11761 351 11819 360
rect 11949 351 12007 360
rect 12805 388 12863 397
rect 13265 388 13323 397
rect 13633 388 13691 397
rect 14093 388 14151 397
rect 14461 388 14519 397
rect 14921 388 14979 397
rect 15289 388 15347 397
rect 15749 388 15807 397
rect 12805 360 15807 388
rect 12805 351 12863 360
rect 13265 351 13323 360
rect 13633 351 13691 360
rect 14093 351 14151 360
rect 14461 351 14519 360
rect 14921 351 14979 360
rect 15289 351 15347 360
rect 15749 351 15807 360
rect 16301 388 16359 397
rect 16945 388 17003 397
rect 17589 388 17647 397
rect 18233 388 18291 397
rect 18877 388 18935 397
rect 19521 388 19579 397
rect 20165 388 20223 397
rect 20809 388 20867 397
rect 16301 360 20867 388
rect 16301 351 16359 360
rect 16945 351 17003 360
rect 17589 351 17647 360
rect 18233 351 18291 360
rect 18877 351 18935 360
rect 19521 351 19579 360
rect 20165 351 20223 360
rect 20809 351 20867 360
rect 21605 388 21663 397
rect 21793 388 21851 397
rect 22953 388 23011 397
rect 23141 388 23199 397
rect 24089 388 24147 397
rect 24277 388 24335 397
rect 25437 388 25495 397
rect 25625 388 25683 397
rect 21605 360 25683 388
rect 21605 351 21663 360
rect 21793 351 21851 360
rect 22953 351 23011 360
rect 23141 351 23199 360
rect 24089 351 24147 360
rect 24277 351 24335 360
rect 25437 351 25495 360
rect 25625 351 25683 360
rect 26329 388 26387 397
rect 26789 388 26847 397
rect 27157 388 27215 397
rect 27617 388 27675 397
rect 27985 388 28043 397
rect 28445 388 28503 397
rect 28813 388 28871 397
rect 29273 388 29331 397
rect 26329 360 29331 388
rect 26329 351 26387 360
rect 26789 351 26847 360
rect 27157 351 27215 360
rect 27617 351 27675 360
rect 27985 351 28043 360
rect 28445 351 28503 360
rect 28813 351 28871 360
rect 29273 351 29331 360
rect 29825 388 29883 397
rect 30469 388 30527 397
rect 31113 388 31171 397
rect 31757 388 31815 397
rect 32401 388 32459 397
rect 33045 388 33103 397
rect 33689 388 33747 397
rect 34333 388 34391 397
rect 29825 360 34391 388
rect 29825 351 29883 360
rect 30469 351 30527 360
rect 31113 351 31171 360
rect 31757 351 31815 360
rect 32401 351 32459 360
rect 33045 351 33103 360
rect 33689 351 33747 360
rect 34333 351 34391 360
rect 35281 388 35339 397
rect 35469 388 35527 397
rect 36417 388 36475 397
rect 36605 388 36663 397
rect 37857 388 37915 397
rect 38045 388 38103 397
rect 38993 388 39051 397
rect 39181 388 39239 397
rect 40525 388 40583 397
rect 40713 388 40771 397
rect 41661 388 41719 397
rect 41849 388 41907 397
rect 43101 388 43159 397
rect 43289 388 43347 397
rect 44237 388 44295 397
rect 44425 388 44483 397
rect 35281 360 44483 388
rect 35281 351 35339 360
rect 35469 351 35527 360
rect 36417 351 36475 360
rect 36605 351 36663 360
rect 37857 351 37915 360
rect 38045 351 38103 360
rect 38993 351 39051 360
rect 39181 351 39239 360
rect 40525 351 40583 360
rect 40713 351 40771 360
rect 41661 351 41719 360
rect 41849 351 41907 360
rect 43101 351 43159 360
rect 43289 351 43347 360
rect 44237 351 44295 360
rect 44425 351 44483 360
rect 0 -48 45080 48
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX -38 -48 45118 1136
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3646992
string GDS_START 3646346
<< end >>
