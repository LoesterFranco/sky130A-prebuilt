magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 2576 561
rect 103 439 157 527
rect 538 428 597 527
rect 17 153 68 335
rect 108 153 164 335
rect 210 153 267 335
rect 719 455 785 527
rect 581 323 617 392
rect 474 215 540 320
rect 581 211 713 323
rect 581 145 620 211
rect 17 17 140 119
rect 365 17 418 109
rect 1189 455 1266 527
rect 538 17 620 111
rect 1412 425 1603 527
rect 1832 447 1898 527
rect 2031 447 2097 527
rect 1328 289 1413 353
rect 725 17 791 109
rect 1776 309 1989 345
rect 1776 285 1827 309
rect 1122 17 1219 93
rect 1341 17 1543 161
rect 2023 17 2073 109
rect 2314 358 2364 527
rect 2407 299 2473 490
rect 2507 299 2559 527
rect 2429 165 2473 299
rect 2314 17 2373 165
rect 2407 51 2473 165
rect 2507 17 2559 177
rect 0 -17 2576 17
<< obsli1 >>
rect 17 405 69 493
rect 191 451 409 493
rect 191 405 225 451
rect 454 417 504 493
rect 17 369 225 405
rect 259 369 339 417
rect 301 323 339 369
rect 301 289 305 323
rect 301 142 339 289
rect 373 354 504 417
rect 651 400 685 465
rect 819 427 888 493
rect 651 398 797 400
rect 373 181 440 354
rect 651 391 799 398
rect 651 366 765 391
rect 747 357 765 366
rect 373 143 504 181
rect 747 177 799 357
rect 301 141 335 142
rect 299 133 335 141
rect 295 132 335 133
rect 295 129 334 132
rect 292 127 333 129
rect 289 126 333 127
rect 288 124 333 126
rect 286 123 332 124
rect 284 122 332 123
rect 281 121 332 122
rect 279 120 332 121
rect 276 119 332 120
rect 174 115 330 119
rect 174 111 328 115
rect 174 51 325 111
rect 452 51 504 143
rect 654 143 799 177
rect 833 284 888 427
rect 923 323 966 493
rect 1007 427 1151 493
rect 1075 357 1083 391
rect 923 318 949 323
rect 932 289 949 318
rect 1041 315 1083 357
rect 833 255 898 284
rect 833 221 857 255
rect 891 221 898 255
rect 833 218 898 221
rect 654 51 691 143
rect 833 117 867 218
rect 932 184 966 289
rect 1117 279 1151 427
rect 1321 421 1364 490
rect 1637 425 1798 492
rect 1185 387 1364 421
rect 1764 413 1798 425
rect 1932 413 1993 490
rect 1185 315 1219 387
rect 1447 357 1512 391
rect 1546 357 1627 391
rect 1447 334 1627 357
rect 1017 255 1295 279
rect 1471 255 1543 265
rect 825 51 867 117
rect 901 51 966 184
rect 1000 245 1543 255
rect 1000 51 1088 245
rect 1129 161 1195 203
rect 1261 195 1543 245
rect 1577 181 1627 334
rect 1685 255 1730 381
rect 1764 379 2097 413
rect 2031 321 2097 379
rect 2131 273 2183 493
rect 1685 221 1696 255
rect 1685 215 1730 221
rect 1764 181 1821 251
rect 1129 127 1307 161
rect 1257 51 1307 127
rect 1577 144 1821 181
rect 1864 239 2183 273
rect 1864 171 1906 239
rect 1942 157 2103 203
rect 1942 109 1982 157
rect 2137 117 2183 239
rect 1693 55 1982 109
rect 2115 51 2183 117
rect 2217 265 2269 493
rect 2217 199 2395 265
rect 2217 51 2269 199
<< obsli1c >>
rect 305 289 339 323
rect 765 357 799 391
rect 1041 357 1075 391
rect 949 289 983 323
rect 857 221 891 255
rect 1512 357 1546 391
rect 1696 221 1730 255
<< metal1 >>
rect 0 496 2576 592
rect 1316 320 1374 329
rect 1776 320 1834 329
rect 1316 292 1834 320
rect 1316 283 1374 292
rect 1776 283 1834 292
rect 109 252 167 261
rect 477 252 535 261
rect 109 224 535 252
rect 109 215 167 224
rect 477 215 535 224
rect 0 -48 2576 48
<< obsm1 >>
rect 753 391 811 397
rect 753 357 765 391
rect 799 388 811 391
rect 1029 391 1087 397
rect 1029 388 1041 391
rect 799 360 1041 388
rect 799 357 811 360
rect 753 351 811 357
rect 1029 357 1041 360
rect 1075 388 1087 391
rect 1500 391 1558 397
rect 1500 388 1512 391
rect 1075 360 1512 388
rect 1075 357 1087 360
rect 1029 351 1087 357
rect 1500 357 1512 360
rect 1546 357 1558 391
rect 1500 351 1558 357
rect 293 323 351 329
rect 293 289 305 323
rect 339 320 351 323
rect 937 323 995 329
rect 937 320 949 323
rect 339 292 949 320
rect 339 289 351 292
rect 293 283 351 289
rect 937 289 949 292
rect 983 289 995 323
rect 937 283 995 289
rect 845 255 903 261
rect 845 221 857 255
rect 891 252 903 255
rect 1684 255 1742 261
rect 1684 252 1696 255
rect 891 224 1696 252
rect 891 221 903 224
rect 845 215 903 221
rect 1684 221 1696 224
rect 1730 221 1742 255
rect 1684 215 1742 221
<< labels >>
rlabel locali s 210 153 267 335 6 D
port 1 nsew signal input
rlabel locali s 2429 165 2473 299 6 Q
port 2 nsew signal output
rlabel locali s 2407 299 2473 490 6 Q
port 2 nsew signal output
rlabel locali s 2407 51 2473 165 6 Q
port 2 nsew signal output
rlabel locali s 17 153 68 335 6 SCD
port 3 nsew signal input
rlabel locali s 108 153 164 335 6 SCE
port 4 nsew signal input
rlabel locali s 474 215 540 320 6 SCE
port 4 nsew signal input
rlabel metal1 s 477 252 535 261 6 SCE
port 4 nsew signal input
rlabel metal1 s 477 215 535 224 6 SCE
port 4 nsew signal input
rlabel metal1 s 109 252 167 261 6 SCE
port 4 nsew signal input
rlabel metal1 s 109 224 535 252 6 SCE
port 4 nsew signal input
rlabel metal1 s 109 215 167 224 6 SCE
port 4 nsew signal input
rlabel locali s 1328 289 1413 353 6 SET_B
port 5 nsew signal input
rlabel locali s 1776 309 1989 345 6 SET_B
port 5 nsew signal input
rlabel locali s 1776 285 1827 309 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1776 320 1834 329 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1776 283 1834 292 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1316 320 1374 329 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1316 292 1834 320 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1316 283 1374 292 6 SET_B
port 5 nsew signal input
rlabel locali s 581 323 617 392 6 CLK
port 6 nsew clock input
rlabel locali s 581 211 713 323 6 CLK
port 6 nsew clock input
rlabel locali s 581 145 620 211 6 CLK
port 6 nsew clock input
rlabel locali s 2507 17 2559 177 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 2314 17 2373 165 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 2023 17 2073 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1341 17 1543 161 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1122 17 1219 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 725 17 791 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 538 17 620 111 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 365 17 418 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 17 17 140 119 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 2576 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 2576 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 2507 299 2559 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 2314 358 2364 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 2031 447 2097 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1832 447 1898 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1412 425 1603 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1189 455 1266 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 719 455 785 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 538 428 597 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 103 439 157 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 2576 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 2576 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2576 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 304536
string GDS_START 284032
<< end >>
