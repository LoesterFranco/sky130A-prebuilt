magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 25 290 178 356
rect 217 294 471 360
rect 1459 287 1703 355
rect 1753 252 1895 355
rect 1945 289 2087 355
rect 2430 260 2567 356
rect 2975 394 3041 596
rect 3165 394 3231 596
rect 2975 360 3335 394
rect 2708 260 2773 310
rect 2430 255 2773 260
rect 2533 226 2773 255
rect 3289 226 3335 360
rect 3013 192 3335 226
rect 3013 70 3063 192
rect 3185 70 3235 192
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3360 683
rect 23 390 73 649
rect 113 428 179 596
rect 219 462 269 649
rect 303 496 369 596
rect 409 530 459 649
rect 505 581 944 615
rect 505 530 572 581
rect 609 496 660 547
rect 303 462 660 496
rect 113 394 539 428
rect 113 390 179 394
rect 505 354 539 394
rect 598 388 660 462
rect 698 388 764 581
rect 804 354 838 547
rect 505 320 838 354
rect 875 384 944 581
rect 505 260 841 286
rect 23 206 274 256
rect 23 17 73 206
rect 109 94 175 172
rect 209 128 274 206
rect 310 252 841 260
rect 310 226 539 252
rect 310 192 360 226
rect 610 192 676 218
rect 394 158 676 192
rect 315 124 428 158
rect 315 94 362 124
rect 109 55 362 94
rect 396 17 462 90
rect 508 85 574 124
rect 610 119 676 158
rect 721 85 755 218
rect 791 119 841 252
rect 875 236 909 384
rect 990 336 1040 596
rect 1080 364 1146 649
rect 1282 581 1630 615
rect 1664 593 1730 649
rect 1878 593 1946 649
rect 1192 407 1242 581
rect 1282 441 1348 581
rect 1596 559 1630 581
rect 1987 559 2053 596
rect 1388 423 1425 547
rect 1462 491 1528 547
rect 1596 525 2053 559
rect 1462 457 1837 491
rect 1987 457 2053 525
rect 2093 457 2127 649
rect 2161 581 2595 615
rect 2161 423 2195 581
rect 1388 407 2195 423
rect 1192 389 2195 407
rect 2229 513 2495 547
rect 1192 373 1425 389
rect 943 307 1040 336
rect 1207 307 1341 339
rect 943 273 1341 307
rect 943 270 1040 273
rect 875 85 943 236
rect 508 51 943 85
rect 989 70 1040 270
rect 1388 253 1425 373
rect 1375 239 1425 253
rect 1075 17 1141 226
rect 1187 205 1425 239
rect 1187 117 1237 205
rect 1273 85 1339 171
rect 1375 153 1425 205
rect 1461 219 1665 253
rect 1461 187 1511 219
rect 1631 218 1665 219
rect 1547 153 1597 185
rect 1631 184 2023 218
rect 1375 119 1597 153
rect 1631 116 1851 150
rect 1631 85 1665 116
rect 1273 51 1665 85
rect 1699 17 1765 82
rect 1801 70 1851 116
rect 1887 17 1937 150
rect 1973 70 2023 184
rect 2059 17 2109 206
rect 2143 85 2177 389
rect 2229 206 2295 513
rect 2211 153 2295 206
rect 2329 221 2395 479
rect 2429 446 2495 513
rect 2529 480 2595 581
rect 2629 446 2695 596
rect 2429 412 2695 446
rect 2429 390 2495 412
rect 2775 378 2841 596
rect 2601 344 2841 378
rect 2875 364 2941 649
rect 3081 428 3131 649
rect 3265 428 3331 649
rect 2601 294 2666 344
rect 2329 192 2499 221
rect 2807 192 2841 344
rect 2329 187 2635 192
rect 2465 158 2635 187
rect 2211 124 2431 153
rect 2211 119 2535 124
rect 2572 119 2635 158
rect 2397 85 2535 119
rect 2669 85 2735 192
rect 2781 119 2841 192
rect 2875 260 3242 326
rect 2875 85 2909 260
rect 2143 51 2363 85
rect 2397 51 2909 85
rect 2943 17 2977 226
rect 3099 17 3149 158
rect 3271 17 3337 158
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3360 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 3199 649 3233 683
rect 3295 649 3329 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
<< metal1 >>
rect 0 683 3360 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3360 683
rect 0 617 3360 649
rect 0 17 3360 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3360 17
rect 0 -49 3360 -17
<< obsm1 >>
rect 883 421 941 430
rect 2323 421 2381 430
rect 883 393 2381 421
rect 883 384 941 393
rect 2323 384 2381 393
<< labels >>
rlabel locali s 217 294 471 360 6 A0
port 1 nsew signal input
rlabel locali s 25 290 178 356 6 A1
port 2 nsew signal input
rlabel locali s 1753 252 1895 355 6 A2
port 3 nsew signal input
rlabel locali s 1945 289 2087 355 6 A3
port 4 nsew signal input
rlabel locali s 1459 287 1703 355 6 S0
port 5 nsew signal input
rlabel locali s 2708 260 2773 310 6 S1
port 6 nsew signal input
rlabel locali s 2533 226 2773 255 6 S1
port 6 nsew signal input
rlabel locali s 2430 260 2567 356 6 S1
port 6 nsew signal input
rlabel locali s 2430 255 2773 260 6 S1
port 6 nsew signal input
rlabel locali s 3289 226 3335 360 6 X
port 7 nsew signal output
rlabel locali s 3185 70 3235 192 6 X
port 7 nsew signal output
rlabel locali s 3165 394 3231 596 6 X
port 7 nsew signal output
rlabel locali s 3013 192 3335 226 6 X
port 7 nsew signal output
rlabel locali s 3013 70 3063 192 6 X
port 7 nsew signal output
rlabel locali s 2975 394 3041 596 6 X
port 7 nsew signal output
rlabel locali s 2975 360 3335 394 6 X
port 7 nsew signal output
rlabel metal1 s 0 -49 3360 49 8 VGND
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 617 3360 715 6 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 3360 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1725522
string GDS_START 1700548
<< end >>
