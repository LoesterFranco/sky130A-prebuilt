magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1104 561
rect 103 441 169 527
rect 85 199 155 339
rect 189 199 247 265
rect 131 17 165 165
rect 559 357 623 475
rect 680 359 730 527
rect 559 290 601 357
rect 775 325 825 493
rect 859 359 909 527
rect 943 325 993 493
rect 1027 359 1077 527
rect 535 199 601 290
rect 647 289 734 323
rect 775 291 1087 325
rect 647 199 681 289
rect 1041 181 1087 291
rect 783 145 1087 181
rect 303 17 369 96
rect 493 17 559 97
rect 671 17 747 97
rect 783 51 833 145
rect 867 17 901 111
rect 935 51 1001 145
rect 1035 17 1069 111
rect 0 -17 1104 17
<< obsli1 >>
rect 17 407 69 491
rect 225 459 489 493
rect 225 407 259 459
rect 17 373 259 407
rect 302 391 421 425
rect 17 165 51 373
rect 198 305 319 339
rect 281 265 319 305
rect 281 199 339 265
rect 281 165 319 199
rect 17 90 80 165
rect 215 131 319 165
rect 387 165 421 391
rect 455 199 489 459
rect 715 215 1007 249
rect 715 165 749 215
rect 387 131 749 165
rect 215 90 249 131
rect 419 61 453 131
rect 593 61 627 131
<< metal1 >>
rect 0 496 1104 592
rect 0 -48 1104 48
<< labels >>
rlabel locali s 647 289 734 323 6 A
port 1 nsew signal input
rlabel locali s 647 199 681 289 6 A
port 1 nsew signal input
rlabel locali s 559 357 623 475 6 B
port 2 nsew signal input
rlabel locali s 559 290 601 357 6 B
port 2 nsew signal input
rlabel locali s 535 199 601 290 6 B
port 2 nsew signal input
rlabel locali s 85 199 155 339 6 C_N
port 3 nsew signal input
rlabel locali s 189 199 247 265 6 D_N
port 4 nsew signal input
rlabel locali s 1041 181 1087 291 6 X
port 5 nsew signal output
rlabel locali s 943 325 993 493 6 X
port 5 nsew signal output
rlabel locali s 935 51 1001 145 6 X
port 5 nsew signal output
rlabel locali s 783 145 1087 181 6 X
port 5 nsew signal output
rlabel locali s 783 51 833 145 6 X
port 5 nsew signal output
rlabel locali s 775 325 825 493 6 X
port 5 nsew signal output
rlabel locali s 775 291 1087 325 6 X
port 5 nsew signal output
rlabel locali s 1035 17 1069 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 867 17 901 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 671 17 747 97 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 493 17 559 97 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 303 17 369 96 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 131 17 165 165 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 1104 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1104 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1027 359 1077 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 859 359 909 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 680 359 730 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 103 441 169 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 1104 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 1104 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1104 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 8888
string GDS_START 130
<< end >>
