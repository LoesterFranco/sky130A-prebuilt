magic
tech sky130A
magscale 1 2
timestamp 1604502697
<< nwell >>
rect -38 261 1326 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 82 47 112 177
rect 186 47 216 177
rect 270 47 300 177
rect 364 47 394 177
rect 570 47 600 177
rect 674 47 704 177
rect 758 47 788 177
rect 869 47 899 177
rect 1057 47 1087 177
rect 1161 47 1191 177
<< pmoshvt >>
rect 84 297 120 497
rect 178 297 214 497
rect 272 297 308 497
rect 366 297 402 497
rect 572 297 608 497
rect 666 297 702 497
rect 760 297 796 497
rect 861 297 897 497
rect 1059 297 1095 497
rect 1153 297 1189 497
<< ndiff >>
rect 27 95 82 177
rect 27 61 38 95
rect 72 61 82 95
rect 27 47 82 61
rect 112 163 186 177
rect 112 129 132 163
rect 166 129 186 163
rect 112 47 186 129
rect 216 163 270 177
rect 216 129 226 163
rect 260 129 270 163
rect 216 95 270 129
rect 216 61 226 95
rect 260 61 270 95
rect 216 47 270 61
rect 300 95 364 177
rect 300 61 320 95
rect 354 61 364 95
rect 300 47 364 61
rect 394 163 460 177
rect 394 129 414 163
rect 448 129 460 163
rect 394 95 460 129
rect 394 61 414 95
rect 448 61 460 95
rect 394 47 460 61
rect 514 163 570 177
rect 514 129 526 163
rect 560 129 570 163
rect 514 95 570 129
rect 514 61 526 95
rect 560 61 570 95
rect 514 47 570 61
rect 600 163 674 177
rect 600 129 620 163
rect 654 129 674 163
rect 600 95 674 129
rect 600 61 620 95
rect 654 61 674 95
rect 600 47 674 61
rect 704 95 758 177
rect 704 61 714 95
rect 748 61 758 95
rect 704 47 758 61
rect 788 163 869 177
rect 788 129 815 163
rect 849 129 869 163
rect 788 95 869 129
rect 788 61 815 95
rect 849 61 869 95
rect 788 47 869 61
rect 899 95 951 177
rect 899 61 909 95
rect 943 61 951 95
rect 899 47 951 61
rect 1005 95 1057 177
rect 1005 61 1013 95
rect 1047 61 1057 95
rect 1005 47 1057 61
rect 1087 163 1161 177
rect 1087 129 1097 163
rect 1131 129 1161 163
rect 1087 47 1161 129
rect 1191 163 1243 177
rect 1191 129 1201 163
rect 1235 129 1243 163
rect 1191 95 1243 129
rect 1191 61 1201 95
rect 1235 61 1243 95
rect 1191 47 1243 61
<< pdiff >>
rect 27 477 84 497
rect 27 443 38 477
rect 72 443 84 477
rect 27 409 84 443
rect 27 375 38 409
rect 72 375 84 409
rect 27 297 84 375
rect 120 477 178 497
rect 120 443 132 477
rect 166 443 178 477
rect 120 297 178 443
rect 214 477 272 497
rect 214 443 226 477
rect 260 443 272 477
rect 214 409 272 443
rect 214 375 226 409
rect 260 375 272 409
rect 214 297 272 375
rect 308 477 366 497
rect 308 443 320 477
rect 354 443 366 477
rect 308 297 366 443
rect 402 477 460 497
rect 402 443 414 477
rect 448 443 460 477
rect 402 409 460 443
rect 402 375 414 409
rect 448 375 460 409
rect 402 297 460 375
rect 514 477 572 497
rect 514 443 526 477
rect 560 443 572 477
rect 514 297 572 443
rect 608 477 666 497
rect 608 443 620 477
rect 654 443 666 477
rect 608 297 666 443
rect 702 477 760 497
rect 702 443 714 477
rect 748 443 760 477
rect 702 297 760 443
rect 796 409 861 497
rect 796 375 815 409
rect 849 375 861 409
rect 796 297 861 375
rect 897 477 951 497
rect 897 443 909 477
rect 943 443 951 477
rect 897 297 951 443
rect 1005 477 1059 497
rect 1005 443 1013 477
rect 1047 443 1059 477
rect 1005 297 1059 443
rect 1095 409 1153 497
rect 1095 375 1107 409
rect 1141 375 1153 409
rect 1095 341 1153 375
rect 1095 307 1107 341
rect 1141 307 1153 341
rect 1095 297 1153 307
rect 1189 477 1247 497
rect 1189 443 1201 477
rect 1235 443 1247 477
rect 1189 409 1247 443
rect 1189 375 1201 409
rect 1235 375 1247 409
rect 1189 297 1247 375
<< ndiffc >>
rect 38 61 72 95
rect 132 129 166 163
rect 226 129 260 163
rect 226 61 260 95
rect 320 61 354 95
rect 414 129 448 163
rect 414 61 448 95
rect 526 129 560 163
rect 526 61 560 95
rect 620 129 654 163
rect 620 61 654 95
rect 714 61 748 95
rect 815 129 849 163
rect 815 61 849 95
rect 909 61 943 95
rect 1013 61 1047 95
rect 1097 129 1131 163
rect 1201 129 1235 163
rect 1201 61 1235 95
<< pdiffc >>
rect 38 443 72 477
rect 38 375 72 409
rect 132 443 166 477
rect 226 443 260 477
rect 226 375 260 409
rect 320 443 354 477
rect 414 443 448 477
rect 414 375 448 409
rect 526 443 560 477
rect 620 443 654 477
rect 714 443 748 477
rect 815 375 849 409
rect 909 443 943 477
rect 1013 443 1047 477
rect 1107 375 1141 409
rect 1107 307 1141 341
rect 1201 443 1235 477
rect 1201 375 1235 409
<< poly >>
rect 84 497 120 523
rect 178 497 214 523
rect 272 497 308 523
rect 366 497 402 523
rect 572 497 608 523
rect 666 497 702 523
rect 760 497 796 523
rect 861 497 897 523
rect 1059 497 1095 523
rect 1153 497 1189 523
rect 84 282 120 297
rect 178 282 214 297
rect 272 282 308 297
rect 366 282 402 297
rect 572 282 608 297
rect 666 282 702 297
rect 760 282 796 297
rect 861 282 897 297
rect 1059 282 1095 297
rect 1153 282 1189 297
rect 82 265 122 282
rect 176 265 216 282
rect 82 249 216 265
rect 82 215 123 249
rect 157 215 216 249
rect 82 199 216 215
rect 82 177 112 199
rect 186 177 216 199
rect 270 265 310 282
rect 364 265 404 282
rect 570 265 610 282
rect 664 265 704 282
rect 270 249 704 265
rect 270 215 287 249
rect 321 215 365 249
rect 399 215 443 249
rect 477 215 515 249
rect 549 215 704 249
rect 270 199 704 215
rect 270 177 300 199
rect 364 177 394 199
rect 570 177 600 199
rect 674 177 704 199
rect 758 265 798 282
rect 859 265 899 282
rect 758 249 899 265
rect 758 215 804 249
rect 838 215 899 249
rect 758 199 899 215
rect 758 177 788 199
rect 869 177 899 199
rect 1057 265 1097 282
rect 1151 265 1191 282
rect 1057 249 1191 265
rect 1057 215 1099 249
rect 1133 215 1191 249
rect 1057 199 1191 215
rect 1057 177 1087 199
rect 1161 177 1191 199
rect 82 21 112 47
rect 186 21 216 47
rect 270 21 300 47
rect 364 21 394 47
rect 570 21 600 47
rect 674 21 704 47
rect 758 21 788 47
rect 869 21 899 47
rect 1057 21 1087 47
rect 1161 21 1191 47
<< polycont >>
rect 123 215 157 249
rect 287 215 321 249
rect 365 215 399 249
rect 443 215 477 249
rect 515 215 549 249
rect 804 215 838 249
rect 1099 215 1133 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 17 477 80 493
rect 17 443 38 477
rect 72 443 80 477
rect 17 409 80 443
rect 124 477 174 527
rect 124 443 132 477
rect 166 443 174 477
rect 124 427 174 443
rect 218 477 268 493
rect 218 443 226 477
rect 260 443 268 477
rect 17 375 38 409
rect 72 393 80 409
rect 218 409 268 443
rect 312 477 362 527
rect 312 443 320 477
rect 354 443 362 477
rect 312 427 362 443
rect 406 477 456 493
rect 406 443 414 477
rect 448 443 456 477
rect 218 393 226 409
rect 72 375 226 393
rect 260 393 268 409
rect 406 409 456 443
rect 518 477 568 493
rect 518 443 526 477
rect 560 459 568 477
rect 518 425 533 443
rect 567 425 568 459
rect 612 477 662 527
rect 612 443 620 477
rect 654 443 662 477
rect 612 427 662 443
rect 706 477 951 493
rect 706 443 714 477
rect 748 459 909 477
rect 706 425 737 443
rect 901 443 909 459
rect 943 443 951 477
rect 901 427 951 443
rect 1005 477 1055 527
rect 1005 443 1013 477
rect 1047 443 1055 477
rect 1005 427 1055 443
rect 1193 477 1268 527
rect 1193 443 1201 477
rect 1235 443 1268 477
rect 406 393 414 409
rect 260 375 414 393
rect 448 391 456 409
rect 815 409 857 425
rect 448 375 756 391
rect 17 357 756 375
rect 849 393 857 409
rect 1099 409 1149 425
rect 1099 393 1107 409
rect 849 375 1107 393
rect 1141 375 1149 409
rect 815 359 1149 375
rect 1193 409 1268 443
rect 1193 375 1201 409
rect 1235 375 1268 409
rect 1193 359 1268 375
rect 17 179 63 357
rect 722 325 756 357
rect 1099 341 1149 359
rect 168 289 670 323
rect 722 291 1041 325
rect 168 257 202 289
rect 97 249 202 257
rect 636 257 670 289
rect 97 215 123 249
rect 157 215 202 249
rect 271 249 581 255
rect 271 215 287 249
rect 321 215 365 249
rect 399 215 443 249
rect 477 215 515 249
rect 549 215 581 249
rect 636 249 861 257
rect 636 215 804 249
rect 838 215 861 249
rect 1007 249 1041 291
rect 1099 307 1107 341
rect 1141 325 1149 341
rect 1141 307 1268 325
rect 1099 283 1268 307
rect 1007 215 1099 249
rect 1133 215 1149 249
rect 17 163 182 179
rect 17 129 132 163
rect 166 129 182 163
rect 226 163 464 181
rect 260 145 414 163
rect 260 129 276 145
rect 226 95 276 129
rect 388 129 414 145
rect 448 129 464 163
rect 21 61 38 95
rect 72 61 226 95
rect 260 61 276 95
rect 21 51 276 61
rect 320 95 354 111
rect 320 17 354 61
rect 388 95 464 129
rect 388 61 414 95
rect 448 61 464 95
rect 388 51 464 61
rect 526 163 560 181
rect 526 95 560 129
rect 526 17 560 61
rect 594 163 1151 181
rect 594 129 620 163
rect 654 145 815 163
rect 654 129 670 145
rect 594 95 670 129
rect 782 129 815 145
rect 849 145 1097 163
rect 849 129 865 145
rect 1081 129 1097 145
rect 1131 129 1151 163
rect 1190 163 1268 283
rect 1190 129 1201 163
rect 1235 129 1268 163
rect 594 61 620 95
rect 654 61 670 95
rect 594 51 670 61
rect 714 95 748 111
rect 714 17 748 61
rect 782 95 865 129
rect 782 61 815 95
rect 849 61 865 95
rect 782 51 865 61
rect 909 95 943 111
rect 1190 95 1268 129
rect 997 61 1013 95
rect 1047 61 1201 95
rect 1235 61 1268 95
rect 909 17 943 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 533 443 560 459
rect 560 443 567 459
rect 533 425 567 443
rect 737 443 748 459
rect 748 443 771 459
rect 737 425 771 443
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 521 459 579 465
rect 521 425 533 459
rect 567 456 579 459
rect 725 459 783 465
rect 725 456 737 459
rect 567 428 737 456
rect 567 425 579 428
rect 521 419 579 425
rect 725 425 737 428
rect 771 425 783 459
rect 725 419 783 425
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew
flabel corelocali s 1222 289 1256 323 0 FreeSans 400 0 0 0 Y
port 7 nsew
flabel corelocali s 397 221 431 255 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 212 289 246 323 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew
rlabel comment s 0 0 0 0 4 xnor2_2
<< properties >>
string FIXED_BBOX 0 0 1288 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 695744
string GDS_START 686584
<< end >>
