magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 590 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 83 47 113 177
rect 187 47 217 177
rect 271 47 301 177
rect 375 47 405 177
<< pmoshvt >>
rect 85 297 121 497
rect 179 297 215 497
rect 273 297 309 497
rect 367 297 403 497
<< ndiff >>
rect 27 163 83 177
rect 27 129 39 163
rect 73 129 83 163
rect 27 95 83 129
rect 27 61 39 95
rect 73 61 83 95
rect 27 47 83 61
rect 113 163 187 177
rect 113 129 133 163
rect 167 129 187 163
rect 113 95 187 129
rect 113 61 133 95
rect 167 61 187 95
rect 113 47 187 61
rect 217 95 271 177
rect 217 61 227 95
rect 261 61 271 95
rect 217 47 271 61
rect 301 163 375 177
rect 301 129 321 163
rect 355 129 375 163
rect 301 95 375 129
rect 301 61 321 95
rect 355 61 375 95
rect 301 47 375 61
rect 405 95 480 177
rect 405 61 438 95
rect 472 61 480 95
rect 405 47 480 61
<< pdiff >>
rect 27 477 85 497
rect 27 443 39 477
rect 73 443 85 477
rect 27 409 85 443
rect 27 375 39 409
rect 73 375 85 409
rect 27 341 85 375
rect 27 307 39 341
rect 73 307 85 341
rect 27 297 85 307
rect 121 485 179 497
rect 121 451 133 485
rect 167 451 179 485
rect 121 417 179 451
rect 121 383 133 417
rect 167 383 179 417
rect 121 297 179 383
rect 215 477 273 497
rect 215 443 227 477
rect 261 443 273 477
rect 215 409 273 443
rect 215 375 227 409
rect 261 375 273 409
rect 215 341 273 375
rect 215 307 227 341
rect 261 307 273 341
rect 215 297 273 307
rect 309 409 367 497
rect 309 375 321 409
rect 355 375 367 409
rect 309 341 367 375
rect 309 307 321 341
rect 355 307 367 341
rect 309 297 367 307
rect 403 485 457 497
rect 403 451 415 485
rect 449 451 457 485
rect 403 417 457 451
rect 403 383 415 417
rect 449 383 457 417
rect 403 297 457 383
<< ndiffc >>
rect 39 129 73 163
rect 39 61 73 95
rect 133 129 167 163
rect 133 61 167 95
rect 227 61 261 95
rect 321 129 355 163
rect 321 61 355 95
rect 438 61 472 95
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 133 451 167 485
rect 133 383 167 417
rect 227 443 261 477
rect 227 375 261 409
rect 227 307 261 341
rect 321 375 355 409
rect 321 307 355 341
rect 415 451 449 485
rect 415 383 449 417
<< poly >>
rect 85 497 121 523
rect 179 497 215 523
rect 273 497 309 523
rect 367 497 403 523
rect 85 282 121 297
rect 179 282 215 297
rect 273 282 309 297
rect 367 282 403 297
rect 83 265 123 282
rect 177 265 217 282
rect 83 249 217 265
rect 83 215 112 249
rect 146 215 217 249
rect 83 199 217 215
rect 83 177 113 199
rect 187 177 217 199
rect 271 265 311 282
rect 365 265 405 282
rect 271 249 405 265
rect 271 215 321 249
rect 355 215 405 249
rect 271 199 405 215
rect 271 177 301 199
rect 375 177 405 199
rect 83 21 113 47
rect 187 21 217 47
rect 271 21 301 47
rect 375 21 405 47
<< polycont >>
rect 112 215 146 249
rect 321 215 355 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 18 477 73 493
rect 18 443 39 477
rect 18 409 73 443
rect 18 375 39 409
rect 18 341 73 375
rect 107 485 183 527
rect 107 451 133 485
rect 167 451 183 485
rect 107 417 183 451
rect 107 383 133 417
rect 167 383 183 417
rect 107 367 183 383
rect 227 485 475 493
rect 227 477 415 485
rect 261 459 415 477
rect 227 409 261 443
rect 449 451 475 485
rect 18 307 39 341
rect 227 341 261 375
rect 73 307 227 333
rect 18 291 261 307
rect 295 409 371 425
rect 295 375 321 409
rect 355 375 371 409
rect 295 341 371 375
rect 415 417 475 451
rect 449 383 475 417
rect 415 367 475 383
rect 295 307 321 341
rect 355 333 371 341
rect 355 307 462 333
rect 295 289 462 307
rect 18 249 172 255
rect 18 215 112 249
rect 146 215 172 249
rect 206 249 380 255
rect 206 215 321 249
rect 355 215 380 249
rect 419 181 462 289
rect 18 163 73 181
rect 18 129 39 163
rect 18 95 73 129
rect 18 61 39 95
rect 18 17 73 61
rect 107 163 462 181
rect 107 129 133 163
rect 167 145 321 163
rect 167 129 183 145
rect 107 95 183 129
rect 295 129 321 145
rect 355 147 462 163
rect 355 129 371 147
rect 107 61 133 95
rect 167 61 183 95
rect 107 51 183 61
rect 227 95 261 111
rect 227 17 261 61
rect 295 95 371 129
rect 295 61 321 95
rect 355 61 371 95
rect 295 51 371 61
rect 428 95 496 111
rect 428 61 438 95
rect 472 61 496 95
rect 428 17 496 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
flabel corelocali s 214 221 248 255 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel corelocali s 307 357 341 391 0 FreeSans 400 0 0 0 Y
port 7 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew
rlabel comment s 0 0 0 0 4 nor2_2
<< properties >>
string FIXED_BBOX 0 0 552 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2390238
string GDS_START 2385208
<< end >>
