magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 828 561
rect 18 425 69 527
rect 18 215 85 391
rect 383 367 439 527
rect 473 391 523 493
rect 557 427 607 527
rect 641 391 691 493
rect 473 357 691 391
rect 725 359 775 527
rect 566 323 691 357
rect 566 289 811 323
rect 326 215 464 255
rect 734 181 811 289
rect 118 17 249 113
rect 396 17 431 181
rect 465 147 811 181
rect 465 58 531 147
rect 565 17 599 110
rect 633 58 699 147
rect 733 17 767 110
rect 0 -17 828 17
<< obsli1 >>
rect 119 265 153 493
rect 198 323 292 493
rect 198 299 532 323
rect 258 289 532 299
rect 119 199 224 265
rect 119 181 169 199
rect 22 147 169 181
rect 258 181 292 289
rect 498 249 532 289
rect 498 215 700 249
rect 258 147 349 181
rect 22 53 84 147
rect 283 61 349 147
<< metal1 >>
rect 0 496 828 592
rect 0 -48 828 48
<< labels >>
rlabel locali s 326 215 464 255 6 A
port 1 nsew signal input
rlabel locali s 18 215 85 391 6 B_N
port 2 nsew signal input
rlabel locali s 734 181 811 289 6 X
port 3 nsew signal output
rlabel locali s 641 391 691 493 6 X
port 3 nsew signal output
rlabel locali s 633 58 699 147 6 X
port 3 nsew signal output
rlabel locali s 566 323 691 357 6 X
port 3 nsew signal output
rlabel locali s 566 289 811 323 6 X
port 3 nsew signal output
rlabel locali s 473 391 523 493 6 X
port 3 nsew signal output
rlabel locali s 473 357 691 391 6 X
port 3 nsew signal output
rlabel locali s 465 147 811 181 6 X
port 3 nsew signal output
rlabel locali s 465 58 531 147 6 X
port 3 nsew signal output
rlabel locali s 733 17 767 110 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 565 17 599 110 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 396 17 431 181 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 118 17 249 113 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 828 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 828 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 725 359 775 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 557 427 607 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 383 367 439 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 18 425 69 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 828 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 828 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1026482
string GDS_START 1019706
<< end >>
