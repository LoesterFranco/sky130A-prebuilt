magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 368 561
rect 112 375 178 527
rect 212 312 263 493
rect 17 197 88 271
rect 229 166 263 312
rect 298 297 350 527
rect 112 17 178 93
rect 212 51 263 166
rect 298 17 350 185
rect 0 -17 368 17
<< obsli1 >>
rect 35 341 69 493
rect 35 307 178 341
rect 144 265 178 307
rect 144 199 195 265
rect 144 161 178 199
rect 35 127 178 161
rect 35 51 69 127
<< metal1 >>
rect 0 496 368 592
rect 0 -48 368 48
<< labels >>
rlabel locali s 17 197 88 271 6 A
port 1 nsew signal input
rlabel locali s 229 166 263 312 6 X
port 2 nsew signal output
rlabel locali s 212 312 263 493 6 X
port 2 nsew signal output
rlabel locali s 212 51 263 166 6 X
port 2 nsew signal output
rlabel locali s 298 17 350 185 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 112 17 178 93 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 0 -17 368 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 368 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 298 297 350 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 112 375 178 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 0 527 368 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 496 368 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 368 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3035940
string GDS_START 3031504
<< end >>
