magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1932 561
rect 104 427 170 527
rect 19 195 89 325
rect 103 17 169 93
rect 376 449 442 527
rect 352 167 386 337
rect 492 271 558 337
rect 746 433 785 527
rect 352 157 398 167
rect 613 157 650 219
rect 706 211 798 331
rect 352 127 650 157
rect 374 123 650 127
rect 1180 367 1214 527
rect 392 17 461 89
rect 495 61 530 123
rect 752 17 792 109
rect 1558 427 1619 527
rect 1775 325 1809 527
rect 1138 17 1212 117
rect 1846 301 1915 479
rect 1543 17 1617 123
rect 1881 164 1915 301
rect 1775 17 1809 139
rect 1846 61 1915 164
rect 0 -17 1932 17
<< obsli1 >>
rect 36 393 70 493
rect 36 391 169 393
rect 36 359 128 391
rect 123 357 128 359
rect 162 357 169 391
rect 123 194 169 357
rect 123 161 162 194
rect 35 127 162 161
rect 204 187 246 493
rect 204 153 208 187
rect 242 153 246 187
rect 204 143 246 153
rect 35 69 69 127
rect 203 69 246 143
rect 284 415 342 489
rect 538 449 712 483
rect 284 372 644 415
rect 284 93 318 372
rect 423 226 458 372
rect 610 327 644 372
rect 678 399 712 449
rect 836 413 884 488
rect 932 438 1146 472
rect 836 399 870 413
rect 678 365 870 399
rect 990 391 1078 402
rect 610 261 654 327
rect 423 192 492 226
rect 836 177 870 365
rect 684 143 870 177
rect 904 207 952 381
rect 990 357 1041 391
rect 1075 357 1078 391
rect 990 331 1078 357
rect 1112 315 1146 438
rect 1248 427 1298 493
rect 1343 433 1520 467
rect 1112 297 1214 315
rect 1054 263 1214 297
rect 904 187 1020 207
rect 904 156 949 187
rect 284 52 358 93
rect 684 89 718 143
rect 836 123 870 143
rect 926 153 949 156
rect 983 153 1020 187
rect 926 141 1020 153
rect 564 55 718 89
rect 836 57 892 123
rect 1054 107 1088 263
rect 1180 249 1214 263
rect 1122 213 1156 219
rect 1248 213 1282 427
rect 1316 391 1354 393
rect 1316 357 1318 391
rect 1352 357 1354 391
rect 1316 249 1354 357
rect 1388 315 1452 381
rect 1122 153 1282 213
rect 1388 207 1426 315
rect 1486 281 1520 433
rect 1687 381 1741 491
rect 1554 315 1741 381
rect 940 73 1088 107
rect 1248 107 1282 153
rect 1316 187 1426 207
rect 1316 153 1326 187
rect 1360 153 1426 187
rect 1316 141 1426 153
rect 1460 265 1520 281
rect 1707 265 1741 315
rect 1460 199 1673 265
rect 1707 199 1847 265
rect 1460 107 1494 199
rect 1707 165 1741 199
rect 1248 73 1340 107
rect 1386 73 1494 107
rect 1671 60 1741 165
<< obsli1c >>
rect 128 357 162 391
rect 208 153 242 187
rect 1041 357 1075 391
rect 949 153 983 187
rect 1318 357 1352 391
rect 1326 153 1360 187
<< metal1 >>
rect 0 496 1932 592
rect 0 -48 1932 48
<< obsm1 >>
rect 116 391 174 397
rect 116 357 128 391
rect 162 388 174 391
rect 1029 391 1087 397
rect 1029 388 1041 391
rect 162 360 1041 388
rect 162 357 174 360
rect 116 351 174 357
rect 1029 357 1041 360
rect 1075 388 1087 391
rect 1306 391 1364 397
rect 1306 388 1318 391
rect 1075 360 1318 388
rect 1075 357 1087 360
rect 1029 351 1087 357
rect 1306 357 1318 360
rect 1352 357 1364 391
rect 1306 351 1364 357
rect 196 187 254 193
rect 196 153 208 187
rect 242 184 254 187
rect 937 187 995 193
rect 937 184 949 187
rect 242 156 949 184
rect 242 153 254 156
rect 196 147 254 153
rect 937 153 949 156
rect 983 184 995 187
rect 1314 187 1372 193
rect 1314 184 1326 187
rect 983 156 1326 184
rect 983 153 995 156
rect 937 147 995 153
rect 1314 153 1326 156
rect 1360 153 1372 187
rect 1314 147 1372 153
<< labels >>
rlabel locali s 492 271 558 337 6 D
port 1 nsew signal input
rlabel locali s 1881 164 1915 301 6 Q
port 2 nsew signal output
rlabel locali s 1846 301 1915 479 6 Q
port 2 nsew signal output
rlabel locali s 1846 61 1915 164 6 Q
port 2 nsew signal output
rlabel locali s 706 211 798 331 6 SCD
port 3 nsew signal input
rlabel locali s 613 157 650 219 6 SCE
port 4 nsew signal input
rlabel locali s 495 61 530 123 6 SCE
port 4 nsew signal input
rlabel locali s 374 123 650 127 6 SCE
port 4 nsew signal input
rlabel locali s 352 167 386 337 6 SCE
port 4 nsew signal input
rlabel locali s 352 157 398 167 6 SCE
port 4 nsew signal input
rlabel locali s 352 127 650 157 6 SCE
port 4 nsew signal input
rlabel locali s 19 195 89 325 6 CLK
port 5 nsew clock input
rlabel locali s 1775 17 1809 139 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1543 17 1617 123 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1138 17 1212 117 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 752 17 792 109 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 392 17 461 89 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 103 17 169 93 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 1932 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1932 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1775 325 1809 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1558 427 1619 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1180 367 1214 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 746 433 785 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 376 449 442 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 104 427 170 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 1932 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 1932 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1932 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 376304
string GDS_START 361098
<< end >>
