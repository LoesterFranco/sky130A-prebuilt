magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 828 561
rect 19 416 85 527
rect 24 153 85 361
rect 197 17 245 177
rect 304 157 343 423
rect 477 439 511 527
rect 632 455 698 527
rect 420 299 735 335
rect 420 249 485 299
rect 419 215 485 249
rect 521 199 643 265
rect 677 259 735 299
rect 677 207 759 259
rect 304 123 612 157
rect 304 51 344 123
rect 388 17 454 89
rect 546 51 612 123
rect 727 17 786 173
rect 0 -17 828 17
<< obsli1 >>
rect 209 457 443 493
rect 119 257 171 453
rect 209 359 270 457
rect 119 214 265 257
rect 119 106 159 214
rect 53 72 159 106
rect 377 405 443 457
rect 562 421 596 493
rect 732 421 784 493
rect 562 405 784 421
rect 377 371 784 405
<< metal1 >>
rect 0 496 828 592
rect 0 -48 828 48
<< labels >>
rlabel locali s 521 199 643 265 6 A1
port 1 nsew signal input
rlabel locali s 677 259 735 299 6 A2
port 2 nsew signal input
rlabel locali s 677 207 759 259 6 A2
port 2 nsew signal input
rlabel locali s 420 299 735 335 6 A2
port 2 nsew signal input
rlabel locali s 420 249 485 299 6 A2
port 2 nsew signal input
rlabel locali s 419 215 485 249 6 A2
port 2 nsew signal input
rlabel locali s 24 153 85 361 6 B1_N
port 3 nsew signal input
rlabel locali s 546 51 612 123 6 Y
port 4 nsew signal output
rlabel locali s 304 157 343 423 6 Y
port 4 nsew signal output
rlabel locali s 304 123 612 157 6 Y
port 4 nsew signal output
rlabel locali s 304 51 344 123 6 Y
port 4 nsew signal output
rlabel locali s 727 17 786 173 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 388 17 454 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 197 17 245 177 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 828 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 828 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 632 455 698 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 477 439 511 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 19 416 85 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 828 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 828 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 4016036
string GDS_START 4009404
<< end >>
