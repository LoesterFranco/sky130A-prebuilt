magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 1478 704
<< pwell >>
rect 0 0 1440 49
<< scnmos >>
rect 84 74 114 202
rect 198 74 228 202
rect 284 74 314 202
rect 384 74 414 202
rect 476 74 506 202
rect 569 74 599 202
rect 805 94 835 222
rect 883 94 913 222
rect 1011 74 1041 222
rect 1126 74 1156 222
rect 1226 74 1256 222
rect 1312 74 1342 222
<< pmoshvt >>
rect 100 392 130 592
rect 190 392 220 592
rect 280 392 310 592
rect 370 392 400 592
rect 572 368 602 536
rect 676 368 706 536
rect 800 368 830 536
rect 890 368 920 536
rect 1014 368 1044 592
rect 1124 368 1154 592
rect 1224 368 1254 592
rect 1315 368 1345 592
<< ndiff >>
rect 27 190 84 202
rect 27 156 39 190
rect 73 156 84 190
rect 27 120 84 156
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 127 198 202
rect 114 93 139 127
rect 173 93 198 127
rect 114 74 198 93
rect 228 190 284 202
rect 228 156 239 190
rect 273 156 284 190
rect 228 120 284 156
rect 228 86 239 120
rect 273 86 284 120
rect 228 74 284 86
rect 314 121 384 202
rect 314 87 339 121
rect 373 87 384 121
rect 314 74 384 87
rect 414 190 476 202
rect 414 156 428 190
rect 462 156 476 190
rect 414 74 476 156
rect 506 121 569 202
rect 506 87 517 121
rect 551 87 569 121
rect 506 74 569 87
rect 599 179 663 202
rect 599 145 617 179
rect 651 145 663 179
rect 599 74 663 145
rect 744 177 805 222
rect 744 143 760 177
rect 794 143 805 177
rect 744 94 805 143
rect 835 94 883 222
rect 913 145 1011 222
rect 913 111 945 145
rect 979 111 1011 145
rect 913 94 1011 111
rect 961 74 1011 94
rect 1041 194 1126 222
rect 1041 160 1067 194
rect 1101 160 1126 194
rect 1041 120 1126 160
rect 1041 86 1067 120
rect 1101 86 1126 120
rect 1041 74 1126 86
rect 1156 124 1226 222
rect 1156 90 1167 124
rect 1201 90 1226 124
rect 1156 74 1226 90
rect 1256 210 1312 222
rect 1256 176 1267 210
rect 1301 176 1312 210
rect 1256 120 1312 176
rect 1256 86 1267 120
rect 1301 86 1312 120
rect 1256 74 1312 86
rect 1342 210 1413 222
rect 1342 176 1367 210
rect 1401 176 1413 210
rect 1342 120 1413 176
rect 1342 86 1367 120
rect 1401 86 1413 120
rect 1342 74 1413 86
<< pdiff >>
rect 724 608 782 620
rect 41 580 100 592
rect 41 546 53 580
rect 87 546 100 580
rect 41 509 100 546
rect 41 475 53 509
rect 87 475 100 509
rect 41 438 100 475
rect 41 404 53 438
rect 87 404 100 438
rect 41 392 100 404
rect 130 580 190 592
rect 130 546 143 580
rect 177 546 190 580
rect 130 508 190 546
rect 130 474 143 508
rect 177 474 190 508
rect 130 392 190 474
rect 220 580 280 592
rect 220 546 233 580
rect 267 546 280 580
rect 220 510 280 546
rect 220 476 233 510
rect 267 476 280 510
rect 220 440 280 476
rect 220 406 233 440
rect 267 406 280 440
rect 220 392 280 406
rect 310 531 370 592
rect 310 497 323 531
rect 357 497 370 531
rect 310 440 370 497
rect 310 406 323 440
rect 357 406 370 440
rect 310 392 370 406
rect 400 580 459 592
rect 400 546 413 580
rect 447 546 459 580
rect 724 574 736 608
rect 770 574 782 608
rect 400 508 459 546
rect 724 536 782 574
rect 938 608 996 620
rect 938 574 950 608
rect 984 592 996 608
rect 984 574 1014 592
rect 938 536 1014 574
rect 400 474 413 508
rect 447 474 459 508
rect 400 392 459 474
rect 513 519 572 536
rect 513 485 525 519
rect 559 485 572 519
rect 513 368 572 485
rect 602 414 676 536
rect 602 380 616 414
rect 650 380 676 414
rect 602 368 676 380
rect 706 368 800 536
rect 830 440 890 536
rect 830 406 843 440
rect 877 406 890 440
rect 830 368 890 406
rect 920 368 1014 536
rect 1044 580 1124 592
rect 1044 546 1067 580
rect 1101 546 1124 580
rect 1044 497 1124 546
rect 1044 463 1067 497
rect 1101 463 1124 497
rect 1044 414 1124 463
rect 1044 380 1067 414
rect 1101 380 1124 414
rect 1044 368 1124 380
rect 1154 582 1224 592
rect 1154 548 1167 582
rect 1201 548 1224 582
rect 1154 514 1224 548
rect 1154 480 1167 514
rect 1201 480 1224 514
rect 1154 446 1224 480
rect 1154 412 1167 446
rect 1201 412 1224 446
rect 1154 368 1224 412
rect 1254 580 1315 592
rect 1254 546 1267 580
rect 1301 546 1315 580
rect 1254 497 1315 546
rect 1254 463 1267 497
rect 1301 463 1315 497
rect 1254 414 1315 463
rect 1254 380 1267 414
rect 1301 380 1315 414
rect 1254 368 1315 380
rect 1345 580 1413 592
rect 1345 546 1367 580
rect 1401 546 1413 580
rect 1345 497 1413 546
rect 1345 463 1367 497
rect 1401 463 1413 497
rect 1345 414 1413 463
rect 1345 380 1367 414
rect 1401 380 1413 414
rect 1345 368 1413 380
<< ndiffc >>
rect 39 156 73 190
rect 39 86 73 120
rect 139 93 173 127
rect 239 156 273 190
rect 239 86 273 120
rect 339 87 373 121
rect 428 156 462 190
rect 517 87 551 121
rect 617 145 651 179
rect 760 143 794 177
rect 945 111 979 145
rect 1067 160 1101 194
rect 1067 86 1101 120
rect 1167 90 1201 124
rect 1267 176 1301 210
rect 1267 86 1301 120
rect 1367 176 1401 210
rect 1367 86 1401 120
<< pdiffc >>
rect 53 546 87 580
rect 53 475 87 509
rect 53 404 87 438
rect 143 546 177 580
rect 143 474 177 508
rect 233 546 267 580
rect 233 476 267 510
rect 233 406 267 440
rect 323 497 357 531
rect 323 406 357 440
rect 413 546 447 580
rect 736 574 770 608
rect 950 574 984 608
rect 413 474 447 508
rect 525 485 559 519
rect 616 380 650 414
rect 843 406 877 440
rect 1067 546 1101 580
rect 1067 463 1101 497
rect 1067 380 1101 414
rect 1167 548 1201 582
rect 1167 480 1201 514
rect 1167 412 1201 446
rect 1267 546 1301 580
rect 1267 463 1301 497
rect 1267 380 1301 414
rect 1367 546 1401 580
rect 1367 463 1401 497
rect 1367 380 1401 414
<< poly >>
rect 100 592 130 618
rect 190 592 220 618
rect 280 592 310 618
rect 370 592 400 618
rect 572 536 602 562
rect 676 536 706 562
rect 1014 592 1044 618
rect 1124 592 1154 618
rect 1224 592 1254 618
rect 1315 592 1345 618
rect 800 536 830 562
rect 890 536 920 562
rect 100 377 130 392
rect 190 377 220 392
rect 280 377 310 392
rect 370 377 400 392
rect 97 318 133 377
rect 187 318 223 377
rect 21 302 223 318
rect 21 268 37 302
rect 71 268 105 302
rect 139 268 173 302
rect 207 282 223 302
rect 277 356 313 377
rect 367 356 403 377
rect 277 340 428 356
rect 572 353 602 368
rect 676 353 706 368
rect 800 353 830 368
rect 890 353 920 368
rect 1014 353 1044 368
rect 1124 353 1154 368
rect 1224 353 1254 368
rect 1315 353 1345 368
rect 277 306 310 340
rect 344 306 378 340
rect 412 306 428 340
rect 569 326 605 353
rect 673 326 706 353
rect 797 336 833 353
rect 887 336 923 353
rect 277 290 428 306
rect 498 310 703 326
rect 498 290 514 310
rect 207 268 228 282
rect 21 252 228 268
rect 84 202 114 252
rect 198 202 228 252
rect 284 202 314 290
rect 384 202 414 290
rect 476 276 514 290
rect 548 276 585 310
rect 619 276 653 310
rect 687 276 703 310
rect 476 260 703 276
rect 769 320 835 336
rect 769 286 785 320
rect 819 286 835 320
rect 769 270 835 286
rect 476 202 506 260
rect 569 202 599 260
rect 805 222 835 270
rect 883 320 949 336
rect 883 286 899 320
rect 933 286 949 320
rect 883 270 949 286
rect 1011 310 1047 353
rect 1121 310 1157 353
rect 1221 310 1257 353
rect 1011 294 1257 310
rect 883 222 913 270
rect 1011 260 1027 294
rect 1061 260 1095 294
rect 1129 260 1163 294
rect 1197 274 1257 294
rect 1312 274 1348 353
rect 1197 260 1348 274
rect 1011 244 1348 260
rect 1011 222 1041 244
rect 1126 222 1156 244
rect 1226 222 1256 244
rect 1312 222 1342 244
rect 84 48 114 74
rect 198 48 228 74
rect 284 48 314 74
rect 384 48 414 74
rect 476 48 506 74
rect 569 48 599 74
rect 805 68 835 94
rect 883 68 913 94
rect 1011 48 1041 74
rect 1126 48 1156 74
rect 1226 48 1256 74
rect 1312 48 1342 74
<< polycont >>
rect 37 268 71 302
rect 105 268 139 302
rect 173 268 207 302
rect 310 306 344 340
rect 378 306 412 340
rect 514 276 548 310
rect 585 276 619 310
rect 653 276 687 310
rect 785 286 819 320
rect 899 286 933 320
rect 1027 260 1061 294
rect 1095 260 1129 294
rect 1163 260 1197 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 37 580 103 596
rect 37 546 53 580
rect 87 546 103 580
rect 37 509 103 546
rect 37 475 53 509
rect 87 475 103 509
rect 37 438 103 475
rect 143 580 177 649
rect 143 508 177 546
rect 143 458 177 474
rect 217 581 463 615
rect 217 580 283 581
rect 217 546 233 580
rect 267 546 283 580
rect 397 580 463 581
rect 217 510 283 546
rect 217 476 233 510
rect 267 476 283 510
rect 37 404 53 438
rect 87 424 103 438
rect 217 440 283 476
rect 217 424 233 440
rect 87 406 233 424
rect 267 406 283 440
rect 87 404 283 406
rect 37 390 283 404
rect 323 531 357 547
rect 323 440 357 497
rect 397 546 413 580
rect 447 546 463 580
rect 397 508 463 546
rect 397 474 413 508
rect 447 474 463 508
rect 397 458 463 474
rect 509 519 575 649
rect 720 608 786 649
rect 720 574 736 608
rect 770 574 786 608
rect 720 558 786 574
rect 934 608 1000 649
rect 934 574 950 608
rect 984 574 1000 608
rect 934 558 1000 574
rect 1051 580 1117 596
rect 1051 546 1067 580
rect 1101 546 1117 580
rect 509 485 525 519
rect 559 485 575 519
rect 509 464 575 485
rect 633 490 1017 524
rect 633 430 667 490
rect 599 424 667 430
rect 357 414 667 424
rect 357 406 616 414
rect 323 390 616 406
rect 37 388 103 390
rect 599 380 616 390
rect 650 380 667 414
rect 599 364 667 380
rect 701 440 893 456
rect 701 406 843 440
rect 877 406 893 440
rect 701 390 893 406
rect 21 302 223 354
rect 21 268 37 302
rect 71 268 105 302
rect 139 268 173 302
rect 207 268 223 302
rect 294 340 455 356
rect 294 306 310 340
rect 344 306 378 340
rect 412 306 455 340
rect 701 326 735 390
rect 294 290 455 306
rect 498 310 735 326
rect 21 252 223 268
rect 498 276 514 310
rect 548 276 585 310
rect 619 276 653 310
rect 687 276 735 310
rect 498 260 735 276
rect 769 320 839 356
rect 769 286 785 320
rect 819 286 839 320
rect 769 270 839 286
rect 883 320 949 356
rect 883 286 899 320
rect 933 286 949 320
rect 883 270 949 286
rect 983 310 1017 490
rect 1051 497 1117 546
rect 1051 463 1067 497
rect 1101 463 1117 497
rect 1051 414 1117 463
rect 1051 380 1067 414
rect 1101 380 1117 414
rect 1151 582 1217 649
rect 1151 548 1167 582
rect 1201 548 1217 582
rect 1151 514 1217 548
rect 1151 480 1167 514
rect 1201 480 1217 514
rect 1151 446 1217 480
rect 1151 412 1167 446
rect 1201 412 1217 446
rect 1251 580 1317 596
rect 1251 546 1267 580
rect 1301 546 1317 580
rect 1251 497 1317 546
rect 1251 463 1267 497
rect 1301 463 1317 497
rect 1251 414 1317 463
rect 1051 378 1117 380
rect 1251 380 1267 414
rect 1301 380 1317 414
rect 1251 378 1317 380
rect 1051 344 1317 378
rect 1351 580 1417 649
rect 1351 546 1367 580
rect 1401 546 1417 580
rect 1351 497 1417 546
rect 1351 463 1367 497
rect 1401 463 1417 497
rect 1351 414 1417 463
rect 1351 380 1367 414
rect 1401 380 1417 414
rect 1351 364 1417 380
rect 983 294 1213 310
rect 701 226 735 260
rect 983 260 1027 294
rect 1061 260 1095 294
rect 1129 260 1163 294
rect 1197 260 1213 294
rect 983 244 1213 260
rect 23 190 667 218
rect 701 192 806 226
rect 983 224 1017 244
rect 23 156 39 190
rect 73 184 239 190
rect 73 156 89 184
rect 23 120 89 156
rect 223 156 239 184
rect 273 156 428 190
rect 462 179 667 190
rect 462 156 617 179
rect 23 86 39 120
rect 73 86 89 120
rect 23 70 89 86
rect 123 127 189 150
rect 123 93 139 127
rect 173 93 189 127
rect 123 17 189 93
rect 223 120 289 156
rect 601 145 617 156
rect 651 145 667 179
rect 223 86 239 120
rect 273 86 289 120
rect 223 70 289 86
rect 323 121 389 122
rect 323 87 339 121
rect 373 87 389 121
rect 323 17 389 87
rect 501 121 567 122
rect 501 87 517 121
rect 551 87 567 121
rect 601 119 667 145
rect 740 177 806 192
rect 740 143 760 177
rect 794 143 806 177
rect 740 127 806 143
rect 840 190 1017 224
rect 1251 210 1317 344
rect 1051 194 1267 210
rect 501 85 567 87
rect 840 85 874 190
rect 1051 160 1067 194
rect 1101 176 1267 194
rect 1301 176 1317 210
rect 1101 162 1317 176
rect 1101 160 1117 162
rect 501 51 874 85
rect 908 145 1016 156
rect 908 111 945 145
rect 979 111 1016 145
rect 908 17 1016 111
rect 1051 120 1117 160
rect 1051 86 1067 120
rect 1101 86 1117 120
rect 1051 70 1117 86
rect 1151 124 1217 128
rect 1151 90 1167 124
rect 1201 90 1217 124
rect 1151 17 1217 90
rect 1251 120 1317 162
rect 1251 86 1267 120
rect 1301 86 1317 120
rect 1251 70 1317 86
rect 1351 210 1417 226
rect 1351 176 1367 210
rect 1401 176 1417 210
rect 1351 120 1417 176
rect 1351 86 1367 120
rect 1401 86 1417 120
rect 1351 17 1417 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 683 1440 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 0 617 1440 649
rect 0 17 1440 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -49 1440 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o2bb2a_4
flabel pwell s 0 0 1440 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nwell s 0 617 1440 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 1440 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 1440 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 1087 168 1121 202 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 1183 168 1217 202 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 A2_N
port 2 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 A1_N
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 1440 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1569982
string GDS_START 1558588
<< end >>
