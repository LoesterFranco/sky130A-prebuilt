magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1472 561
rect 35 367 69 527
rect 203 367 237 527
rect 371 367 405 527
rect 455 323 489 493
rect 523 367 589 527
rect 623 323 657 493
rect 691 367 757 527
rect 791 323 825 493
rect 859 367 925 527
rect 959 323 993 493
rect 1027 367 1093 527
rect 1127 323 1161 493
rect 1195 367 1261 527
rect 1295 323 1329 493
rect 455 289 1329 323
rect 1363 297 1429 527
rect 27 215 332 255
rect 942 181 1329 289
rect 455 147 1329 181
rect 19 17 85 113
rect 187 17 253 113
rect 355 17 421 113
rect 455 51 489 147
rect 523 17 589 113
rect 623 51 657 147
rect 691 17 757 113
rect 791 51 825 147
rect 859 17 925 113
rect 959 51 993 147
rect 1027 17 1093 113
rect 1127 51 1161 147
rect 1195 17 1261 113
rect 1295 51 1329 147
rect 1363 17 1429 177
rect 0 -17 1472 17
<< obsli1 >>
rect 103 323 169 493
rect 271 323 337 493
rect 103 289 403 323
rect 368 249 403 289
rect 368 215 893 249
rect 368 181 403 215
rect 119 147 403 181
rect 119 51 153 147
rect 287 52 321 147
<< metal1 >>
rect 0 496 1472 592
rect 0 -48 1472 48
<< labels >>
rlabel locali s 27 215 332 255 6 A
port 1 nsew signal input
rlabel locali s 1295 323 1329 493 6 X
port 2 nsew signal output
rlabel locali s 1295 51 1329 147 6 X
port 2 nsew signal output
rlabel locali s 1127 323 1161 493 6 X
port 2 nsew signal output
rlabel locali s 1127 51 1161 147 6 X
port 2 nsew signal output
rlabel locali s 959 323 993 493 6 X
port 2 nsew signal output
rlabel locali s 959 51 993 147 6 X
port 2 nsew signal output
rlabel locali s 942 181 1329 289 6 X
port 2 nsew signal output
rlabel locali s 791 323 825 493 6 X
port 2 nsew signal output
rlabel locali s 791 51 825 147 6 X
port 2 nsew signal output
rlabel locali s 623 323 657 493 6 X
port 2 nsew signal output
rlabel locali s 623 51 657 147 6 X
port 2 nsew signal output
rlabel locali s 455 323 489 493 6 X
port 2 nsew signal output
rlabel locali s 455 289 1329 323 6 X
port 2 nsew signal output
rlabel locali s 455 147 1329 181 6 X
port 2 nsew signal output
rlabel locali s 455 51 489 147 6 X
port 2 nsew signal output
rlabel locali s 1363 17 1429 177 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1195 17 1261 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1027 17 1093 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 859 17 925 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 691 17 757 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 523 17 589 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 355 17 421 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 187 17 253 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 19 17 85 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 0 -17 1472 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1472 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1363 297 1429 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1195 367 1261 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1027 367 1093 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 859 367 925 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 691 367 757 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 523 367 589 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 371 367 405 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 203 367 237 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 35 367 69 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 0 527 1472 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 496 1472 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1472 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3015918
string GDS_START 3004784
<< end >>
