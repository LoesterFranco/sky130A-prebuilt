magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 518 704
<< pwell >>
rect 0 0 480 49
<< scnmos >>
rect 125 112 155 222
rect 250 112 280 222
rect 366 74 396 222
<< pmoshvt >>
rect 122 368 152 536
rect 206 368 236 536
rect 364 368 394 592
<< ndiff >>
rect 27 183 125 222
rect 27 149 80 183
rect 114 149 125 183
rect 27 112 125 149
rect 155 181 250 222
rect 155 147 198 181
rect 232 147 250 181
rect 155 112 250 147
rect 280 152 366 222
rect 280 118 307 152
rect 341 118 366 152
rect 280 112 366 118
rect 295 74 366 112
rect 396 210 453 222
rect 396 176 407 210
rect 441 176 453 210
rect 396 120 453 176
rect 396 86 407 120
rect 441 86 453 120
rect 396 74 453 86
<< pdiff >>
rect 270 580 364 592
rect 270 546 317 580
rect 351 546 364 580
rect 270 536 364 546
rect 63 524 122 536
rect 63 490 75 524
rect 109 490 122 524
rect 63 414 122 490
rect 63 380 75 414
rect 109 380 122 414
rect 63 368 122 380
rect 152 368 206 536
rect 236 508 364 536
rect 236 492 317 508
rect 236 458 249 492
rect 283 474 317 492
rect 351 474 364 508
rect 283 458 364 474
rect 236 368 364 458
rect 394 580 453 592
rect 394 546 407 580
rect 441 546 453 580
rect 394 497 453 546
rect 394 463 407 497
rect 441 463 453 497
rect 394 414 453 463
rect 394 380 407 414
rect 441 380 453 414
rect 394 368 453 380
<< ndiffc >>
rect 80 149 114 183
rect 198 147 232 181
rect 307 118 341 152
rect 407 176 441 210
rect 407 86 441 120
<< pdiffc >>
rect 317 546 351 580
rect 75 490 109 524
rect 75 380 109 414
rect 249 458 283 492
rect 317 474 351 508
rect 407 546 441 580
rect 407 463 441 497
rect 407 380 441 414
<< poly >>
rect 364 592 394 618
rect 122 536 152 562
rect 206 536 236 562
rect 122 353 152 368
rect 206 353 236 368
rect 364 353 394 368
rect 119 310 155 353
rect 21 294 155 310
rect 203 336 239 353
rect 203 320 280 336
rect 361 326 397 353
rect 203 306 225 320
rect 21 260 37 294
rect 71 260 105 294
rect 139 260 155 294
rect 209 286 225 306
rect 259 286 280 320
rect 209 270 280 286
rect 21 244 155 260
rect 125 222 155 244
rect 250 222 280 270
rect 328 310 397 326
rect 328 276 344 310
rect 378 276 397 310
rect 328 260 397 276
rect 366 222 396 260
rect 125 86 155 112
rect 250 86 280 112
rect 366 48 396 74
<< polycont >>
rect 37 260 71 294
rect 105 260 139 294
rect 225 286 259 320
rect 344 276 378 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 233 580 357 649
rect 233 546 317 580
rect 351 546 357 580
rect 59 524 125 540
rect 59 490 75 524
rect 109 490 125 524
rect 59 424 125 490
rect 233 508 357 546
rect 233 492 317 508
rect 233 458 249 492
rect 283 474 317 492
rect 351 474 357 508
rect 283 458 357 474
rect 391 580 462 596
rect 391 546 407 580
rect 441 546 462 580
rect 391 497 462 546
rect 391 463 407 497
rect 441 463 462 497
rect 59 414 357 424
rect 59 380 75 414
rect 109 390 357 414
rect 109 380 125 390
rect 59 364 125 380
rect 209 320 275 356
rect 21 294 155 310
rect 21 260 37 294
rect 71 260 105 294
rect 139 260 155 294
rect 209 286 225 320
rect 259 286 275 320
rect 209 270 275 286
rect 323 326 357 390
rect 391 414 462 463
rect 391 380 407 414
rect 441 380 462 414
rect 391 364 462 380
rect 323 310 394 326
rect 323 276 344 310
rect 378 276 394 310
rect 21 236 155 260
rect 323 260 394 276
rect 323 236 357 260
rect 189 202 357 236
rect 428 226 462 364
rect 391 210 462 226
rect 59 183 130 199
rect 59 149 80 183
rect 114 149 130 183
rect 59 17 130 149
rect 189 181 248 202
rect 189 147 198 181
rect 232 147 248 181
rect 391 176 407 210
rect 441 176 462 210
rect 189 108 248 147
rect 291 152 357 168
rect 291 118 307 152
rect 341 118 357 152
rect 291 17 357 118
rect 391 120 462 176
rect 391 86 407 120
rect 441 86 462 120
rect 391 70 462 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< metal1 >>
rect 0 683 480 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 0 617 480 649
rect 0 17 480 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
rect 0 -49 480 -17
<< labels >>
rlabel comment s 0 0 0 0 4 or2_1
flabel pwell s 0 0 480 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 0 617 480 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 0 617 480 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 480 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 415 390 449 424 0 FreeSans 340 0 0 0 X
port 7 nsew
flabel corelocali s 415 464 449 498 0 FreeSans 340 0 0 0 X
port 7 nsew
flabel corelocali s 415 538 449 572 0 FreeSans 340 0 0 0 X
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 480 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1026914
string GDS_START 1022144
<< end >>
