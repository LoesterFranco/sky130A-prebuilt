magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 710 704
<< pwell >>
rect 0 0 672 49
<< scnmos >>
rect 185 112 215 222
rect 321 74 351 222
rect 407 74 437 222
rect 501 74 531 222
<< pmoshvt >>
rect 84 424 114 592
rect 318 368 348 592
rect 408 368 438 592
rect 504 368 534 592
<< ndiff >>
rect 132 176 185 222
rect 132 142 140 176
rect 174 142 185 176
rect 132 112 185 142
rect 215 204 321 222
rect 215 170 240 204
rect 274 170 321 204
rect 215 136 321 170
rect 215 112 276 136
rect 268 102 276 112
rect 310 102 321 136
rect 268 74 321 102
rect 351 210 407 222
rect 351 176 362 210
rect 396 176 407 210
rect 351 120 407 176
rect 351 86 362 120
rect 396 86 407 120
rect 351 74 407 86
rect 437 74 501 222
rect 531 197 588 222
rect 531 163 542 197
rect 576 163 588 197
rect 531 120 588 163
rect 531 86 542 120
rect 576 86 588 120
rect 531 74 588 86
<< pdiff >>
rect 29 580 84 592
rect 29 546 37 580
rect 71 546 84 580
rect 29 470 84 546
rect 29 436 37 470
rect 71 436 84 470
rect 29 424 84 436
rect 114 580 169 592
rect 114 546 127 580
rect 161 546 169 580
rect 114 473 169 546
rect 114 439 127 473
rect 161 439 169 473
rect 114 424 169 439
rect 263 580 318 592
rect 263 546 271 580
rect 305 546 318 580
rect 263 497 318 546
rect 263 463 271 497
rect 305 463 318 497
rect 263 414 318 463
rect 263 380 271 414
rect 305 380 318 414
rect 263 368 318 380
rect 348 580 408 592
rect 348 546 361 580
rect 395 546 408 580
rect 348 462 408 546
rect 348 428 361 462
rect 395 428 408 462
rect 348 368 408 428
rect 438 582 504 592
rect 438 548 454 582
rect 488 548 504 582
rect 438 514 504 548
rect 438 480 454 514
rect 488 480 504 514
rect 438 368 504 480
rect 534 580 589 592
rect 534 546 547 580
rect 581 546 589 580
rect 534 497 589 546
rect 534 463 547 497
rect 581 463 589 497
rect 534 414 589 463
rect 534 380 547 414
rect 581 380 589 414
rect 534 368 589 380
<< ndiffc >>
rect 140 142 174 176
rect 240 170 274 204
rect 276 102 310 136
rect 362 176 396 210
rect 362 86 396 120
rect 542 163 576 197
rect 542 86 576 120
<< pdiffc >>
rect 37 546 71 580
rect 37 436 71 470
rect 127 546 161 580
rect 127 439 161 473
rect 271 546 305 580
rect 271 463 305 497
rect 271 380 305 414
rect 361 546 395 580
rect 361 428 395 462
rect 454 548 488 582
rect 454 480 488 514
rect 547 546 581 580
rect 547 463 581 497
rect 547 380 581 414
<< poly >>
rect 84 592 114 618
rect 318 592 348 618
rect 408 592 438 618
rect 504 592 534 618
rect 84 409 114 424
rect 81 321 117 409
rect 318 353 348 368
rect 408 353 438 368
rect 504 353 534 368
rect 24 305 111 321
rect 315 310 351 353
rect 405 336 441 353
rect 24 271 40 305
rect 74 271 111 305
rect 24 267 111 271
rect 257 294 351 310
rect 24 237 215 267
rect 257 260 273 294
rect 307 260 351 294
rect 393 320 459 336
rect 393 286 409 320
rect 443 286 459 320
rect 393 270 459 286
rect 501 310 537 353
rect 501 294 567 310
rect 257 244 351 260
rect 24 203 40 237
rect 74 203 111 237
rect 185 222 215 237
rect 321 222 351 244
rect 407 222 437 270
rect 501 260 517 294
rect 551 260 567 294
rect 501 244 567 260
rect 501 222 531 244
rect 24 169 111 203
rect 24 135 40 169
rect 74 135 111 169
rect 24 101 111 135
rect 24 67 40 101
rect 74 67 111 101
rect 185 86 215 112
rect 24 51 111 67
rect 321 48 351 74
rect 407 48 437 74
rect 501 48 531 74
<< polycont >>
rect 40 271 74 305
rect 273 260 307 294
rect 409 286 443 320
rect 40 203 74 237
rect 517 260 551 294
rect 40 135 74 169
rect 40 67 74 101
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 21 580 87 596
rect 21 546 37 580
rect 71 546 87 580
rect 21 470 87 546
rect 21 436 37 470
rect 71 436 87 470
rect 21 389 87 436
rect 127 580 177 649
rect 161 546 177 580
rect 127 473 177 546
rect 161 439 177 473
rect 127 423 177 439
rect 217 580 305 596
rect 217 546 271 580
rect 217 497 305 546
rect 217 463 271 497
rect 217 414 305 463
rect 21 355 183 389
rect 217 384 271 414
rect 24 305 90 321
rect 24 271 40 305
rect 74 271 90 305
rect 24 237 90 271
rect 24 203 40 237
rect 74 203 90 237
rect 149 310 183 355
rect 255 380 271 384
rect 345 580 404 596
rect 345 546 361 580
rect 395 546 404 580
rect 345 462 404 546
rect 438 582 504 649
rect 438 548 454 582
rect 488 548 504 582
rect 438 514 504 548
rect 438 480 454 514
rect 488 480 504 514
rect 538 580 597 596
rect 538 546 547 580
rect 581 546 597 580
rect 538 497 597 546
rect 345 428 361 462
rect 395 446 404 462
rect 538 463 547 497
rect 581 463 597 497
rect 538 446 597 463
rect 395 428 597 446
rect 345 414 597 428
rect 345 412 547 414
rect 255 378 305 380
rect 531 380 547 412
rect 581 380 597 414
rect 255 344 375 378
rect 531 364 597 380
rect 149 294 307 310
rect 149 260 273 294
rect 149 244 307 260
rect 149 210 190 244
rect 341 236 375 344
rect 409 320 459 356
rect 443 286 459 320
rect 409 270 459 286
rect 501 294 647 310
rect 501 260 517 294
rect 551 260 647 294
rect 501 236 647 260
rect 341 210 412 236
rect 24 169 90 203
rect 24 135 40 169
rect 74 135 90 169
rect 24 101 90 135
rect 124 176 190 210
rect 124 142 140 176
rect 174 142 190 176
rect 124 108 190 142
rect 224 204 290 210
rect 224 170 240 204
rect 274 170 290 204
rect 341 202 362 210
rect 224 152 290 170
rect 396 176 412 210
rect 224 136 326 152
rect 24 67 40 101
rect 74 67 90 101
rect 24 51 90 67
rect 224 102 276 136
rect 310 102 326 136
rect 224 17 326 102
rect 362 120 412 176
rect 396 86 412 120
rect 362 70 412 86
rect 526 197 592 202
rect 526 163 542 197
rect 576 163 592 197
rect 526 120 592 163
rect 526 86 542 120
rect 576 86 592 120
rect 526 17 592 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a21boi_1
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 31 94 65 128 0 FreeSans 340 0 0 0 B1_N
port 3 nsew
flabel corelocali s 31 168 65 202 0 FreeSans 340 0 0 0 B1_N
port 3 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 B1_N
port 3 nsew
flabel corelocali s 223 390 257 424 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 223 464 257 498 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 223 538 257 572 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 511 242 545 276 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 607 242 641 276 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 672 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3988470
string GDS_START 3981668
<< end >>
