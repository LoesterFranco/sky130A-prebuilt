magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 576 289 1363 323
rect 576 255 620 289
rect 1319 255 1363 289
rect 85 215 620 255
rect 654 221 1268 255
rect 654 215 1100 221
rect 1319 215 1624 255
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 17 401 80 493
rect 124 435 174 527
rect 218 401 268 493
rect 312 435 362 527
rect 406 459 832 493
rect 406 401 456 459
rect 594 425 644 459
rect 17 357 456 401
rect 500 391 550 425
rect 688 391 738 425
rect 500 357 738 391
rect 782 359 832 459
rect 886 401 936 493
rect 980 435 1030 527
rect 1074 401 1124 493
rect 1168 435 1218 527
rect 1262 401 1312 493
rect 1356 435 1406 527
rect 1450 401 1500 493
rect 1544 435 1594 527
rect 1638 459 2076 493
rect 1638 401 1688 459
rect 886 357 1688 401
rect 500 323 534 357
rect 17 289 534 323
rect 1450 291 1500 357
rect 1736 333 1794 425
rect 1838 367 1888 459
rect 1932 333 1982 425
rect 2026 359 2076 459
rect 1736 325 1982 333
rect 2110 325 2191 493
rect 1602 289 1702 323
rect 1736 289 2191 325
rect 17 181 51 289
rect 1668 255 1702 289
rect 1668 215 2026 255
rect 1130 181 1226 187
rect 2127 181 2191 289
rect 17 147 746 181
rect 913 179 1226 181
rect 106 145 746 147
rect 17 17 72 113
rect 106 51 182 145
rect 226 17 260 111
rect 294 51 370 145
rect 414 17 448 111
rect 482 51 558 145
rect 602 17 636 111
rect 670 51 746 145
rect 790 17 844 179
rect 913 145 1141 179
rect 1175 145 1226 179
rect 913 129 1226 145
rect 1270 145 1696 181
rect 1730 179 2191 181
rect 1730 145 1753 179
rect 1787 147 2191 179
rect 1787 145 1896 147
rect 1270 95 1320 145
rect 878 51 1320 95
rect 1364 17 1398 111
rect 1432 51 1508 145
rect 1552 17 1586 111
rect 1620 51 1696 145
rect 1752 17 1786 111
rect 1820 51 1896 145
rect 1940 17 1974 111
rect 2008 51 2084 147
rect 2128 17 2162 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 1141 145 1175 179
rect 1753 145 1787 179
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
<< metal1 >>
rect 0 561 2208 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 0 496 2208 527
rect 1129 179 1799 185
rect 1129 145 1141 179
rect 1175 156 1753 179
rect 1175 145 1187 156
rect 1129 139 1187 145
rect 1741 145 1753 156
rect 1787 145 1799 179
rect 1741 139 1799 145
rect 0 17 2208 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
rect 0 -48 2208 -17
<< obsm1 >>
rect 425 320 483 329
rect 1649 320 1707 329
rect 425 292 1707 320
rect 425 283 483 292
rect 1649 283 1707 292
<< labels >>
rlabel locali s 1319 255 1363 289 6 A
port 1 nsew signal input
rlabel locali s 1319 215 1624 255 6 A
port 1 nsew signal input
rlabel locali s 576 289 1363 323 6 A
port 1 nsew signal input
rlabel locali s 576 255 620 289 6 A
port 1 nsew signal input
rlabel locali s 85 215 620 255 6 A
port 1 nsew signal input
rlabel locali s 654 221 1268 255 6 B
port 2 nsew signal input
rlabel locali s 654 215 1100 221 6 B
port 2 nsew signal input
rlabel metal1 s 1741 139 1799 156 6 X
port 3 nsew signal output
rlabel metal1 s 1129 156 1799 185 6 X
port 3 nsew signal output
rlabel metal1 s 1129 139 1187 156 6 X
port 3 nsew signal output
rlabel metal1 s 0 -48 2208 48 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 496 2208 592 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2208 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 780560
string GDS_START 765290
<< end >>
