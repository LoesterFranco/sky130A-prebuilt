magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1012 561
rect 17 427 73 527
rect 21 199 89 391
rect 17 17 69 165
rect 359 324 431 475
rect 467 357 527 475
rect 584 359 634 527
rect 359 199 393 324
rect 467 290 505 357
rect 679 325 729 493
rect 763 359 813 527
rect 847 325 897 493
rect 931 359 981 527
rect 439 199 505 290
rect 551 289 638 323
rect 679 291 993 325
rect 551 199 585 289
rect 945 181 993 291
rect 687 145 993 181
rect 207 17 257 117
rect 397 17 463 97
rect 575 17 651 97
rect 687 51 737 145
rect 771 17 805 111
rect 839 51 905 145
rect 939 17 973 111
rect 0 -17 1012 17
<< obsli1 >>
rect 119 413 157 491
rect 123 265 157 413
rect 207 349 273 490
rect 207 315 325 349
rect 123 199 243 265
rect 123 181 157 199
rect 119 87 157 181
rect 291 165 325 315
rect 619 215 911 249
rect 619 165 653 215
rect 291 131 653 165
rect 323 61 357 131
rect 497 61 531 131
<< metal1 >>
rect 0 496 1012 592
rect 0 -48 1012 48
<< labels >>
rlabel locali s 551 289 638 323 6 A
port 1 nsew signal input
rlabel locali s 551 199 585 289 6 A
port 1 nsew signal input
rlabel locali s 467 357 527 475 6 B
port 2 nsew signal input
rlabel locali s 467 290 505 357 6 B
port 2 nsew signal input
rlabel locali s 439 199 505 290 6 B
port 2 nsew signal input
rlabel locali s 359 324 431 475 6 C
port 3 nsew signal input
rlabel locali s 359 199 393 324 6 C
port 3 nsew signal input
rlabel locali s 21 199 89 391 6 D_N
port 4 nsew signal input
rlabel locali s 945 181 993 291 6 X
port 5 nsew signal output
rlabel locali s 847 325 897 493 6 X
port 5 nsew signal output
rlabel locali s 839 51 905 145 6 X
port 5 nsew signal output
rlabel locali s 687 145 993 181 6 X
port 5 nsew signal output
rlabel locali s 687 51 737 145 6 X
port 5 nsew signal output
rlabel locali s 679 325 729 493 6 X
port 5 nsew signal output
rlabel locali s 679 291 993 325 6 X
port 5 nsew signal output
rlabel locali s 939 17 973 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 771 17 805 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 575 17 651 97 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 397 17 463 97 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 207 17 257 117 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 17 17 69 165 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 1012 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1012 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 931 359 981 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 763 359 813 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 584 359 634 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 17 427 73 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 1012 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 1012 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1012 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1105282
string GDS_START 1096850
<< end >>
