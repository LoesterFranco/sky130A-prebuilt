magic
tech sky130A
magscale 1 2
timestamp 1601050088
<< locali >>
rect 21 260 87 356
rect 121 260 217 356
rect 319 378 369 596
rect 319 344 402 378
rect 368 204 402 344
rect 325 170 402 204
rect 325 158 359 170
rect 293 70 359 158
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 22 390 88 649
rect 128 424 178 596
rect 212 458 278 649
rect 128 390 285 424
rect 251 310 285 390
rect 409 412 459 649
rect 251 244 334 310
rect 251 226 285 244
rect 27 192 285 226
rect 27 70 93 192
rect 191 17 257 158
rect 395 17 457 136
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< metal1 >>
rect 0 683 480 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 0 617 480 649
rect 0 17 480 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
rect 0 -49 480 -17
<< labels >>
rlabel locali s 21 260 87 356 6 A
port 1 nsew signal input
rlabel locali s 121 260 217 356 6 B
port 2 nsew signal input
rlabel locali s 368 204 402 344 6 X
port 3 nsew signal output
rlabel locali s 325 170 402 204 6 X
port 3 nsew signal output
rlabel locali s 325 158 359 170 6 X
port 3 nsew signal output
rlabel locali s 319 378 369 596 6 X
port 3 nsew signal output
rlabel locali s 319 344 402 378 6 X
port 3 nsew signal output
rlabel locali s 293 70 359 158 6 X
port 3 nsew signal output
rlabel metal1 s 0 -49 480 49 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 617 480 715 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 480 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3114526
string GDS_START 3109452
<< end >>
