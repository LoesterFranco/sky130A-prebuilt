magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 25 260 99 356
rect 385 236 551 302
rect 2137 270 2203 356
rect 2315 364 2385 596
rect 2351 230 2385 364
rect 2311 81 2385 230
rect 2601 70 2668 596
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2688 683
rect 21 424 87 596
rect 127 458 161 649
rect 201 581 425 615
rect 21 390 167 424
rect 133 326 167 390
rect 201 364 283 581
rect 133 260 215 326
rect 133 226 167 260
rect 249 226 283 364
rect 23 192 167 226
rect 23 70 73 192
rect 109 17 175 158
rect 211 70 283 226
rect 317 481 357 547
rect 317 202 351 481
rect 391 371 425 581
rect 459 505 493 649
rect 527 581 906 615
rect 527 471 561 581
rect 618 513 716 547
rect 474 405 561 471
rect 595 371 648 471
rect 391 337 648 371
rect 595 291 648 337
rect 682 359 716 513
rect 750 427 800 547
rect 840 498 906 581
rect 1008 532 1074 649
rect 1114 498 1164 596
rect 1204 532 1270 649
rect 840 464 1290 498
rect 840 461 963 464
rect 750 393 895 427
rect 682 325 827 359
rect 595 225 693 291
rect 727 279 827 325
rect 317 168 550 202
rect 727 191 761 279
rect 861 233 895 393
rect 317 115 373 168
rect 409 17 482 134
rect 516 85 550 168
rect 590 157 761 191
rect 795 199 895 233
rect 929 233 963 461
rect 1087 424 1127 430
rect 1121 392 1127 424
rect 1121 390 1170 392
rect 1087 335 1170 390
rect 1224 335 1290 464
rect 1372 420 1483 596
rect 1581 594 1654 649
rect 1700 560 1766 596
rect 1807 594 1873 649
rect 1998 560 2064 596
rect 997 301 1053 333
rect 1342 312 1415 386
rect 1449 380 1483 420
rect 1578 526 2064 560
rect 2209 526 2275 649
rect 1578 414 1644 526
rect 1998 492 2064 526
rect 1678 458 1880 492
rect 1998 458 2277 492
rect 1678 380 1712 458
rect 1846 424 1880 458
rect 1449 346 1712 380
rect 1746 390 1759 424
rect 1793 390 1812 424
rect 1846 390 2034 424
rect 997 267 1297 301
rect 929 199 1029 233
rect 590 119 656 157
rect 795 123 829 199
rect 692 85 829 123
rect 516 51 829 85
rect 863 85 929 165
rect 963 143 1029 199
rect 1063 85 1129 207
rect 863 51 1129 85
rect 1163 17 1229 207
rect 1263 102 1297 267
rect 1342 236 1573 312
rect 1607 202 1641 346
rect 1746 255 1812 390
rect 1860 221 1926 312
rect 1968 284 2034 390
rect 2069 390 2170 424
rect 2069 221 2103 390
rect 2243 330 2277 458
rect 2243 264 2317 330
rect 1344 136 1641 202
rect 1675 187 2178 221
rect 1675 102 1709 187
rect 2243 153 2277 264
rect 1263 68 1709 102
rect 1743 17 1777 153
rect 1813 85 1863 153
rect 1899 119 2277 153
rect 1813 51 2072 85
rect 2211 17 2277 85
rect 2422 317 2472 582
rect 2511 364 2561 649
rect 2422 251 2567 317
rect 2422 70 2472 251
rect 2516 17 2566 162
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2688 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 1087 390 1121 424
rect 1759 390 1793 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
<< metal1 >>
rect 0 683 2688 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2688 683
rect 0 617 2688 649
rect 1075 424 1133 430
rect 1075 390 1087 424
rect 1121 421 1133 424
rect 1747 424 1805 430
rect 1747 421 1759 424
rect 1121 393 1759 421
rect 1121 390 1133 393
rect 1075 384 1133 390
rect 1747 390 1759 393
rect 1793 390 1805 424
rect 1747 384 1805 390
rect 0 17 2688 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2688 17
rect 0 -49 2688 -17
<< obsm1 >>
rect 595 273 653 282
rect 1363 273 1421 282
rect 595 245 1421 273
rect 595 236 653 245
rect 1363 236 1421 245
<< labels >>
rlabel locali s 385 236 551 302 6 D
port 1 nsew signal input
rlabel locali s 2601 70 2668 596 6 Q
port 2 nsew signal output
rlabel locali s 2351 230 2385 364 6 Q_N
port 3 nsew signal output
rlabel locali s 2315 364 2385 596 6 Q_N
port 3 nsew signal output
rlabel locali s 2311 81 2385 230 6 Q_N
port 3 nsew signal output
rlabel locali s 2137 270 2203 356 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 1747 421 1805 430 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1747 384 1805 393 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1075 421 1133 430 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1075 393 1805 421 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1075 384 1133 393 6 SET_B
port 5 nsew signal input
rlabel locali s 25 260 99 356 6 CLK_N
port 6 nsew clock input
rlabel metal1 s 0 -49 2688 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 617 2688 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2688 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 2774134
string GDS_START 2753522
<< end >>
