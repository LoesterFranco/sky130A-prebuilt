magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 95 47 125 177
rect 192 93 222 177
rect 430 47 460 177
rect 526 47 556 177
rect 610 47 640 177
<< pmoshvt >>
rect 81 297 117 497
rect 194 297 230 381
rect 422 297 458 497
rect 518 297 554 497
rect 612 297 648 497
<< ndiff >>
rect 43 149 95 177
rect 43 115 51 149
rect 85 115 95 149
rect 43 47 95 115
rect 125 149 192 177
rect 125 115 135 149
rect 169 115 192 149
rect 125 93 192 115
rect 222 149 284 177
rect 222 115 242 149
rect 276 115 284 149
rect 222 93 284 115
rect 370 131 430 177
rect 370 97 378 131
rect 412 97 430 131
rect 125 47 177 93
rect 370 47 430 97
rect 460 163 526 177
rect 460 129 472 163
rect 506 129 526 163
rect 460 95 526 129
rect 460 61 472 95
rect 506 61 526 95
rect 460 47 526 61
rect 556 95 610 177
rect 556 61 566 95
rect 600 61 610 95
rect 556 47 610 61
rect 640 163 706 177
rect 640 129 663 163
rect 697 129 706 163
rect 640 95 706 129
rect 640 61 663 95
rect 697 61 706 95
rect 640 47 706 61
<< pdiff >>
rect 27 482 81 497
rect 27 448 35 482
rect 69 448 81 482
rect 27 414 81 448
rect 27 380 35 414
rect 69 380 81 414
rect 27 346 81 380
rect 27 312 35 346
rect 69 312 81 346
rect 27 297 81 312
rect 117 475 177 497
rect 117 441 135 475
rect 169 441 177 475
rect 117 381 177 441
rect 362 477 422 497
rect 362 443 370 477
rect 404 443 422 477
rect 117 297 194 381
rect 230 339 288 381
rect 230 305 242 339
rect 276 305 288 339
rect 230 297 288 305
rect 362 297 422 443
rect 458 477 518 497
rect 458 443 472 477
rect 506 443 518 477
rect 458 409 518 443
rect 458 375 472 409
rect 506 375 518 409
rect 458 341 518 375
rect 458 307 472 341
rect 506 307 518 341
rect 458 297 518 307
rect 554 297 612 497
rect 648 477 706 497
rect 648 443 660 477
rect 694 443 706 477
rect 648 409 706 443
rect 648 375 660 409
rect 694 375 706 409
rect 648 341 706 375
rect 648 307 660 341
rect 694 307 706 341
rect 648 297 706 307
<< ndiffc >>
rect 51 115 85 149
rect 135 115 169 149
rect 242 115 276 149
rect 378 97 412 131
rect 472 129 506 163
rect 472 61 506 95
rect 566 61 600 95
rect 663 129 697 163
rect 663 61 697 95
<< pdiffc >>
rect 35 448 69 482
rect 35 380 69 414
rect 35 312 69 346
rect 135 441 169 475
rect 370 443 404 477
rect 242 305 276 339
rect 472 443 506 477
rect 472 375 506 409
rect 472 307 506 341
rect 660 443 694 477
rect 660 375 694 409
rect 660 307 694 341
<< poly >>
rect 81 497 117 523
rect 422 497 458 523
rect 518 497 554 523
rect 612 497 648 523
rect 194 381 230 407
rect 81 282 117 297
rect 194 282 230 297
rect 422 282 458 297
rect 518 282 554 297
rect 612 282 648 297
rect 79 265 119 282
rect 192 265 232 282
rect 420 265 460 282
rect 516 265 556 282
rect 79 249 146 265
rect 79 215 102 249
rect 136 215 146 249
rect 79 199 146 215
rect 192 249 254 265
rect 192 215 210 249
rect 244 215 254 249
rect 192 199 254 215
rect 300 249 460 265
rect 300 215 310 249
rect 344 215 460 249
rect 300 199 460 215
rect 502 249 556 265
rect 502 215 512 249
rect 546 215 556 249
rect 502 199 556 215
rect 95 177 125 199
rect 192 177 222 199
rect 430 177 460 199
rect 526 177 556 199
rect 610 265 650 282
rect 610 249 664 265
rect 610 215 620 249
rect 654 215 664 249
rect 610 199 664 215
rect 610 177 640 199
rect 192 67 222 93
rect 95 21 125 47
rect 430 21 460 47
rect 526 21 556 47
rect 610 21 640 47
<< polycont >>
rect 102 215 136 249
rect 210 215 244 249
rect 310 215 344 249
rect 512 215 546 249
rect 620 215 654 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 17 482 85 493
rect 17 448 35 482
rect 69 448 85 482
rect 17 414 85 448
rect 119 475 201 527
rect 119 441 135 475
rect 169 441 201 475
rect 354 477 420 527
rect 354 443 370 477
rect 404 443 420 477
rect 456 477 517 493
rect 456 443 472 477
rect 506 443 517 477
rect 17 380 35 414
rect 69 380 85 414
rect 456 409 517 443
rect 456 407 472 409
rect 17 346 85 380
rect 17 312 35 346
rect 69 312 85 346
rect 17 296 85 312
rect 129 375 472 407
rect 506 375 517 409
rect 129 373 517 375
rect 17 165 68 296
rect 129 265 172 373
rect 378 341 517 373
rect 215 305 242 339
rect 276 305 344 339
rect 102 249 172 265
rect 136 215 172 249
rect 102 199 172 215
rect 206 249 276 265
rect 206 215 210 249
rect 244 215 276 249
rect 206 199 276 215
rect 310 249 344 305
rect 310 165 344 215
rect 17 149 89 165
rect 17 115 51 149
rect 85 115 89 149
rect 17 90 89 115
rect 135 149 169 165
rect 135 17 169 115
rect 242 149 344 165
rect 276 131 344 149
rect 378 307 472 341
rect 506 307 517 341
rect 634 477 710 527
rect 634 443 660 477
rect 694 443 710 477
rect 634 409 710 443
rect 634 375 660 409
rect 694 375 710 409
rect 634 341 710 375
rect 634 307 660 341
rect 694 307 710 341
rect 378 291 517 307
rect 378 131 412 291
rect 446 249 570 257
rect 446 215 512 249
rect 546 215 570 249
rect 604 249 714 257
rect 604 215 620 249
rect 654 215 714 249
rect 242 90 276 115
rect 378 51 412 97
rect 456 163 713 181
rect 456 129 472 163
rect 506 147 663 163
rect 506 129 522 147
rect 456 95 522 129
rect 647 129 663 147
rect 697 129 713 163
rect 456 61 472 95
rect 506 61 522 95
rect 456 51 522 61
rect 566 95 600 111
rect 566 17 600 61
rect 647 95 713 129
rect 647 61 663 95
rect 697 61 713 95
rect 647 54 713 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel corelocali s 213 221 247 255 0 FreeSans 400 0 0 0 B1_N
port 3 nsew
flabel corelocali s 674 238 674 238 0 FreeSans 400 0 0 0 A1
port 1 nsew
flabel corelocali s 29 425 63 459 0 FreeSans 400 0 0 0 X
port 8 nsew
flabel corelocali s 490 238 490 238 0 FreeSans 400 0 0 0 A2
port 2 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
rlabel comment s 0 0 0 0 4 o21ba_1
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 994076
string GDS_START 987844
<< end >>
