magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 2852 561
rect 103 427 169 527
rect 17 195 87 325
rect 286 377 357 527
rect 662 443 728 527
rect 103 17 169 93
rect 283 205 339 337
rect 387 230 431 339
rect 765 335 812 475
rect 387 163 463 230
rect 755 315 812 335
rect 755 281 821 315
rect 286 17 341 127
rect 387 69 431 163
rect 1141 441 1217 527
rect 1435 383 1501 527
rect 1924 451 2000 527
rect 1174 193 1243 213
rect 1174 147 1259 193
rect 2188 451 2466 527
rect 645 17 711 89
rect 1167 17 1201 105
rect 1951 147 2026 213
rect 2500 326 2557 493
rect 2307 219 2398 265
rect 1524 17 1595 93
rect 1912 17 1964 105
rect 2400 17 2466 161
rect 2521 143 2557 326
rect 2500 51 2557 143
rect 2691 353 2748 527
rect 2783 294 2835 493
rect 2793 157 2835 294
rect 2691 17 2749 109
rect 2783 51 2835 157
rect 0 -17 2852 17
<< obsli1 >>
rect 19 393 69 493
rect 19 359 167 393
rect 121 187 167 359
rect 19 153 121 161
rect 155 153 167 187
rect 19 127 167 153
rect 203 391 247 493
rect 203 357 213 391
rect 443 375 515 477
rect 594 381 628 493
rect 19 69 69 127
rect 203 69 247 357
rect 481 301 515 375
rect 552 349 628 381
rect 552 315 721 349
rect 846 427 889 493
rect 927 450 1093 484
rect 481 293 521 301
rect 481 286 526 293
rect 481 281 534 286
rect 481 259 615 281
rect 492 255 615 259
rect 492 251 581 255
rect 497 221 581 251
rect 497 215 615 221
rect 686 219 721 315
rect 855 261 889 427
rect 849 255 889 261
rect 845 247 846 255
rect 790 221 846 247
rect 880 235 889 255
rect 923 357 949 391
rect 983 357 1025 391
rect 923 315 1025 357
rect 880 221 882 235
rect 497 119 531 215
rect 686 159 754 219
rect 465 53 531 119
rect 574 153 754 159
rect 790 213 880 221
rect 574 125 729 153
rect 574 61 608 125
rect 790 119 824 213
rect 923 207 958 315
rect 1059 281 1093 450
rect 1277 407 1311 475
rect 1127 357 1397 407
rect 1710 450 1876 484
rect 1672 391 1719 397
rect 1127 315 1177 357
rect 1279 281 1329 297
rect 1059 247 1329 281
rect 1059 239 1134 247
rect 914 141 958 207
rect 1000 187 1066 203
rect 1000 153 1031 187
rect 1065 153 1066 187
rect 1000 147 1066 153
rect 1100 131 1134 239
rect 1285 231 1329 247
rect 1363 213 1397 357
rect 1672 357 1685 391
rect 1431 323 1632 331
rect 1431 289 1593 323
rect 1627 289 1632 323
rect 1672 315 1719 357
rect 1431 283 1632 289
rect 1431 247 1497 283
rect 1767 261 1808 381
rect 1684 255 1808 261
rect 1559 213 1625 247
rect 1363 212 1625 213
rect 1362 179 1625 212
rect 1684 221 1685 255
rect 1719 225 1808 255
rect 1842 281 1876 450
rect 2048 417 2082 475
rect 1910 383 2466 417
rect 1910 315 1960 383
rect 1842 247 2112 281
rect 1719 221 1741 225
rect 1362 156 1402 179
rect 790 85 866 119
rect 1097 117 1134 131
rect 1336 122 1402 156
rect 1097 93 1131 117
rect 832 53 866 85
rect 911 53 1131 93
rect 1252 85 1318 93
rect 1436 85 1470 143
rect 1684 141 1741 221
rect 1842 93 1876 247
rect 2068 215 2112 247
rect 2146 156 2181 383
rect 2115 119 2181 156
rect 2216 323 2371 349
rect 2216 289 2237 323
rect 2271 315 2371 323
rect 2216 185 2271 289
rect 2432 265 2466 383
rect 2432 199 2485 265
rect 2216 151 2355 185
rect 1252 51 1470 85
rect 1723 53 1876 93
rect 2016 85 2082 109
rect 2215 85 2250 117
rect 2016 51 2250 85
rect 2313 53 2355 151
rect 2592 265 2655 483
rect 2592 199 2759 265
rect 2592 51 2655 199
<< obsli1c >>
rect 121 153 155 187
rect 213 357 247 391
rect 581 221 615 255
rect 846 221 880 255
rect 949 357 983 391
rect 1031 153 1065 187
rect 1685 357 1719 391
rect 1593 289 1627 323
rect 1685 221 1719 255
rect 2237 289 2271 323
<< metal1 >>
rect 0 496 2852 592
rect 1213 184 1271 193
rect 1949 184 2007 193
rect 1213 156 2007 184
rect 1213 147 1271 156
rect 1949 147 2007 156
rect 0 -48 2852 48
<< obsm1 >>
rect 201 391 259 397
rect 201 357 213 391
rect 247 388 259 391
rect 937 391 995 397
rect 937 388 949 391
rect 247 360 949 388
rect 247 357 259 360
rect 201 351 259 357
rect 937 357 949 360
rect 983 388 995 391
rect 1673 391 1731 397
rect 1673 388 1685 391
rect 983 360 1685 388
rect 983 357 995 360
rect 937 351 995 357
rect 1673 357 1685 360
rect 1719 357 1731 391
rect 1673 351 1731 357
rect 1581 323 1639 329
rect 1581 289 1593 323
rect 1627 320 1639 323
rect 2225 323 2283 329
rect 2225 320 2237 323
rect 1627 292 2237 320
rect 1627 289 1639 292
rect 1581 283 1639 289
rect 2225 289 2237 292
rect 2271 289 2283 323
rect 2225 283 2283 289
rect 569 255 627 261
rect 569 221 581 255
rect 615 252 627 255
rect 834 255 892 261
rect 834 252 846 255
rect 615 224 846 252
rect 615 221 627 224
rect 569 215 627 221
rect 834 221 846 224
rect 880 221 892 255
rect 1673 255 1731 261
rect 1673 252 1685 255
rect 834 215 892 221
rect 1034 224 1685 252
rect 1034 193 1077 224
rect 1673 221 1685 224
rect 1719 221 1731 255
rect 1673 215 1731 221
rect 109 187 167 193
rect 109 153 121 187
rect 155 184 167 187
rect 1019 187 1077 193
rect 1019 184 1031 187
rect 155 156 1031 184
rect 155 153 167 156
rect 109 147 167 153
rect 1019 153 1031 156
rect 1065 153 1077 187
rect 1019 147 1077 153
<< labels >>
rlabel locali s 765 335 812 475 6 D
port 1 nsew signal input
rlabel locali s 755 315 812 335 6 D
port 1 nsew signal input
rlabel locali s 755 281 821 315 6 D
port 1 nsew signal input
rlabel locali s 2793 157 2835 294 6 Q
port 2 nsew signal output
rlabel locali s 2783 294 2835 493 6 Q
port 2 nsew signal output
rlabel locali s 2783 51 2835 157 6 Q
port 2 nsew signal output
rlabel locali s 2521 143 2557 326 6 Q_N
port 3 nsew signal output
rlabel locali s 2500 326 2557 493 6 Q_N
port 3 nsew signal output
rlabel locali s 2500 51 2557 143 6 Q_N
port 3 nsew signal output
rlabel locali s 2307 219 2398 265 6 RESET_B
port 4 nsew signal input
rlabel locali s 283 205 339 337 6 SCD
port 5 nsew signal input
rlabel locali s 387 230 431 339 6 SCE
port 6 nsew signal input
rlabel locali s 387 163 463 230 6 SCE
port 6 nsew signal input
rlabel locali s 387 69 431 163 6 SCE
port 6 nsew signal input
rlabel locali s 1174 193 1243 213 6 SET_B
port 7 nsew signal input
rlabel locali s 1174 147 1259 193 6 SET_B
port 7 nsew signal input
rlabel locali s 1951 147 2026 213 6 SET_B
port 7 nsew signal input
rlabel metal1 s 1949 184 2007 193 6 SET_B
port 7 nsew signal input
rlabel metal1 s 1949 147 2007 156 6 SET_B
port 7 nsew signal input
rlabel metal1 s 1213 184 1271 193 6 SET_B
port 7 nsew signal input
rlabel metal1 s 1213 156 2007 184 6 SET_B
port 7 nsew signal input
rlabel metal1 s 1213 147 1271 156 6 SET_B
port 7 nsew signal input
rlabel locali s 17 195 87 325 6 CLK_N
port 8 nsew clock input
rlabel locali s 2691 17 2749 109 6 VGND
port 9 nsew ground bidirectional abutment
rlabel locali s 2400 17 2466 161 6 VGND
port 9 nsew ground bidirectional abutment
rlabel locali s 1912 17 1964 105 6 VGND
port 9 nsew ground bidirectional abutment
rlabel locali s 1524 17 1595 93 6 VGND
port 9 nsew ground bidirectional abutment
rlabel locali s 1167 17 1201 105 6 VGND
port 9 nsew ground bidirectional abutment
rlabel locali s 645 17 711 89 6 VGND
port 9 nsew ground bidirectional abutment
rlabel locali s 286 17 341 127 6 VGND
port 9 nsew ground bidirectional abutment
rlabel locali s 103 17 169 93 6 VGND
port 9 nsew ground bidirectional abutment
rlabel locali s 0 -17 2852 17 8 VGND
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 2852 48 8 VGND
port 9 nsew ground bidirectional abutment
rlabel locali s 2691 353 2748 527 6 VPWR
port 10 nsew power bidirectional abutment
rlabel locali s 2188 451 2466 527 6 VPWR
port 10 nsew power bidirectional abutment
rlabel locali s 1924 451 2000 527 6 VPWR
port 10 nsew power bidirectional abutment
rlabel locali s 1435 383 1501 527 6 VPWR
port 10 nsew power bidirectional abutment
rlabel locali s 1141 441 1217 527 6 VPWR
port 10 nsew power bidirectional abutment
rlabel locali s 662 443 728 527 6 VPWR
port 10 nsew power bidirectional abutment
rlabel locali s 286 377 357 527 6 VPWR
port 10 nsew power bidirectional abutment
rlabel locali s 103 427 169 527 6 VPWR
port 10 nsew power bidirectional abutment
rlabel locali s 0 527 2852 561 6 VPWR
port 10 nsew power bidirectional abutment
rlabel metal1 s 0 496 2852 592 6 VPWR
port 10 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2852 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 54774
string GDS_START 31832
<< end >>
