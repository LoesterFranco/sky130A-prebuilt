magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 1353 325 1403 425
rect 1541 325 1591 425
rect 1353 291 1591 325
rect 79 215 401 257
rect 455 215 830 257
rect 877 215 1257 257
rect 1353 181 1450 291
rect 1771 215 1910 257
rect 103 145 1599 181
rect 103 51 179 145
rect 291 51 367 145
rect 479 51 555 145
rect 667 51 743 145
rect 959 51 1035 145
rect 1147 51 1223 145
rect 1335 51 1411 145
rect 1523 51 1599 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 19 325 85 493
rect 129 359 171 527
rect 215 325 265 493
rect 309 359 359 527
rect 403 459 829 493
rect 403 325 453 459
rect 19 291 453 325
rect 497 325 547 425
rect 591 359 641 459
rect 685 325 735 425
rect 779 359 829 459
rect 883 459 1685 493
rect 883 359 933 459
rect 977 325 1027 425
rect 1071 359 1121 459
rect 1165 325 1215 425
rect 497 291 1215 325
rect 1259 291 1309 459
rect 1447 359 1497 459
rect 1635 359 1685 459
rect 1730 325 1797 493
rect 1654 291 1797 325
rect 1841 291 1887 527
rect 1654 257 1688 291
rect 1484 215 1688 257
rect 1654 181 1688 215
rect 35 17 69 179
rect 1654 147 1797 181
rect 223 17 257 111
rect 411 17 445 111
rect 599 17 633 111
rect 787 17 925 111
rect 1079 17 1113 111
rect 1267 17 1301 111
rect 1455 17 1489 111
rect 1643 17 1677 111
rect 1722 51 1797 147
rect 1841 17 1887 181
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< labels >>
rlabel locali s 79 215 401 257 6 A
port 1 nsew signal input
rlabel locali s 455 215 830 257 6 B
port 2 nsew signal input
rlabel locali s 877 215 1257 257 6 C
port 3 nsew signal input
rlabel locali s 1771 215 1910 257 6 D_N
port 4 nsew signal input
rlabel locali s 1541 325 1591 425 6 Y
port 5 nsew signal output
rlabel locali s 1523 51 1599 145 6 Y
port 5 nsew signal output
rlabel locali s 1353 325 1403 425 6 Y
port 5 nsew signal output
rlabel locali s 1353 291 1591 325 6 Y
port 5 nsew signal output
rlabel locali s 1353 181 1450 291 6 Y
port 5 nsew signal output
rlabel locali s 1335 51 1411 145 6 Y
port 5 nsew signal output
rlabel locali s 1147 51 1223 145 6 Y
port 5 nsew signal output
rlabel locali s 959 51 1035 145 6 Y
port 5 nsew signal output
rlabel locali s 667 51 743 145 6 Y
port 5 nsew signal output
rlabel locali s 479 51 555 145 6 Y
port 5 nsew signal output
rlabel locali s 291 51 367 145 6 Y
port 5 nsew signal output
rlabel locali s 103 145 1599 181 6 Y
port 5 nsew signal output
rlabel locali s 103 51 179 145 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -48 1932 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 1932 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1932 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2530600
string GDS_START 2516274
<< end >>
