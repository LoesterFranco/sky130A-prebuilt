magic
tech sky130A
magscale 1 2
timestamp 1604502729
<< locali >>
rect 95 196 161 398
rect 263 236 355 310
rect 2235 416 2291 596
rect 2425 430 2471 596
rect 2425 416 2567 430
rect 2235 364 2567 416
rect 2521 230 2567 364
rect 2136 196 2567 230
rect 2136 70 2202 196
rect 2403 70 2469 196
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2592 683
rect 23 482 73 592
rect 113 516 179 649
rect 315 516 381 649
rect 421 581 759 615
rect 421 482 455 581
rect 23 448 359 482
rect 489 459 589 547
rect 623 459 691 547
rect 489 448 523 459
rect 23 162 57 448
rect 325 414 523 448
rect 195 378 291 414
rect 195 344 455 378
rect 195 202 229 344
rect 389 270 455 344
rect 23 70 73 162
rect 109 17 159 162
rect 195 68 287 202
rect 323 17 373 202
rect 409 85 443 226
rect 489 185 523 414
rect 557 291 623 425
rect 489 119 555 185
rect 589 85 623 291
rect 409 51 623 85
rect 657 260 691 459
rect 725 467 759 581
rect 797 551 831 649
rect 903 581 1102 615
rect 797 501 869 551
rect 903 467 937 581
rect 725 433 937 467
rect 971 459 1034 547
rect 725 294 759 433
rect 971 399 1005 459
rect 1068 453 1102 581
rect 1136 487 1188 649
rect 1318 530 1453 596
rect 1577 530 1611 649
rect 1334 496 1543 530
rect 1651 496 1717 596
rect 1756 530 1806 649
rect 1846 530 1912 596
rect 1068 419 1295 453
rect 823 348 1005 399
rect 1039 350 1127 385
rect 1039 316 1087 350
rect 1121 316 1127 350
rect 793 280 1005 314
rect 1039 310 1127 316
rect 793 260 827 280
rect 657 226 827 260
rect 954 274 1005 280
rect 1161 274 1227 298
rect 657 70 707 226
rect 861 190 918 246
rect 954 240 1227 274
rect 1261 290 1295 419
rect 1334 358 1368 496
rect 1509 462 1822 496
rect 1409 404 1475 462
rect 1334 324 1407 358
rect 954 224 1005 240
rect 1261 224 1339 290
rect 861 156 1010 190
rect 918 124 1010 156
rect 805 17 884 120
rect 1134 17 1200 206
rect 1261 85 1295 224
rect 1373 185 1407 324
rect 1329 119 1407 185
rect 1441 85 1475 404
rect 1637 350 1703 370
rect 1509 202 1575 331
rect 1637 316 1663 350
rect 1697 316 1703 350
rect 1637 236 1703 316
rect 1756 274 1822 462
rect 1856 202 1890 530
rect 1951 364 2001 649
rect 2041 330 2107 540
rect 2145 364 2201 649
rect 2325 450 2391 649
rect 2505 464 2571 649
rect 2041 298 2399 330
rect 1509 168 1890 202
rect 1261 51 1475 85
rect 1587 17 1790 134
rect 1824 84 1890 168
rect 1936 264 2399 298
rect 1936 70 2002 264
rect 2036 17 2102 226
rect 2236 17 2369 160
rect 2503 17 2569 162
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2592 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 1087 316 1121 350
rect 1663 316 1697 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
<< metal1 >>
rect 0 683 2592 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2592 683
rect 0 617 2592 649
rect 1075 350 1133 356
rect 1075 316 1087 350
rect 1121 347 1133 350
rect 1651 350 1709 356
rect 1651 347 1663 350
rect 1121 319 1663 347
rect 1121 316 1133 319
rect 1075 310 1133 316
rect 1651 316 1663 319
rect 1697 316 1709 350
rect 1651 310 1709 316
rect 0 17 2592 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2592 17
rect 0 -49 2592 -17
<< labels >>
rlabel locali s 95 196 161 398 6 D
port 1 nsew signal input
rlabel locali s 2521 230 2567 364 6 Q
port 2 nsew signal output
rlabel locali s 2425 430 2471 596 6 Q
port 2 nsew signal output
rlabel locali s 2425 416 2567 430 6 Q
port 2 nsew signal output
rlabel locali s 2403 70 2469 196 6 Q
port 2 nsew signal output
rlabel locali s 2235 416 2291 596 6 Q
port 2 nsew signal output
rlabel locali s 2235 364 2567 416 6 Q
port 2 nsew signal output
rlabel locali s 2136 196 2567 230 6 Q
port 2 nsew signal output
rlabel locali s 2136 70 2202 196 6 Q
port 2 nsew signal output
rlabel metal1 s 1651 347 1709 356 6 SET_B
port 3 nsew signal input
rlabel metal1 s 1651 310 1709 319 6 SET_B
port 3 nsew signal input
rlabel metal1 s 1075 347 1133 356 6 SET_B
port 3 nsew signal input
rlabel metal1 s 1075 319 1709 347 6 SET_B
port 3 nsew signal input
rlabel metal1 s 1075 310 1133 319 6 SET_B
port 3 nsew signal input
rlabel locali s 263 236 355 310 6 CLK
port 4 nsew clock input
rlabel metal1 s 0 -49 2592 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 617 2592 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2592 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 2835402
string GDS_START 2816604
<< end >>
