magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 106 357 306 493
rect 18 137 72 265
rect 106 165 150 357
rect 184 199 261 323
rect 295 199 349 323
rect 383 199 441 493
rect 479 199 598 265
rect 106 131 179 165
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 18 299 72 527
rect 557 299 627 527
rect 213 131 511 165
rect 213 97 288 131
rect 17 51 288 97
rect 329 17 395 97
rect 477 75 511 131
rect 545 17 619 165
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 479 199 598 265 6 A1
port 1 nsew signal input
rlabel locali s 383 199 441 493 6 A2
port 2 nsew signal input
rlabel locali s 295 199 349 323 6 A3
port 3 nsew signal input
rlabel locali s 18 137 72 265 6 B1
port 4 nsew signal input
rlabel locali s 184 199 261 323 6 B2
port 5 nsew signal input
rlabel locali s 106 357 306 493 6 Y
port 6 nsew signal output
rlabel locali s 106 165 150 357 6 Y
port 6 nsew signal output
rlabel locali s 106 131 179 165 6 Y
port 6 nsew signal output
rlabel metal1 s 0 -48 644 48 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 580764
string GDS_START 574152
<< end >>
