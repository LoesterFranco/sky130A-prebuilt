magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 2438 704
rect 193 322 1343 332
rect 1135 305 1343 322
<< pwell >>
rect 0 0 2400 49
<< scnmos >>
rect 84 80 114 164
rect 282 74 312 222
rect 368 74 398 222
rect 566 81 596 165
rect 718 81 748 165
rect 796 81 826 165
rect 1031 74 1061 158
rect 1109 74 1139 158
rect 1232 74 1262 202
rect 1330 74 1360 202
rect 1432 74 1462 158
rect 1510 74 1540 158
rect 1588 74 1618 158
rect 1760 74 1790 158
rect 1972 74 2002 222
rect 2170 74 2200 184
rect 2286 74 2316 222
<< pmoshvt >>
rect 86 508 116 592
rect 288 358 318 582
rect 378 358 408 582
rect 598 463 628 547
rect 698 463 728 547
rect 782 463 812 547
rect 963 463 993 547
rect 1065 463 1095 547
rect 1224 341 1254 541
rect 1325 377 1355 577
rect 1487 508 1517 592
rect 1571 508 1601 592
rect 1661 508 1691 592
rect 1880 508 1910 592
rect 1981 368 2011 592
rect 2183 403 2213 571
rect 2284 368 2314 592
<< ndiff >>
rect 225 197 282 222
rect 27 139 84 164
rect 27 105 39 139
rect 73 105 84 139
rect 27 80 84 105
rect 114 139 171 164
rect 114 105 125 139
rect 159 105 171 139
rect 114 80 171 105
rect 225 163 237 197
rect 271 163 282 197
rect 225 120 282 163
rect 225 86 237 120
rect 271 86 282 120
rect 225 74 282 86
rect 312 186 368 222
rect 312 152 323 186
rect 357 152 368 186
rect 312 118 368 152
rect 312 84 323 118
rect 357 84 368 118
rect 312 74 368 84
rect 398 210 455 222
rect 398 176 409 210
rect 443 176 455 210
rect 398 120 455 176
rect 398 86 409 120
rect 443 86 455 120
rect 398 74 455 86
rect 509 153 566 165
rect 509 119 521 153
rect 555 119 566 153
rect 509 81 566 119
rect 596 140 718 165
rect 596 106 673 140
rect 707 106 718 140
rect 596 81 718 106
rect 748 81 796 165
rect 826 127 883 165
rect 1175 189 1232 202
rect 1175 158 1187 189
rect 826 93 837 127
rect 871 93 883 127
rect 826 81 883 93
rect 978 137 1031 158
rect 978 103 986 137
rect 1020 103 1031 137
rect 978 74 1031 103
rect 1061 74 1109 158
rect 1139 155 1187 158
rect 1221 155 1232 189
rect 1139 116 1232 155
rect 1139 82 1187 116
rect 1221 82 1232 116
rect 1139 74 1232 82
rect 1262 74 1330 202
rect 1360 169 1417 202
rect 1360 135 1371 169
rect 1405 158 1417 169
rect 1405 135 1432 158
rect 1360 74 1432 135
rect 1462 74 1510 158
rect 1540 74 1588 158
rect 1618 128 1760 158
rect 1618 94 1629 128
rect 1663 94 1701 128
rect 1735 94 1760 128
rect 1618 74 1760 94
rect 1790 133 1847 158
rect 1790 99 1801 133
rect 1835 99 1847 133
rect 1790 74 1847 99
rect 1901 127 1972 222
rect 1901 93 1913 127
rect 1947 93 1972 127
rect 1901 74 1972 93
rect 2002 210 2059 222
rect 2002 176 2013 210
rect 2047 176 2059 210
rect 2215 184 2286 222
rect 2002 120 2059 176
rect 2002 86 2013 120
rect 2047 86 2059 120
rect 2002 74 2059 86
rect 2113 146 2170 184
rect 2113 112 2125 146
rect 2159 112 2170 146
rect 2113 74 2170 112
rect 2200 150 2227 184
rect 2261 150 2286 184
rect 2200 116 2286 150
rect 2200 82 2227 116
rect 2261 82 2286 116
rect 2200 74 2286 82
rect 2316 194 2373 222
rect 2316 160 2327 194
rect 2361 160 2373 194
rect 2316 120 2373 160
rect 2316 86 2327 120
rect 2361 86 2373 120
rect 2316 74 2373 86
<< pdiff >>
rect 27 567 86 592
rect 27 533 39 567
rect 73 533 86 567
rect 27 508 86 533
rect 116 568 175 592
rect 116 534 129 568
rect 163 534 175 568
rect 116 508 175 534
rect 229 404 288 582
rect 229 370 241 404
rect 275 370 288 404
rect 229 358 288 370
rect 318 556 378 582
rect 318 522 331 556
rect 365 522 378 556
rect 318 358 378 522
rect 408 530 467 582
rect 408 496 421 530
rect 455 496 467 530
rect 408 358 467 496
rect 1434 577 1487 592
rect 1130 547 1206 555
rect 539 520 598 547
rect 539 486 551 520
rect 585 486 598 520
rect 539 463 598 486
rect 628 520 698 547
rect 628 486 651 520
rect 685 486 698 520
rect 628 463 698 486
rect 728 463 782 547
rect 812 535 963 547
rect 812 501 831 535
rect 865 501 963 535
rect 812 463 963 501
rect 993 520 1065 547
rect 993 486 1006 520
rect 1040 486 1065 520
rect 993 463 1065 486
rect 1095 543 1206 547
rect 1095 509 1151 543
rect 1185 541 1206 543
rect 1272 541 1325 577
rect 1185 509 1224 541
rect 1095 463 1224 509
rect 1171 341 1224 463
rect 1254 377 1325 541
rect 1355 565 1487 577
rect 1355 531 1368 565
rect 1402 531 1440 565
rect 1474 531 1487 565
rect 1355 508 1487 531
rect 1517 508 1571 592
rect 1601 580 1661 592
rect 1601 546 1614 580
rect 1648 546 1661 580
rect 1601 508 1661 546
rect 1691 567 1750 592
rect 1691 533 1704 567
rect 1738 533 1750 567
rect 1691 508 1750 533
rect 1804 567 1880 592
rect 1804 533 1816 567
rect 1850 533 1880 567
rect 1804 508 1880 533
rect 1910 580 1981 592
rect 1910 546 1930 580
rect 1964 546 1981 580
rect 1910 508 1981 546
rect 1355 469 1414 508
rect 1355 435 1368 469
rect 1402 435 1414 469
rect 1355 377 1414 435
rect 1254 341 1307 377
rect 1928 368 1981 508
rect 2011 580 2070 592
rect 2011 546 2024 580
rect 2058 546 2070 580
rect 2231 571 2284 592
rect 2011 497 2070 546
rect 2011 463 2024 497
rect 2058 463 2070 497
rect 2011 414 2070 463
rect 2011 380 2024 414
rect 2058 380 2070 414
rect 2124 559 2183 571
rect 2124 525 2136 559
rect 2170 525 2183 559
rect 2124 449 2183 525
rect 2124 415 2136 449
rect 2170 415 2183 449
rect 2124 403 2183 415
rect 2213 559 2284 571
rect 2213 525 2226 559
rect 2260 525 2284 559
rect 2213 449 2284 525
rect 2213 415 2226 449
rect 2260 415 2284 449
rect 2213 403 2284 415
rect 2011 368 2070 380
rect 2231 368 2284 403
rect 2314 580 2373 592
rect 2314 546 2327 580
rect 2361 546 2373 580
rect 2314 497 2373 546
rect 2314 463 2327 497
rect 2361 463 2373 497
rect 2314 414 2373 463
rect 2314 380 2327 414
rect 2361 380 2373 414
rect 2314 368 2373 380
<< ndiffc >>
rect 39 105 73 139
rect 125 105 159 139
rect 237 163 271 197
rect 237 86 271 120
rect 323 152 357 186
rect 323 84 357 118
rect 409 176 443 210
rect 409 86 443 120
rect 521 119 555 153
rect 673 106 707 140
rect 837 93 871 127
rect 986 103 1020 137
rect 1187 155 1221 189
rect 1187 82 1221 116
rect 1371 135 1405 169
rect 1629 94 1663 128
rect 1701 94 1735 128
rect 1801 99 1835 133
rect 1913 93 1947 127
rect 2013 176 2047 210
rect 2013 86 2047 120
rect 2125 112 2159 146
rect 2227 150 2261 184
rect 2227 82 2261 116
rect 2327 160 2361 194
rect 2327 86 2361 120
<< pdiffc >>
rect 39 533 73 567
rect 129 534 163 568
rect 241 370 275 404
rect 331 522 365 556
rect 421 496 455 530
rect 551 486 585 520
rect 651 486 685 520
rect 831 501 865 535
rect 1006 486 1040 520
rect 1151 509 1185 543
rect 1368 531 1402 565
rect 1440 531 1474 565
rect 1614 546 1648 580
rect 1704 533 1738 567
rect 1816 533 1850 567
rect 1930 546 1964 580
rect 1368 435 1402 469
rect 2024 546 2058 580
rect 2024 463 2058 497
rect 2024 380 2058 414
rect 2136 525 2170 559
rect 2136 415 2170 449
rect 2226 525 2260 559
rect 2226 415 2260 449
rect 2327 546 2361 580
rect 2327 463 2361 497
rect 2327 380 2361 414
<< poly >>
rect 86 592 116 618
rect 482 615 1358 645
rect 288 582 318 608
rect 378 582 408 608
rect 86 493 116 508
rect 83 404 119 493
rect 83 388 161 404
rect 83 354 111 388
rect 145 354 161 388
rect 83 320 161 354
rect 288 343 318 358
rect 378 343 408 358
rect 83 286 111 320
rect 145 286 161 320
rect 285 310 321 343
rect 375 326 411 343
rect 482 326 512 615
rect 598 547 628 573
rect 695 562 731 615
rect 1322 592 1358 615
rect 1487 592 1517 618
rect 1571 592 1601 618
rect 1661 592 1691 618
rect 1880 592 1910 618
rect 1981 592 2011 618
rect 1325 577 1355 592
rect 698 547 728 562
rect 782 547 812 573
rect 963 547 993 573
rect 1065 547 1095 573
rect 1224 541 1254 567
rect 598 448 628 463
rect 595 421 631 448
rect 698 437 728 463
rect 782 448 812 463
rect 963 448 993 463
rect 1065 448 1095 463
rect 375 310 512 326
rect 83 252 161 286
rect 83 218 111 252
rect 145 218 161 252
rect 260 294 326 310
rect 260 260 276 294
rect 310 260 326 294
rect 375 290 421 310
rect 260 244 326 260
rect 368 276 421 290
rect 455 276 512 310
rect 573 405 639 421
rect 573 371 589 405
rect 623 371 639 405
rect 779 410 815 448
rect 779 394 912 410
rect 779 380 862 394
rect 573 338 639 371
rect 846 360 862 380
rect 896 360 912 394
rect 846 344 912 360
rect 573 337 798 338
rect 573 303 589 337
rect 623 322 798 337
rect 623 303 748 322
rect 573 288 748 303
rect 782 288 798 322
rect 573 287 798 288
rect 368 260 512 276
rect 282 222 312 244
rect 368 222 398 260
rect 482 239 512 260
rect 718 272 798 287
rect 83 202 161 218
rect 84 164 114 202
rect 84 54 114 80
rect 482 209 596 239
rect 566 165 596 209
rect 718 165 748 272
rect 882 253 912 344
rect 960 344 996 448
rect 1062 391 1098 448
rect 1062 375 1139 391
rect 960 314 1020 344
rect 1062 341 1089 375
rect 1123 341 1139 375
rect 1487 493 1517 508
rect 1571 493 1601 508
rect 1661 493 1691 508
rect 1880 493 1910 508
rect 1484 470 1520 493
rect 1446 454 1520 470
rect 1446 420 1462 454
rect 1496 440 1520 454
rect 1496 420 1512 440
rect 1446 404 1512 420
rect 1568 383 1604 493
rect 1658 461 1694 493
rect 1658 431 1698 461
rect 1877 444 1913 493
rect 1325 362 1355 377
rect 1554 367 1620 383
rect 1062 325 1139 341
rect 1224 326 1254 341
rect 1322 332 1462 362
rect 1554 347 1570 367
rect 990 277 1020 314
rect 990 261 1061 277
rect 882 237 948 253
rect 882 217 898 237
rect 796 203 898 217
rect 932 203 948 237
rect 990 227 1006 261
rect 1040 227 1061 261
rect 990 211 1061 227
rect 796 187 948 203
rect 796 165 826 187
rect 1031 158 1061 211
rect 1109 158 1139 325
rect 1221 290 1257 326
rect 1187 274 1262 290
rect 1187 240 1203 274
rect 1237 240 1262 274
rect 1187 224 1262 240
rect 1310 274 1376 290
rect 1310 240 1326 274
rect 1360 240 1376 274
rect 1310 224 1376 240
rect 1232 202 1262 224
rect 1330 202 1360 224
rect 282 48 312 74
rect 368 48 398 74
rect 566 55 596 81
rect 718 55 748 81
rect 796 55 826 81
rect 1432 158 1462 332
rect 1510 333 1570 347
rect 1604 333 1620 367
rect 1510 317 1620 333
rect 1510 158 1540 317
rect 1668 311 1698 431
rect 1813 428 1907 444
rect 1813 394 1829 428
rect 1863 394 1907 428
rect 1813 360 1907 394
rect 2183 571 2213 597
rect 2284 592 2314 618
rect 2183 388 2213 403
rect 1813 326 1829 360
rect 1863 326 1907 360
rect 1981 353 2011 368
rect 2170 358 2216 388
rect 1813 322 1907 326
rect 1978 322 2014 353
rect 2170 322 2200 358
rect 2284 353 2314 368
rect 1668 295 1734 311
rect 1668 275 1684 295
rect 1588 261 1684 275
rect 1718 261 1734 295
rect 1588 245 1734 261
rect 1813 292 2200 322
rect 2281 310 2317 353
rect 1813 258 1829 292
rect 1863 258 2200 292
rect 1588 158 1618 245
rect 1813 242 2200 258
rect 2251 294 2317 310
rect 2251 260 2267 294
rect 2301 260 2317 294
rect 2251 244 2317 260
rect 1813 203 1843 242
rect 1972 222 2002 242
rect 1760 173 1843 203
rect 1760 158 1790 173
rect 2170 184 2200 242
rect 2286 222 2316 244
rect 1031 48 1061 74
rect 1109 48 1139 74
rect 1232 48 1262 74
rect 1330 48 1360 74
rect 1432 48 1462 74
rect 1510 48 1540 74
rect 1588 48 1618 74
rect 1760 48 1790 74
rect 1972 48 2002 74
rect 2170 48 2200 74
rect 2286 48 2316 74
<< polycont >>
rect 111 354 145 388
rect 111 286 145 320
rect 111 218 145 252
rect 276 260 310 294
rect 421 276 455 310
rect 589 371 623 405
rect 862 360 896 394
rect 589 303 623 337
rect 748 288 782 322
rect 1089 341 1123 375
rect 1462 420 1496 454
rect 898 203 932 237
rect 1006 227 1040 261
rect 1203 240 1237 274
rect 1326 240 1360 274
rect 1570 333 1604 367
rect 1829 394 1863 428
rect 1829 326 1863 360
rect 1684 261 1718 295
rect 1829 258 1863 292
rect 2267 260 2301 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2400 683
rect 23 567 73 596
rect 23 533 39 567
rect 23 472 73 533
rect 113 568 179 649
rect 113 534 129 568
rect 163 534 179 568
rect 113 518 179 534
rect 315 556 381 649
rect 315 522 331 556
rect 365 522 381 556
rect 315 506 381 522
rect 421 581 775 615
rect 421 530 471 581
rect 455 496 471 530
rect 421 480 471 496
rect 505 520 601 547
rect 505 486 551 520
rect 585 486 601 520
rect 23 446 359 472
rect 505 459 601 486
rect 635 520 707 547
rect 635 486 651 520
rect 685 486 707 520
rect 635 459 707 486
rect 505 446 539 459
rect 23 438 539 446
rect 23 168 57 438
rect 325 412 539 438
rect 95 388 161 404
rect 95 354 111 388
rect 145 354 161 388
rect 95 320 161 354
rect 95 286 111 320
rect 145 286 161 320
rect 95 252 161 286
rect 95 218 111 252
rect 145 218 161 252
rect 95 202 161 218
rect 195 370 241 404
rect 275 378 291 404
rect 275 370 471 378
rect 195 344 471 370
rect 195 202 229 344
rect 405 310 471 344
rect 263 294 359 310
rect 263 260 276 294
rect 310 260 359 294
rect 405 276 421 310
rect 455 276 471 310
rect 405 260 471 276
rect 263 236 359 260
rect 409 210 459 226
rect 195 197 287 202
rect 23 139 73 168
rect 23 105 39 139
rect 23 76 73 105
rect 109 139 159 168
rect 109 105 125 139
rect 109 17 159 105
rect 195 163 237 197
rect 271 163 287 197
rect 195 120 287 163
rect 195 86 237 120
rect 271 86 287 120
rect 195 70 287 86
rect 321 186 373 202
rect 321 152 323 186
rect 357 152 373 186
rect 321 118 373 152
rect 321 84 323 118
rect 357 84 373 118
rect 321 17 373 84
rect 443 176 459 210
rect 409 120 459 176
rect 443 86 459 120
rect 505 169 539 412
rect 573 405 639 421
rect 573 371 589 405
rect 623 371 639 405
rect 573 337 639 371
rect 573 303 589 337
rect 623 303 639 337
rect 573 287 639 303
rect 505 153 571 169
rect 505 119 521 153
rect 555 119 571 153
rect 409 85 459 86
rect 605 85 639 287
rect 409 51 639 85
rect 673 211 707 459
rect 741 467 775 581
rect 809 535 888 649
rect 809 501 831 535
rect 865 501 888 535
rect 922 581 1108 615
rect 922 467 956 581
rect 741 433 956 467
rect 990 520 1040 547
rect 990 486 1006 520
rect 741 322 789 433
rect 990 399 1040 486
rect 1074 459 1108 581
rect 1142 543 1210 649
rect 1142 509 1151 543
rect 1185 509 1210 543
rect 1142 493 1210 509
rect 1352 565 1490 581
rect 1352 531 1368 565
rect 1402 531 1440 565
rect 1474 531 1490 565
rect 1352 530 1490 531
rect 1614 580 1648 649
rect 1614 530 1648 546
rect 1688 567 1754 596
rect 1688 533 1704 567
rect 1738 533 1754 567
rect 1352 496 1580 530
rect 1688 496 1754 533
rect 1352 469 1402 496
rect 1074 425 1207 459
rect 846 394 1040 399
rect 846 360 862 394
rect 896 360 1040 394
rect 846 355 1040 360
rect 1081 375 1139 391
rect 741 288 748 322
rect 782 288 789 322
rect 1081 350 1089 375
rect 741 272 789 288
rect 823 287 1047 321
rect 1081 316 1087 350
rect 1123 341 1139 375
rect 1121 316 1139 341
rect 1173 358 1207 425
rect 1352 435 1368 469
rect 1352 392 1402 435
rect 1446 454 1512 462
rect 1446 420 1462 454
rect 1496 420 1512 454
rect 1446 404 1512 420
rect 1546 444 1754 496
rect 1800 567 1866 596
rect 1800 533 1816 567
rect 1850 533 1866 567
rect 1912 580 1982 649
rect 1912 546 1930 580
rect 1964 546 1982 580
rect 2024 580 2087 596
rect 2058 546 2087 580
rect 1800 512 1866 533
rect 1800 478 1947 512
rect 1546 428 1879 444
rect 1546 410 1829 428
rect 1368 370 1402 392
rect 1173 324 1321 358
rect 1368 336 1444 370
rect 1081 310 1139 316
rect 1287 290 1321 324
rect 823 211 857 287
rect 990 261 1047 287
rect 673 177 857 211
rect 891 237 955 253
rect 891 203 898 237
rect 932 203 955 237
rect 990 227 1006 261
rect 1040 258 1047 261
rect 1187 274 1253 290
rect 1187 258 1203 274
rect 1040 240 1203 258
rect 1237 240 1253 274
rect 1040 227 1253 240
rect 990 224 1253 227
rect 1287 274 1376 290
rect 1287 240 1326 274
rect 1360 240 1376 274
rect 1287 224 1376 240
rect 990 211 1047 224
rect 891 177 955 203
rect 1171 189 1237 190
rect 673 140 723 177
rect 707 106 723 140
rect 673 77 723 106
rect 821 127 887 143
rect 821 93 837 127
rect 871 93 887 127
rect 821 17 887 93
rect 921 137 1036 177
rect 921 103 986 137
rect 1020 103 1036 137
rect 921 87 1036 103
rect 1171 155 1187 189
rect 1221 155 1237 189
rect 1171 116 1237 155
rect 1171 82 1187 116
rect 1221 82 1237 116
rect 1171 17 1237 82
rect 1287 85 1321 224
rect 1410 185 1444 336
rect 1355 169 1444 185
rect 1355 135 1371 169
rect 1405 135 1444 169
rect 1355 119 1444 135
rect 1478 85 1512 404
rect 1813 394 1829 410
rect 1863 394 1879 428
rect 1554 367 1620 376
rect 1554 333 1570 367
rect 1604 333 1620 367
rect 1813 360 1879 394
rect 1554 202 1620 333
rect 1657 350 1734 356
rect 1657 316 1663 350
rect 1697 316 1734 350
rect 1657 295 1734 316
rect 1657 261 1684 295
rect 1718 261 1734 295
rect 1657 236 1734 261
rect 1813 326 1829 360
rect 1863 326 1879 360
rect 1813 292 1879 326
rect 1813 258 1829 292
rect 1863 258 1879 292
rect 1813 242 1879 258
rect 1913 202 1947 478
rect 2024 497 2087 546
rect 2058 463 2087 497
rect 2024 414 2087 463
rect 2058 380 2087 414
rect 2024 236 2087 380
rect 2136 559 2170 575
rect 2136 449 2170 525
rect 2136 310 2170 415
rect 2210 559 2276 649
rect 2210 525 2226 559
rect 2260 525 2276 559
rect 2210 449 2276 525
rect 2210 415 2226 449
rect 2260 415 2276 449
rect 2210 399 2276 415
rect 2311 580 2377 596
rect 2311 546 2327 580
rect 2361 546 2377 580
rect 2311 497 2377 546
rect 2311 463 2327 497
rect 2361 463 2377 497
rect 2311 414 2377 463
rect 2311 380 2327 414
rect 2361 380 2377 414
rect 2311 364 2377 380
rect 2136 294 2308 310
rect 2136 260 2267 294
rect 2301 260 2308 294
rect 2136 244 2308 260
rect 2024 226 2063 236
rect 1554 168 1947 202
rect 1997 210 2063 226
rect 1997 176 2013 210
rect 2047 176 2063 210
rect 2136 188 2175 244
rect 2343 210 2377 364
rect 2311 194 2377 210
rect 1287 51 1512 85
rect 1613 128 1751 134
rect 1613 94 1629 128
rect 1663 94 1701 128
rect 1735 94 1751 128
rect 1613 17 1751 94
rect 1785 133 1851 168
rect 1785 99 1801 133
rect 1835 99 1851 133
rect 1785 83 1851 99
rect 1897 127 1963 134
rect 1897 93 1913 127
rect 1947 93 1963 127
rect 1897 17 1963 93
rect 1997 120 2063 176
rect 1997 86 2013 120
rect 2047 86 2063 120
rect 1997 70 2063 86
rect 2109 146 2175 188
rect 2109 112 2125 146
rect 2159 112 2175 146
rect 2109 70 2175 112
rect 2211 184 2277 188
rect 2211 150 2227 184
rect 2261 150 2277 184
rect 2211 116 2277 150
rect 2211 82 2227 116
rect 2261 82 2277 116
rect 2211 17 2277 82
rect 2311 160 2327 194
rect 2361 160 2377 194
rect 2311 120 2377 160
rect 2311 86 2327 120
rect 2361 86 2377 120
rect 2311 70 2377 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2400 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 1087 341 1089 350
rect 1089 341 1121 350
rect 1087 316 1121 341
rect 1663 316 1697 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
<< metal1 >>
rect 0 683 2400 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2400 683
rect 0 617 2400 649
rect 1075 350 1133 356
rect 1075 316 1087 350
rect 1121 347 1133 350
rect 1651 350 1709 356
rect 1651 347 1663 350
rect 1121 319 1663 347
rect 1121 316 1133 319
rect 1075 310 1133 316
rect 1651 316 1663 319
rect 1697 316 1709 350
rect 1651 310 1709 316
rect 0 17 2400 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2400 17
rect 0 -49 2400 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dfsbp_1
flabel comment s 898 276 898 276 0 FreeSans 200 0 0 0 no_jumper_check
flabel comment s 657 309 657 309 0 FreeSans 200 0 0 0 no_jumper_check
flabel pwell s 0 0 2400 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 2400 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 1663 316 1697 350 0 FreeSans 340 0 0 0 SET_B
port 3 nsew
flabel metal1 s 0 617 2400 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 2400 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 2335 390 2369 424 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 2335 464 2369 498 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 2335 538 2369 572 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 2047 242 2081 276 0 FreeSans 340 0 0 0 Q_N
port 9 nsew
flabel corelocali s 2047 316 2081 350 0 FreeSans 340 0 0 0 Q_N
port 9 nsew
flabel corelocali s 2047 390 2081 424 0 FreeSans 340 0 0 0 Q_N
port 9 nsew
flabel corelocali s 2047 464 2081 498 0 FreeSans 340 0 0 0 Q_N
port 9 nsew
flabel corelocali s 2047 538 2081 572 0 FreeSans 340 0 0 0 Q_N
port 9 nsew
flabel corelocali s 127 242 161 276 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 319 242 353 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 2400 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2787538
string GDS_START 2769364
<< end >>
