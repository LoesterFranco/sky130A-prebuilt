magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 368 561
rect 19 337 74 491
rect 208 439 247 527
rect 19 299 136 337
rect 19 135 67 265
rect 101 165 136 299
rect 170 199 253 265
rect 289 199 348 265
rect 101 129 167 165
rect 22 17 88 95
rect 122 53 167 129
rect 207 75 253 199
rect 289 17 349 163
rect 0 -17 368 17
<< obsli1 >>
rect 108 405 174 491
rect 283 405 349 491
rect 108 371 349 405
rect 170 305 349 371
<< metal1 >>
rect 0 496 368 592
rect 0 -48 368 48
<< labels >>
rlabel locali s 207 75 253 199 6 A1
port 1 nsew signal input
rlabel locali s 170 199 253 265 6 A1
port 1 nsew signal input
rlabel locali s 289 199 348 265 6 A2
port 2 nsew signal input
rlabel locali s 19 135 67 265 6 B1
port 3 nsew signal input
rlabel locali s 122 53 167 129 6 Y
port 4 nsew signal output
rlabel locali s 101 165 136 299 6 Y
port 4 nsew signal output
rlabel locali s 101 129 167 165 6 Y
port 4 nsew signal output
rlabel locali s 19 337 74 491 6 Y
port 4 nsew signal output
rlabel locali s 19 299 136 337 6 Y
port 4 nsew signal output
rlabel locali s 289 17 349 163 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 22 17 88 95 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 368 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 368 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 208 439 247 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 368 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 368 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 368 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 4020762
string GDS_START 4016092
<< end >>
