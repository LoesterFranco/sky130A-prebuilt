magic
tech sky130A
magscale 1 2
timestamp 1604502697
<< nwell >>
rect -38 261 406 582
<< pwell >>
rect 233 -17 267 17
<< scnmos >>
rect 89 47 119 151
rect 249 47 279 151
<< pmoshvt >>
rect 81 339 117 497
rect 251 339 287 497
<< ndiff >>
rect 27 123 89 151
rect 27 89 35 123
rect 69 89 89 123
rect 27 47 89 89
rect 119 93 249 151
rect 119 59 131 93
rect 165 59 199 93
rect 233 59 249 93
rect 119 47 249 59
rect 279 106 333 151
rect 279 72 291 106
rect 325 72 333 106
rect 279 47 333 72
<< pdiff >>
rect 27 477 81 497
rect 27 443 35 477
rect 69 443 81 477
rect 27 396 81 443
rect 27 362 35 396
rect 69 362 81 396
rect 27 339 81 362
rect 117 477 251 497
rect 117 375 131 477
rect 233 375 251 477
rect 117 339 251 375
rect 287 477 341 497
rect 287 443 299 477
rect 333 443 341 477
rect 287 409 341 443
rect 287 375 299 409
rect 333 375 341 409
rect 287 339 341 375
<< ndiffc >>
rect 35 89 69 123
rect 131 59 165 93
rect 199 59 233 93
rect 291 72 325 106
<< pdiffc >>
rect 35 443 69 477
rect 35 362 69 396
rect 131 375 233 477
rect 299 443 333 477
rect 299 375 333 409
<< poly >>
rect 81 497 117 523
rect 251 497 287 523
rect 81 324 117 339
rect 251 324 287 339
rect 79 278 119 324
rect 75 262 139 278
rect 75 228 85 262
rect 119 228 139 262
rect 75 212 139 228
rect 249 265 289 324
rect 249 249 343 265
rect 249 215 299 249
rect 333 215 343 249
rect 89 151 119 212
rect 249 199 343 215
rect 249 151 279 199
rect 89 21 119 47
rect 249 21 279 47
<< polycont >>
rect 85 228 119 262
rect 299 215 333 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 17 477 71 493
rect 17 443 35 477
rect 69 443 71 477
rect 17 396 71 443
rect 17 362 35 396
rect 69 362 71 396
rect 105 477 255 527
rect 105 375 131 477
rect 233 375 255 477
rect 299 477 333 493
rect 299 409 333 443
rect 17 312 71 362
rect 299 341 333 375
rect 17 152 51 312
rect 108 307 333 341
rect 108 278 152 307
rect 85 262 152 278
rect 119 228 152 262
rect 85 212 152 228
rect 108 161 152 212
rect 273 249 349 271
rect 273 215 299 249
rect 333 215 349 249
rect 273 197 349 215
rect 17 123 69 152
rect 108 127 325 161
rect 17 89 35 123
rect 291 106 325 127
rect 17 51 69 89
rect 105 59 131 93
rect 165 59 199 93
rect 233 59 255 93
rect 105 17 255 59
rect 291 51 325 72
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
<< metal1 >>
rect 0 561 368 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 0 496 368 527
rect 0 17 368 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
rect 0 -48 368 -17
<< labels >>
flabel metal1 s 230 0 230 0 0 FreeSans 200 180 0 0 VGND
port 2 nsew
flabel metal1 s 230 544 230 544 0 FreeSans 200 180 0 0 VPWR
port 5 nsew
flabel corelocali s 29 85 63 119 0 FreeSans 200 180 0 0 X
port 6 nsew
flabel corelocali s 29 357 63 391 0 FreeSans 200 180 0 0 X
port 6 nsew
flabel corelocali s 29 425 63 459 0 FreeSans 200 180 0 0 X
port 6 nsew
flabel corelocali s 286 221 320 255 0 FreeSans 200 180 0 0 A
port 1 nsew
flabel nbase s 230 544 230 544 0 FreeSans 200 180 0 0 VPB
port 4 nsew
flabel pwell s 230 0 230 0 0 FreeSans 200 180 0 0 VNB
port 3 nsew
rlabel comment s 0 0 0 0 4 clkbuf_1
<< properties >>
string FIXED_BBOX 0 0 368 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1747334
string GDS_START 1743232
<< end >>
