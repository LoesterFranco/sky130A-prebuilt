magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 644 561
rect 115 365 165 527
rect 96 213 184 255
rect 283 179 333 425
rect 555 429 605 527
rect 582 255 625 393
rect 520 213 625 255
rect 17 17 73 179
rect 107 145 341 179
rect 107 51 173 145
rect 207 17 241 111
rect 275 51 341 145
rect 375 17 409 179
rect 555 17 606 169
rect 0 -17 644 17
<< obsli1 >>
rect 17 331 81 493
rect 199 459 425 493
rect 199 331 249 459
rect 17 289 249 331
rect 367 378 425 459
rect 367 289 418 378
rect 479 323 513 492
rect 452 289 513 323
rect 452 249 486 289
rect 375 215 486 249
rect 443 179 486 215
rect 443 145 513 179
rect 479 89 513 145
<< metal1 >>
rect 0 496 644 592
rect 0 -48 644 48
<< labels >>
rlabel locali s 96 213 184 255 6 A
port 1 nsew signal input
rlabel locali s 582 255 625 393 6 B_N
port 2 nsew signal input
rlabel locali s 520 213 625 255 6 B_N
port 2 nsew signal input
rlabel locali s 283 179 333 425 6 Y
port 3 nsew signal output
rlabel locali s 275 51 341 145 6 Y
port 3 nsew signal output
rlabel locali s 107 145 341 179 6 Y
port 3 nsew signal output
rlabel locali s 107 51 173 145 6 Y
port 3 nsew signal output
rlabel locali s 555 17 606 169 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 375 17 409 179 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 207 17 241 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 17 17 73 179 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 644 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 644 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 555 429 605 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 115 365 165 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 644 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 644 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1959814
string GDS_START 1953884
<< end >>
