magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 1357 325 1407 425
rect 1545 325 1595 425
rect 1357 291 1726 325
rect 36 215 405 257
rect 459 215 894 257
rect 939 215 1261 257
rect 1295 215 1609 257
rect 1672 181 1726 291
rect 107 145 1726 181
rect 107 51 183 145
rect 295 51 371 145
rect 483 51 559 145
rect 671 51 747 145
rect 963 51 1039 145
rect 1151 51 1227 145
rect 1339 51 1415 145
rect 1527 51 1603 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 18 325 81 493
rect 125 359 175 527
rect 219 325 269 493
rect 313 359 363 527
rect 407 459 844 493
rect 407 325 457 459
rect 18 291 457 325
rect 501 325 551 425
rect 595 359 645 459
rect 689 325 739 425
rect 783 359 844 459
rect 881 459 1689 493
rect 881 359 937 459
rect 981 325 1031 425
rect 1075 359 1125 459
rect 1169 325 1219 425
rect 1263 359 1313 459
rect 501 291 1219 325
rect 1451 359 1501 459
rect 1639 359 1689 459
rect 18 17 73 181
rect 227 17 261 111
rect 415 17 449 111
rect 603 17 637 111
rect 791 17 929 111
rect 1083 17 1117 111
rect 1271 17 1305 111
rect 1459 17 1493 111
rect 1647 17 1681 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
<< metal1 >>
rect 0 561 1748 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 0 496 1748 527
rect 0 17 1748 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
rect 0 -48 1748 -17
<< labels >>
rlabel locali s 36 215 405 257 6 A
port 1 nsew signal input
rlabel locali s 459 215 894 257 6 B
port 2 nsew signal input
rlabel locali s 939 215 1261 257 6 C
port 3 nsew signal input
rlabel locali s 1295 215 1609 257 6 D
port 4 nsew signal input
rlabel locali s 1672 181 1726 291 6 Y
port 5 nsew signal output
rlabel locali s 1545 325 1595 425 6 Y
port 5 nsew signal output
rlabel locali s 1527 51 1603 145 6 Y
port 5 nsew signal output
rlabel locali s 1357 325 1407 425 6 Y
port 5 nsew signal output
rlabel locali s 1357 291 1726 325 6 Y
port 5 nsew signal output
rlabel locali s 1339 51 1415 145 6 Y
port 5 nsew signal output
rlabel locali s 1151 51 1227 145 6 Y
port 5 nsew signal output
rlabel locali s 963 51 1039 145 6 Y
port 5 nsew signal output
rlabel locali s 671 51 747 145 6 Y
port 5 nsew signal output
rlabel locali s 483 51 559 145 6 Y
port 5 nsew signal output
rlabel locali s 295 51 371 145 6 Y
port 5 nsew signal output
rlabel locali s 107 145 1726 181 6 Y
port 5 nsew signal output
rlabel locali s 107 51 183 145 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -48 1748 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 1748 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1748 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2500888
string GDS_START 2487770
<< end >>
