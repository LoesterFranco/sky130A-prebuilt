magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 90 243 164 356
rect 198 243 264 356
rect 600 243 666 430
rect 700 243 774 430
rect 1170 289 1236 356
rect 1844 512 1897 578
rect 1641 270 1707 356
rect 1849 236 1897 512
rect 1816 80 1897 236
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 22 390 111 576
rect 145 390 211 649
rect 406 501 510 545
rect 653 535 719 649
rect 759 581 1110 615
rect 759 501 804 581
rect 406 467 804 501
rect 22 206 56 390
rect 406 337 510 467
rect 861 433 1033 547
rect 1070 501 1110 581
rect 1146 535 1212 649
rect 1258 501 1324 596
rect 1070 467 1324 501
rect 306 240 372 306
rect 306 206 340 240
rect 406 206 440 337
rect 22 172 340 206
rect 22 70 89 172
rect 140 17 218 136
rect 306 85 340 172
rect 375 119 440 206
rect 492 209 558 290
rect 861 399 1136 433
rect 816 209 882 290
rect 916 289 1068 355
rect 916 209 950 289
rect 1102 255 1136 399
rect 1258 390 1324 467
rect 1358 581 1704 615
rect 492 175 950 209
rect 984 221 1247 255
rect 492 85 526 175
rect 984 141 1018 221
rect 306 51 526 85
rect 625 17 743 136
rect 842 75 1018 141
rect 1052 17 1118 187
rect 1197 89 1247 221
rect 1281 157 1315 390
rect 1358 257 1424 581
rect 1349 223 1424 257
rect 1458 389 1524 547
rect 1570 390 1636 547
rect 1670 424 1704 581
rect 1738 458 1804 649
rect 1670 390 1783 424
rect 1458 255 1492 389
rect 1570 355 1607 390
rect 1526 289 1607 355
rect 1349 191 1385 223
rect 1458 221 1539 255
rect 1421 157 1471 187
rect 1281 123 1471 157
rect 1421 121 1471 123
rect 1197 87 1297 89
rect 1505 87 1539 221
rect 1573 236 1607 289
rect 1749 336 1783 390
rect 1749 270 1815 336
rect 1573 100 1682 236
rect 1197 53 1539 87
rect 1716 17 1782 236
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
<< metal1 >>
rect 0 683 1920 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 0 617 1920 649
rect 0 17 1920 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
rect 0 -49 1920 -17
<< labels >>
rlabel locali s 198 243 264 356 6 A0
port 1 nsew signal input
rlabel locali s 600 243 666 430 6 A1
port 2 nsew signal input
rlabel locali s 700 243 774 430 6 A2
port 3 nsew signal input
rlabel locali s 1170 289 1236 356 6 A3
port 4 nsew signal input
rlabel locali s 90 243 164 356 6 S0
port 5 nsew signal input
rlabel locali s 1641 270 1707 356 6 S1
port 6 nsew signal input
rlabel locali s 1849 236 1897 512 6 X
port 7 nsew signal output
rlabel locali s 1844 512 1897 578 6 X
port 7 nsew signal output
rlabel locali s 1816 80 1897 236 6 X
port 7 nsew signal output
rlabel metal1 s 0 -49 1920 49 8 VGND
port 8 nsew ground bidirectional
rlabel metal1 s 0 617 1920 715 6 VPWR
port 9 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1920 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1990768
string GDS_START 1976338
<< end >>
