magic
tech sky130A
magscale 1 2
timestamp 1601050047
<< nwell >>
rect -38 332 2918 704
rect 1624 311 1956 332
<< pwell >>
rect 0 0 2880 49
<< scpmos >>
rect 86 464 116 592
rect 310 464 340 592
rect 394 464 424 592
rect 484 464 514 592
rect 592 464 622 592
rect 706 464 736 592
rect 914 368 944 592
rect 1004 368 1034 592
rect 1212 457 1242 541
rect 1302 457 1332 541
rect 1386 457 1416 541
rect 1511 457 1541 541
rect 1713 347 1743 547
rect 1837 366 1867 566
rect 2007 508 2037 592
rect 2085 508 2115 592
rect 2255 508 2285 592
rect 2345 508 2375 592
rect 2462 392 2492 592
rect 2664 368 2694 592
rect 2754 368 2784 592
<< nmoslvt >>
rect 84 74 114 158
rect 282 81 312 165
rect 360 81 390 165
rect 517 81 547 165
rect 595 81 625 165
rect 704 81 734 165
rect 923 74 953 222
rect 1023 74 1053 222
rect 1224 138 1254 222
rect 1324 138 1354 222
rect 1402 138 1432 222
rect 1480 138 1510 222
rect 1693 74 1723 222
rect 1794 74 1824 222
rect 2048 74 2078 158
rect 2126 74 2156 158
rect 2212 74 2242 158
rect 2284 74 2314 158
rect 2482 74 2512 202
rect 2680 74 2710 222
rect 2766 74 2796 222
<< ndiff >>
rect 866 202 923 222
rect 866 168 878 202
rect 912 168 923 202
rect 27 133 84 158
rect 27 99 39 133
rect 73 99 84 133
rect 27 74 84 99
rect 114 128 171 158
rect 114 94 125 128
rect 159 94 171 128
rect 114 74 171 94
rect 225 127 282 165
rect 225 93 237 127
rect 271 93 282 127
rect 225 81 282 93
rect 312 81 360 165
rect 390 153 517 165
rect 390 119 471 153
rect 505 119 517 153
rect 390 81 517 119
rect 547 81 595 165
rect 625 140 704 165
rect 625 106 659 140
rect 693 106 704 140
rect 625 81 704 106
rect 734 140 805 165
rect 734 106 759 140
rect 793 106 805 140
rect 734 81 805 106
rect 866 120 923 168
rect 866 86 878 120
rect 912 86 923 120
rect 866 74 923 86
rect 953 127 1023 222
rect 953 93 964 127
rect 998 93 1023 127
rect 953 74 1023 93
rect 1053 209 1110 222
rect 1053 175 1064 209
rect 1098 175 1110 209
rect 1053 120 1110 175
rect 1167 197 1224 222
rect 1167 163 1179 197
rect 1213 163 1224 197
rect 1167 138 1224 163
rect 1254 196 1324 222
rect 1254 162 1279 196
rect 1313 162 1324 196
rect 1254 138 1324 162
rect 1354 138 1402 222
rect 1432 138 1480 222
rect 1510 138 1693 222
rect 1053 86 1064 120
rect 1098 86 1110 120
rect 1053 74 1110 86
rect 1525 82 1693 138
rect 1525 48 1551 82
rect 1585 74 1693 82
rect 1723 189 1794 222
rect 1723 155 1734 189
rect 1768 155 1794 189
rect 1723 74 1794 155
rect 1824 158 1874 222
rect 2623 210 2680 222
rect 1824 146 2048 158
rect 1824 112 1902 146
rect 1936 112 2003 146
rect 2037 112 2048 146
rect 1824 74 2048 112
rect 2078 74 2126 158
rect 2156 133 2212 158
rect 2156 99 2167 133
rect 2201 99 2212 133
rect 2156 74 2212 99
rect 2242 74 2284 158
rect 2314 133 2371 158
rect 2314 99 2325 133
rect 2359 99 2371 133
rect 2314 74 2371 99
rect 2425 120 2482 202
rect 2425 86 2437 120
rect 2471 86 2482 120
rect 2425 74 2482 86
rect 2512 190 2569 202
rect 2512 156 2523 190
rect 2557 156 2569 190
rect 2512 120 2569 156
rect 2512 86 2523 120
rect 2557 86 2569 120
rect 2512 74 2569 86
rect 2623 176 2635 210
rect 2669 176 2680 210
rect 2623 120 2680 176
rect 2623 86 2635 120
rect 2669 86 2680 120
rect 2623 74 2680 86
rect 2710 210 2766 222
rect 2710 176 2721 210
rect 2755 176 2766 210
rect 2710 120 2766 176
rect 2710 86 2721 120
rect 2755 86 2766 120
rect 2710 74 2766 86
rect 2796 210 2853 222
rect 2796 176 2807 210
rect 2841 176 2853 210
rect 2796 120 2853 176
rect 2796 86 2807 120
rect 2841 86 2853 120
rect 2796 74 2853 86
rect 1585 48 1612 74
rect 1525 36 1612 48
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 510 86 546
rect 27 476 39 510
rect 73 476 86 510
rect 27 464 86 476
rect 116 580 310 592
rect 116 546 139 580
rect 173 546 263 580
rect 297 546 310 580
rect 116 510 310 546
rect 116 476 139 510
rect 173 476 263 510
rect 297 476 310 510
rect 116 464 310 476
rect 340 464 394 592
rect 424 580 484 592
rect 424 546 437 580
rect 471 546 484 580
rect 424 510 484 546
rect 424 476 437 510
rect 471 476 484 510
rect 424 464 484 476
rect 514 464 592 592
rect 622 575 706 592
rect 622 541 635 575
rect 669 541 706 575
rect 622 464 706 541
rect 736 580 795 592
rect 736 546 749 580
rect 783 546 795 580
rect 736 510 795 546
rect 736 476 749 510
rect 783 476 795 510
rect 736 464 795 476
rect 855 421 914 592
rect 855 387 867 421
rect 901 387 914 421
rect 855 368 914 387
rect 944 580 1004 592
rect 944 546 957 580
rect 991 546 1004 580
rect 944 368 1004 546
rect 1034 429 1093 592
rect 1034 395 1047 429
rect 1081 395 1093 429
rect 1034 368 1093 395
rect 1434 582 1493 594
rect 1434 548 1446 582
rect 1480 548 1493 582
rect 1434 541 1493 548
rect 1948 566 2007 592
rect 1761 547 1837 566
rect 1153 516 1212 541
rect 1153 482 1165 516
rect 1199 482 1212 516
rect 1153 457 1212 482
rect 1242 529 1302 541
rect 1242 495 1255 529
rect 1289 495 1302 529
rect 1242 457 1302 495
rect 1332 457 1386 541
rect 1416 457 1511 541
rect 1541 521 1600 541
rect 1541 487 1554 521
rect 1588 487 1600 521
rect 1541 457 1600 487
rect 1654 524 1713 547
rect 1654 490 1666 524
rect 1700 490 1713 524
rect 1654 468 1713 490
rect 1660 347 1713 468
rect 1743 535 1837 547
rect 1743 501 1773 535
rect 1807 501 1837 535
rect 1743 464 1837 501
rect 1743 430 1773 464
rect 1807 430 1837 464
rect 1743 393 1837 430
rect 1743 359 1773 393
rect 1807 366 1837 393
rect 1867 554 2007 566
rect 1867 520 1880 554
rect 1914 520 1960 554
rect 1994 520 2007 554
rect 1867 508 2007 520
rect 2037 508 2085 592
rect 2115 580 2255 592
rect 2115 546 2128 580
rect 2162 546 2198 580
rect 2232 546 2255 580
rect 2115 508 2255 546
rect 2285 567 2345 592
rect 2285 533 2298 567
rect 2332 533 2345 567
rect 2285 508 2345 533
rect 2375 580 2462 592
rect 2375 546 2405 580
rect 2439 546 2462 580
rect 2375 509 2462 546
rect 2375 508 2405 509
rect 1867 486 1925 508
rect 1867 452 1880 486
rect 1914 452 1925 486
rect 1867 418 1925 452
rect 1867 384 1880 418
rect 1914 384 1925 418
rect 1867 366 1925 384
rect 1807 359 1819 366
rect 1743 347 1819 359
rect 2393 475 2405 508
rect 2439 475 2462 509
rect 2393 438 2462 475
rect 2393 404 2405 438
rect 2439 404 2462 438
rect 2393 392 2462 404
rect 2492 580 2551 592
rect 2492 546 2505 580
rect 2539 546 2551 580
rect 2492 509 2551 546
rect 2492 475 2505 509
rect 2539 475 2551 509
rect 2492 438 2551 475
rect 2492 404 2505 438
rect 2539 404 2551 438
rect 2492 392 2551 404
rect 2605 580 2664 592
rect 2605 546 2617 580
rect 2651 546 2664 580
rect 2605 497 2664 546
rect 2605 463 2617 497
rect 2651 463 2664 497
rect 2605 414 2664 463
rect 2605 380 2617 414
rect 2651 380 2664 414
rect 2605 368 2664 380
rect 2694 580 2754 592
rect 2694 546 2707 580
rect 2741 546 2754 580
rect 2694 497 2754 546
rect 2694 463 2707 497
rect 2741 463 2754 497
rect 2694 414 2754 463
rect 2694 380 2707 414
rect 2741 380 2754 414
rect 2694 368 2754 380
rect 2784 580 2853 592
rect 2784 546 2807 580
rect 2841 546 2853 580
rect 2784 497 2853 546
rect 2784 463 2807 497
rect 2841 463 2853 497
rect 2784 414 2853 463
rect 2784 380 2807 414
rect 2841 380 2853 414
rect 2784 368 2853 380
<< ndiffc >>
rect 878 168 912 202
rect 39 99 73 133
rect 125 94 159 128
rect 237 93 271 127
rect 471 119 505 153
rect 659 106 693 140
rect 759 106 793 140
rect 878 86 912 120
rect 964 93 998 127
rect 1064 175 1098 209
rect 1179 163 1213 197
rect 1279 162 1313 196
rect 1064 86 1098 120
rect 1551 48 1585 82
rect 1734 155 1768 189
rect 1902 112 1936 146
rect 2003 112 2037 146
rect 2167 99 2201 133
rect 2325 99 2359 133
rect 2437 86 2471 120
rect 2523 156 2557 190
rect 2523 86 2557 120
rect 2635 176 2669 210
rect 2635 86 2669 120
rect 2721 176 2755 210
rect 2721 86 2755 120
rect 2807 176 2841 210
rect 2807 86 2841 120
<< pdiffc >>
rect 39 546 73 580
rect 39 476 73 510
rect 139 546 173 580
rect 263 546 297 580
rect 139 476 173 510
rect 263 476 297 510
rect 437 546 471 580
rect 437 476 471 510
rect 635 541 669 575
rect 749 546 783 580
rect 749 476 783 510
rect 867 387 901 421
rect 957 546 991 580
rect 1047 395 1081 429
rect 1446 548 1480 582
rect 1165 482 1199 516
rect 1255 495 1289 529
rect 1554 487 1588 521
rect 1666 490 1700 524
rect 1773 501 1807 535
rect 1773 430 1807 464
rect 1773 359 1807 393
rect 1880 520 1914 554
rect 1960 520 1994 554
rect 2128 546 2162 580
rect 2198 546 2232 580
rect 2298 533 2332 567
rect 2405 546 2439 580
rect 1880 452 1914 486
rect 1880 384 1914 418
rect 2405 475 2439 509
rect 2405 404 2439 438
rect 2505 546 2539 580
rect 2505 475 2539 509
rect 2505 404 2539 438
rect 2617 546 2651 580
rect 2617 463 2651 497
rect 2617 380 2651 414
rect 2707 546 2741 580
rect 2707 463 2741 497
rect 2707 380 2741 414
rect 2807 546 2841 580
rect 2807 463 2841 497
rect 2807 380 2841 414
<< poly >>
rect 86 592 116 618
rect 310 592 340 618
rect 394 592 424 618
rect 484 592 514 618
rect 592 592 622 618
rect 706 592 736 618
rect 914 592 944 618
rect 1004 592 1034 618
rect 1108 615 1870 645
rect 86 449 116 464
rect 310 449 340 464
rect 394 449 424 464
rect 484 449 514 464
rect 592 449 622 464
rect 706 449 736 464
rect 83 367 119 449
rect 307 367 343 449
rect 83 351 343 367
rect 83 317 137 351
rect 171 317 205 351
rect 239 317 273 351
rect 307 317 343 351
rect 83 301 343 317
rect 84 158 114 301
rect 391 253 427 449
rect 481 432 517 449
rect 475 416 541 432
rect 475 382 491 416
rect 525 382 541 416
rect 475 366 541 382
rect 589 430 625 449
rect 703 432 739 449
rect 589 414 655 430
rect 589 380 605 414
rect 639 380 655 414
rect 589 346 655 380
rect 703 416 823 432
rect 703 382 773 416
rect 807 382 823 416
rect 703 366 823 382
rect 162 237 228 253
rect 162 203 178 237
rect 212 217 228 237
rect 354 237 427 253
rect 475 302 547 318
rect 475 268 491 302
rect 525 268 547 302
rect 589 312 605 346
rect 639 312 655 346
rect 589 296 655 312
rect 475 252 547 268
rect 212 203 312 217
rect 162 187 312 203
rect 354 203 370 237
rect 404 203 427 237
rect 354 187 427 203
rect 282 165 312 187
rect 360 165 390 187
rect 517 165 547 252
rect 595 165 625 296
rect 704 165 734 366
rect 914 353 944 368
rect 1004 353 1034 368
rect 911 318 947 353
rect 1001 325 1037 353
rect 795 302 953 318
rect 795 268 811 302
rect 845 268 879 302
rect 913 268 953 302
rect 795 252 953 268
rect 923 222 953 252
rect 995 309 1061 325
rect 995 275 1011 309
rect 1045 279 1061 309
rect 1108 279 1138 615
rect 1212 541 1242 567
rect 1299 556 1335 615
rect 1302 541 1332 556
rect 1386 541 1416 567
rect 1834 581 1870 615
rect 2007 592 2037 618
rect 2085 592 2115 618
rect 2255 592 2285 618
rect 2345 592 2375 618
rect 2462 592 2492 618
rect 2664 592 2694 618
rect 2754 592 2784 618
rect 1511 541 1541 567
rect 1713 547 1743 573
rect 1837 566 1867 581
rect 1212 442 1242 457
rect 1209 393 1245 442
rect 1302 431 1332 457
rect 1386 442 1416 457
rect 1511 442 1541 457
rect 1383 415 1419 442
rect 1508 425 1544 442
rect 1383 399 1466 415
rect 1180 377 1246 393
rect 1180 343 1196 377
rect 1230 357 1246 377
rect 1383 365 1416 399
rect 1450 365 1466 399
rect 1230 343 1332 357
rect 1383 349 1466 365
rect 1508 409 1628 425
rect 1508 375 1578 409
rect 1612 375 1628 409
rect 1508 359 1628 375
rect 1180 327 1332 343
rect 1302 301 1332 327
rect 1045 275 1254 279
rect 995 249 1254 275
rect 1302 271 1354 301
rect 1023 222 1053 249
rect 1224 222 1254 249
rect 1324 222 1354 271
rect 1402 222 1432 349
rect 1514 267 1544 359
rect 2007 493 2037 508
rect 2085 493 2115 508
rect 2255 493 2285 508
rect 2345 493 2375 508
rect 2004 466 2040 493
rect 1957 450 2040 466
rect 1957 416 1973 450
rect 2007 416 2040 450
rect 2082 476 2118 493
rect 2082 460 2170 476
rect 2082 446 2120 460
rect 1957 400 2040 416
rect 2088 426 2120 446
rect 2154 426 2170 460
rect 2252 447 2288 493
rect 2088 392 2170 426
rect 2222 431 2288 447
rect 2222 411 2238 431
rect 1837 351 1867 366
rect 2088 358 2120 392
rect 2154 358 2170 392
rect 1713 332 1743 347
rect 1834 345 1870 351
rect 1710 315 1746 332
rect 1834 315 2040 345
rect 1480 237 1544 267
rect 1618 299 1746 315
rect 1618 265 1634 299
rect 1668 285 1746 299
rect 1668 265 1723 285
rect 1618 249 1723 265
rect 1480 222 1510 237
rect 1693 222 1723 249
rect 1794 251 1962 267
rect 1794 237 1912 251
rect 1794 222 1824 237
rect 84 48 114 74
rect 282 55 312 81
rect 360 55 390 81
rect 517 55 547 81
rect 595 55 625 81
rect 704 55 734 81
rect 1224 112 1254 138
rect 1324 112 1354 138
rect 1402 112 1432 138
rect 1480 112 1510 138
rect 923 48 953 74
rect 1023 48 1053 74
rect 1896 217 1912 237
rect 1946 217 1962 251
rect 1896 201 1962 217
rect 2010 226 2040 315
rect 2088 324 2170 358
rect 2088 290 2120 324
rect 2154 290 2170 324
rect 2088 274 2170 290
rect 2212 397 2238 411
rect 2272 397 2288 431
rect 2212 381 2288 397
rect 2010 196 2078 226
rect 2048 158 2078 196
rect 2126 158 2156 274
rect 2212 158 2242 381
rect 2342 333 2378 493
rect 2462 377 2492 392
rect 2348 285 2378 333
rect 2459 285 2495 377
rect 2664 353 2694 368
rect 2754 353 2784 368
rect 2661 326 2697 353
rect 2751 326 2787 353
rect 2312 269 2495 285
rect 2312 249 2328 269
rect 2284 235 2328 249
rect 2362 249 2495 269
rect 2605 310 2787 326
rect 2605 276 2621 310
rect 2655 290 2787 310
rect 2655 276 2796 290
rect 2605 260 2796 276
rect 2362 235 2512 249
rect 2284 219 2512 235
rect 2680 222 2710 260
rect 2766 222 2796 260
rect 2284 158 2314 219
rect 2482 202 2512 219
rect 1693 48 1723 74
rect 1794 48 1824 74
rect 2048 48 2078 74
rect 2126 48 2156 74
rect 2212 48 2242 74
rect 2284 48 2314 74
rect 2482 48 2512 74
rect 2680 48 2710 74
rect 2766 48 2796 74
<< polycont >>
rect 137 317 171 351
rect 205 317 239 351
rect 273 317 307 351
rect 491 382 525 416
rect 605 380 639 414
rect 773 382 807 416
rect 178 203 212 237
rect 491 268 525 302
rect 605 312 639 346
rect 370 203 404 237
rect 811 268 845 302
rect 879 268 913 302
rect 1011 275 1045 309
rect 1196 343 1230 377
rect 1416 365 1450 399
rect 1578 375 1612 409
rect 1973 416 2007 450
rect 2120 426 2154 460
rect 2120 358 2154 392
rect 1634 265 1668 299
rect 1912 217 1946 251
rect 2120 290 2154 324
rect 2238 397 2272 431
rect 2328 235 2362 269
rect 2621 276 2655 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2880 683
rect 23 580 89 596
rect 23 546 39 580
rect 73 546 89 580
rect 23 510 89 546
rect 23 476 39 510
rect 73 476 89 510
rect 23 435 89 476
rect 123 580 313 649
rect 123 546 139 580
rect 173 546 263 580
rect 297 546 313 580
rect 123 510 313 546
rect 123 476 139 510
rect 173 476 263 510
rect 297 476 313 510
rect 123 469 313 476
rect 421 580 487 596
rect 421 546 437 580
rect 471 546 487 580
rect 421 510 487 546
rect 619 575 685 649
rect 619 541 635 575
rect 669 541 685 575
rect 619 537 685 541
rect 723 580 799 596
rect 723 546 749 580
rect 783 546 799 580
rect 941 580 1007 649
rect 941 546 957 580
rect 991 546 1007 580
rect 1430 582 1497 649
rect 1430 548 1446 582
rect 1480 548 1497 582
rect 421 476 437 510
rect 471 503 487 510
rect 723 512 799 546
rect 1149 516 1199 545
rect 1149 512 1165 516
rect 723 510 1165 512
rect 723 503 749 510
rect 471 476 749 503
rect 783 482 1165 510
rect 1239 529 1374 545
rect 1430 532 1497 548
rect 1239 495 1255 529
rect 1289 498 1374 529
rect 1538 521 1604 545
rect 1538 498 1554 521
rect 1289 495 1554 498
rect 783 478 1199 482
rect 783 476 799 478
rect 421 469 799 476
rect 689 466 799 469
rect 23 416 541 435
rect 23 401 491 416
rect 23 253 57 401
rect 475 382 491 401
rect 525 382 541 416
rect 121 351 359 367
rect 475 366 541 382
rect 589 414 655 430
rect 589 380 605 414
rect 639 380 655 414
rect 121 317 137 351
rect 171 317 205 351
rect 239 317 273 351
rect 307 332 359 351
rect 589 346 655 380
rect 307 317 541 332
rect 121 302 541 317
rect 121 298 491 302
rect 475 268 491 298
rect 525 268 541 302
rect 589 312 605 346
rect 639 312 655 346
rect 589 296 655 312
rect 23 237 228 253
rect 23 203 178 237
rect 212 203 228 237
rect 23 187 228 203
rect 313 237 420 253
rect 475 252 541 268
rect 689 262 723 466
rect 1149 461 1199 478
rect 1340 487 1554 495
rect 1588 487 1604 521
rect 1340 464 1604 487
rect 1650 524 1716 649
rect 2112 580 2248 649
rect 1864 554 2078 570
rect 1650 490 1666 524
rect 1700 490 1716 524
rect 1650 464 1716 490
rect 1750 535 1823 551
rect 1750 501 1773 535
rect 1807 501 1823 535
rect 1750 464 1823 501
rect 757 424 833 432
rect 757 416 799 424
rect 757 382 773 416
rect 807 382 833 390
rect 757 366 833 382
rect 867 421 917 444
rect 901 398 917 421
rect 1031 429 1097 444
rect 901 387 997 398
rect 867 364 997 387
rect 963 325 997 364
rect 1031 395 1047 429
rect 1081 395 1097 429
rect 1149 427 1306 461
rect 1031 393 1097 395
rect 1031 377 1238 393
rect 1031 359 1196 377
rect 1095 343 1196 359
rect 1230 343 1238 377
rect 1095 327 1238 343
rect 313 203 370 237
rect 404 203 420 237
rect 23 133 73 187
rect 313 162 420 203
rect 575 228 723 262
rect 793 302 929 318
rect 793 268 811 302
rect 845 268 879 302
rect 913 268 929 302
rect 793 252 929 268
rect 963 309 1061 325
rect 963 275 1011 309
rect 1045 275 1061 309
rect 963 259 1061 275
rect 793 236 839 252
rect 575 169 609 228
rect 963 218 997 259
rect 1095 225 1129 327
rect 1272 293 1306 427
rect 878 202 997 218
rect 454 153 609 169
rect 23 99 39 133
rect 23 70 73 99
rect 109 128 175 153
rect 109 94 125 128
rect 159 94 175 128
rect 109 17 175 94
rect 221 127 287 128
rect 221 93 237 127
rect 271 93 287 127
rect 454 119 471 153
rect 505 119 609 153
rect 643 140 709 169
rect 221 85 287 93
rect 643 106 659 140
rect 693 106 709 140
rect 643 85 709 106
rect 221 51 709 85
rect 743 140 809 169
rect 743 106 759 140
rect 793 106 809 140
rect 743 17 809 106
rect 912 184 997 202
rect 1048 209 1129 225
rect 878 120 912 168
rect 1048 175 1064 209
rect 1098 175 1129 209
rect 878 70 912 86
rect 948 127 1014 150
rect 948 93 964 127
rect 998 93 1014 127
rect 948 17 1014 93
rect 1048 120 1129 175
rect 1163 259 1306 293
rect 1163 197 1229 259
rect 1340 225 1374 464
rect 1163 163 1179 197
rect 1213 163 1229 197
rect 1163 134 1229 163
rect 1263 196 1374 225
rect 1263 162 1279 196
rect 1313 191 1374 196
rect 1408 399 1463 415
rect 1408 365 1416 399
rect 1450 365 1463 399
rect 1408 218 1463 365
rect 1497 315 1531 464
rect 1750 430 1773 464
rect 1807 430 1823 464
rect 1565 424 1703 430
rect 1565 409 1663 424
rect 1565 375 1578 409
rect 1612 390 1663 409
rect 1697 390 1703 424
rect 1612 375 1703 390
rect 1565 359 1703 375
rect 1750 393 1823 430
rect 1750 359 1773 393
rect 1807 359 1823 393
rect 1864 520 1880 554
rect 1914 520 1960 554
rect 1994 520 2078 554
rect 2112 546 2128 580
rect 2162 546 2198 580
rect 2232 546 2248 580
rect 2282 567 2348 596
rect 1864 504 2078 520
rect 2282 533 2298 567
rect 2332 533 2348 567
rect 2282 512 2348 533
rect 1864 486 1920 504
rect 1864 452 1880 486
rect 1914 452 1920 486
rect 1864 418 1920 452
rect 1864 384 1880 418
rect 1914 384 1920 418
rect 1864 368 1920 384
rect 1957 450 2010 466
rect 1957 416 1973 450
rect 2007 416 2010 450
rect 1750 343 1823 359
rect 1497 299 1684 315
rect 1497 265 1634 299
rect 1668 265 1684 299
rect 1497 252 1684 265
rect 1750 226 1784 343
rect 1957 267 2010 416
rect 1718 218 1784 226
rect 1313 162 1329 191
rect 1408 189 1784 218
rect 1408 184 1734 189
rect 1263 134 1329 162
rect 1718 155 1734 184
rect 1768 155 1784 189
rect 1048 86 1064 120
rect 1098 100 1129 120
rect 1408 116 1684 150
rect 1718 119 1784 155
rect 1818 251 2010 267
rect 1818 217 1912 251
rect 1946 217 2010 251
rect 1818 201 2010 217
rect 2044 240 2078 504
rect 2112 478 2348 512
rect 2389 580 2455 649
rect 2389 546 2405 580
rect 2439 546 2455 580
rect 2389 509 2455 546
rect 2112 460 2170 478
rect 2112 426 2120 460
rect 2154 426 2170 460
rect 2389 475 2405 509
rect 2439 475 2455 509
rect 2112 392 2170 426
rect 2112 358 2120 392
rect 2154 358 2170 392
rect 2222 431 2288 444
rect 2222 397 2238 431
rect 2272 424 2288 431
rect 2222 390 2239 397
rect 2273 390 2288 424
rect 2222 384 2288 390
rect 2389 438 2455 475
rect 2389 404 2405 438
rect 2439 404 2455 438
rect 2389 388 2455 404
rect 2489 580 2555 596
rect 2489 546 2505 580
rect 2539 546 2555 580
rect 2489 509 2555 546
rect 2489 475 2505 509
rect 2539 475 2555 509
rect 2489 438 2555 475
rect 2489 404 2505 438
rect 2539 404 2555 438
rect 2489 388 2555 404
rect 2112 350 2170 358
rect 2112 324 2446 350
rect 2112 290 2120 324
rect 2154 316 2446 324
rect 2154 290 2170 316
rect 2112 274 2170 290
rect 2204 269 2378 282
rect 2204 240 2328 269
rect 2044 235 2328 240
rect 2362 235 2378 269
rect 2044 222 2378 235
rect 2044 206 2238 222
rect 1408 100 1442 116
rect 1098 86 1442 100
rect 1048 66 1442 86
rect 1650 85 1684 116
rect 1818 85 1852 201
rect 2044 162 2078 206
rect 2412 188 2446 316
rect 1886 146 2078 162
rect 1886 112 1902 146
rect 1936 112 2003 146
rect 2037 112 2078 146
rect 1886 96 2078 112
rect 2151 133 2217 162
rect 2151 99 2167 133
rect 2201 99 2217 133
rect 1521 48 1551 82
rect 1585 48 1616 82
rect 1650 51 1852 85
rect 1521 17 1616 48
rect 2151 17 2217 99
rect 2309 154 2446 188
rect 2521 326 2555 388
rect 2601 580 2667 649
rect 2601 546 2617 580
rect 2651 546 2667 580
rect 2601 497 2667 546
rect 2601 463 2617 497
rect 2651 463 2667 497
rect 2601 414 2667 463
rect 2601 380 2617 414
rect 2651 380 2667 414
rect 2601 364 2667 380
rect 2705 580 2757 596
rect 2705 546 2707 580
rect 2741 546 2757 580
rect 2705 497 2757 546
rect 2705 463 2707 497
rect 2741 463 2757 497
rect 2705 414 2757 463
rect 2705 380 2707 414
rect 2741 380 2757 414
rect 2521 310 2671 326
rect 2521 276 2621 310
rect 2655 276 2671 310
rect 2521 260 2671 276
rect 2705 282 2757 380
rect 2791 580 2857 649
rect 2791 546 2807 580
rect 2841 546 2857 580
rect 2791 497 2857 546
rect 2791 463 2807 497
rect 2841 463 2857 497
rect 2791 414 2857 463
rect 2791 380 2807 414
rect 2841 380 2857 414
rect 2791 364 2857 380
rect 2521 190 2573 260
rect 2521 156 2523 190
rect 2557 156 2573 190
rect 2309 133 2375 154
rect 2309 99 2325 133
rect 2359 99 2375 133
rect 2521 120 2573 156
rect 2309 70 2375 99
rect 2421 86 2437 120
rect 2471 86 2487 120
rect 2421 17 2487 86
rect 2521 86 2523 120
rect 2557 86 2573 120
rect 2521 70 2573 86
rect 2619 210 2669 226
rect 2619 176 2635 210
rect 2619 120 2669 176
rect 2619 86 2635 120
rect 2619 17 2669 86
rect 2705 210 2771 282
rect 2705 176 2721 210
rect 2755 176 2771 210
rect 2705 120 2771 176
rect 2705 86 2721 120
rect 2755 86 2771 120
rect 2705 70 2771 86
rect 2807 210 2857 226
rect 2841 176 2857 210
rect 2807 120 2857 176
rect 2841 86 2857 120
rect 2807 17 2857 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2880 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 799 416 833 424
rect 799 390 807 416
rect 807 390 833 416
rect 1663 390 1697 424
rect 2239 397 2272 424
rect 2272 397 2273 424
rect 2239 390 2273 397
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
<< metal1 >>
rect 0 683 2880 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2880 683
rect 0 617 2880 649
rect 787 424 845 430
rect 787 390 799 424
rect 833 421 845 424
rect 1651 424 1709 430
rect 1651 421 1663 424
rect 833 393 1663 421
rect 833 390 845 393
rect 787 384 845 390
rect 1651 390 1663 393
rect 1697 421 1709 424
rect 2227 424 2285 430
rect 2227 421 2239 424
rect 1697 393 2239 421
rect 1697 390 1709 393
rect 1651 384 1709 390
rect 2227 390 2239 393
rect 2273 390 2285 424
rect 2227 384 2285 390
rect 0 17 2880 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2880 17
rect 0 -49 2880 -17
<< labels >>
rlabel comment s 0 0 0 0 4 sdfrtp_2
flabel pwell s 0 0 2880 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 0 617 2880 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 2239 390 2273 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew
flabel metal1 s 0 617 2880 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 2880 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 319 168 353 202 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 SCD
port 4 nsew
flabel corelocali s 607 390 641 424 0 FreeSans 340 0 0 0 SCD
port 4 nsew
flabel corelocali s 799 242 833 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 2719 94 2753 128 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2719 168 2753 202 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2719 242 2753 276 0 FreeSans 340 0 0 0 Q
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 2880 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 214974
string GDS_START 193972
<< end >>
