magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 644 561
rect 212 367 246 527
rect 288 401 354 493
rect 388 435 422 527
rect 456 401 522 493
rect 288 367 522 401
rect 556 367 590 527
rect 456 333 522 367
rect 456 299 627 333
rect 18 153 69 265
rect 173 199 248 265
rect 558 181 627 299
rect 21 17 69 119
rect 212 17 246 165
rect 288 147 627 181
rect 288 53 354 147
rect 388 17 422 113
rect 456 53 522 147
rect 556 17 590 113
rect 0 -17 644 17
<< obsli1 >>
rect 31 333 103 493
rect 31 299 323 333
rect 103 165 139 299
rect 282 249 323 299
rect 282 215 524 249
rect 103 58 169 165
<< metal1 >>
rect 0 496 644 592
rect 0 -48 644 48
<< labels >>
rlabel locali s 173 199 248 265 6 A
port 1 nsew signal input
rlabel locali s 18 153 69 265 6 B
port 2 nsew signal input
rlabel locali s 558 181 627 299 6 X
port 3 nsew signal output
rlabel locali s 456 401 522 493 6 X
port 3 nsew signal output
rlabel locali s 456 333 522 367 6 X
port 3 nsew signal output
rlabel locali s 456 299 627 333 6 X
port 3 nsew signal output
rlabel locali s 456 53 522 147 6 X
port 3 nsew signal output
rlabel locali s 288 401 354 493 6 X
port 3 nsew signal output
rlabel locali s 288 367 522 401 6 X
port 3 nsew signal output
rlabel locali s 288 147 627 181 6 X
port 3 nsew signal output
rlabel locali s 288 53 354 147 6 X
port 3 nsew signal output
rlabel locali s 556 17 590 113 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 388 17 422 113 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 212 17 246 165 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 21 17 69 119 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 644 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 644 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 556 367 590 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 388 435 422 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 212 367 246 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 644 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 644 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1009186
string GDS_START 1003484
<< end >>
