magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1104 561
rect 19 299 69 527
rect 187 383 253 527
rect 357 383 427 527
rect 529 383 595 527
rect 932 383 1001 417
rect 932 349 998 383
rect 932 336 1001 349
rect 852 315 1001 336
rect 852 302 998 315
rect 27 199 160 265
rect 211 199 361 265
rect 400 199 623 265
rect 679 199 811 265
rect 852 165 895 302
rect 1035 259 1082 325
rect 946 215 1082 259
rect 459 131 1069 165
rect 103 17 169 93
rect 647 51 681 131
rect 717 17 783 93
rect 817 51 851 131
rect 935 17 1001 93
rect 1035 51 1069 131
rect 0 -17 1104 17
<< obsli1 >>
rect 119 349 153 493
rect 287 349 321 493
rect 461 349 495 493
rect 822 485 888 493
rect 1035 485 1069 493
rect 629 451 1069 485
rect 717 349 783 417
rect 822 383 888 451
rect 119 315 783 349
rect 1035 359 1069 451
rect 35 131 421 165
rect 35 51 69 131
rect 203 51 237 131
rect 271 61 609 95
<< metal1 >>
rect 0 496 1104 592
rect 0 -48 1104 48
<< labels >>
rlabel locali s 400 199 623 265 6 A1
port 1 nsew signal input
rlabel locali s 211 199 361 265 6 A2
port 2 nsew signal input
rlabel locali s 27 199 160 265 6 A3
port 3 nsew signal input
rlabel locali s 679 199 811 265 6 B1
port 4 nsew signal input
rlabel locali s 1035 259 1082 325 6 C1
port 5 nsew signal input
rlabel locali s 946 215 1082 259 6 C1
port 5 nsew signal input
rlabel locali s 1035 51 1069 131 6 Y
port 6 nsew signal output
rlabel locali s 932 383 1001 417 6 Y
port 6 nsew signal output
rlabel locali s 932 349 998 383 6 Y
port 6 nsew signal output
rlabel locali s 932 336 1001 349 6 Y
port 6 nsew signal output
rlabel locali s 852 315 1001 336 6 Y
port 6 nsew signal output
rlabel locali s 852 302 998 315 6 Y
port 6 nsew signal output
rlabel locali s 852 165 895 302 6 Y
port 6 nsew signal output
rlabel locali s 817 51 851 131 6 Y
port 6 nsew signal output
rlabel locali s 647 51 681 131 6 Y
port 6 nsew signal output
rlabel locali s 459 131 1069 165 6 Y
port 6 nsew signal output
rlabel locali s 935 17 1001 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 717 17 783 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 103 17 169 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 1104 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1104 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 529 383 595 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 357 383 427 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 187 383 253 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 19 299 69 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 1104 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 1104 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1104 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3595280
string GDS_START 3584962
<< end >>
