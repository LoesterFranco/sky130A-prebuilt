magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1564 561
rect 115 359 165 527
rect 283 359 333 527
rect 1227 325 1277 425
rect 1395 325 1445 425
rect 1227 291 1547 325
rect 36 215 365 257
rect 419 215 814 257
rect 859 215 1141 257
rect 1175 215 1459 257
rect 1493 181 1547 291
rect 18 17 73 181
rect 107 145 1547 181
rect 107 51 173 145
rect 207 17 241 111
rect 275 51 341 145
rect 375 17 409 111
rect 443 51 509 145
rect 543 17 577 111
rect 611 51 677 145
rect 711 17 849 111
rect 883 51 949 145
rect 983 17 1017 111
rect 1051 51 1117 145
rect 1151 17 1185 111
rect 1219 51 1285 145
rect 1319 17 1353 111
rect 1387 51 1453 145
rect 1487 17 1521 111
rect 0 -17 1564 17
<< obsli1 >>
rect 18 325 81 493
rect 199 325 249 493
rect 367 459 764 493
rect 367 325 417 459
rect 18 291 417 325
rect 451 325 501 425
rect 535 359 585 459
rect 619 325 669 425
rect 703 359 764 459
rect 801 459 1529 493
rect 801 359 857 459
rect 891 325 941 425
rect 975 359 1025 459
rect 1059 325 1109 425
rect 1143 359 1193 459
rect 451 291 1109 325
rect 1311 359 1361 459
rect 1479 359 1529 459
<< metal1 >>
rect 0 496 1564 592
rect 0 -48 1564 48
<< labels >>
rlabel locali s 36 215 365 257 6 A
port 1 nsew signal input
rlabel locali s 419 215 814 257 6 B
port 2 nsew signal input
rlabel locali s 859 215 1141 257 6 C
port 3 nsew signal input
rlabel locali s 1175 215 1459 257 6 D
port 4 nsew signal input
rlabel locali s 1493 181 1547 291 6 Y
port 5 nsew signal output
rlabel locali s 1395 325 1445 425 6 Y
port 5 nsew signal output
rlabel locali s 1387 51 1453 145 6 Y
port 5 nsew signal output
rlabel locali s 1227 325 1277 425 6 Y
port 5 nsew signal output
rlabel locali s 1227 291 1547 325 6 Y
port 5 nsew signal output
rlabel locali s 1219 51 1285 145 6 Y
port 5 nsew signal output
rlabel locali s 1051 51 1117 145 6 Y
port 5 nsew signal output
rlabel locali s 883 51 949 145 6 Y
port 5 nsew signal output
rlabel locali s 611 51 677 145 6 Y
port 5 nsew signal output
rlabel locali s 443 51 509 145 6 Y
port 5 nsew signal output
rlabel locali s 275 51 341 145 6 Y
port 5 nsew signal output
rlabel locali s 107 145 1547 181 6 Y
port 5 nsew signal output
rlabel locali s 107 51 173 145 6 Y
port 5 nsew signal output
rlabel locali s 1487 17 1521 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1319 17 1353 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1151 17 1185 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 983 17 1017 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 711 17 849 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 543 17 577 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 375 17 409 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 207 17 241 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 18 17 73 181 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 1564 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1564 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 283 359 333 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 115 359 165 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 1564 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 1564 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1564 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1162934
string GDS_START 1150616
<< end >>
