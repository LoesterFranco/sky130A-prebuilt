magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 107 297 183 493
rect 19 211 86 265
rect 130 177 164 297
rect 198 215 275 265
rect 130 51 279 177
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 17 299 73 527
rect 227 299 279 527
rect 17 17 79 177
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
<< metal1 >>
rect 0 561 368 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 0 496 368 527
rect 0 17 368 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
rect 0 -48 368 -17
<< labels >>
rlabel locali s 198 215 275 265 6 A
port 1 nsew signal input
rlabel locali s 19 211 86 265 6 B
port 2 nsew signal input
rlabel locali s 130 177 164 297 6 Y
port 3 nsew signal output
rlabel locali s 130 51 279 177 6 Y
port 3 nsew signal output
rlabel locali s 107 297 183 493 6 Y
port 3 nsew signal output
rlabel metal1 s 0 -48 368 48 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 496 368 592 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 368 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2191256
string GDS_START 2187140
<< end >>
