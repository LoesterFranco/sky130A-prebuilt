magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 1326 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 79 47 109 177
rect 183 47 213 177
rect 267 47 297 177
rect 371 47 401 177
rect 455 47 485 177
rect 559 47 589 177
rect 643 47 673 177
rect 737 47 767 177
rect 831 47 861 177
rect 935 47 965 177
rect 1019 47 1049 177
rect 1123 47 1153 177
<< pmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 457 297 493 497
rect 551 297 587 497
rect 645 297 681 497
rect 739 297 775 497
rect 833 297 869 497
rect 927 297 963 497
rect 1021 297 1057 497
rect 1115 297 1151 497
<< ndiff >>
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 93 183 177
rect 109 59 129 93
rect 163 59 183 93
rect 109 47 183 59
rect 213 161 267 177
rect 213 127 223 161
rect 257 127 267 161
rect 213 93 267 127
rect 213 59 223 93
rect 257 59 267 93
rect 213 47 267 59
rect 297 93 371 177
rect 297 59 317 93
rect 351 59 371 93
rect 297 47 371 59
rect 401 161 455 177
rect 401 127 411 161
rect 445 127 455 161
rect 401 93 455 127
rect 401 59 411 93
rect 445 59 455 93
rect 401 47 455 59
rect 485 93 559 177
rect 485 59 505 93
rect 539 59 559 93
rect 485 47 559 59
rect 589 161 643 177
rect 589 127 599 161
rect 633 127 643 161
rect 589 93 643 127
rect 589 59 599 93
rect 633 59 643 93
rect 589 47 643 59
rect 673 161 737 177
rect 673 127 693 161
rect 727 127 737 161
rect 673 47 737 127
rect 767 93 831 177
rect 767 59 787 93
rect 821 59 831 93
rect 767 47 831 59
rect 861 161 935 177
rect 861 127 881 161
rect 915 127 935 161
rect 861 47 935 127
rect 965 93 1019 177
rect 965 59 975 93
rect 1009 59 1019 93
rect 965 47 1019 59
rect 1049 161 1123 177
rect 1049 127 1069 161
rect 1103 127 1123 161
rect 1049 47 1123 127
rect 1153 161 1205 177
rect 1153 127 1163 161
rect 1197 127 1205 161
rect 1153 93 1205 127
rect 1153 59 1163 93
rect 1197 59 1205 93
rect 1153 47 1205 59
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 485 175 497
rect 117 451 129 485
rect 163 451 175 485
rect 117 417 175 451
rect 117 383 129 417
rect 163 383 175 417
rect 117 349 175 383
rect 117 315 129 349
rect 163 315 175 349
rect 117 297 175 315
rect 211 485 269 497
rect 211 451 223 485
rect 257 451 269 485
rect 211 417 269 451
rect 211 383 223 417
rect 257 383 269 417
rect 211 297 269 383
rect 305 485 363 497
rect 305 451 317 485
rect 351 451 363 485
rect 305 417 363 451
rect 305 383 317 417
rect 351 383 363 417
rect 305 349 363 383
rect 305 315 317 349
rect 351 315 363 349
rect 305 297 363 315
rect 399 485 457 497
rect 399 451 411 485
rect 445 451 457 485
rect 399 417 457 451
rect 399 383 411 417
rect 445 383 457 417
rect 399 297 457 383
rect 493 485 551 497
rect 493 451 505 485
rect 539 451 551 485
rect 493 417 551 451
rect 493 383 505 417
rect 539 383 551 417
rect 493 349 551 383
rect 493 315 505 349
rect 539 315 551 349
rect 493 297 551 315
rect 587 485 645 497
rect 587 451 599 485
rect 633 451 645 485
rect 587 417 645 451
rect 587 383 599 417
rect 633 383 645 417
rect 587 297 645 383
rect 681 485 739 497
rect 681 451 693 485
rect 727 451 739 485
rect 681 417 739 451
rect 681 383 693 417
rect 727 383 739 417
rect 681 349 739 383
rect 681 315 693 349
rect 727 315 739 349
rect 681 297 739 315
rect 775 485 833 497
rect 775 451 787 485
rect 821 451 833 485
rect 775 417 833 451
rect 775 383 787 417
rect 821 383 833 417
rect 775 297 833 383
rect 869 485 927 497
rect 869 451 881 485
rect 915 451 927 485
rect 869 417 927 451
rect 869 383 881 417
rect 915 383 927 417
rect 869 349 927 383
rect 869 315 881 349
rect 915 315 927 349
rect 869 297 927 315
rect 963 485 1021 497
rect 963 451 975 485
rect 1009 451 1021 485
rect 963 417 1021 451
rect 963 383 975 417
rect 1009 383 1021 417
rect 963 297 1021 383
rect 1057 485 1115 497
rect 1057 451 1069 485
rect 1103 451 1115 485
rect 1057 417 1115 451
rect 1057 383 1069 417
rect 1103 383 1115 417
rect 1057 349 1115 383
rect 1057 315 1069 349
rect 1103 315 1115 349
rect 1057 297 1115 315
rect 1151 485 1205 497
rect 1151 451 1163 485
rect 1197 451 1205 485
rect 1151 417 1205 451
rect 1151 383 1163 417
rect 1197 383 1205 417
rect 1151 349 1205 383
rect 1151 315 1163 349
rect 1197 315 1205 349
rect 1151 297 1205 315
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 129 59 163 93
rect 223 127 257 161
rect 223 59 257 93
rect 317 59 351 93
rect 411 127 445 161
rect 411 59 445 93
rect 505 59 539 93
rect 599 127 633 161
rect 599 59 633 93
rect 693 127 727 161
rect 787 59 821 93
rect 881 127 915 161
rect 975 59 1009 93
rect 1069 127 1103 161
rect 1163 127 1197 161
rect 1163 59 1197 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 451 163 485
rect 129 383 163 417
rect 129 315 163 349
rect 223 451 257 485
rect 223 383 257 417
rect 317 451 351 485
rect 317 383 351 417
rect 317 315 351 349
rect 411 451 445 485
rect 411 383 445 417
rect 505 451 539 485
rect 505 383 539 417
rect 505 315 539 349
rect 599 451 633 485
rect 599 383 633 417
rect 693 451 727 485
rect 693 383 727 417
rect 693 315 727 349
rect 787 451 821 485
rect 787 383 821 417
rect 881 451 915 485
rect 881 383 915 417
rect 881 315 915 349
rect 975 451 1009 485
rect 975 383 1009 417
rect 1069 451 1103 485
rect 1069 383 1103 417
rect 1069 315 1103 349
rect 1163 451 1197 485
rect 1163 383 1197 417
rect 1163 315 1197 349
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 457 497 493 523
rect 551 497 587 523
rect 645 497 681 523
rect 739 497 775 523
rect 833 497 869 523
rect 927 497 963 523
rect 1021 497 1057 523
rect 1115 497 1151 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 457 282 493 297
rect 551 282 587 297
rect 645 282 681 297
rect 739 282 775 297
rect 833 282 869 297
rect 927 282 963 297
rect 1021 282 1057 297
rect 1115 282 1151 297
rect 79 265 119 282
rect 173 265 213 282
rect 267 265 307 282
rect 361 265 401 282
rect 455 265 495 282
rect 549 265 589 282
rect 79 249 589 265
rect 79 215 95 249
rect 129 215 163 249
rect 197 215 231 249
rect 265 215 299 249
rect 333 215 367 249
rect 401 215 435 249
rect 469 215 503 249
rect 537 215 589 249
rect 79 199 589 215
rect 79 177 109 199
rect 183 177 213 199
rect 267 177 297 199
rect 371 177 401 199
rect 455 177 485 199
rect 559 177 589 199
rect 643 265 683 282
rect 737 265 777 282
rect 831 265 871 282
rect 925 265 965 282
rect 1019 265 1059 282
rect 1113 265 1153 282
rect 643 249 1153 265
rect 643 215 777 249
rect 811 215 845 249
rect 879 215 913 249
rect 947 215 981 249
rect 1015 215 1153 249
rect 643 199 1153 215
rect 643 177 673 199
rect 737 177 767 199
rect 831 177 861 199
rect 935 177 965 199
rect 1019 177 1049 199
rect 1123 177 1153 199
rect 79 21 109 47
rect 183 21 213 47
rect 267 21 297 47
rect 371 21 401 47
rect 455 21 485 47
rect 559 21 589 47
rect 643 21 673 47
rect 737 21 767 47
rect 831 21 861 47
rect 935 21 965 47
rect 1019 21 1049 47
rect 1123 21 1153 47
<< polycont >>
rect 95 215 129 249
rect 163 215 197 249
rect 231 215 265 249
rect 299 215 333 249
rect 367 215 401 249
rect 435 215 469 249
rect 503 215 537 249
rect 777 215 811 249
rect 845 215 879 249
rect 913 215 947 249
rect 981 215 1015 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 25 485 79 527
rect 25 451 35 485
rect 69 451 79 485
rect 25 417 79 451
rect 25 383 35 417
rect 69 383 79 417
rect 25 349 79 383
rect 25 315 35 349
rect 69 315 79 349
rect 25 299 79 315
rect 113 485 179 493
rect 113 451 129 485
rect 163 451 179 485
rect 113 417 179 451
rect 113 383 129 417
rect 163 383 179 417
rect 113 349 179 383
rect 213 485 267 527
rect 213 451 223 485
rect 257 451 267 485
rect 213 417 267 451
rect 213 383 223 417
rect 257 383 267 417
rect 213 367 267 383
rect 301 485 367 493
rect 301 451 317 485
rect 351 451 367 485
rect 301 417 367 451
rect 301 383 317 417
rect 351 383 367 417
rect 113 315 129 349
rect 163 333 179 349
rect 301 349 367 383
rect 401 485 455 527
rect 401 451 411 485
rect 445 451 455 485
rect 401 417 455 451
rect 401 383 411 417
rect 445 383 455 417
rect 401 367 455 383
rect 489 485 555 493
rect 489 451 505 485
rect 539 451 555 485
rect 489 417 555 451
rect 489 383 505 417
rect 539 383 555 417
rect 301 333 317 349
rect 163 315 317 333
rect 351 333 367 349
rect 489 349 555 383
rect 589 485 643 527
rect 589 451 599 485
rect 633 451 643 485
rect 589 417 643 451
rect 589 383 599 417
rect 633 383 643 417
rect 589 367 643 383
rect 677 485 743 493
rect 677 451 693 485
rect 727 451 743 485
rect 677 417 743 451
rect 677 383 693 417
rect 727 383 743 417
rect 489 333 505 349
rect 351 315 505 333
rect 539 333 555 349
rect 677 349 743 383
rect 777 485 831 527
rect 777 451 787 485
rect 821 451 831 485
rect 777 417 831 451
rect 777 383 787 417
rect 821 383 831 417
rect 777 367 831 383
rect 865 485 931 493
rect 865 451 881 485
rect 915 451 931 485
rect 865 417 931 451
rect 865 383 881 417
rect 915 383 931 417
rect 677 333 693 349
rect 539 315 693 333
rect 727 333 743 349
rect 865 349 931 383
rect 965 485 1019 527
rect 965 451 975 485
rect 1009 451 1019 485
rect 965 417 1019 451
rect 965 383 975 417
rect 1009 383 1019 417
rect 965 367 1019 383
rect 1053 485 1119 493
rect 1053 451 1069 485
rect 1103 451 1119 485
rect 1053 417 1119 451
rect 1053 383 1069 417
rect 1103 383 1119 417
rect 865 333 881 349
rect 727 315 881 333
rect 915 333 931 349
rect 1053 349 1119 383
rect 1053 333 1069 349
rect 915 315 1069 333
rect 1103 315 1119 349
rect 113 299 1119 315
rect 1153 485 1207 527
rect 1153 451 1163 485
rect 1197 451 1207 485
rect 1153 417 1207 451
rect 1153 383 1163 417
rect 1197 383 1207 417
rect 1153 349 1207 383
rect 1153 315 1163 349
rect 1197 315 1207 349
rect 1153 299 1207 315
rect 79 249 553 265
rect 79 215 95 249
rect 129 215 163 249
rect 197 215 231 249
rect 265 215 299 249
rect 333 215 367 249
rect 401 215 435 249
rect 469 215 503 249
rect 537 215 553 249
rect 79 211 553 215
rect 667 177 727 299
rect 1065 265 1119 299
rect 761 249 1031 265
rect 761 215 777 249
rect 811 215 845 249
rect 879 215 913 249
rect 947 215 981 249
rect 1015 215 1031 249
rect 761 211 1031 215
rect 1065 211 1183 265
rect 1065 177 1119 211
rect 18 161 633 177
rect 18 127 35 161
rect 69 143 223 161
rect 69 127 85 143
rect 18 93 85 127
rect 207 127 223 143
rect 257 143 411 161
rect 257 127 273 143
rect 18 59 35 93
rect 69 59 85 93
rect 18 51 85 59
rect 119 93 173 109
rect 119 59 129 93
rect 163 59 173 93
rect 119 17 173 59
rect 207 93 273 127
rect 395 127 411 143
rect 445 143 599 161
rect 445 127 461 143
rect 207 59 223 93
rect 257 59 273 93
rect 207 51 273 59
rect 307 93 361 109
rect 307 59 317 93
rect 351 59 361 93
rect 307 17 361 59
rect 395 93 461 127
rect 583 127 599 143
rect 667 161 1119 177
rect 667 127 693 161
rect 727 127 881 161
rect 915 127 1069 161
rect 1103 127 1119 161
rect 1153 161 1213 177
rect 1153 127 1163 161
rect 1197 127 1213 161
rect 395 59 411 93
rect 445 59 461 93
rect 395 51 461 59
rect 495 93 549 109
rect 495 59 505 93
rect 539 59 549 93
rect 495 17 549 59
rect 583 93 633 127
rect 1153 93 1213 127
rect 583 59 599 93
rect 633 59 787 93
rect 821 59 975 93
rect 1009 59 1163 93
rect 1197 59 1213 93
rect 583 51 1213 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
flabel corelocali s 673 221 707 255 0 FreeSans 250 0 0 0 Y
port 7 nsew
flabel corelocali s 857 221 891 255 0 FreeSans 250 0 0 0 A
port 1 nsew
flabel corelocali s 305 221 339 255 0 FreeSans 250 0 0 0 B
port 2 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew
rlabel comment s 0 0 0 0 4 nand2_6
<< properties >>
string FIXED_BBOX 0 0 1288 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3440178
string GDS_START 3430442
<< end >>
