magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 920 561
rect 18 299 69 527
rect 103 333 169 493
rect 203 367 237 527
rect 271 333 337 493
rect 371 367 437 527
rect 471 333 537 493
rect 599 367 665 527
rect 719 333 785 493
rect 103 289 785 333
rect 819 289 885 527
rect 22 215 169 255
rect 214 215 340 255
rect 447 215 616 255
rect 674 211 785 289
rect 833 215 899 255
rect 119 17 153 109
rect 719 127 785 211
rect 0 -17 920 17
<< obsli1 >>
rect 18 147 237 181
rect 18 51 85 147
rect 187 93 237 147
rect 271 127 617 181
rect 651 93 685 177
rect 819 93 885 181
rect 187 51 425 93
rect 463 51 885 93
<< metal1 >>
rect 0 496 920 592
rect 0 -48 920 48
<< labels >>
rlabel locali s 833 215 899 255 6 A
port 1 nsew signal input
rlabel locali s 447 215 616 255 6 B
port 2 nsew signal input
rlabel locali s 214 215 340 255 6 C
port 3 nsew signal input
rlabel locali s 22 215 169 255 6 D
port 4 nsew signal input
rlabel locali s 719 333 785 493 6 Y
port 5 nsew signal output
rlabel locali s 719 127 785 211 6 Y
port 5 nsew signal output
rlabel locali s 674 211 785 289 6 Y
port 5 nsew signal output
rlabel locali s 471 333 537 493 6 Y
port 5 nsew signal output
rlabel locali s 271 333 337 493 6 Y
port 5 nsew signal output
rlabel locali s 103 333 169 493 6 Y
port 5 nsew signal output
rlabel locali s 103 289 785 333 6 Y
port 5 nsew signal output
rlabel locali s 119 17 153 109 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 920 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 920 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 819 289 885 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 599 367 665 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 371 367 437 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 203 367 237 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 18 299 69 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 920 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 920 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 920 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1850160
string GDS_START 1841432
<< end >>
