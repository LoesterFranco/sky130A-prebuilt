magic
tech sky130A
magscale 1 2
timestamp 1604502701
<< nwell >>
rect -38 332 902 704
<< pwell >>
rect 0 0 864 49
<< scpmos >>
rect 125 368 155 568
rect 279 368 309 592
rect 369 368 399 592
rect 477 368 507 592
rect 567 368 597 592
rect 657 368 687 592
rect 748 368 778 592
<< nmoslvt >>
rect 84 74 114 202
rect 282 74 312 222
rect 368 74 398 222
rect 468 74 498 222
rect 574 74 604 222
rect 660 74 690 222
rect 746 74 776 222
<< ndiff >>
rect 27 190 84 202
rect 27 156 39 190
rect 73 156 84 190
rect 27 120 84 156
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 152 171 202
rect 114 118 125 152
rect 159 118 171 152
rect 114 74 171 118
rect 225 152 282 222
rect 225 118 237 152
rect 271 118 282 152
rect 225 74 282 118
rect 312 177 368 222
rect 312 143 323 177
rect 357 143 368 177
rect 312 74 368 143
rect 398 210 468 222
rect 398 176 423 210
rect 457 176 468 210
rect 398 120 468 176
rect 398 86 423 120
rect 457 86 468 120
rect 398 74 468 86
rect 498 152 574 222
rect 498 118 523 152
rect 557 118 574 152
rect 498 74 574 118
rect 604 210 660 222
rect 604 176 615 210
rect 649 176 660 210
rect 604 120 660 176
rect 604 86 615 120
rect 649 86 660 120
rect 604 74 660 86
rect 690 146 746 222
rect 690 112 701 146
rect 735 112 746 146
rect 690 74 746 112
rect 776 210 833 222
rect 776 176 787 210
rect 821 176 833 210
rect 776 120 833 176
rect 776 86 787 120
rect 821 86 833 120
rect 776 74 833 86
<< pdiff >>
rect 191 580 279 592
rect 191 568 217 580
rect 64 560 125 568
rect 64 526 78 560
rect 112 526 125 560
rect 64 492 125 526
rect 64 458 78 492
rect 112 458 125 492
rect 64 424 125 458
rect 64 390 78 424
rect 112 390 125 424
rect 64 368 125 390
rect 155 546 217 568
rect 251 546 279 580
rect 155 497 279 546
rect 155 463 217 497
rect 251 463 279 497
rect 155 414 279 463
rect 155 380 217 414
rect 251 380 279 414
rect 155 368 279 380
rect 309 580 369 592
rect 309 546 322 580
rect 356 546 369 580
rect 309 497 369 546
rect 309 463 322 497
rect 356 463 369 497
rect 309 414 369 463
rect 309 380 322 414
rect 356 380 369 414
rect 309 368 369 380
rect 399 580 477 592
rect 399 546 416 580
rect 450 546 477 580
rect 399 368 477 546
rect 507 578 567 592
rect 507 544 520 578
rect 554 544 567 578
rect 507 368 567 544
rect 597 519 657 592
rect 597 485 610 519
rect 644 485 657 519
rect 597 368 657 485
rect 687 580 748 592
rect 687 546 700 580
rect 734 546 748 580
rect 687 492 748 546
rect 687 458 700 492
rect 734 458 748 492
rect 687 368 748 458
rect 778 580 837 592
rect 778 546 791 580
rect 825 546 837 580
rect 778 497 837 546
rect 778 463 791 497
rect 825 463 837 497
rect 778 414 837 463
rect 778 380 791 414
rect 825 380 837 414
rect 778 368 837 380
<< ndiffc >>
rect 39 156 73 190
rect 39 86 73 120
rect 125 118 159 152
rect 237 118 271 152
rect 323 143 357 177
rect 423 176 457 210
rect 423 86 457 120
rect 523 118 557 152
rect 615 176 649 210
rect 615 86 649 120
rect 701 112 735 146
rect 787 176 821 210
rect 787 86 821 120
<< pdiffc >>
rect 78 526 112 560
rect 78 458 112 492
rect 78 390 112 424
rect 217 546 251 580
rect 217 463 251 497
rect 217 380 251 414
rect 322 546 356 580
rect 322 463 356 497
rect 322 380 356 414
rect 416 546 450 580
rect 520 544 554 578
rect 610 485 644 519
rect 700 546 734 580
rect 700 458 734 492
rect 791 546 825 580
rect 791 463 825 497
rect 791 380 825 414
<< poly >>
rect 125 568 155 594
rect 279 592 309 618
rect 369 592 399 618
rect 477 592 507 618
rect 567 592 597 618
rect 657 592 687 618
rect 748 592 778 618
rect 125 353 155 368
rect 279 353 309 368
rect 369 353 399 368
rect 477 353 507 368
rect 567 353 597 368
rect 657 353 687 368
rect 748 353 778 368
rect 122 336 158 353
rect 84 320 158 336
rect 84 286 108 320
rect 142 286 158 320
rect 276 310 312 353
rect 84 270 158 286
rect 206 305 312 310
rect 366 305 402 353
rect 474 336 510 353
rect 564 336 600 353
rect 654 336 690 353
rect 206 294 402 305
rect 84 202 114 270
rect 206 260 222 294
rect 256 274 402 294
rect 450 320 516 336
rect 450 286 466 320
rect 500 286 516 320
rect 256 260 398 274
rect 450 270 516 286
rect 564 320 690 336
rect 564 286 589 320
rect 623 286 690 320
rect 564 270 690 286
rect 206 244 398 260
rect 282 222 312 244
rect 368 222 398 244
rect 468 222 498 270
rect 574 222 604 270
rect 660 222 690 270
rect 745 330 781 353
rect 745 314 811 330
rect 745 280 761 314
rect 795 280 811 314
rect 745 264 811 280
rect 746 222 776 264
rect 84 48 114 74
rect 282 48 312 74
rect 368 48 398 74
rect 468 48 498 74
rect 574 48 604 74
rect 660 48 690 74
rect 746 48 776 74
<< polycont >>
rect 108 286 142 320
rect 222 260 256 294
rect 466 286 500 320
rect 589 286 623 320
rect 761 280 795 314
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 201 580 267 649
rect 23 560 128 572
rect 23 526 78 560
rect 112 526 128 560
rect 23 492 128 526
rect 23 458 78 492
rect 112 458 128 492
rect 23 424 128 458
rect 23 390 78 424
rect 112 390 128 424
rect 201 546 217 580
rect 251 546 267 580
rect 201 497 267 546
rect 201 463 217 497
rect 251 463 267 497
rect 201 414 267 463
rect 23 236 57 390
rect 201 380 217 414
rect 251 380 267 414
rect 201 364 267 380
rect 306 580 356 596
rect 306 546 322 580
rect 306 497 356 546
rect 396 580 470 649
rect 396 546 416 580
rect 450 546 470 580
rect 396 530 470 546
rect 504 581 751 615
rect 504 578 570 581
rect 504 544 520 578
rect 554 544 570 578
rect 684 580 751 581
rect 504 526 570 544
rect 306 463 322 497
rect 610 519 644 547
rect 356 485 610 492
rect 356 463 644 485
rect 306 458 644 463
rect 684 546 700 580
rect 734 546 751 580
rect 684 492 751 546
rect 684 458 700 492
rect 734 458 751 492
rect 791 580 841 649
rect 825 546 841 580
rect 791 497 841 546
rect 825 463 841 497
rect 306 414 373 458
rect 306 380 322 414
rect 356 380 373 414
rect 92 320 167 356
rect 92 286 108 320
rect 142 286 167 320
rect 92 270 167 286
rect 206 294 272 310
rect 206 260 222 294
rect 256 260 272 294
rect 206 236 272 260
rect 306 236 373 380
rect 450 390 743 424
rect 450 320 516 390
rect 450 286 466 320
rect 500 286 516 320
rect 450 270 516 286
rect 564 320 647 356
rect 564 286 589 320
rect 623 286 647 320
rect 564 270 647 286
rect 697 330 743 390
rect 791 414 841 463
rect 825 380 841 414
rect 791 364 841 380
rect 697 314 811 330
rect 697 280 761 314
rect 795 280 811 314
rect 697 264 811 280
rect 23 202 272 236
rect 23 190 73 202
rect 23 156 39 190
rect 323 177 373 236
rect 23 120 73 156
rect 23 86 39 120
rect 23 70 73 86
rect 109 152 175 168
rect 109 118 125 152
rect 159 118 175 152
rect 109 17 175 118
rect 221 152 287 168
rect 221 118 237 152
rect 271 118 287 152
rect 357 143 373 177
rect 323 123 373 143
rect 407 230 649 236
rect 407 210 837 230
rect 407 176 423 210
rect 457 202 615 210
rect 457 176 473 202
rect 221 85 287 118
rect 407 120 473 176
rect 649 196 787 210
rect 407 86 423 120
rect 457 86 473 120
rect 407 85 473 86
rect 221 51 473 85
rect 507 152 573 168
rect 507 118 523 152
rect 557 118 573 152
rect 507 17 573 118
rect 615 120 649 176
rect 821 176 837 210
rect 615 70 649 86
rect 685 146 751 162
rect 685 112 701 146
rect 735 112 751 146
rect 685 17 751 112
rect 787 120 837 176
rect 821 86 837 120
rect 787 70 837 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o21bai_2
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 B1_N
port 3 nsew
flabel corelocali s 319 242 353 276 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 319 390 353 424 0 FreeSans 340 0 0 0 Y
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 864 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1143252
string GDS_START 1135664
<< end >>
