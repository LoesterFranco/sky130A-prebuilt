magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 736 561
rect 17 312 85 527
rect 122 425 532 483
rect 566 367 622 527
rect 17 151 85 265
rect 304 199 452 323
rect 664 299 719 493
rect 486 199 562 265
rect 17 17 85 117
rect 685 152 719 299
rect 207 17 273 117
rect 382 17 448 97
rect 550 17 626 97
rect 664 83 719 152
rect 0 -17 736 17
<< obsli1 >>
rect 119 265 167 384
rect 206 357 532 391
rect 206 299 270 357
rect 498 333 532 357
rect 119 199 250 265
rect 498 299 630 333
rect 596 265 630 299
rect 596 199 651 265
rect 119 61 168 199
rect 596 165 630 199
rect 313 131 630 165
rect 313 61 347 131
rect 482 61 516 131
<< metal1 >>
rect 0 496 736 592
rect 0 -48 736 48
<< labels >>
rlabel locali s 486 199 562 265 6 A
port 1 nsew signal input
rlabel locali s 122 425 532 483 6 B
port 2 nsew signal input
rlabel locali s 304 199 452 323 6 C
port 3 nsew signal input
rlabel locali s 17 151 85 265 6 D_N
port 4 nsew signal input
rlabel locali s 685 152 719 299 6 X
port 5 nsew signal output
rlabel locali s 664 299 719 493 6 X
port 5 nsew signal output
rlabel locali s 664 83 719 152 6 X
port 5 nsew signal output
rlabel locali s 550 17 626 97 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 382 17 448 97 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 207 17 273 117 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 17 17 85 117 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 736 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 736 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 566 367 622 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 17 312 85 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 736 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 736 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1090244
string GDS_START 1083020
<< end >>
