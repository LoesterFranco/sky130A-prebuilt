magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2300 561
rect 22 261 66 393
rect 103 349 179 417
rect 291 349 367 417
rect 435 349 555 417
rect 667 349 743 417
rect 103 315 743 349
rect 859 383 935 527
rect 1064 383 1208 527
rect 1373 383 1449 527
rect 1561 383 1637 527
rect 1853 383 1929 527
rect 2041 383 2117 527
rect 22 215 380 261
rect 435 198 523 315
rect 567 199 791 265
rect 835 215 1213 257
rect 1349 215 1709 260
rect 1829 215 2207 256
rect 479 161 523 198
rect 479 127 1233 161
rect 2151 151 2207 215
rect 103 17 179 93
rect 291 17 367 93
rect 1769 17 1835 93
rect 1947 17 2023 93
rect 2137 17 2215 93
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2300 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
<< obsli1 >>
rect 19 451 821 485
rect 787 349 821 451
rect 979 349 1013 493
rect 1258 349 1292 493
rect 1493 349 1527 493
rect 1681 349 1715 493
rect 1973 349 2007 493
rect 2161 349 2195 493
rect 787 315 2195 349
rect 35 127 445 161
rect 1373 127 2101 161
rect 35 51 69 127
rect 223 51 257 127
rect 411 93 445 127
rect 411 59 837 93
rect 885 59 1731 93
rect 1879 51 1913 127
rect 2067 51 2101 127
<< metal1 >>
rect 0 561 2300 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2300 561
rect 0 496 2300 527
rect 0 17 2300 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2300 17
rect 0 -48 2300 -17
<< labels >>
rlabel locali s 835 215 1213 257 6 A1
port 1 nsew signal input
rlabel locali s 1349 215 1709 260 6 A2
port 2 nsew signal input
rlabel locali s 2151 151 2207 215 6 A3
port 3 nsew signal input
rlabel locali s 1829 215 2207 256 6 A3
port 3 nsew signal input
rlabel locali s 567 199 791 265 6 B1
port 4 nsew signal input
rlabel locali s 22 261 66 393 6 B2
port 5 nsew signal input
rlabel locali s 22 215 380 261 6 B2
port 5 nsew signal input
rlabel locali s 667 349 743 417 6 Y
port 6 nsew signal output
rlabel locali s 479 161 523 198 6 Y
port 6 nsew signal output
rlabel locali s 479 127 1233 161 6 Y
port 6 nsew signal output
rlabel locali s 435 349 555 417 6 Y
port 6 nsew signal output
rlabel locali s 435 198 523 315 6 Y
port 6 nsew signal output
rlabel locali s 291 349 367 417 6 Y
port 6 nsew signal output
rlabel locali s 103 349 179 417 6 Y
port 6 nsew signal output
rlabel locali s 103 315 743 349 6 Y
port 6 nsew signal output
rlabel viali s 2145 -17 2179 17 8 VGND
port 7 nsew ground bidirectional
rlabel viali s 2053 -17 2087 17 8 VGND
port 7 nsew ground bidirectional
rlabel viali s 1961 -17 1995 17 8 VGND
port 7 nsew ground bidirectional
rlabel viali s 1869 -17 1903 17 8 VGND
port 7 nsew ground bidirectional
rlabel viali s 1777 -17 1811 17 8 VGND
port 7 nsew ground bidirectional
rlabel viali s 1685 -17 1719 17 8 VGND
port 7 nsew ground bidirectional
rlabel viali s 1593 -17 1627 17 8 VGND
port 7 nsew ground bidirectional
rlabel viali s 1501 -17 1535 17 8 VGND
port 7 nsew ground bidirectional
rlabel viali s 1409 -17 1443 17 8 VGND
port 7 nsew ground bidirectional
rlabel viali s 1317 -17 1351 17 8 VGND
port 7 nsew ground bidirectional
rlabel viali s 1225 -17 1259 17 8 VGND
port 7 nsew ground bidirectional
rlabel viali s 1133 -17 1167 17 8 VGND
port 7 nsew ground bidirectional
rlabel viali s 1041 -17 1075 17 8 VGND
port 7 nsew ground bidirectional
rlabel viali s 949 -17 983 17 8 VGND
port 7 nsew ground bidirectional
rlabel viali s 857 -17 891 17 8 VGND
port 7 nsew ground bidirectional
rlabel viali s 765 -17 799 17 8 VGND
port 7 nsew ground bidirectional
rlabel viali s 673 -17 707 17 8 VGND
port 7 nsew ground bidirectional
rlabel viali s 581 -17 615 17 8 VGND
port 7 nsew ground bidirectional
rlabel viali s 489 -17 523 17 8 VGND
port 7 nsew ground bidirectional
rlabel viali s 397 -17 431 17 8 VGND
port 7 nsew ground bidirectional
rlabel viali s 305 -17 339 17 8 VGND
port 7 nsew ground bidirectional
rlabel viali s 213 -17 247 17 8 VGND
port 7 nsew ground bidirectional
rlabel viali s 121 -17 155 17 8 VGND
port 7 nsew ground bidirectional
rlabel viali s 29 -17 63 17 8 VGND
port 7 nsew ground bidirectional
rlabel locali s 2137 17 2215 93 6 VGND
port 7 nsew ground bidirectional
rlabel locali s 1947 17 2023 93 6 VGND
port 7 nsew ground bidirectional
rlabel locali s 1769 17 1835 93 6 VGND
port 7 nsew ground bidirectional
rlabel locali s 291 17 367 93 6 VGND
port 7 nsew ground bidirectional
rlabel locali s 103 17 179 93 6 VGND
port 7 nsew ground bidirectional
rlabel locali s 0 -17 2300 17 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 -48 2300 48 8 VGND
port 7 nsew ground bidirectional
rlabel viali s 2145 527 2179 561 6 VPWR
port 8 nsew power bidirectional
rlabel viali s 2053 527 2087 561 6 VPWR
port 8 nsew power bidirectional
rlabel viali s 1961 527 1995 561 6 VPWR
port 8 nsew power bidirectional
rlabel viali s 1869 527 1903 561 6 VPWR
port 8 nsew power bidirectional
rlabel viali s 1777 527 1811 561 6 VPWR
port 8 nsew power bidirectional
rlabel viali s 1685 527 1719 561 6 VPWR
port 8 nsew power bidirectional
rlabel viali s 1593 527 1627 561 6 VPWR
port 8 nsew power bidirectional
rlabel viali s 1501 527 1535 561 6 VPWR
port 8 nsew power bidirectional
rlabel viali s 1409 527 1443 561 6 VPWR
port 8 nsew power bidirectional
rlabel viali s 1317 527 1351 561 6 VPWR
port 8 nsew power bidirectional
rlabel viali s 1225 527 1259 561 6 VPWR
port 8 nsew power bidirectional
rlabel viali s 1133 527 1167 561 6 VPWR
port 8 nsew power bidirectional
rlabel viali s 1041 527 1075 561 6 VPWR
port 8 nsew power bidirectional
rlabel viali s 949 527 983 561 6 VPWR
port 8 nsew power bidirectional
rlabel viali s 857 527 891 561 6 VPWR
port 8 nsew power bidirectional
rlabel viali s 765 527 799 561 6 VPWR
port 8 nsew power bidirectional
rlabel viali s 673 527 707 561 6 VPWR
port 8 nsew power bidirectional
rlabel viali s 581 527 615 561 6 VPWR
port 8 nsew power bidirectional
rlabel viali s 489 527 523 561 6 VPWR
port 8 nsew power bidirectional
rlabel viali s 397 527 431 561 6 VPWR
port 8 nsew power bidirectional
rlabel viali s 305 527 339 561 6 VPWR
port 8 nsew power bidirectional
rlabel viali s 213 527 247 561 6 VPWR
port 8 nsew power bidirectional
rlabel viali s 121 527 155 561 6 VPWR
port 8 nsew power bidirectional
rlabel viali s 29 527 63 561 6 VPWR
port 8 nsew power bidirectional
rlabel locali s 2041 383 2117 527 6 VPWR
port 8 nsew power bidirectional
rlabel locali s 1853 383 1929 527 6 VPWR
port 8 nsew power bidirectional
rlabel locali s 1561 383 1637 527 6 VPWR
port 8 nsew power bidirectional
rlabel locali s 1373 383 1449 527 6 VPWR
port 8 nsew power bidirectional
rlabel locali s 1064 383 1208 527 6 VPWR
port 8 nsew power bidirectional
rlabel locali s 859 383 935 527 6 VPWR
port 8 nsew power bidirectional
rlabel locali s 0 527 2300 561 6 VPWR
port 8 nsew power bidirectional
rlabel metal1 s 0 496 2300 592 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2300 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1478552
string GDS_START 1461808
<< end >>
