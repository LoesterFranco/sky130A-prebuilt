magic
tech sky130A
magscale 1 2
timestamp 1601050088
<< obsli1 >>
rect 0 649 31 683
rect 65 649 96 683
rect 18 572 78 613
rect 18 538 31 572
rect 65 538 78 572
rect 18 378 78 538
rect 18 17 78 288
rect 0 -17 31 17
rect 65 -17 96 17
<< obsli1c >>
rect 31 649 65 683
rect 31 538 65 572
rect 31 -17 65 17
<< metal1 >>
rect 0 683 96 715
rect 0 649 31 683
rect 65 649 96 683
rect 0 617 96 649
rect 16 572 80 581
rect 16 538 31 572
rect 65 538 80 572
rect 16 529 80 538
rect 0 17 96 49
rect 0 -17 31 17
rect 65 -17 96 17
rect 0 -49 96 -17
<< labels >>
rlabel metal1 s 0 -49 96 49 8 VGND
port 1 nsew ground bidirectional
rlabel metal1 s 16 529 80 581 6 VPB
port 2 nsew power bidirectional
rlabel metal1 s 0 617 96 715 6 VPWR
port 3 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE WELLTAP
string FIXED_BBOX 0 0 96 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 460178
string GDS_START 458274
<< end >>
