magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 17 435 73 596
rect 213 435 265 547
rect 399 435 493 547
rect 17 401 493 435
rect 17 384 73 401
rect 17 199 51 384
rect 121 333 425 367
rect 121 299 167 333
rect 85 233 167 299
rect 201 233 267 299
rect 359 226 425 333
rect 459 260 493 401
rect 613 390 855 424
rect 989 390 1211 424
rect 613 360 647 390
rect 535 294 647 360
rect 821 356 855 390
rect 989 356 1023 390
rect 1177 356 1211 390
rect 459 226 568 260
rect 681 252 747 356
rect 821 290 895 356
rect 937 290 1023 356
rect 1061 290 1127 356
rect 1177 290 1291 356
rect 502 218 568 226
rect 890 222 1316 256
rect 890 218 943 222
rect 17 165 284 199
rect 218 156 284 165
rect 502 184 943 218
rect 502 70 568 184
rect 890 70 943 184
rect 1264 70 1316 222
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 113 596 667 615
rect 113 581 865 596
rect 113 469 179 581
rect 299 469 365 581
rect 527 492 561 547
rect 601 530 865 581
rect 601 526 667 530
rect 900 496 943 596
rect 979 530 1051 649
rect 1085 496 1131 596
rect 1165 530 1231 649
rect 1267 496 1321 600
rect 900 492 1321 496
rect 527 458 1321 492
rect 527 394 561 458
rect 889 390 955 458
rect 1255 390 1321 458
rect 23 17 96 131
rect 318 122 356 177
rect 132 70 356 122
rect 390 17 456 188
rect 604 116 854 150
rect 604 70 654 116
rect 690 17 768 82
rect 804 70 854 116
rect 977 154 1230 188
rect 977 70 1043 154
rect 1077 17 1143 120
rect 1180 66 1230 154
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
<< metal1 >>
rect 0 683 1344 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 0 617 1344 649
rect 0 17 1344 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
rect 0 -49 1344 -17
<< labels >>
rlabel locali s 1177 356 1211 390 6 A1
port 1 nsew signal input
rlabel locali s 1177 290 1291 356 6 A1
port 1 nsew signal input
rlabel locali s 989 390 1211 424 6 A1
port 1 nsew signal input
rlabel locali s 989 356 1023 390 6 A1
port 1 nsew signal input
rlabel locali s 937 290 1023 356 6 A1
port 1 nsew signal input
rlabel locali s 1061 290 1127 356 6 A2
port 2 nsew signal input
rlabel locali s 821 356 855 390 6 B1
port 3 nsew signal input
rlabel locali s 821 290 895 356 6 B1
port 3 nsew signal input
rlabel locali s 613 390 855 424 6 B1
port 3 nsew signal input
rlabel locali s 613 360 647 390 6 B1
port 3 nsew signal input
rlabel locali s 535 294 647 360 6 B1
port 3 nsew signal input
rlabel locali s 681 252 747 356 6 B2
port 4 nsew signal input
rlabel locali s 201 233 267 299 6 C1
port 5 nsew signal input
rlabel locali s 359 226 425 333 6 C2
port 6 nsew signal input
rlabel locali s 121 333 425 367 6 C2
port 6 nsew signal input
rlabel locali s 121 299 167 333 6 C2
port 6 nsew signal input
rlabel locali s 85 233 167 299 6 C2
port 6 nsew signal input
rlabel locali s 1264 70 1316 222 6 Y
port 7 nsew signal output
rlabel locali s 890 222 1316 256 6 Y
port 7 nsew signal output
rlabel locali s 890 218 943 222 6 Y
port 7 nsew signal output
rlabel locali s 890 70 943 184 6 Y
port 7 nsew signal output
rlabel locali s 502 218 568 226 6 Y
port 7 nsew signal output
rlabel locali s 502 184 943 218 6 Y
port 7 nsew signal output
rlabel locali s 502 70 568 184 6 Y
port 7 nsew signal output
rlabel locali s 459 260 493 401 6 Y
port 7 nsew signal output
rlabel locali s 459 226 568 260 6 Y
port 7 nsew signal output
rlabel locali s 399 435 493 547 6 Y
port 7 nsew signal output
rlabel locali s 218 156 284 165 6 Y
port 7 nsew signal output
rlabel locali s 213 435 265 547 6 Y
port 7 nsew signal output
rlabel locali s 17 435 73 596 6 Y
port 7 nsew signal output
rlabel locali s 17 401 493 435 6 Y
port 7 nsew signal output
rlabel locali s 17 384 73 401 6 Y
port 7 nsew signal output
rlabel locali s 17 199 51 384 6 Y
port 7 nsew signal output
rlabel locali s 17 165 284 199 6 Y
port 7 nsew signal output
rlabel metal1 s 0 -49 1344 49 8 VGND
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1344 715 6 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1344 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3475432
string GDS_START 3463852
<< end >>
