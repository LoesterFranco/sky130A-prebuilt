magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 121 424 363 596
rect 106 390 363 424
rect 21 236 72 356
rect 106 226 140 390
rect 174 260 263 356
rect 297 260 363 356
rect 106 176 361 226
rect 123 73 161 176
rect 295 70 361 176
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 384 683
rect 21 465 87 649
rect 21 390 71 465
rect 23 142 72 202
rect 23 17 89 142
rect 195 17 261 142
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 384 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
<< metal1 >>
rect 0 683 384 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 384 683
rect 0 617 384 649
rect 0 17 384 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 384 17
rect 0 -49 384 -17
<< labels >>
rlabel locali s 21 236 72 356 6 A
port 1 nsew signal input
rlabel locali s 174 260 263 356 6 B
port 2 nsew signal input
rlabel locali s 297 260 363 356 6 C
port 3 nsew signal input
rlabel locali s 295 70 361 176 6 Y
port 4 nsew signal output
rlabel locali s 123 73 161 176 6 Y
port 4 nsew signal output
rlabel locali s 121 424 363 596 6 Y
port 4 nsew signal output
rlabel locali s 106 390 363 424 6 Y
port 4 nsew signal output
rlabel locali s 106 226 140 390 6 Y
port 4 nsew signal output
rlabel locali s 106 176 361 226 6 Y
port 4 nsew signal output
rlabel metal1 s 0 -49 384 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 617 384 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 384 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1579262
string GDS_START 1574480
<< end >>
