magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 17 197 66 325
rect 295 191 378 265
rect 1119 299 1179 491
rect 1142 265 1179 299
rect 1307 265 1361 491
rect 1142 199 1447 265
rect 1142 149 1179 199
rect 1119 83 1179 149
rect 1307 77 1361 199
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 35 393 69 493
rect 103 427 179 527
rect 35 359 178 393
rect 132 314 178 359
rect 166 280 178 314
rect 132 161 178 280
rect 35 127 178 161
rect 223 388 257 493
rect 35 69 69 127
rect 103 17 179 93
rect 223 69 257 354
rect 311 333 377 483
rect 421 367 484 527
rect 605 451 790 485
rect 534 388 591 401
rect 568 354 591 388
rect 311 299 458 333
rect 424 219 458 299
rect 534 271 591 354
rect 635 314 713 399
rect 669 283 713 314
rect 424 157 508 219
rect 635 207 669 280
rect 327 153 508 157
rect 327 123 458 153
rect 583 141 669 207
rect 756 265 790 451
rect 824 427 858 527
rect 928 373 972 487
rect 828 307 972 373
rect 934 265 972 307
rect 1018 299 1075 527
rect 1213 299 1263 527
rect 1401 299 1435 527
rect 756 199 900 265
rect 934 199 1098 265
rect 327 69 361 123
rect 756 107 790 199
rect 395 17 471 89
rect 618 73 790 107
rect 824 17 858 122
rect 934 83 972 199
rect 1018 17 1075 143
rect 1213 17 1263 165
rect 1401 17 1435 143
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 132 280 166 314
rect 223 354 257 388
rect 534 354 568 388
rect 635 280 669 314
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< obsm1 >>
rect 211 388 269 394
rect 522 388 580 394
rect 211 354 223 388
rect 257 360 534 388
rect 257 354 269 360
rect 211 348 269 354
rect 522 354 534 360
rect 568 354 580 388
rect 522 348 580 354
rect 120 314 682 320
rect 120 280 132 314
rect 166 292 635 314
rect 166 280 178 292
rect 120 274 178 280
rect 623 280 635 292
rect 669 280 682 314
rect 623 274 682 280
<< labels >>
rlabel locali s 295 191 378 265 6 D
port 1 nsew signal input
rlabel locali s 17 197 66 325 6 GATE_N
port 2 nsew signal input
rlabel locali s 1307 265 1361 491 6 Q
port 3 nsew signal output
rlabel locali s 1307 77 1361 199 6 Q
port 3 nsew signal output
rlabel locali s 1142 265 1179 299 6 Q
port 3 nsew signal output
rlabel locali s 1142 199 1447 265 6 Q
port 3 nsew signal output
rlabel locali s 1142 149 1179 199 6 Q
port 3 nsew signal output
rlabel locali s 1119 299 1179 491 6 Q
port 3 nsew signal output
rlabel locali s 1119 83 1179 149 6 Q
port 3 nsew signal output
rlabel metal1 s 0 -48 1472 48 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 496 1472 592 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1472 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1960880
string GDS_START 1948756
<< end >>
