magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1564 561
rect 119 325 161 425
rect 279 325 329 425
rect 447 325 497 425
rect 615 325 665 425
rect 119 289 665 325
rect 887 359 937 527
rect 1055 359 1105 527
rect 1223 359 1273 527
rect 1391 359 1441 527
rect 18 215 379 255
rect 119 17 153 111
rect 287 17 321 111
rect 439 177 489 289
rect 523 215 808 255
rect 855 215 1137 257
rect 1182 215 1547 257
rect 439 129 1113 177
rect 1231 17 1265 111
rect 1399 17 1433 111
rect 0 -17 1564 17
<< obsli1 >>
rect 18 459 853 493
rect 18 291 85 459
rect 195 359 245 459
rect 363 359 413 459
rect 531 359 581 459
rect 699 325 853 459
rect 971 325 1021 493
rect 1139 325 1189 493
rect 1307 325 1357 493
rect 1475 325 1525 493
rect 699 291 1525 325
rect 19 145 405 181
rect 19 51 85 145
rect 187 51 253 145
rect 355 95 405 145
rect 1147 145 1533 181
rect 1147 95 1197 145
rect 355 51 757 95
rect 795 51 1197 95
rect 1299 51 1365 145
rect 1467 51 1533 145
<< metal1 >>
rect 0 496 1564 592
rect 0 -48 1564 48
<< labels >>
rlabel locali s 855 215 1137 257 6 A1
port 1 nsew signal input
rlabel locali s 1182 215 1547 257 6 A2
port 2 nsew signal input
rlabel locali s 523 215 808 255 6 B1
port 3 nsew signal input
rlabel locali s 18 215 379 255 6 B2
port 4 nsew signal input
rlabel locali s 615 325 665 425 6 Y
port 5 nsew signal output
rlabel locali s 447 325 497 425 6 Y
port 5 nsew signal output
rlabel locali s 439 177 489 289 6 Y
port 5 nsew signal output
rlabel locali s 439 129 1113 177 6 Y
port 5 nsew signal output
rlabel locali s 279 325 329 425 6 Y
port 5 nsew signal output
rlabel locali s 119 325 161 425 6 Y
port 5 nsew signal output
rlabel locali s 119 289 665 325 6 Y
port 5 nsew signal output
rlabel locali s 1399 17 1433 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1231 17 1265 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 287 17 321 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 119 17 153 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 1564 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1564 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1391 359 1441 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1223 359 1273 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1055 359 1105 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 887 359 937 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 1564 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 1564 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1564 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3448538
string GDS_START 3436546
<< end >>
