magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 644 561
rect 131 435 185 527
rect 17 211 125 323
rect 415 435 480 527
rect 514 299 627 493
rect 131 17 185 109
rect 535 165 627 299
rect 415 17 480 109
rect 514 51 627 165
rect 0 -17 644 17
<< obsli1 >>
rect 17 401 97 493
rect 231 427 285 493
rect 17 357 206 401
rect 159 265 206 357
rect 251 323 285 427
rect 323 401 375 493
rect 323 357 480 401
rect 159 199 217 265
rect 251 211 406 323
rect 440 265 480 357
rect 159 177 206 199
rect 17 143 206 177
rect 17 51 97 143
rect 251 117 285 211
rect 440 199 501 265
rect 440 177 480 199
rect 231 51 285 117
rect 323 143 480 177
rect 323 51 375 143
<< metal1 >>
rect 0 496 644 592
rect 0 -48 644 48
<< labels >>
rlabel locali s 17 211 125 323 6 A
port 1 nsew signal input
rlabel locali s 535 165 627 299 6 X
port 2 nsew signal output
rlabel locali s 514 299 627 493 6 X
port 2 nsew signal output
rlabel locali s 514 51 627 165 6 X
port 2 nsew signal output
rlabel locali s 415 17 480 109 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 131 17 185 109 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 0 -17 644 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 644 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 415 435 480 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 131 435 185 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 0 527 644 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 496 644 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2817530
string GDS_START 2811670
<< end >>
