magic
tech sky130A
magscale 1 2
timestamp 1599588244
<< locali >>
rect 25 256 167 310
rect 201 290 267 356
rect 341 256 407 310
rect 25 222 407 256
rect 1082 430 1138 596
rect 1272 430 1318 596
rect 1082 364 1415 430
rect 889 236 963 310
rect 1273 294 1331 364
rect 1265 260 1331 294
rect 1265 230 1315 260
rect 1065 196 1315 230
rect 1065 70 1131 196
rect 1265 70 1315 196
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 23 424 89 596
rect 129 492 163 596
rect 203 526 269 649
rect 303 492 369 596
rect 129 458 369 492
rect 403 506 469 596
rect 503 540 749 596
rect 789 506 839 596
rect 403 472 839 506
rect 403 424 469 472
rect 23 390 469 424
rect 579 404 659 438
rect 789 412 839 472
rect 23 388 89 390
rect 449 276 545 356
rect 449 242 511 276
rect 449 236 545 242
rect 579 226 613 404
rect 885 378 951 572
rect 693 360 951 378
rect 992 364 1042 649
rect 1172 464 1238 649
rect 1352 464 1418 649
rect 647 344 951 360
rect 647 294 727 344
rect 773 276 839 302
rect 773 242 799 276
rect 833 242 839 276
rect 773 236 839 242
rect 997 264 1231 330
rect 579 202 654 226
rect 997 202 1031 264
rect 579 188 1031 202
rect 23 168 1031 188
rect 23 154 654 168
rect 23 70 89 154
rect 123 17 189 120
rect 223 70 440 154
rect 474 17 545 120
rect 579 70 654 154
rect 688 68 913 134
rect 965 17 1031 134
rect 1165 17 1231 162
rect 1351 17 1417 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 511 242 545 276
rect 799 242 833 276
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 683 1440 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 0 617 1440 649
rect 0 616 50 617
rect 499 276 557 282
rect 499 242 511 276
rect 545 273 557 276
rect 787 276 845 282
rect 787 273 799 276
rect 545 245 799 273
rect 545 242 557 245
rect 499 236 557 242
rect 787 242 799 245
rect 833 242 845 276
rect 787 236 845 242
rect 0 49 50 50
rect 0 17 1440 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -49 1440 -17
<< labels >>
rlabel locali s 201 290 267 356 6 A
port 1 nsew signal input
rlabel locali s 341 256 407 310 6 B
port 2 nsew signal input
rlabel locali s 25 256 167 310 6 B
port 2 nsew signal input
rlabel locali s 25 222 407 256 6 B
port 2 nsew signal input
rlabel metal1 s 787 273 845 282 6 C
port 3 nsew signal input
rlabel metal1 s 787 236 845 245 6 C
port 3 nsew signal input
rlabel metal1 s 499 273 557 282 6 C
port 3 nsew signal input
rlabel metal1 s 499 245 845 273 6 C
port 3 nsew signal input
rlabel metal1 s 499 236 557 245 6 C
port 3 nsew signal input
rlabel locali s 889 236 963 310 6 D_N
port 4 nsew signal input
rlabel locali s 1273 294 1331 364 6 X
port 5 nsew signal output
rlabel locali s 1272 430 1318 596 6 X
port 5 nsew signal output
rlabel locali s 1265 260 1331 294 6 X
port 5 nsew signal output
rlabel locali s 1265 230 1315 260 6 X
port 5 nsew signal output
rlabel locali s 1265 70 1315 196 6 X
port 5 nsew signal output
rlabel locali s 1082 430 1138 596 6 X
port 5 nsew signal output
rlabel locali s 1082 364 1415 430 6 X
port 5 nsew signal output
rlabel locali s 1065 196 1315 230 6 X
port 5 nsew signal output
rlabel locali s 1065 70 1131 196 6 X
port 5 nsew signal output
rlabel metal1 s 0 -49 1440 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 7 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 617 1440 715 6 VPWR
port 9 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1440 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 888762
string GDS_START 876798
<< end >>
