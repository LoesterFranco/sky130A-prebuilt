magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 85 290 161 356
rect 195 290 258 356
rect 1509 426 1575 596
rect 1709 426 1775 596
rect 1509 394 1775 426
rect 1509 392 1895 394
rect 1709 360 1895 392
rect 1264 224 1511 290
rect 1849 226 1895 360
rect 1587 192 1895 226
rect 1587 72 1625 192
rect 1759 160 1895 192
rect 1759 72 1797 160
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 17 390 95 566
rect 129 390 195 649
rect 451 588 517 649
rect 229 554 326 566
rect 229 520 840 554
rect 918 526 1064 649
rect 229 390 326 520
rect 17 250 51 390
rect 292 350 326 390
rect 360 418 441 486
rect 636 452 740 486
rect 360 384 672 418
rect 292 284 373 350
rect 292 250 326 284
rect 407 250 441 384
rect 17 166 89 250
rect 227 200 326 250
rect 360 200 441 250
rect 498 166 564 334
rect 606 304 672 384
rect 706 372 740 452
rect 774 406 840 520
rect 1098 472 1164 592
rect 888 406 1164 472
rect 1198 416 1264 649
rect 706 338 1044 372
rect 606 238 852 304
rect 963 224 1044 338
rect 1098 358 1164 406
rect 1298 358 1364 592
rect 1409 416 1475 649
rect 1609 460 1675 649
rect 1809 428 1875 649
rect 1098 326 1579 358
rect 1098 324 1815 326
rect 963 204 997 224
rect 17 132 564 166
rect 748 170 997 204
rect 125 17 191 98
rect 462 17 625 98
rect 748 80 814 170
rect 919 17 985 136
rect 1031 85 1097 190
rect 1133 119 1167 324
rect 1545 260 1815 324
rect 1203 154 1441 190
rect 1203 85 1253 154
rect 1031 51 1253 85
rect 1289 17 1355 120
rect 1389 71 1441 154
rect 1487 17 1553 190
rect 1659 17 1725 158
rect 1831 17 1897 126
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
<< metal1 >>
rect 0 683 1920 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 0 617 1920 649
rect 0 17 1920 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
rect 0 -49 1920 -17
<< labels >>
rlabel locali s 85 290 161 356 6 D
port 1 nsew signal input
rlabel locali s 1849 226 1895 360 6 Q
port 2 nsew signal output
rlabel locali s 1759 160 1895 192 6 Q
port 2 nsew signal output
rlabel locali s 1759 72 1797 160 6 Q
port 2 nsew signal output
rlabel locali s 1709 426 1775 596 6 Q
port 2 nsew signal output
rlabel locali s 1709 360 1895 392 6 Q
port 2 nsew signal output
rlabel locali s 1587 192 1895 226 6 Q
port 2 nsew signal output
rlabel locali s 1587 72 1625 192 6 Q
port 2 nsew signal output
rlabel locali s 1509 426 1575 596 6 Q
port 2 nsew signal output
rlabel locali s 1509 394 1775 426 6 Q
port 2 nsew signal output
rlabel locali s 1509 392 1895 394 6 Q
port 2 nsew signal output
rlabel locali s 1264 224 1511 290 6 RESET_B
port 3 nsew signal input
rlabel locali s 195 290 258 356 6 GATE_N
port 4 nsew clock input
rlabel metal1 s 0 -49 1920 49 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1920 715 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1920 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3020568
string GDS_START 3006388
<< end >>
