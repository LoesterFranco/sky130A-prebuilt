magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1196 561
rect 114 427 164 527
rect 554 427 604 527
rect 722 427 783 527
rect 1005 325 1055 425
rect 141 289 376 323
rect 141 255 175 289
rect 342 255 376 289
rect 109 215 175 255
rect 209 215 308 255
rect 342 215 646 255
rect 684 215 818 255
rect 1005 283 1179 325
rect 1097 181 1179 283
rect 38 17 72 111
rect 206 17 240 111
rect 374 17 408 111
rect 562 17 596 111
rect 725 145 1179 181
rect 725 129 791 145
rect 997 129 1063 145
rect 929 17 963 111
rect 1097 17 1131 111
rect 0 -17 1196 17
<< obsli1 >>
rect 24 459 80 493
rect 24 427 29 459
rect 63 427 80 459
rect 198 459 416 493
rect 198 427 213 459
rect 247 427 248 459
rect 366 427 416 459
rect 457 425 520 493
rect 282 391 332 425
rect 478 391 520 425
rect 638 391 688 493
rect 817 459 1139 493
rect 817 391 971 459
rect 24 357 444 391
rect 478 357 971 391
rect 24 181 58 357
rect 410 323 444 357
rect 1089 359 1139 459
rect 410 289 957 323
rect 923 249 957 289
rect 923 215 1055 249
rect 24 145 340 181
rect 106 51 172 145
rect 274 51 340 145
rect 462 145 680 181
rect 462 51 528 145
rect 630 95 680 145
rect 630 51 876 95
<< obsli1c >>
rect 29 425 63 459
rect 213 425 247 459
<< metal1 >>
rect 0 496 1196 592
rect 201 252 259 261
rect 753 252 811 261
rect 201 224 811 252
rect 201 215 259 224
rect 753 215 811 224
rect 0 -48 1196 48
<< obsm1 >>
rect 17 459 75 465
rect 17 425 29 459
rect 63 456 75 459
rect 201 459 259 465
rect 201 456 213 459
rect 63 428 213 456
rect 63 425 75 428
rect 17 419 75 425
rect 201 425 213 428
rect 247 425 259 459
rect 201 419 259 425
<< labels >>
rlabel locali s 342 255 376 289 6 A
port 1 nsew signal input
rlabel locali s 342 215 646 255 6 A
port 1 nsew signal input
rlabel locali s 141 289 376 323 6 A
port 1 nsew signal input
rlabel locali s 141 255 175 289 6 A
port 1 nsew signal input
rlabel locali s 109 215 175 255 6 A
port 1 nsew signal input
rlabel locali s 209 215 308 255 6 B
port 2 nsew signal input
rlabel locali s 684 215 818 255 6 B
port 2 nsew signal input
rlabel metal1 s 753 252 811 261 6 B
port 2 nsew signal input
rlabel metal1 s 753 215 811 224 6 B
port 2 nsew signal input
rlabel metal1 s 201 252 259 261 6 B
port 2 nsew signal input
rlabel metal1 s 201 224 811 252 6 B
port 2 nsew signal input
rlabel metal1 s 201 215 259 224 6 B
port 2 nsew signal input
rlabel locali s 1097 181 1179 283 6 X
port 3 nsew signal output
rlabel locali s 1005 325 1055 425 6 X
port 3 nsew signal output
rlabel locali s 1005 283 1179 325 6 X
port 3 nsew signal output
rlabel locali s 997 129 1063 145 6 X
port 3 nsew signal output
rlabel locali s 725 145 1179 181 6 X
port 3 nsew signal output
rlabel locali s 725 129 791 145 6 X
port 3 nsew signal output
rlabel locali s 1097 17 1131 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 929 17 963 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 562 17 596 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 374 17 408 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 206 17 240 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 38 17 72 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 1196 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1196 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 722 427 783 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 554 427 604 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 114 427 164 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 1196 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 1196 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 646902
string GDS_START 637824
<< end >>
