magic
tech sky130A
magscale 1 2
timestamp 1604502701
<< nwell >>
rect -38 332 710 704
<< pwell >>
rect 0 0 672 49
<< scpmos >>
rect 120 392 150 592
rect 204 392 234 592
rect 318 392 348 592
rect 440 368 470 592
rect 530 368 560 592
<< nmoslvt >>
rect 84 74 114 202
rect 215 74 245 202
rect 315 74 345 202
rect 458 74 488 222
rect 544 74 574 222
<< ndiff >>
rect 408 202 458 222
rect 27 147 84 202
rect 27 113 39 147
rect 73 113 84 147
rect 27 74 84 113
rect 114 120 215 202
rect 114 86 147 120
rect 181 86 215 120
rect 114 74 215 86
rect 245 148 315 202
rect 245 114 256 148
rect 290 114 315 148
rect 245 74 315 114
rect 345 120 458 202
rect 345 86 377 120
rect 411 86 458 120
rect 345 74 458 86
rect 488 210 544 222
rect 488 176 499 210
rect 533 176 544 210
rect 488 120 544 176
rect 488 86 499 120
rect 533 86 544 120
rect 488 74 544 86
rect 574 131 645 222
rect 574 97 599 131
rect 633 97 645 131
rect 574 74 645 97
<< pdiff >>
rect 61 580 120 592
rect 61 546 73 580
rect 107 546 120 580
rect 61 511 120 546
rect 61 477 73 511
rect 107 477 120 511
rect 61 442 120 477
rect 61 408 73 442
rect 107 408 120 442
rect 61 392 120 408
rect 150 392 204 592
rect 234 392 318 592
rect 348 580 440 592
rect 348 546 361 580
rect 395 546 440 580
rect 348 509 440 546
rect 348 475 361 509
rect 395 475 440 509
rect 348 438 440 475
rect 348 404 361 438
rect 395 404 440 438
rect 348 392 440 404
rect 387 368 440 392
rect 470 580 530 592
rect 470 546 483 580
rect 517 546 530 580
rect 470 497 530 546
rect 470 463 483 497
rect 517 463 530 497
rect 470 414 530 463
rect 470 380 483 414
rect 517 380 530 414
rect 470 368 530 380
rect 560 580 629 592
rect 560 546 583 580
rect 617 546 629 580
rect 560 462 629 546
rect 560 428 583 462
rect 617 428 629 462
rect 560 368 629 428
<< ndiffc >>
rect 39 113 73 147
rect 147 86 181 120
rect 256 114 290 148
rect 377 86 411 120
rect 499 176 533 210
rect 499 86 533 120
rect 599 97 633 131
<< pdiffc >>
rect 73 546 107 580
rect 73 477 107 511
rect 73 408 107 442
rect 361 546 395 580
rect 361 475 395 509
rect 361 404 395 438
rect 483 546 517 580
rect 483 463 517 497
rect 483 380 517 414
rect 583 546 617 580
rect 583 428 617 462
<< poly >>
rect 120 592 150 618
rect 204 592 234 618
rect 318 592 348 618
rect 440 592 470 618
rect 530 592 560 618
rect 120 377 150 392
rect 204 377 234 392
rect 318 377 348 392
rect 117 358 153 377
rect 84 342 153 358
rect 84 308 103 342
rect 137 308 153 342
rect 84 274 153 308
rect 84 240 103 274
rect 137 240 153 274
rect 84 224 153 240
rect 201 360 237 377
rect 201 344 267 360
rect 201 310 217 344
rect 251 310 267 344
rect 201 276 267 310
rect 201 242 217 276
rect 251 242 267 276
rect 201 226 267 242
rect 315 310 351 377
rect 440 353 470 368
rect 530 353 560 368
rect 437 326 473 353
rect 527 326 563 353
rect 429 310 563 326
rect 315 294 381 310
rect 315 260 331 294
rect 365 260 381 294
rect 429 276 445 310
rect 479 276 513 310
rect 547 290 563 310
rect 547 276 574 290
rect 429 260 574 276
rect 315 244 381 260
rect 84 202 114 224
rect 215 202 245 226
rect 315 202 345 244
rect 458 222 488 260
rect 544 222 574 260
rect 84 48 114 74
rect 215 48 245 74
rect 315 48 345 74
rect 458 48 488 74
rect 544 48 574 74
<< polycont >>
rect 103 308 137 342
rect 103 240 137 274
rect 217 310 251 344
rect 217 242 251 276
rect 331 260 365 294
rect 445 276 479 310
rect 513 276 547 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 57 580 123 596
rect 57 546 73 580
rect 107 546 123 580
rect 345 580 411 649
rect 57 511 123 546
rect 57 477 73 511
rect 107 477 123 511
rect 57 442 123 477
rect 57 426 73 442
rect 19 408 73 426
rect 107 408 123 442
rect 19 392 123 408
rect 19 190 53 392
rect 87 342 167 358
rect 87 308 103 342
rect 137 308 167 342
rect 87 274 167 308
rect 87 240 103 274
rect 137 240 167 274
rect 87 224 167 240
rect 201 344 267 578
rect 345 546 361 580
rect 395 546 411 580
rect 345 509 411 546
rect 345 475 361 509
rect 395 475 411 509
rect 345 438 411 475
rect 345 404 361 438
rect 395 404 411 438
rect 345 388 411 404
rect 467 580 533 596
rect 467 546 483 580
rect 517 546 533 580
rect 467 497 533 546
rect 467 463 483 497
rect 517 463 533 497
rect 467 414 533 463
rect 567 580 633 649
rect 567 546 583 580
rect 617 546 633 580
rect 567 462 633 546
rect 567 428 583 462
rect 617 428 633 462
rect 467 380 483 414
rect 517 394 533 414
rect 517 380 647 394
rect 467 360 647 380
rect 201 310 217 344
rect 251 310 267 344
rect 415 310 563 326
rect 201 276 267 310
rect 201 242 217 276
rect 251 242 267 276
rect 201 226 267 242
rect 313 294 381 310
rect 313 260 331 294
rect 365 260 381 294
rect 313 236 381 260
rect 415 276 445 310
rect 479 276 513 310
rect 547 276 563 310
rect 415 260 563 276
rect 415 192 449 260
rect 601 226 647 360
rect 240 190 449 192
rect 19 158 449 190
rect 483 210 647 226
rect 483 176 499 210
rect 533 192 647 210
rect 533 176 549 192
rect 19 156 306 158
rect 19 147 89 156
rect 19 113 39 147
rect 73 113 89 147
rect 240 148 306 156
rect 19 70 89 113
rect 123 86 147 120
rect 181 86 206 120
rect 123 17 206 86
rect 240 114 256 148
rect 290 114 306 148
rect 483 120 549 176
rect 240 70 306 114
rect 340 86 377 120
rect 411 86 449 120
rect 340 17 449 86
rect 483 86 499 120
rect 533 86 549 120
rect 483 70 549 86
rect 583 131 649 158
rect 583 97 599 131
rect 633 97 649 131
rect 583 17 649 97
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel comment s 0 0 0 0 4 or3_2
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 607 242 641 276 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 127 242 161 276 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 319 242 353 276 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 223 390 257 424 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 223 464 257 498 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 223 538 257 572 0 FreeSans 340 0 0 0 B
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 672 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 885666
string GDS_START 879174
<< end >>
