magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 460 561
rect 175 371 241 527
rect 331 370 443 493
rect 20 145 65 265
rect 192 213 265 265
rect 407 179 443 370
rect 171 17 213 179
rect 247 145 443 179
rect 247 51 313 145
rect 347 17 424 111
rect 0 -17 460 17
<< obsli1 >>
rect 83 336 135 381
rect 83 302 341 336
rect 99 109 135 302
rect 307 249 341 302
rect 307 215 373 249
rect 66 74 135 109
<< metal1 >>
rect 0 496 460 592
rect 0 -48 460 48
<< labels >>
rlabel locali s 192 213 265 265 6 A
port 1 nsew signal input
rlabel locali s 20 145 65 265 6 B_N
port 2 nsew signal input
rlabel locali s 407 179 443 370 6 Y
port 3 nsew signal output
rlabel locali s 331 370 443 493 6 Y
port 3 nsew signal output
rlabel locali s 247 145 443 179 6 Y
port 3 nsew signal output
rlabel locali s 247 51 313 145 6 Y
port 3 nsew signal output
rlabel locali s 347 17 424 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 171 17 213 179 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 460 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 460 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 175 371 241 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 460 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 460 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 460 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1953828
string GDS_START 1949574
<< end >>
