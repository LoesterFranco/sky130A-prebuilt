magic
tech sky130A
magscale 1 2
timestamp 1604502697
<< nwell >>
rect -38 261 1694 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 95 47 125 177
rect 189 47 219 177
rect 283 47 313 177
rect 367 47 397 177
rect 461 47 491 177
rect 555 47 585 177
rect 659 47 689 177
rect 753 47 783 177
rect 847 47 877 177
rect 941 47 971 177
rect 1045 47 1075 177
rect 1129 47 1159 177
rect 1223 47 1253 177
rect 1317 47 1347 177
rect 1421 47 1451 177
rect 1515 47 1545 177
<< pmoshvt >>
rect 87 297 123 497
rect 181 297 217 497
rect 275 297 311 497
rect 369 297 405 497
rect 463 297 499 497
rect 557 297 593 497
rect 651 297 687 497
rect 745 297 781 497
rect 849 297 885 497
rect 943 297 979 497
rect 1037 297 1073 497
rect 1131 297 1167 497
rect 1225 297 1261 497
rect 1319 297 1355 497
rect 1413 297 1449 497
rect 1507 297 1543 497
<< ndiff >>
rect 33 163 95 177
rect 33 129 41 163
rect 75 129 95 163
rect 33 95 95 129
rect 33 61 41 95
rect 75 61 95 95
rect 33 47 95 61
rect 125 95 189 177
rect 125 61 135 95
rect 169 61 189 95
rect 125 47 189 61
rect 219 163 283 177
rect 219 129 229 163
rect 263 129 283 163
rect 219 95 283 129
rect 219 61 229 95
rect 263 61 283 95
rect 219 47 283 61
rect 313 95 367 177
rect 313 61 323 95
rect 357 61 367 95
rect 313 47 367 61
rect 397 163 461 177
rect 397 129 417 163
rect 451 129 461 163
rect 397 95 461 129
rect 397 61 417 95
rect 451 61 461 95
rect 397 47 461 61
rect 491 95 555 177
rect 491 61 511 95
rect 545 61 555 95
rect 491 47 555 61
rect 585 163 659 177
rect 585 129 605 163
rect 639 129 659 163
rect 585 95 659 129
rect 585 61 605 95
rect 639 61 659 95
rect 585 47 659 61
rect 689 95 753 177
rect 689 61 699 95
rect 733 61 753 95
rect 689 47 753 61
rect 783 163 847 177
rect 783 129 793 163
rect 827 129 847 163
rect 783 95 847 129
rect 783 61 793 95
rect 827 61 847 95
rect 783 47 847 61
rect 877 163 941 177
rect 877 129 897 163
rect 931 129 941 163
rect 877 47 941 129
rect 971 95 1045 177
rect 971 61 991 95
rect 1025 61 1045 95
rect 971 47 1045 61
rect 1075 163 1129 177
rect 1075 129 1085 163
rect 1119 129 1129 163
rect 1075 47 1129 129
rect 1159 95 1223 177
rect 1159 61 1179 95
rect 1213 61 1223 95
rect 1159 47 1223 61
rect 1253 163 1317 177
rect 1253 129 1273 163
rect 1307 129 1317 163
rect 1253 47 1317 129
rect 1347 95 1421 177
rect 1347 61 1367 95
rect 1401 61 1421 95
rect 1347 47 1421 61
rect 1451 163 1515 177
rect 1451 129 1461 163
rect 1495 129 1515 163
rect 1451 47 1515 129
rect 1545 95 1597 177
rect 1545 61 1555 95
rect 1589 61 1597 95
rect 1545 47 1597 61
<< pdiff >>
rect 27 477 87 497
rect 27 443 41 477
rect 75 443 87 477
rect 27 409 87 443
rect 27 375 41 409
rect 75 375 87 409
rect 27 341 87 375
rect 27 307 41 341
rect 75 307 87 341
rect 27 297 87 307
rect 123 477 181 497
rect 123 443 135 477
rect 169 443 181 477
rect 123 409 181 443
rect 123 375 135 409
rect 169 375 181 409
rect 123 341 181 375
rect 123 307 135 341
rect 169 307 181 341
rect 123 297 181 307
rect 217 477 275 497
rect 217 443 229 477
rect 263 443 275 477
rect 217 297 275 443
rect 311 477 369 497
rect 311 443 323 477
rect 357 443 369 477
rect 311 409 369 443
rect 311 375 323 409
rect 357 375 369 409
rect 311 297 369 375
rect 405 409 463 497
rect 405 375 417 409
rect 451 375 463 409
rect 405 297 463 375
rect 499 477 557 497
rect 499 443 511 477
rect 545 443 557 477
rect 499 297 557 443
rect 593 409 651 497
rect 593 375 605 409
rect 639 375 651 409
rect 593 297 651 375
rect 687 477 745 497
rect 687 443 699 477
rect 733 443 745 477
rect 687 297 745 443
rect 781 477 849 497
rect 781 443 801 477
rect 835 443 849 477
rect 781 297 849 443
rect 885 477 943 497
rect 885 443 897 477
rect 931 443 943 477
rect 885 297 943 443
rect 979 477 1037 497
rect 979 443 991 477
rect 1025 443 1037 477
rect 979 297 1037 443
rect 1073 477 1131 497
rect 1073 443 1085 477
rect 1119 443 1131 477
rect 1073 409 1131 443
rect 1073 375 1085 409
rect 1119 375 1131 409
rect 1073 297 1131 375
rect 1167 409 1225 497
rect 1167 375 1179 409
rect 1213 375 1225 409
rect 1167 297 1225 375
rect 1261 477 1319 497
rect 1261 443 1273 477
rect 1307 443 1319 477
rect 1261 297 1319 443
rect 1355 409 1413 497
rect 1355 375 1367 409
rect 1401 375 1413 409
rect 1355 297 1413 375
rect 1449 477 1507 497
rect 1449 443 1461 477
rect 1495 443 1507 477
rect 1449 297 1507 443
rect 1543 477 1597 497
rect 1543 443 1555 477
rect 1589 443 1597 477
rect 1543 297 1597 443
<< ndiffc >>
rect 41 129 75 163
rect 41 61 75 95
rect 135 61 169 95
rect 229 129 263 163
rect 229 61 263 95
rect 323 61 357 95
rect 417 129 451 163
rect 417 61 451 95
rect 511 61 545 95
rect 605 129 639 163
rect 605 61 639 95
rect 699 61 733 95
rect 793 129 827 163
rect 793 61 827 95
rect 897 129 931 163
rect 991 61 1025 95
rect 1085 129 1119 163
rect 1179 61 1213 95
rect 1273 129 1307 163
rect 1367 61 1401 95
rect 1461 129 1495 163
rect 1555 61 1589 95
<< pdiffc >>
rect 41 443 75 477
rect 41 375 75 409
rect 41 307 75 341
rect 135 443 169 477
rect 135 375 169 409
rect 135 307 169 341
rect 229 443 263 477
rect 323 443 357 477
rect 323 375 357 409
rect 417 375 451 409
rect 511 443 545 477
rect 605 375 639 409
rect 699 443 733 477
rect 801 443 835 477
rect 897 443 931 477
rect 991 443 1025 477
rect 1085 443 1119 477
rect 1085 375 1119 409
rect 1179 375 1213 409
rect 1273 443 1307 477
rect 1367 375 1401 409
rect 1461 443 1495 477
rect 1555 443 1589 477
<< poly >>
rect 87 497 123 523
rect 181 497 217 523
rect 275 497 311 523
rect 369 497 405 523
rect 463 497 499 523
rect 557 497 593 523
rect 651 497 687 523
rect 745 497 781 523
rect 849 497 885 523
rect 943 497 979 523
rect 1037 497 1073 523
rect 1131 497 1167 523
rect 1225 497 1261 523
rect 1319 497 1355 523
rect 1413 497 1449 523
rect 1507 497 1543 523
rect 87 282 123 297
rect 181 282 217 297
rect 275 282 311 297
rect 369 282 405 297
rect 463 282 499 297
rect 557 282 593 297
rect 651 282 687 297
rect 745 282 781 297
rect 849 282 885 297
rect 943 282 979 297
rect 1037 282 1073 297
rect 1131 282 1167 297
rect 1225 282 1261 297
rect 1319 282 1355 297
rect 1413 282 1449 297
rect 1507 282 1543 297
rect 85 265 125 282
rect 179 265 219 282
rect 273 265 313 282
rect 76 249 313 265
rect 76 215 97 249
rect 131 215 175 249
rect 209 215 253 249
rect 287 215 313 249
rect 76 199 313 215
rect 95 177 125 199
rect 189 177 219 199
rect 283 177 313 199
rect 367 265 407 282
rect 461 265 501 282
rect 555 265 595 282
rect 649 265 689 282
rect 743 265 783 282
rect 847 265 887 282
rect 941 265 981 282
rect 1035 265 1075 282
rect 1129 265 1169 282
rect 1223 265 1263 282
rect 1317 265 1357 282
rect 1411 265 1451 282
rect 1505 265 1545 282
rect 367 249 689 265
rect 367 215 395 249
rect 429 215 473 249
rect 507 215 551 249
rect 585 215 629 249
rect 663 215 689 249
rect 367 199 689 215
rect 731 249 795 265
rect 731 215 741 249
rect 775 215 795 249
rect 731 199 795 215
rect 847 249 1087 265
rect 847 215 949 249
rect 983 215 1027 249
rect 1061 215 1087 249
rect 847 199 1087 215
rect 1129 249 1451 265
rect 1129 215 1148 249
rect 1182 215 1226 249
rect 1260 215 1304 249
rect 1338 215 1382 249
rect 1416 215 1451 249
rect 1129 199 1451 215
rect 1493 249 1563 265
rect 1493 215 1503 249
rect 1537 215 1563 249
rect 1493 199 1563 215
rect 367 177 397 199
rect 461 177 491 199
rect 555 177 585 199
rect 659 177 689 199
rect 753 177 783 199
rect 847 177 877 199
rect 941 177 971 199
rect 1045 177 1075 199
rect 1129 177 1159 199
rect 1223 177 1253 199
rect 1317 177 1347 199
rect 1421 177 1451 199
rect 1515 177 1545 199
rect 95 21 125 47
rect 189 21 219 47
rect 283 21 313 47
rect 367 21 397 47
rect 461 21 491 47
rect 555 21 585 47
rect 659 21 689 47
rect 753 21 783 47
rect 847 21 877 47
rect 941 21 971 47
rect 1045 21 1075 47
rect 1129 21 1159 47
rect 1223 21 1253 47
rect 1317 21 1347 47
rect 1421 21 1451 47
rect 1515 21 1545 47
<< polycont >>
rect 97 215 131 249
rect 175 215 209 249
rect 253 215 287 249
rect 395 215 429 249
rect 473 215 507 249
rect 551 215 585 249
rect 629 215 663 249
rect 741 215 775 249
rect 949 215 983 249
rect 1027 215 1061 249
rect 1148 215 1182 249
rect 1226 215 1260 249
rect 1304 215 1338 249
rect 1382 215 1416 249
rect 1503 215 1537 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 33 477 83 527
rect 33 443 41 477
rect 75 443 83 477
rect 33 409 83 443
rect 33 375 41 409
rect 75 375 83 409
rect 33 341 83 375
rect 33 307 41 341
rect 75 307 83 341
rect 33 289 83 307
rect 127 477 177 493
rect 127 443 135 477
rect 169 443 177 477
rect 127 409 177 443
rect 221 477 271 527
rect 221 443 229 477
rect 263 443 271 477
rect 221 425 271 443
rect 315 477 749 493
rect 315 443 323 477
rect 357 459 511 477
rect 127 375 135 409
rect 169 391 177 409
rect 315 409 357 443
rect 503 443 511 459
rect 545 459 699 477
rect 545 443 553 459
rect 503 425 553 443
rect 691 443 699 459
rect 733 443 749 477
rect 691 425 749 443
rect 793 477 837 527
rect 793 443 801 477
rect 835 443 837 477
rect 793 425 837 443
rect 871 477 942 493
rect 871 443 897 477
rect 931 443 942 477
rect 871 425 942 443
rect 985 477 1033 527
rect 985 443 991 477
rect 1025 443 1033 477
rect 985 425 1033 443
rect 1077 477 1503 493
rect 1077 443 1085 477
rect 1119 459 1273 477
rect 1119 443 1127 459
rect 315 391 323 409
rect 169 375 323 391
rect 127 357 357 375
rect 391 409 459 425
rect 391 375 417 409
rect 451 391 459 409
rect 597 409 647 425
rect 597 391 605 409
rect 451 375 605 391
rect 639 391 647 409
rect 908 391 942 425
rect 1077 409 1127 443
rect 1265 443 1273 459
rect 1307 459 1461 477
rect 1307 443 1315 459
rect 1265 425 1315 443
rect 1453 443 1461 459
rect 1495 443 1503 477
rect 1453 427 1503 443
rect 1547 477 1603 527
rect 1547 443 1555 477
rect 1589 443 1603 477
rect 1547 425 1603 443
rect 1077 391 1085 409
rect 639 375 874 391
rect 391 357 874 375
rect 908 375 1085 391
rect 1119 375 1127 409
rect 908 357 1127 375
rect 1171 409 1221 425
rect 1171 375 1179 409
rect 1213 391 1221 409
rect 1359 409 1409 425
rect 1359 391 1367 409
rect 1213 375 1367 391
rect 1401 391 1409 409
rect 1401 375 1634 391
rect 1171 357 1634 375
rect 127 341 177 357
rect 127 307 135 341
rect 169 307 177 341
rect 840 323 874 357
rect 127 289 177 307
rect 250 289 806 323
rect 840 289 915 323
rect 250 255 313 289
rect 17 249 313 255
rect 17 215 97 249
rect 131 215 175 249
rect 209 215 253 249
rect 287 215 313 249
rect 367 249 689 255
rect 367 215 395 249
rect 429 215 473 249
rect 507 215 551 249
rect 585 215 629 249
rect 663 215 689 249
rect 725 249 806 289
rect 725 215 741 249
rect 775 215 806 249
rect 25 163 837 181
rect 25 129 41 163
rect 75 145 229 163
rect 75 129 91 145
rect 25 95 91 129
rect 203 129 229 145
rect 263 147 417 163
rect 263 129 279 147
rect 25 61 41 95
rect 75 61 91 95
rect 25 51 91 61
rect 135 95 169 111
rect 135 17 169 61
rect 203 95 279 129
rect 391 129 417 147
rect 451 145 605 163
rect 451 129 467 145
rect 203 61 229 95
rect 263 61 279 95
rect 203 51 279 61
rect 323 95 357 111
rect 323 17 357 61
rect 391 95 467 129
rect 579 129 605 145
rect 639 147 793 163
rect 639 129 655 147
rect 391 61 417 95
rect 451 61 467 95
rect 391 51 467 61
rect 511 95 545 111
rect 511 17 545 61
rect 579 95 655 129
rect 767 129 793 147
rect 827 129 837 163
rect 871 164 915 289
rect 949 289 1547 323
rect 949 249 1098 289
rect 983 215 1027 249
rect 1061 215 1098 249
rect 1132 249 1432 255
rect 1132 215 1148 249
rect 1182 215 1226 249
rect 1260 215 1304 249
rect 1338 215 1382 249
rect 1416 215 1432 249
rect 1493 249 1547 289
rect 1493 215 1503 249
rect 1537 215 1547 249
rect 949 199 1098 215
rect 1493 199 1547 215
rect 1581 164 1634 357
rect 871 163 1634 164
rect 871 129 897 163
rect 931 129 1085 163
rect 1119 129 1273 163
rect 1307 129 1461 163
rect 1495 129 1634 163
rect 579 61 605 95
rect 639 61 655 95
rect 579 51 655 61
rect 699 95 733 111
rect 699 17 733 61
rect 767 95 837 129
rect 767 61 793 95
rect 827 61 991 95
rect 1025 61 1179 95
rect 1213 61 1367 95
rect 1401 61 1555 95
rect 1589 61 1609 95
rect 767 51 1609 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
<< metal1 >>
rect 0 561 1656 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 0 496 1656 527
rect 0 17 1656 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
rect 0 -48 1656 -17
<< labels >>
flabel corelocali s 230 238 230 238 0 FreeSans 400 0 0 0 A1
port 1 nsew
flabel corelocali s 641 357 675 391 0 FreeSans 400 0 0 0 Y
port 9 nsew
flabel corelocali s 506 238 506 238 0 FreeSans 400 0 0 0 A2
port 2 nsew
flabel corelocali s 966 238 966 238 0 FreeSans 400 180 0 0 B1
port 3 nsew
flabel corelocali s 1242 238 1242 238 0 FreeSans 400 180 0 0 B2
port 4 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
rlabel comment s 0 0 0 0 4 o22ai_4
<< properties >>
string FIXED_BBOX 0 0 1656 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 950120
string GDS_START 938732
<< end >>
