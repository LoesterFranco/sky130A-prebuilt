magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 828 561
rect 117 375 183 527
rect 17 199 105 265
rect 217 323 251 493
rect 294 359 344 527
rect 481 323 530 425
rect 217 289 530 323
rect 641 367 707 527
rect 305 181 356 289
rect 390 215 618 255
rect 652 215 811 255
rect 36 17 70 165
rect 305 129 371 181
rect 489 17 523 111
rect 657 17 691 111
rect 0 -17 828 17
<< obsli1 >>
rect 36 333 70 383
rect 36 299 173 333
rect 139 249 173 299
rect 391 459 607 493
rect 391 359 447 459
rect 573 333 607 459
rect 741 333 796 493
rect 573 291 796 333
rect 139 215 267 249
rect 139 165 173 215
rect 120 89 173 165
rect 215 95 271 181
rect 405 145 796 181
rect 405 95 455 145
rect 215 51 455 95
rect 557 51 623 145
rect 725 53 796 145
<< metal1 >>
rect 0 496 828 592
rect 0 -48 828 48
<< labels >>
rlabel locali s 652 215 811 255 6 A1
port 1 nsew signal input
rlabel locali s 390 215 618 255 6 A2
port 2 nsew signal input
rlabel locali s 17 199 105 265 6 B1_N
port 3 nsew signal input
rlabel locali s 481 323 530 425 6 Y
port 4 nsew signal output
rlabel locali s 305 181 356 289 6 Y
port 4 nsew signal output
rlabel locali s 305 129 371 181 6 Y
port 4 nsew signal output
rlabel locali s 217 323 251 493 6 Y
port 4 nsew signal output
rlabel locali s 217 289 530 323 6 Y
port 4 nsew signal output
rlabel locali s 657 17 691 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 489 17 523 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 36 17 70 165 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 828 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 828 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 641 367 707 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 294 359 344 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 117 375 183 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 828 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 828 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1401524
string GDS_START 1394468
<< end >>
