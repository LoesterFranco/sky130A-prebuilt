magic
tech sky130A
magscale 1 2
timestamp 1599588201
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 268 47 298 131
rect 354 47 384 131
rect 440 47 470 131
rect 526 47 556 131
rect 612 47 642 131
rect 698 47 728 131
rect 784 47 814 131
rect 870 47 900 131
<< pmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 248 297 278 497
rect 332 297 362 497
rect 416 297 446 497
rect 500 297 530 497
rect 584 297 614 497
rect 668 297 698 497
rect 752 297 782 497
rect 836 297 866 497
rect 920 297 950 497
rect 1004 297 1034 497
<< ndiff >>
rect 215 95 268 131
rect 215 61 223 95
rect 257 61 268 95
rect 215 47 268 61
rect 298 106 354 131
rect 298 72 309 106
rect 343 72 354 106
rect 298 47 354 72
rect 384 95 440 131
rect 384 61 395 95
rect 429 61 440 95
rect 384 47 440 61
rect 470 106 526 131
rect 470 72 481 106
rect 515 72 526 106
rect 470 47 526 72
rect 556 95 612 131
rect 556 61 567 95
rect 601 61 612 95
rect 556 47 612 61
rect 642 106 698 131
rect 642 72 653 106
rect 687 72 698 106
rect 642 47 698 72
rect 728 95 784 131
rect 728 61 739 95
rect 773 61 784 95
rect 728 47 784 61
rect 814 106 870 131
rect 814 72 825 106
rect 859 72 870 106
rect 814 47 870 72
rect 900 95 953 131
rect 900 61 911 95
rect 945 61 953 95
rect 900 47 953 61
<< pdiff >>
rect 27 478 79 497
rect 27 444 35 478
rect 69 444 79 478
rect 27 410 79 444
rect 27 376 35 410
rect 69 376 79 410
rect 27 297 79 376
rect 109 471 163 497
rect 109 437 119 471
rect 153 437 163 471
rect 109 403 163 437
rect 109 369 119 403
rect 153 369 163 403
rect 109 297 163 369
rect 193 478 248 497
rect 193 444 204 478
rect 238 444 248 478
rect 193 410 248 444
rect 193 376 204 410
rect 238 376 248 410
rect 193 297 248 376
rect 278 471 332 497
rect 278 437 288 471
rect 322 437 332 471
rect 278 383 332 437
rect 278 349 288 383
rect 322 349 332 383
rect 278 297 332 349
rect 362 478 416 497
rect 362 444 372 478
rect 406 444 416 478
rect 362 410 416 444
rect 362 376 372 410
rect 406 376 416 410
rect 362 297 416 376
rect 446 471 500 497
rect 446 437 456 471
rect 490 437 500 471
rect 446 383 500 437
rect 446 349 456 383
rect 490 349 500 383
rect 446 297 500 349
rect 530 478 584 497
rect 530 444 540 478
rect 574 444 584 478
rect 530 410 584 444
rect 530 376 540 410
rect 574 376 584 410
rect 530 297 584 376
rect 614 471 668 497
rect 614 437 624 471
rect 658 437 668 471
rect 614 383 668 437
rect 614 349 624 383
rect 658 349 668 383
rect 614 297 668 349
rect 698 478 752 497
rect 698 444 708 478
rect 742 444 752 478
rect 698 410 752 444
rect 698 376 708 410
rect 742 376 752 410
rect 698 297 752 376
rect 782 471 836 497
rect 782 437 792 471
rect 826 437 836 471
rect 782 383 836 437
rect 782 349 792 383
rect 826 349 836 383
rect 782 297 836 349
rect 866 478 920 497
rect 866 444 876 478
rect 910 444 920 478
rect 866 410 920 444
rect 866 376 876 410
rect 910 376 920 410
rect 866 297 920 376
rect 950 471 1004 497
rect 950 437 960 471
rect 994 437 1004 471
rect 950 383 1004 437
rect 950 349 960 383
rect 994 349 1004 383
rect 950 297 1004 349
rect 1034 478 1086 497
rect 1034 444 1044 478
rect 1078 444 1086 478
rect 1034 410 1086 444
rect 1034 376 1044 410
rect 1078 376 1086 410
rect 1034 297 1086 376
<< ndiffc >>
rect 223 61 257 95
rect 309 72 343 106
rect 395 61 429 95
rect 481 72 515 106
rect 567 61 601 95
rect 653 72 687 106
rect 739 61 773 95
rect 825 72 859 106
rect 911 61 945 95
<< pdiffc >>
rect 35 444 69 478
rect 35 376 69 410
rect 119 437 153 471
rect 119 369 153 403
rect 204 444 238 478
rect 204 376 238 410
rect 288 437 322 471
rect 288 349 322 383
rect 372 444 406 478
rect 372 376 406 410
rect 456 437 490 471
rect 456 349 490 383
rect 540 444 574 478
rect 540 376 574 410
rect 624 437 658 471
rect 624 349 658 383
rect 708 444 742 478
rect 708 376 742 410
rect 792 437 826 471
rect 792 349 826 383
rect 876 444 910 478
rect 876 376 910 410
rect 960 437 994 471
rect 960 349 994 383
rect 1044 444 1078 478
rect 1044 376 1078 410
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 248 497 278 523
rect 332 497 362 523
rect 416 497 446 523
rect 500 497 530 523
rect 584 497 614 523
rect 668 497 698 523
rect 752 497 782 523
rect 836 497 866 523
rect 920 497 950 523
rect 1004 497 1034 523
rect 79 277 109 297
rect 163 277 193 297
rect 248 277 278 297
rect 332 277 362 297
rect 416 277 446 297
rect 500 277 530 297
rect 584 277 614 297
rect 668 277 698 297
rect 752 277 782 297
rect 836 277 866 297
rect 920 277 950 297
rect 1004 277 1034 297
rect 79 249 1034 277
rect 79 215 107 249
rect 141 215 175 249
rect 209 215 243 249
rect 277 215 311 249
rect 345 215 379 249
rect 413 215 447 249
rect 481 215 515 249
rect 549 215 583 249
rect 617 215 651 249
rect 685 215 719 249
rect 753 215 787 249
rect 821 215 855 249
rect 889 215 923 249
rect 957 215 1034 249
rect 79 162 1034 215
rect 268 131 298 162
rect 354 131 384 162
rect 440 131 470 162
rect 526 131 556 162
rect 612 131 642 162
rect 698 131 728 162
rect 784 131 814 162
rect 870 131 900 162
rect 268 21 298 47
rect 354 21 384 47
rect 440 21 470 47
rect 526 21 556 47
rect 612 21 642 47
rect 698 21 728 47
rect 784 21 814 47
rect 870 21 900 47
<< polycont >>
rect 107 215 141 249
rect 175 215 209 249
rect 243 215 277 249
rect 311 215 345 249
rect 379 215 413 249
rect 447 215 481 249
rect 515 215 549 249
rect 583 215 617 249
rect 651 215 685 249
rect 719 215 753 249
rect 787 215 821 249
rect 855 215 889 249
rect 923 215 957 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 19 478 85 493
rect 19 459 35 478
rect 19 425 26 459
rect 69 444 85 478
rect 60 425 85 444
rect 19 410 85 425
rect 19 376 35 410
rect 69 376 85 410
rect 19 360 85 376
rect 119 471 153 487
rect 119 403 153 437
rect 119 326 153 369
rect 188 478 254 493
rect 188 459 204 478
rect 188 425 198 459
rect 238 444 254 478
rect 232 425 254 444
rect 188 410 254 425
rect 188 376 204 410
rect 238 376 254 410
rect 188 360 254 376
rect 288 471 322 487
rect 288 383 322 437
rect 356 478 422 493
rect 356 444 372 478
rect 406 459 422 478
rect 356 425 378 444
rect 412 425 422 459
rect 356 410 422 425
rect 356 376 372 410
rect 406 376 422 410
rect 356 360 422 376
rect 456 471 490 487
rect 456 383 490 437
rect 288 326 322 349
rect 524 478 590 493
rect 524 444 540 478
rect 574 459 590 478
rect 524 425 554 444
rect 588 425 590 459
rect 524 410 590 425
rect 524 376 540 410
rect 574 376 590 410
rect 524 360 590 376
rect 624 471 658 487
rect 624 383 658 437
rect 456 326 490 349
rect 692 478 758 493
rect 692 459 708 478
rect 692 425 699 459
rect 742 444 758 478
rect 733 425 758 444
rect 692 410 758 425
rect 692 376 708 410
rect 742 376 758 410
rect 692 360 758 376
rect 792 471 826 487
rect 792 383 826 437
rect 624 326 658 349
rect 860 478 926 493
rect 860 459 876 478
rect 860 425 871 459
rect 910 444 926 478
rect 905 425 926 444
rect 860 410 926 425
rect 860 376 876 410
rect 910 376 926 410
rect 860 360 926 376
rect 960 471 994 487
rect 960 383 994 437
rect 792 326 826 349
rect 1028 478 1094 493
rect 1028 444 1044 478
rect 1078 459 1094 478
rect 1028 425 1051 444
rect 1085 425 1094 459
rect 1028 410 1094 425
rect 1028 376 1044 410
rect 1078 376 1094 410
rect 1028 360 1094 376
rect 960 326 994 349
rect 23 292 1088 326
rect 23 173 57 292
rect 91 249 973 258
rect 91 215 107 249
rect 141 215 175 249
rect 209 215 243 249
rect 277 215 311 249
rect 345 215 379 249
rect 413 215 447 249
rect 481 215 515 249
rect 549 215 583 249
rect 617 215 651 249
rect 685 215 719 249
rect 753 215 787 249
rect 821 215 855 249
rect 889 215 923 249
rect 957 215 973 249
rect 91 207 973 215
rect 1034 173 1088 292
rect 23 139 1088 173
rect 307 106 345 139
rect 207 95 273 105
rect 207 61 223 95
rect 257 61 273 95
rect 207 17 273 61
rect 307 72 309 106
rect 343 72 345 106
rect 479 106 517 139
rect 307 56 345 72
rect 379 95 445 105
rect 379 61 395 95
rect 429 61 445 95
rect 379 17 445 61
rect 479 72 481 106
rect 515 72 517 106
rect 651 106 689 139
rect 479 56 517 72
rect 551 95 617 105
rect 551 61 567 95
rect 601 61 617 95
rect 551 17 617 61
rect 651 72 653 106
rect 687 72 689 106
rect 823 106 861 139
rect 651 56 689 72
rect 723 95 789 105
rect 723 61 739 95
rect 773 61 789 95
rect 723 17 789 61
rect 823 72 825 106
rect 859 72 861 106
rect 823 56 861 72
rect 895 95 961 105
rect 895 61 911 95
rect 945 61 961 95
rect 895 17 961 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 26 444 35 459
rect 35 444 60 459
rect 26 425 60 444
rect 198 444 204 459
rect 204 444 232 459
rect 198 425 232 444
rect 378 444 406 459
rect 406 444 412 459
rect 378 425 412 444
rect 554 444 574 459
rect 574 444 588 459
rect 554 425 588 444
rect 699 444 708 459
rect 708 444 733 459
rect 699 425 733 444
rect 871 444 876 459
rect 876 444 905 459
rect 871 425 905 444
rect 1051 444 1078 459
rect 1078 444 1085 459
rect 1051 425 1085 444
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 14 459 1182 468
rect 14 425 26 459
rect 60 428 198 459
rect 60 425 72 428
rect 14 416 72 425
rect 186 425 198 428
rect 232 428 378 459
rect 232 425 244 428
rect 186 416 244 425
rect 366 425 378 428
rect 412 428 554 459
rect 412 425 424 428
rect 366 416 424 425
rect 542 425 554 428
rect 588 428 699 459
rect 588 425 600 428
rect 542 416 600 425
rect 687 425 699 428
rect 733 428 871 459
rect 733 425 745 428
rect 687 416 745 425
rect 859 425 871 428
rect 905 428 1051 459
rect 905 425 917 428
rect 859 416 917 425
rect 1039 425 1051 428
rect 1085 428 1182 459
rect 1085 425 1097 428
rect 1039 416 1097 425
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
flabel corelocali s 1042 289 1076 323 0 FreeSans 400 0 0 0 Y
port 7 nsew
flabel corelocali s 1042 221 1076 255 0 FreeSans 400 0 0 0 Y
port 7 nsew
flabel corelocali s 1042 153 1076 187 0 FreeSans 400 0 0 0 Y
port 7 nsew
flabel corelocali s 490 221 524 255 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 398 221 432 255 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 306 221 340 255 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 214 221 248 255 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 858 221 892 255 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 766 221 800 255 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 674 221 708 255 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 582 221 616 255 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 122 221 156 255 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 34 432 72 466 0 FreeSans 200 0 0 0 KAPWR
port 2 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew
rlabel comment s 0 0 0 0 4 lpflow_clkinvkapwr_8
<< properties >>
string FIXED_BBOX 0 0 1196 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2272554
string GDS_START 2262086
string path 0.000 0.000 29.900 0.000 
<< end >>
