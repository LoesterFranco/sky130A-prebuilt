magic
tech sky130A
magscale 1 2
timestamp 1601050088
<< locali >>
rect 217 364 469 444
rect 217 310 263 364
rect 85 236 167 310
rect 229 224 263 310
rect 835 290 935 356
rect 969 290 1223 356
rect 229 190 442 224
rect 229 70 268 190
rect 392 70 442 190
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 17 512 89 596
rect 123 546 199 649
rect 313 546 379 649
rect 493 546 641 649
rect 17 478 664 512
rect 17 364 89 478
rect 630 392 664 478
rect 698 460 748 596
rect 789 494 855 649
rect 889 581 1135 615
rect 889 494 955 581
rect 995 460 1029 547
rect 698 426 1029 460
rect 17 202 51 364
rect 630 326 698 392
rect 732 390 1029 426
rect 1069 390 1135 581
rect 1175 390 1225 649
rect 297 292 596 324
rect 732 292 766 390
rect 297 258 766 292
rect 17 70 95 202
rect 129 17 195 202
rect 306 17 356 156
rect 478 17 528 224
rect 562 85 596 258
rect 800 224 1225 256
rect 630 222 1225 224
rect 630 190 866 222
rect 630 119 664 190
rect 700 85 766 156
rect 800 121 866 190
rect 562 51 766 85
rect 900 17 950 188
rect 986 121 1036 222
rect 1072 17 1122 188
rect 1158 121 1225 222
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
<< metal1 >>
rect 0 683 1248 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 0 617 1248 649
rect 0 17 1248 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
rect 0 -49 1248 -17
<< labels >>
rlabel locali s 835 290 935 356 6 A1
port 1 nsew signal input
rlabel locali s 969 290 1223 356 6 A2
port 2 nsew signal input
rlabel locali s 85 236 167 310 6 B1_N
port 3 nsew signal input
rlabel locali s 392 70 442 190 6 X
port 4 nsew signal output
rlabel locali s 229 224 263 310 6 X
port 4 nsew signal output
rlabel locali s 229 190 442 224 6 X
port 4 nsew signal output
rlabel locali s 229 70 268 190 6 X
port 4 nsew signal output
rlabel locali s 217 364 469 444 6 X
port 4 nsew signal output
rlabel locali s 217 310 263 364 6 X
port 4 nsew signal output
rlabel metal1 s 0 -49 1248 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 617 1248 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1248 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1101342
string GDS_START 1091676
<< end >>
