magic
tech sky130A
magscale 1 2
timestamp 1601050082
<< locali >>
rect 25 260 101 356
rect 374 405 450 471
rect 394 225 450 405
rect 1543 406 1615 596
rect 1581 226 1615 406
rect 1543 70 1615 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 23 424 89 596
rect 129 458 163 649
rect 203 559 269 596
rect 315 593 382 649
rect 760 593 826 649
rect 416 559 692 593
rect 956 581 1168 615
rect 956 559 990 581
rect 203 525 450 559
rect 658 525 990 559
rect 23 390 169 424
rect 135 310 169 390
rect 203 364 295 525
rect 261 336 295 364
rect 135 226 227 310
rect 23 192 227 226
rect 23 70 73 192
rect 109 17 159 158
rect 193 85 227 192
rect 261 270 352 336
rect 261 119 295 270
rect 484 248 518 525
rect 552 491 624 525
rect 552 457 828 491
rect 552 316 586 457
rect 620 350 752 416
rect 552 282 684 316
rect 484 214 595 248
rect 329 146 531 180
rect 329 85 363 146
rect 193 51 363 85
rect 397 17 463 112
rect 497 89 531 146
rect 631 123 684 282
rect 718 172 752 350
rect 794 391 828 457
rect 867 425 922 491
rect 794 325 854 391
rect 786 240 852 283
rect 888 240 922 425
rect 956 308 990 525
rect 1024 376 1058 547
rect 1102 410 1168 581
rect 1240 504 1306 649
rect 1024 342 1164 376
rect 956 274 1096 308
rect 786 206 1000 240
rect 1034 230 1096 274
rect 1130 280 1164 342
rect 1210 372 1276 448
rect 1352 372 1402 540
rect 1442 406 1508 649
rect 1210 338 1547 372
rect 1210 314 1276 338
rect 1375 280 1441 304
rect 1130 246 1441 280
rect 718 138 932 172
rect 718 89 752 138
rect 497 55 752 89
rect 814 17 864 104
rect 898 85 932 138
rect 966 119 1000 206
rect 1130 196 1164 246
rect 1375 238 1441 246
rect 1475 270 1547 338
rect 1044 146 1164 196
rect 1113 85 1179 102
rect 898 51 1179 85
rect 1246 17 1312 212
rect 1475 204 1509 270
rect 1358 170 1509 204
rect 1358 70 1408 170
rect 1444 17 1507 136
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
rlabel locali s 394 225 450 405 6 D
port 1 nsew signal input
rlabel locali s 374 405 450 471 6 D
port 1 nsew signal input
rlabel locali s 1581 226 1615 406 6 Q
port 2 nsew signal output
rlabel locali s 1543 406 1615 596 6 Q
port 2 nsew signal output
rlabel locali s 1543 70 1615 226 6 Q
port 2 nsew signal output
rlabel locali s 25 260 101 356 6 CLK
port 3 nsew clock input
rlabel metal1 s 0 -49 1632 49 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1632 715 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2664938
string GDS_START 2652306
<< end >>
