magic
tech sky130A
magscale 1 2
timestamp 1601050047
<< nwell >>
rect -38 332 1190 704
<< pwell >>
rect 0 0 1152 49
<< scpmos >>
rect 219 368 249 536
rect 309 368 339 536
rect 416 368 446 592
rect 582 368 612 592
rect 932 368 962 592
rect 1026 368 1056 592
<< nmoslvt >>
rect 88 74 118 222
rect 300 74 330 222
rect 386 74 416 222
rect 472 74 502 222
rect 585 74 615 222
rect 671 74 701 222
rect 771 74 801 222
rect 857 74 887 222
rect 1038 74 1068 222
<< ndiff >>
rect 31 210 88 222
rect 31 176 43 210
rect 77 176 88 210
rect 31 120 88 176
rect 31 86 43 120
rect 77 86 88 120
rect 31 74 88 86
rect 118 131 175 222
rect 118 97 129 131
rect 163 97 175 131
rect 118 74 175 97
rect 243 131 300 222
rect 243 97 255 131
rect 289 97 300 131
rect 243 74 300 97
rect 330 181 386 222
rect 330 147 341 181
rect 375 147 386 181
rect 330 74 386 147
rect 416 184 472 222
rect 416 150 427 184
rect 461 150 472 184
rect 416 116 472 150
rect 416 82 427 116
rect 461 82 472 116
rect 416 74 472 82
rect 502 181 585 222
rect 502 147 528 181
rect 562 147 585 181
rect 502 74 585 147
rect 615 184 671 222
rect 615 150 626 184
rect 660 150 671 184
rect 615 116 671 150
rect 615 82 626 116
rect 660 82 671 116
rect 615 74 671 82
rect 701 116 771 222
rect 701 82 726 116
rect 760 82 771 116
rect 701 74 771 82
rect 801 205 857 222
rect 801 171 812 205
rect 846 171 857 205
rect 801 116 857 171
rect 801 82 812 116
rect 846 82 857 116
rect 801 74 857 82
rect 887 142 1038 222
rect 887 108 898 142
rect 932 108 993 142
rect 1027 108 1038 142
rect 887 74 1038 108
rect 1068 210 1125 222
rect 1068 176 1079 210
rect 1113 176 1125 210
rect 1068 120 1125 176
rect 1068 86 1079 120
rect 1113 86 1125 120
rect 1068 74 1125 86
<< pdiff >>
rect 357 580 416 592
rect 357 546 369 580
rect 403 546 416 580
rect 357 536 416 546
rect 91 524 219 536
rect 91 490 103 524
rect 137 490 171 524
rect 205 490 219 524
rect 91 440 219 490
rect 91 406 103 440
rect 137 406 171 440
rect 205 406 219 440
rect 91 368 219 406
rect 249 524 309 536
rect 249 490 262 524
rect 296 490 309 524
rect 249 440 309 490
rect 249 406 262 440
rect 296 406 309 440
rect 249 368 309 406
rect 339 500 416 536
rect 339 466 369 500
rect 403 466 416 500
rect 339 420 416 466
rect 339 386 369 420
rect 403 386 416 420
rect 339 368 416 386
rect 446 580 582 592
rect 446 546 459 580
rect 493 546 535 580
rect 569 546 582 580
rect 446 500 582 546
rect 446 466 459 500
rect 493 466 535 500
rect 569 466 582 500
rect 446 420 582 466
rect 446 386 459 420
rect 493 386 535 420
rect 569 386 582 420
rect 446 368 582 386
rect 612 580 932 592
rect 612 546 625 580
rect 659 546 709 580
rect 743 546 795 580
rect 829 546 879 580
rect 913 546 932 580
rect 612 498 932 546
rect 612 464 625 498
rect 659 464 709 498
rect 743 464 795 498
rect 829 464 879 498
rect 913 464 932 498
rect 612 368 932 464
rect 962 580 1026 592
rect 962 546 979 580
rect 1013 546 1026 580
rect 962 510 1026 546
rect 962 476 979 510
rect 1013 476 1026 510
rect 962 440 1026 476
rect 962 406 979 440
rect 1013 406 1026 440
rect 962 368 1026 406
rect 1056 580 1116 592
rect 1056 546 1070 580
rect 1104 546 1116 580
rect 1056 510 1116 546
rect 1056 476 1070 510
rect 1104 476 1116 510
rect 1056 440 1116 476
rect 1056 406 1070 440
rect 1104 406 1116 440
rect 1056 368 1116 406
<< ndiffc >>
rect 43 176 77 210
rect 43 86 77 120
rect 129 97 163 131
rect 255 97 289 131
rect 341 147 375 181
rect 427 150 461 184
rect 427 82 461 116
rect 528 147 562 181
rect 626 150 660 184
rect 626 82 660 116
rect 726 82 760 116
rect 812 171 846 205
rect 812 82 846 116
rect 898 108 932 142
rect 993 108 1027 142
rect 1079 176 1113 210
rect 1079 86 1113 120
<< pdiffc >>
rect 369 546 403 580
rect 103 490 137 524
rect 171 490 205 524
rect 103 406 137 440
rect 171 406 205 440
rect 262 490 296 524
rect 262 406 296 440
rect 369 466 403 500
rect 369 386 403 420
rect 459 546 493 580
rect 535 546 569 580
rect 459 466 493 500
rect 535 466 569 500
rect 459 386 493 420
rect 535 386 569 420
rect 625 546 659 580
rect 709 546 743 580
rect 795 546 829 580
rect 879 546 913 580
rect 625 464 659 498
rect 709 464 743 498
rect 795 464 829 498
rect 879 464 913 498
rect 979 546 1013 580
rect 979 476 1013 510
rect 979 406 1013 440
rect 1070 546 1104 580
rect 1070 476 1104 510
rect 1070 406 1104 440
<< poly >>
rect 416 592 446 618
rect 582 592 612 618
rect 932 592 962 618
rect 1026 592 1056 618
rect 219 536 249 562
rect 309 536 339 562
rect 219 353 249 368
rect 309 353 339 368
rect 416 353 446 368
rect 582 353 612 368
rect 932 353 962 368
rect 1026 353 1056 368
rect 216 345 252 353
rect 306 345 342 353
rect 21 315 342 345
rect 413 336 449 353
rect 579 336 615 353
rect 413 320 615 336
rect 929 326 965 353
rect 1023 326 1059 353
rect 21 310 252 315
rect 21 276 37 310
rect 71 276 105 310
rect 139 276 173 310
rect 207 276 252 310
rect 21 260 252 276
rect 413 286 429 320
rect 463 286 497 320
rect 531 286 565 320
rect 599 286 615 320
rect 413 267 615 286
rect 88 222 118 260
rect 300 237 615 267
rect 300 222 330 237
rect 386 222 416 237
rect 472 222 502 237
rect 585 222 615 237
rect 671 310 1107 326
rect 671 276 785 310
rect 819 276 853 310
rect 887 276 921 310
rect 955 276 989 310
rect 1023 276 1057 310
rect 1091 276 1107 310
rect 671 260 1107 276
rect 671 222 701 260
rect 771 222 801 260
rect 857 222 887 260
rect 1038 222 1068 260
rect 88 48 118 74
rect 300 48 330 74
rect 386 48 416 74
rect 472 48 502 74
rect 585 48 615 74
rect 671 48 701 74
rect 771 48 801 74
rect 857 48 887 74
rect 1038 48 1068 74
<< polycont >>
rect 37 276 71 310
rect 105 276 139 310
rect 173 276 207 310
rect 429 286 463 320
rect 497 286 531 320
rect 565 286 599 320
rect 785 276 819 310
rect 853 276 887 310
rect 921 276 955 310
rect 989 276 1023 310
rect 1057 276 1091 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 87 524 212 649
rect 353 580 419 649
rect 353 546 369 580
rect 403 546 419 580
rect 87 490 103 524
rect 137 490 171 524
rect 205 490 212 524
rect 87 440 212 490
rect 87 406 103 440
rect 137 406 171 440
rect 205 406 212 440
rect 87 390 212 406
rect 246 524 312 540
rect 246 490 262 524
rect 296 490 312 524
rect 246 440 312 490
rect 246 406 262 440
rect 296 406 312 440
rect 246 390 312 406
rect 353 500 419 546
rect 353 466 369 500
rect 403 466 419 500
rect 353 420 419 466
rect 21 310 223 356
rect 21 276 37 310
rect 71 276 105 310
rect 139 276 173 310
rect 207 276 223 310
rect 21 260 223 276
rect 257 336 291 390
rect 353 386 369 420
rect 403 386 419 420
rect 353 370 419 386
rect 453 580 575 596
rect 453 546 459 580
rect 493 546 535 580
rect 569 546 575 580
rect 453 500 575 546
rect 453 466 459 500
rect 493 466 535 500
rect 569 466 575 500
rect 453 430 575 466
rect 609 580 929 649
rect 609 546 625 580
rect 659 546 709 580
rect 743 546 795 580
rect 829 546 879 580
rect 913 546 929 580
rect 609 498 929 546
rect 609 464 625 498
rect 659 464 709 498
rect 743 464 795 498
rect 829 464 879 498
rect 913 464 929 498
rect 963 580 1029 596
rect 963 546 979 580
rect 1013 546 1029 580
rect 963 510 1029 546
rect 963 476 979 510
rect 1013 476 1029 510
rect 963 440 1029 476
rect 963 430 979 440
rect 453 420 979 430
rect 453 386 459 420
rect 493 386 535 420
rect 569 406 979 420
rect 1013 406 1029 440
rect 569 390 1029 406
rect 1063 580 1120 649
rect 1063 546 1070 580
rect 1104 546 1120 580
rect 1063 510 1120 546
rect 1063 476 1070 510
rect 1104 476 1120 510
rect 1063 440 1120 476
rect 1063 406 1070 440
rect 1104 406 1120 440
rect 1063 390 1120 406
rect 569 386 839 390
rect 453 370 839 386
rect 257 320 615 336
rect 257 286 429 320
rect 463 286 497 320
rect 531 286 565 320
rect 599 286 615 320
rect 257 226 291 286
rect 657 252 731 370
rect 889 326 1131 356
rect 769 310 1131 326
rect 769 276 785 310
rect 819 276 853 310
rect 887 276 921 310
rect 955 276 989 310
rect 1023 276 1057 310
rect 1091 276 1131 310
rect 769 260 1131 276
rect 27 210 291 226
rect 27 176 43 210
rect 77 192 291 210
rect 325 218 731 252
rect 27 120 77 176
rect 325 181 377 218
rect 27 86 43 120
rect 27 70 77 86
rect 113 131 179 158
rect 113 97 129 131
rect 163 97 179 131
rect 113 17 179 97
rect 239 131 291 158
rect 239 97 255 131
rect 289 97 291 131
rect 325 147 341 181
rect 375 147 377 181
rect 325 127 377 147
rect 411 150 427 184
rect 461 150 477 184
rect 239 85 291 97
rect 411 116 477 150
rect 511 181 576 218
rect 796 210 1129 226
rect 796 205 1079 210
rect 796 184 812 205
rect 511 147 528 181
rect 562 147 576 181
rect 511 127 576 147
rect 610 150 626 184
rect 660 171 812 184
rect 846 192 1079 205
rect 846 171 862 192
rect 660 150 862 171
rect 1063 176 1079 192
rect 1113 176 1129 210
rect 411 85 427 116
rect 239 82 427 85
rect 461 85 477 116
rect 610 116 676 150
rect 810 116 862 150
rect 610 85 626 116
rect 461 82 626 85
rect 660 82 676 116
rect 239 51 676 82
rect 710 82 726 116
rect 760 82 776 116
rect 710 17 776 82
rect 810 82 812 116
rect 846 82 862 116
rect 810 66 862 82
rect 896 142 1029 158
rect 896 108 898 142
rect 932 108 993 142
rect 1027 108 1029 142
rect 896 17 1029 108
rect 1063 120 1129 176
rect 1063 86 1079 120
rect 1113 86 1129 120
rect 1063 70 1129 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
rlabel comment s 0 0 0 0 4 nand2b_4
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew
flabel corelocali s 703 390 737 424 0 FreeSans 340 0 0 0 Y
port 7 nsew
flabel corelocali s 799 390 833 424 0 FreeSans 340 0 0 0 Y
port 7 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 1087 316 1121 350 0 FreeSans 340 0 0 0 B
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 1152 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 2052084
string GDS_START 2042736
<< end >>
