magic
tech sky130A
magscale 1 2
timestamp 1601050058
<< locali >>
rect 507 359 557 493
rect 25 153 66 331
rect 168 199 249 265
rect 178 84 249 199
rect 283 85 340 265
rect 381 187 415 265
rect 523 331 557 359
rect 675 349 709 493
rect 675 331 810 349
rect 523 297 810 331
rect 381 146 431 187
rect 760 162 810 297
rect 507 128 810 162
rect 507 51 541 128
rect 675 51 709 128
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 21 367 77 527
rect 111 333 153 493
rect 191 387 257 527
rect 291 333 329 493
rect 405 371 471 527
rect 591 367 641 527
rect 100 299 483 333
rect 100 117 134 299
rect 35 51 134 117
rect 449 261 483 299
rect 743 383 809 527
rect 449 221 717 261
rect 515 215 717 221
rect 405 17 467 110
rect 575 17 641 94
rect 743 17 809 94
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
rlabel locali s 25 153 66 331 6 A
port 1 nsew signal input
rlabel locali s 178 84 249 199 6 B
port 2 nsew signal input
rlabel locali s 168 199 249 265 6 B
port 2 nsew signal input
rlabel locali s 283 85 340 265 6 C
port 3 nsew signal input
rlabel locali s 381 187 415 265 6 D
port 4 nsew signal input
rlabel locali s 381 146 431 187 6 D
port 4 nsew signal input
rlabel locali s 760 162 810 297 6 X
port 5 nsew signal output
rlabel locali s 675 349 709 493 6 X
port 5 nsew signal output
rlabel locali s 675 331 810 349 6 X
port 5 nsew signal output
rlabel locali s 675 51 709 128 6 X
port 5 nsew signal output
rlabel locali s 523 331 557 359 6 X
port 5 nsew signal output
rlabel locali s 523 297 810 331 6 X
port 5 nsew signal output
rlabel locali s 507 359 557 493 6 X
port 5 nsew signal output
rlabel locali s 507 128 810 162 6 X
port 5 nsew signal output
rlabel locali s 507 51 541 128 6 X
port 5 nsew signal output
rlabel metal1 s 0 -48 828 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 828 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3835332
string GDS_START 3827942
<< end >>
