magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 103 333 179 493
rect 291 333 367 493
rect 479 337 555 493
rect 479 333 653 337
rect 103 299 653 333
rect 57 215 539 265
rect 573 181 653 299
rect 129 145 653 181
rect 129 51 163 145
rect 317 51 351 145
rect 505 51 539 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 35 299 69 527
rect 223 367 257 527
rect 411 367 445 527
rect 599 435 633 527
rect 26 17 79 109
rect 223 17 257 109
rect 411 17 445 109
rect 573 17 633 110
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel locali s 57 215 539 265 6 A
port 1 nsew signal input
rlabel locali s 573 181 653 299 6 Y
port 2 nsew signal output
rlabel locali s 505 51 539 145 6 Y
port 2 nsew signal output
rlabel locali s 479 337 555 493 6 Y
port 2 nsew signal output
rlabel locali s 479 333 653 337 6 Y
port 2 nsew signal output
rlabel locali s 317 51 351 145 6 Y
port 2 nsew signal output
rlabel locali s 291 333 367 493 6 Y
port 2 nsew signal output
rlabel locali s 129 145 653 181 6 Y
port 2 nsew signal output
rlabel locali s 129 51 163 145 6 Y
port 2 nsew signal output
rlabel locali s 103 333 179 493 6 Y
port 2 nsew signal output
rlabel locali s 103 299 653 333 6 Y
port 2 nsew signal output
rlabel metal1 s 0 -48 736 48 8 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 496 736 592 6 VPWR
port 4 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2113776
string GDS_START 2107410
<< end >>
