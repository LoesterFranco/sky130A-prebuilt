magic
tech sky130A
magscale 1 2
timestamp 1604502729
<< locali >>
rect 25 270 114 356
rect 329 390 559 440
rect 329 364 455 390
rect 409 278 455 364
rect 340 244 455 278
rect 489 270 555 356
rect 340 126 374 244
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 23 424 89 572
rect 145 458 219 649
rect 403 542 469 649
rect 583 542 649 649
rect 261 474 649 508
rect 23 390 195 424
rect 161 294 195 390
rect 161 236 227 294
rect 23 228 227 236
rect 23 202 195 228
rect 23 70 89 202
rect 261 194 295 474
rect 123 17 175 168
rect 238 85 304 194
rect 615 226 649 474
rect 410 85 476 210
rect 238 51 476 85
rect 512 17 546 226
rect 583 70 649 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel locali s 25 270 114 356 6 A_N
port 1 nsew signal input
rlabel locali s 489 270 555 356 6 B
port 2 nsew signal input
rlabel locali s 409 278 455 364 6 Y
port 3 nsew signal output
rlabel locali s 340 244 455 278 6 Y
port 3 nsew signal output
rlabel locali s 340 126 374 244 6 Y
port 3 nsew signal output
rlabel locali s 329 390 559 440 6 Y
port 3 nsew signal output
rlabel locali s 329 364 455 390 6 Y
port 3 nsew signal output
rlabel metal1 s 0 -49 672 49 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 617 672 715 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 2057990
string GDS_START 2052142
<< end >>
