magic
tech sky130A
magscale 1 2
timestamp 1601050047
<< nwell >>
rect -38 332 518 704
<< pwell >>
rect 0 0 480 49
<< scpmos >>
rect 93 368 123 592
rect 183 368 213 592
rect 273 368 303 592
rect 363 368 393 592
<< nmoslvt >>
rect 90 74 120 222
rect 184 74 214 222
rect 280 74 310 222
rect 366 74 396 222
<< ndiff >>
rect 27 210 90 222
rect 27 176 39 210
rect 73 176 90 210
rect 27 120 90 176
rect 27 86 39 120
rect 73 86 90 120
rect 27 74 90 86
rect 120 210 184 222
rect 120 176 139 210
rect 173 176 184 210
rect 120 120 184 176
rect 120 86 139 120
rect 173 86 184 120
rect 120 74 184 86
rect 214 136 280 222
rect 214 102 225 136
rect 259 102 280 136
rect 214 74 280 102
rect 310 210 366 222
rect 310 176 321 210
rect 355 176 366 210
rect 310 120 366 176
rect 310 86 321 120
rect 355 86 366 120
rect 310 74 366 86
rect 396 136 453 222
rect 396 102 407 136
rect 441 102 453 136
rect 396 74 453 102
<< pdiff >>
rect 34 580 93 592
rect 34 546 46 580
rect 80 546 93 580
rect 34 510 93 546
rect 34 476 46 510
rect 80 476 93 510
rect 34 440 93 476
rect 34 406 46 440
rect 80 406 93 440
rect 34 368 93 406
rect 123 580 183 592
rect 123 546 136 580
rect 170 546 183 580
rect 123 510 183 546
rect 123 476 136 510
rect 170 476 183 510
rect 123 440 183 476
rect 123 406 136 440
rect 170 406 183 440
rect 123 368 183 406
rect 213 580 273 592
rect 213 546 226 580
rect 260 546 273 580
rect 213 508 273 546
rect 213 474 226 508
rect 260 474 273 508
rect 213 368 273 474
rect 303 580 363 592
rect 303 546 316 580
rect 350 546 363 580
rect 303 510 363 546
rect 303 476 316 510
rect 350 476 363 510
rect 303 440 363 476
rect 303 406 316 440
rect 350 406 363 440
rect 303 368 363 406
rect 393 580 452 592
rect 393 546 406 580
rect 440 546 452 580
rect 393 508 452 546
rect 393 474 406 508
rect 440 474 452 508
rect 393 368 452 474
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 139 176 173 210
rect 139 86 173 120
rect 225 102 259 136
rect 321 176 355 210
rect 321 86 355 120
rect 407 102 441 136
<< pdiffc >>
rect 46 546 80 580
rect 46 476 80 510
rect 46 406 80 440
rect 136 546 170 580
rect 136 476 170 510
rect 136 406 170 440
rect 226 546 260 580
rect 226 474 260 508
rect 316 546 350 580
rect 316 476 350 510
rect 316 406 350 440
rect 406 546 440 580
rect 406 474 440 508
<< poly >>
rect 93 592 123 618
rect 183 592 213 618
rect 273 592 303 618
rect 363 592 393 618
rect 93 353 123 368
rect 183 353 213 368
rect 273 353 303 368
rect 363 353 393 368
rect 90 336 126 353
rect 180 336 216 353
rect 270 336 306 353
rect 360 336 396 353
rect 90 320 396 336
rect 90 286 106 320
rect 140 286 174 320
rect 208 286 242 320
rect 276 286 310 320
rect 344 286 396 320
rect 90 270 396 286
rect 90 222 120 270
rect 184 222 214 270
rect 280 222 310 270
rect 366 222 396 270
rect 90 48 120 74
rect 184 48 214 74
rect 280 48 310 74
rect 366 48 396 74
<< polycont >>
rect 106 286 140 320
rect 174 286 208 320
rect 242 286 276 320
rect 310 286 344 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 30 580 80 649
rect 30 546 46 580
rect 30 510 80 546
rect 30 476 46 510
rect 30 440 80 476
rect 30 406 46 440
rect 30 390 80 406
rect 120 580 186 596
rect 120 546 136 580
rect 170 546 186 580
rect 120 510 186 546
rect 120 476 136 510
rect 170 476 186 510
rect 120 440 186 476
rect 226 580 260 649
rect 226 508 260 546
rect 226 458 260 474
rect 300 580 366 596
rect 300 546 316 580
rect 350 546 366 580
rect 300 510 366 546
rect 300 476 316 510
rect 350 476 366 510
rect 120 406 136 440
rect 170 424 186 440
rect 300 440 366 476
rect 406 580 456 649
rect 440 546 456 580
rect 406 508 456 546
rect 440 474 456 508
rect 406 458 456 474
rect 300 424 316 440
rect 170 406 316 424
rect 350 424 366 440
rect 350 406 455 424
rect 120 390 455 406
rect 25 320 360 356
rect 25 286 106 320
rect 140 286 174 320
rect 208 286 242 320
rect 276 286 310 320
rect 344 286 360 320
rect 25 270 360 286
rect 409 236 455 390
rect 23 210 89 226
rect 23 176 39 210
rect 73 176 89 210
rect 23 120 89 176
rect 23 86 39 120
rect 73 86 89 120
rect 23 17 89 86
rect 123 210 455 236
rect 123 176 139 210
rect 173 202 321 210
rect 123 120 173 176
rect 355 202 455 210
rect 123 86 139 120
rect 123 70 173 86
rect 209 136 275 168
rect 209 102 225 136
rect 259 102 275 136
rect 209 17 275 102
rect 321 120 355 176
rect 321 70 355 86
rect 391 136 457 168
rect 391 102 407 136
rect 441 102 457 136
rect 391 17 457 102
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< metal1 >>
rect 0 683 480 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 0 617 480 649
rect 0 17 480 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
rect 0 -49 480 -17
<< labels >>
rlabel comment s 0 0 0 0 4 inv_4
flabel pwell s 0 0 480 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew
flabel nbase s 0 617 480 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew
flabel metal1 s 0 617 480 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew
flabel metal1 s 0 0 480 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew
flabel corelocali s 415 242 449 276 0 FreeSans 340 0 0 0 Y
port 6 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 480 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1861282
string GDS_START 1856128
<< end >>
