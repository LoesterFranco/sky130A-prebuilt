magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 1326 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 95 47 125 177
rect 191 47 221 177
rect 287 47 317 177
rect 373 47 403 177
rect 469 47 499 177
rect 565 47 595 177
rect 671 47 701 177
rect 775 47 805 177
rect 861 47 891 177
rect 957 47 987 177
rect 1053 47 1083 177
rect 1159 47 1189 177
<< pmoshvt >>
rect 87 297 123 497
rect 183 297 219 497
rect 279 297 315 497
rect 375 297 411 497
rect 471 297 507 497
rect 567 297 603 497
rect 663 297 699 497
rect 759 297 795 497
rect 863 297 899 497
rect 959 297 995 497
rect 1055 297 1091 497
rect 1151 297 1187 497
<< ndiff >>
rect 32 157 95 177
rect 32 123 40 157
rect 74 123 95 157
rect 32 47 95 123
rect 125 89 191 177
rect 125 55 136 89
rect 170 55 191 89
rect 125 47 191 55
rect 221 157 287 177
rect 221 123 232 157
rect 266 123 287 157
rect 221 47 287 123
rect 317 89 373 177
rect 317 55 328 89
rect 362 55 373 89
rect 317 47 373 55
rect 403 157 469 177
rect 403 123 424 157
rect 458 123 469 157
rect 403 47 469 123
rect 499 89 565 177
rect 499 55 520 89
rect 554 55 565 89
rect 499 47 565 55
rect 595 157 671 177
rect 595 123 616 157
rect 650 123 671 157
rect 595 47 671 123
rect 701 89 775 177
rect 701 55 712 89
rect 746 55 775 89
rect 701 47 775 55
rect 805 125 861 177
rect 805 91 816 125
rect 850 91 861 125
rect 805 47 861 91
rect 891 157 957 177
rect 891 123 912 157
rect 946 123 957 157
rect 891 47 957 123
rect 987 89 1053 177
rect 987 55 1008 89
rect 1042 55 1053 89
rect 987 47 1053 55
rect 1083 157 1159 177
rect 1083 123 1104 157
rect 1138 123 1159 157
rect 1083 47 1159 123
rect 1189 89 1246 177
rect 1189 55 1200 89
rect 1234 55 1246 89
rect 1189 47 1246 55
<< pdiff >>
rect 32 485 87 497
rect 32 451 40 485
rect 74 451 87 485
rect 32 417 87 451
rect 32 383 40 417
rect 74 383 87 417
rect 32 297 87 383
rect 123 477 183 497
rect 123 443 136 477
rect 170 443 183 477
rect 123 297 183 443
rect 219 485 279 497
rect 219 451 232 485
rect 266 451 279 485
rect 219 297 279 451
rect 315 477 375 497
rect 315 443 328 477
rect 362 443 375 477
rect 315 297 375 443
rect 411 405 471 497
rect 411 371 424 405
rect 458 371 471 405
rect 411 297 471 371
rect 507 489 567 497
rect 507 455 520 489
rect 554 455 567 489
rect 507 297 567 455
rect 603 405 663 497
rect 603 371 616 405
rect 650 371 663 405
rect 603 297 663 371
rect 699 489 759 497
rect 699 455 712 489
rect 746 455 759 489
rect 699 297 759 455
rect 795 489 863 497
rect 795 455 812 489
rect 846 455 863 489
rect 795 297 863 455
rect 899 477 959 497
rect 899 443 912 477
rect 946 443 959 477
rect 899 382 959 443
rect 899 348 912 382
rect 946 348 959 382
rect 899 297 959 348
rect 995 485 1055 497
rect 995 451 1008 485
rect 1042 451 1055 485
rect 995 297 1055 451
rect 1091 477 1151 497
rect 1091 443 1104 477
rect 1138 443 1151 477
rect 1091 382 1151 443
rect 1091 348 1104 382
rect 1138 348 1151 382
rect 1091 297 1151 348
rect 1187 485 1242 497
rect 1187 451 1200 485
rect 1234 451 1242 485
rect 1187 410 1242 451
rect 1187 376 1200 410
rect 1234 376 1242 410
rect 1187 297 1242 376
<< ndiffc >>
rect 40 123 74 157
rect 136 55 170 89
rect 232 123 266 157
rect 328 55 362 89
rect 424 123 458 157
rect 520 55 554 89
rect 616 123 650 157
rect 712 55 746 89
rect 816 91 850 125
rect 912 123 946 157
rect 1008 55 1042 89
rect 1104 123 1138 157
rect 1200 55 1234 89
<< pdiffc >>
rect 40 451 74 485
rect 40 383 74 417
rect 136 443 170 477
rect 232 451 266 485
rect 328 443 362 477
rect 424 371 458 405
rect 520 455 554 489
rect 616 371 650 405
rect 712 455 746 489
rect 812 455 846 489
rect 912 443 946 477
rect 912 348 946 382
rect 1008 451 1042 485
rect 1104 443 1138 477
rect 1104 348 1138 382
rect 1200 451 1234 485
rect 1200 376 1234 410
<< poly >>
rect 87 497 123 523
rect 183 497 219 523
rect 279 497 315 523
rect 375 497 411 523
rect 471 497 507 523
rect 567 497 603 523
rect 663 497 699 523
rect 759 497 795 523
rect 863 497 899 523
rect 959 497 995 523
rect 1055 497 1091 523
rect 1151 497 1187 523
rect 87 282 123 297
rect 183 282 219 297
rect 279 282 315 297
rect 375 282 411 297
rect 471 282 507 297
rect 567 282 603 297
rect 663 282 699 297
rect 759 282 795 297
rect 863 282 899 297
rect 959 282 995 297
rect 1055 282 1091 297
rect 1151 282 1187 297
rect 85 265 125 282
rect 181 265 221 282
rect 277 265 317 282
rect 373 265 413 282
rect 469 265 509 282
rect 565 265 605 282
rect 661 265 701 282
rect 757 265 797 282
rect 861 265 901 282
rect 957 265 997 282
rect 1053 265 1093 282
rect 1149 265 1189 282
rect 25 249 325 265
rect 25 215 41 249
rect 75 215 109 249
rect 143 215 187 249
rect 221 215 265 249
rect 299 215 325 249
rect 25 199 325 215
rect 373 249 701 265
rect 373 215 455 249
rect 489 215 551 249
rect 585 215 641 249
rect 675 215 701 249
rect 373 199 701 215
rect 743 249 819 265
rect 743 215 759 249
rect 793 215 819 249
rect 743 199 819 215
rect 861 249 1189 265
rect 861 215 877 249
rect 911 215 955 249
rect 989 215 1033 249
rect 1067 215 1189 249
rect 861 199 1189 215
rect 95 177 125 199
rect 191 177 221 199
rect 287 177 317 199
rect 373 177 403 199
rect 469 177 499 199
rect 565 177 595 199
rect 671 177 701 199
rect 775 177 805 199
rect 861 177 891 199
rect 957 177 987 199
rect 1053 177 1083 199
rect 1159 177 1189 199
rect 95 21 125 47
rect 191 21 221 47
rect 287 21 317 47
rect 373 21 403 47
rect 469 21 499 47
rect 565 21 595 47
rect 671 21 701 47
rect 775 21 805 47
rect 861 21 891 47
rect 957 21 987 47
rect 1053 21 1083 47
rect 1159 21 1189 47
<< polycont >>
rect 41 215 75 249
rect 109 215 143 249
rect 187 215 221 249
rect 265 215 299 249
rect 455 215 489 249
rect 551 215 585 249
rect 641 215 675 249
rect 759 215 793 249
rect 877 215 911 249
rect 955 215 989 249
rect 1033 215 1067 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 24 485 81 527
rect 24 451 40 485
rect 74 451 81 485
rect 24 417 81 451
rect 24 383 40 417
rect 74 383 81 417
rect 125 477 172 493
rect 125 443 136 477
rect 170 443 172 477
rect 206 485 282 527
rect 206 451 232 485
rect 266 451 282 485
rect 326 489 762 493
rect 326 477 520 489
rect 125 417 172 443
rect 326 443 328 477
rect 362 455 520 477
rect 554 455 712 489
rect 746 455 762 489
rect 806 489 862 527
rect 806 455 812 489
rect 846 455 862 489
rect 362 443 364 455
rect 326 417 364 443
rect 806 439 862 455
rect 906 477 948 493
rect 906 443 912 477
rect 946 443 948 477
rect 982 485 1058 527
rect 982 451 1008 485
rect 1042 451 1058 485
rect 1102 477 1140 493
rect 125 383 364 417
rect 906 417 948 443
rect 1102 443 1104 477
rect 1138 443 1140 477
rect 1102 417 1140 443
rect 906 405 1140 417
rect 24 364 81 383
rect 398 371 424 405
rect 458 371 616 405
rect 650 382 1140 405
rect 650 371 912 382
rect 867 348 912 371
rect 946 348 1104 382
rect 1138 348 1140 382
rect 1174 485 1250 527
rect 1174 451 1200 485
rect 1234 451 1250 485
rect 1174 410 1250 451
rect 1174 376 1200 410
rect 1234 376 1250 410
rect 867 340 1140 348
rect 125 303 819 337
rect 125 264 325 303
rect 25 249 325 264
rect 25 215 41 249
rect 75 215 109 249
rect 143 215 187 249
rect 221 215 265 249
rect 299 215 325 249
rect 25 203 325 215
rect 437 249 725 269
rect 437 215 455 249
rect 489 215 551 249
rect 585 215 641 249
rect 675 215 725 249
rect 437 214 725 215
rect 759 249 819 303
rect 867 289 1266 340
rect 793 215 819 249
rect 759 198 819 215
rect 861 249 1120 255
rect 861 215 877 249
rect 911 215 955 249
rect 989 215 1033 249
rect 1067 215 1120 249
rect 861 203 1120 215
rect 1184 169 1266 289
rect 24 157 852 164
rect 24 123 40 157
rect 74 123 232 157
rect 266 123 424 157
rect 458 123 616 157
rect 650 125 852 157
rect 650 123 816 125
rect 806 91 816 123
rect 850 91 852 125
rect 886 157 1266 169
rect 886 123 912 157
rect 946 123 1104 157
rect 1138 123 1266 157
rect 806 89 852 91
rect 110 55 136 89
rect 170 55 186 89
rect 110 17 186 55
rect 302 55 328 89
rect 362 55 378 89
rect 302 17 378 55
rect 494 55 520 89
rect 554 55 570 89
rect 494 17 570 55
rect 686 55 712 89
rect 746 55 762 89
rect 686 17 762 55
rect 806 55 1008 89
rect 1042 55 1200 89
rect 1234 55 1250 89
rect 806 51 1250 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
flabel corelocali s 1232 153 1266 187 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 947 221 981 255 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 472 238 472 238 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 230 306 230 306 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
rlabel comment s 0 0 0 0 4 o21ai_4
<< properties >>
string FIXED_BBOX 0 0 1288 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1002668
string GDS_START 994134
<< end >>
