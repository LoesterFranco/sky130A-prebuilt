magic
tech sky130A
magscale 1 2
timestamp 1599588238
<< locali >>
rect 25 270 110 356
rect 212 370 278 420
rect 212 236 246 370
rect 697 294 785 360
rect 212 88 263 236
rect 887 260 939 356
rect 697 114 743 134
rect 630 51 743 114
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 21 488 87 596
rect 121 522 187 649
rect 302 522 368 649
rect 410 556 476 596
rect 410 522 521 556
rect 21 454 453 488
rect 21 420 178 454
rect 144 236 178 420
rect 24 202 178 236
rect 280 270 346 336
rect 394 294 453 454
rect 312 260 346 270
rect 487 260 521 522
rect 764 462 830 649
rect 872 428 938 564
rect 555 394 938 428
rect 555 294 614 394
rect 819 390 938 394
rect 24 134 90 202
rect 126 17 176 168
rect 312 226 747 260
rect 315 17 407 182
rect 462 116 528 226
rect 562 148 639 192
rect 681 168 747 226
rect 819 226 853 390
rect 819 192 937 226
rect 562 17 596 148
rect 785 17 851 158
rect 887 87 937 192
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
rlabel locali s 697 294 785 360 6 A
port 1 nsew signal input
rlabel locali s 697 114 743 134 6 B
port 2 nsew signal input
rlabel locali s 630 51 743 114 6 B
port 2 nsew signal input
rlabel locali s 887 260 939 356 6 C_N
port 3 nsew signal input
rlabel locali s 25 270 110 356 6 D_N
port 4 nsew signal input
rlabel locali s 212 370 278 420 6 X
port 5 nsew signal output
rlabel locali s 212 236 246 370 6 X
port 5 nsew signal output
rlabel locali s 212 88 263 236 6 X
port 5 nsew signal output
rlabel metal1 s 0 -49 960 49 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 617 960 715 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1136710
string GDS_START 1128688
<< end >>
