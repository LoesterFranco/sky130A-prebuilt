magic
tech sky130A
magscale 1 2
timestamp 1604502701
<< nwell >>
rect -38 332 1574 704
<< pwell >>
rect 0 0 1536 49
<< scpmos >>
rect 86 368 116 592
rect 176 368 206 592
rect 266 368 296 592
rect 356 368 386 592
rect 446 368 476 592
rect 536 368 566 592
rect 626 368 656 592
rect 716 368 746 592
rect 806 368 836 592
rect 896 368 926 592
rect 986 368 1016 592
rect 1076 368 1106 592
rect 1270 424 1300 592
rect 1360 424 1390 592
<< nmoslvt >>
rect 99 74 129 222
rect 185 74 215 222
rect 271 74 301 222
rect 357 74 387 222
rect 443 74 473 222
rect 529 74 559 222
rect 615 74 645 222
rect 701 74 731 222
rect 897 74 927 222
rect 983 74 1013 222
rect 1069 74 1099 222
rect 1155 74 1185 222
rect 1241 74 1271 222
<< ndiff >>
rect 46 210 99 222
rect 46 176 54 210
rect 88 176 99 210
rect 46 120 99 176
rect 46 86 54 120
rect 88 86 99 120
rect 46 74 99 86
rect 129 207 185 222
rect 129 173 140 207
rect 174 173 185 207
rect 129 74 185 173
rect 215 120 271 222
rect 215 86 226 120
rect 260 86 271 120
rect 215 74 271 86
rect 301 207 357 222
rect 301 173 312 207
rect 346 173 357 207
rect 301 74 357 173
rect 387 162 443 222
rect 387 128 398 162
rect 432 128 443 162
rect 387 74 443 128
rect 473 116 529 222
rect 473 82 484 116
rect 518 82 529 116
rect 473 74 529 82
rect 559 162 615 222
rect 559 128 570 162
rect 604 128 615 162
rect 559 74 615 128
rect 645 116 701 222
rect 645 82 656 116
rect 690 82 701 116
rect 645 74 701 82
rect 731 162 784 222
rect 731 128 742 162
rect 776 128 784 162
rect 731 74 784 128
rect 844 160 897 222
rect 844 126 852 160
rect 886 126 897 160
rect 844 74 897 126
rect 927 210 983 222
rect 927 176 938 210
rect 972 176 983 210
rect 927 120 983 176
rect 927 86 938 120
rect 972 86 983 120
rect 927 74 983 86
rect 1013 146 1069 222
rect 1013 112 1024 146
rect 1058 112 1069 146
rect 1013 74 1069 112
rect 1099 210 1155 222
rect 1099 176 1110 210
rect 1144 176 1155 210
rect 1099 120 1155 176
rect 1099 86 1110 120
rect 1144 86 1155 120
rect 1099 74 1155 86
rect 1185 191 1241 222
rect 1185 157 1196 191
rect 1230 157 1241 191
rect 1185 116 1241 157
rect 1185 82 1196 116
rect 1230 82 1241 116
rect 1185 74 1241 82
rect 1271 210 1324 222
rect 1271 176 1282 210
rect 1316 176 1324 210
rect 1271 120 1324 176
rect 1271 86 1282 120
rect 1316 86 1324 120
rect 1271 74 1324 86
<< pdiff >>
rect 31 580 86 592
rect 31 546 39 580
rect 73 546 86 580
rect 31 510 86 546
rect 31 476 39 510
rect 73 476 86 510
rect 31 440 86 476
rect 31 406 39 440
rect 73 406 86 440
rect 31 368 86 406
rect 116 580 176 592
rect 116 546 129 580
rect 163 546 176 580
rect 116 508 176 546
rect 116 474 129 508
rect 163 474 176 508
rect 116 368 176 474
rect 206 580 266 592
rect 206 546 219 580
rect 253 546 266 580
rect 206 510 266 546
rect 206 476 219 510
rect 253 476 266 510
rect 206 440 266 476
rect 206 406 219 440
rect 253 406 266 440
rect 206 368 266 406
rect 296 580 356 592
rect 296 546 309 580
rect 343 546 356 580
rect 296 508 356 546
rect 296 474 309 508
rect 343 474 356 508
rect 296 368 356 474
rect 386 580 446 592
rect 386 546 399 580
rect 433 546 446 580
rect 386 497 446 546
rect 386 463 399 497
rect 433 463 446 497
rect 386 414 446 463
rect 386 380 399 414
rect 433 380 446 414
rect 386 368 446 380
rect 476 580 536 592
rect 476 546 489 580
rect 523 546 536 580
rect 476 508 536 546
rect 476 474 489 508
rect 523 474 536 508
rect 476 368 536 474
rect 566 580 626 592
rect 566 546 579 580
rect 613 546 626 580
rect 566 510 626 546
rect 566 476 579 510
rect 613 476 626 510
rect 566 440 626 476
rect 566 406 579 440
rect 613 406 626 440
rect 566 368 626 406
rect 656 580 716 592
rect 656 546 669 580
rect 703 546 716 580
rect 656 508 716 546
rect 656 474 669 508
rect 703 474 716 508
rect 656 368 716 474
rect 746 580 806 592
rect 746 546 759 580
rect 793 546 806 580
rect 746 510 806 546
rect 746 476 759 510
rect 793 476 806 510
rect 746 440 806 476
rect 746 406 759 440
rect 793 406 806 440
rect 746 368 806 406
rect 836 547 896 592
rect 836 513 849 547
rect 883 513 896 547
rect 836 479 896 513
rect 836 445 849 479
rect 883 445 896 479
rect 836 411 896 445
rect 836 377 849 411
rect 883 377 896 411
rect 836 368 896 377
rect 926 580 986 592
rect 926 546 939 580
rect 973 546 986 580
rect 926 482 986 546
rect 926 448 939 482
rect 973 448 986 482
rect 926 368 986 448
rect 1016 547 1076 592
rect 1016 513 1029 547
rect 1063 513 1076 547
rect 1016 479 1076 513
rect 1016 445 1029 479
rect 1063 445 1076 479
rect 1016 411 1076 445
rect 1016 377 1029 411
rect 1063 377 1076 411
rect 1016 368 1076 377
rect 1106 580 1161 592
rect 1106 546 1119 580
rect 1153 546 1161 580
rect 1106 497 1161 546
rect 1106 463 1119 497
rect 1153 463 1161 497
rect 1106 414 1161 463
rect 1215 574 1270 592
rect 1215 540 1223 574
rect 1257 540 1270 574
rect 1215 506 1270 540
rect 1215 472 1223 506
rect 1257 472 1270 506
rect 1215 424 1270 472
rect 1300 580 1360 592
rect 1300 546 1313 580
rect 1347 546 1360 580
rect 1300 470 1360 546
rect 1300 436 1313 470
rect 1347 436 1360 470
rect 1300 424 1360 436
rect 1390 580 1445 592
rect 1390 546 1403 580
rect 1437 546 1445 580
rect 1390 470 1445 546
rect 1390 436 1403 470
rect 1437 436 1445 470
rect 1390 424 1445 436
rect 1106 380 1119 414
rect 1153 380 1161 414
rect 1106 368 1161 380
<< ndiffc >>
rect 54 176 88 210
rect 54 86 88 120
rect 140 173 174 207
rect 226 86 260 120
rect 312 173 346 207
rect 398 128 432 162
rect 484 82 518 116
rect 570 128 604 162
rect 656 82 690 116
rect 742 128 776 162
rect 852 126 886 160
rect 938 176 972 210
rect 938 86 972 120
rect 1024 112 1058 146
rect 1110 176 1144 210
rect 1110 86 1144 120
rect 1196 157 1230 191
rect 1196 82 1230 116
rect 1282 176 1316 210
rect 1282 86 1316 120
<< pdiffc >>
rect 39 546 73 580
rect 39 476 73 510
rect 39 406 73 440
rect 129 546 163 580
rect 129 474 163 508
rect 219 546 253 580
rect 219 476 253 510
rect 219 406 253 440
rect 309 546 343 580
rect 309 474 343 508
rect 399 546 433 580
rect 399 463 433 497
rect 399 380 433 414
rect 489 546 523 580
rect 489 474 523 508
rect 579 546 613 580
rect 579 476 613 510
rect 579 406 613 440
rect 669 546 703 580
rect 669 474 703 508
rect 759 546 793 580
rect 759 476 793 510
rect 759 406 793 440
rect 849 513 883 547
rect 849 445 883 479
rect 849 377 883 411
rect 939 546 973 580
rect 939 448 973 482
rect 1029 513 1063 547
rect 1029 445 1063 479
rect 1029 377 1063 411
rect 1119 546 1153 580
rect 1119 463 1153 497
rect 1223 540 1257 574
rect 1223 472 1257 506
rect 1313 546 1347 580
rect 1313 436 1347 470
rect 1403 546 1437 580
rect 1403 436 1437 470
rect 1119 380 1153 414
<< poly >>
rect 86 592 116 618
rect 176 592 206 618
rect 266 592 296 618
rect 356 592 386 618
rect 446 592 476 618
rect 536 592 566 618
rect 626 592 656 618
rect 716 592 746 618
rect 806 592 836 618
rect 896 592 926 618
rect 986 592 1016 618
rect 1076 592 1106 618
rect 1270 592 1300 618
rect 1360 592 1390 618
rect 1270 409 1300 424
rect 1360 409 1390 424
rect 86 353 116 368
rect 176 353 206 368
rect 266 353 296 368
rect 356 353 386 368
rect 446 353 476 368
rect 536 353 566 368
rect 626 353 656 368
rect 716 353 746 368
rect 806 353 836 368
rect 896 353 926 368
rect 986 353 1016 368
rect 1076 353 1106 368
rect 1267 364 1303 409
rect 1357 364 1393 409
rect 83 336 119 353
rect 173 336 209 353
rect 263 336 299 353
rect 353 336 389 353
rect 83 320 389 336
rect 83 286 99 320
rect 133 286 167 320
rect 201 286 235 320
rect 269 286 303 320
rect 337 286 389 320
rect 83 270 389 286
rect 443 336 479 353
rect 533 336 569 353
rect 623 336 659 353
rect 713 336 746 353
rect 443 320 743 336
rect 803 330 929 353
rect 983 330 1019 353
rect 1073 330 1109 353
rect 1267 348 1393 364
rect 803 323 1185 330
rect 1267 328 1289 348
rect 443 286 489 320
rect 523 286 557 320
rect 591 286 625 320
rect 659 286 693 320
rect 727 286 743 320
rect 443 270 743 286
rect 897 314 1185 323
rect 897 300 999 314
rect 99 222 129 270
rect 185 222 215 270
rect 271 222 301 270
rect 357 222 387 270
rect 443 222 473 270
rect 529 222 559 270
rect 615 222 645 270
rect 701 222 731 270
rect 897 222 927 300
rect 983 280 999 300
rect 1033 280 1067 314
rect 1101 280 1135 314
rect 1169 280 1185 314
rect 983 264 1185 280
rect 983 222 1013 264
rect 1069 222 1099 264
rect 1155 222 1185 264
rect 1241 314 1289 328
rect 1323 314 1393 348
rect 1241 298 1393 314
rect 1241 222 1271 298
rect 99 48 129 74
rect 185 48 215 74
rect 271 48 301 74
rect 357 48 387 74
rect 443 48 473 74
rect 529 48 559 74
rect 615 48 645 74
rect 701 48 731 74
rect 897 48 927 74
rect 983 48 1013 74
rect 1069 48 1099 74
rect 1155 48 1185 74
rect 1241 48 1271 74
<< polycont >>
rect 99 286 133 320
rect 167 286 201 320
rect 235 286 269 320
rect 303 286 337 320
rect 489 286 523 320
rect 557 286 591 320
rect 625 286 659 320
rect 693 286 727 320
rect 999 280 1033 314
rect 1067 280 1101 314
rect 1135 280 1169 314
rect 1289 314 1323 348
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 23 580 73 596
rect 23 546 39 580
rect 23 510 73 546
rect 23 476 39 510
rect 23 440 73 476
rect 113 580 179 649
rect 113 546 129 580
rect 163 546 179 580
rect 113 508 179 546
rect 113 474 129 508
rect 163 474 179 508
rect 113 458 179 474
rect 219 580 253 596
rect 219 510 253 546
rect 23 406 39 440
rect 219 440 253 476
rect 293 580 359 649
rect 293 546 309 580
rect 343 546 359 580
rect 293 508 359 546
rect 293 474 309 508
rect 343 474 359 508
rect 293 458 359 474
rect 399 580 433 596
rect 399 497 433 546
rect 73 406 219 424
rect 399 424 433 463
rect 473 580 523 649
rect 473 546 489 580
rect 473 508 523 546
rect 473 474 489 508
rect 473 458 523 474
rect 563 580 629 596
rect 563 546 579 580
rect 613 546 629 580
rect 563 510 629 546
rect 563 476 579 510
rect 613 476 629 510
rect 563 440 629 476
rect 669 580 703 649
rect 669 508 703 546
rect 669 458 703 474
rect 743 581 1169 615
rect 743 580 799 581
rect 743 546 759 580
rect 793 546 799 580
rect 933 580 979 581
rect 743 510 799 546
rect 743 476 759 510
rect 793 476 799 510
rect 563 424 579 440
rect 253 414 579 424
rect 253 406 399 414
rect 23 390 399 406
rect 433 406 579 414
rect 613 424 629 440
rect 743 440 799 476
rect 743 424 759 440
rect 613 406 759 424
rect 793 406 799 440
rect 433 390 799 406
rect 833 513 849 547
rect 883 513 899 547
rect 833 479 899 513
rect 833 445 849 479
rect 883 445 899 479
rect 833 411 899 445
rect 933 546 939 580
rect 973 546 979 580
rect 1113 580 1169 581
rect 933 482 979 546
rect 933 448 939 482
rect 973 448 979 482
rect 933 432 979 448
rect 1013 513 1029 547
rect 1063 513 1079 547
rect 1013 479 1079 513
rect 1013 445 1029 479
rect 1063 445 1079 479
rect 399 364 433 380
rect 833 377 849 411
rect 883 398 899 411
rect 1013 411 1079 445
rect 1013 398 1029 411
rect 883 377 1029 398
rect 1063 377 1079 411
rect 833 364 1079 377
rect 1113 546 1119 580
rect 1153 546 1169 580
rect 1113 497 1169 546
rect 1113 463 1119 497
rect 1153 463 1169 497
rect 1207 574 1273 649
rect 1207 540 1223 574
rect 1257 540 1273 574
rect 1207 506 1273 540
rect 1207 472 1223 506
rect 1257 472 1273 506
rect 1207 466 1273 472
rect 1307 580 1363 596
rect 1307 546 1313 580
rect 1347 546 1363 580
rect 1307 470 1363 546
rect 1113 414 1169 463
rect 1307 436 1313 470
rect 1347 436 1363 470
rect 1307 432 1363 436
rect 1113 380 1119 414
rect 1153 380 1169 414
rect 1113 364 1169 380
rect 1205 398 1363 432
rect 1403 580 1453 649
rect 1437 546 1453 580
rect 1403 470 1453 546
rect 1437 436 1453 470
rect 1403 420 1453 436
rect 833 356 949 364
rect 25 320 359 356
rect 25 286 99 320
rect 133 286 167 320
rect 201 286 235 320
rect 269 286 303 320
rect 337 286 359 320
rect 473 320 743 356
rect 473 286 489 320
rect 523 286 557 320
rect 591 286 625 320
rect 659 286 693 320
rect 727 286 743 320
rect 793 252 949 356
rect 1205 330 1239 398
rect 983 314 1239 330
rect 983 280 999 314
rect 1033 280 1067 314
rect 1101 280 1135 314
rect 1169 280 1239 314
rect 1273 348 1511 364
rect 1273 314 1289 348
rect 1323 314 1511 348
rect 1273 298 1511 314
rect 983 264 1239 280
rect 296 230 949 252
rect 1205 230 1332 264
rect 38 210 104 226
rect 38 176 54 210
rect 88 176 104 210
rect 38 120 104 176
rect 140 207 190 226
rect 174 188 190 207
rect 296 218 1144 230
rect 296 207 362 218
rect 296 188 312 207
rect 174 173 312 188
rect 346 173 362 207
rect 915 210 1144 218
rect 915 196 938 210
rect 140 154 362 173
rect 398 162 792 184
rect 922 176 938 196
rect 972 196 1110 210
rect 432 150 570 162
rect 398 120 432 128
rect 38 86 54 120
rect 88 86 226 120
rect 260 86 432 120
rect 604 150 742 162
rect 38 70 432 86
rect 468 82 484 116
rect 518 82 534 116
rect 570 102 604 128
rect 776 128 792 162
rect 468 17 534 82
rect 640 82 656 116
rect 690 82 706 116
rect 742 102 792 128
rect 836 160 886 176
rect 836 126 852 160
rect 640 17 706 82
rect 836 17 886 126
rect 922 120 972 176
rect 1094 176 1110 196
rect 1280 210 1332 230
rect 922 86 938 120
rect 922 70 972 86
rect 1008 146 1058 162
rect 1008 112 1024 146
rect 1008 17 1058 112
rect 1094 120 1144 176
rect 1094 86 1110 120
rect 1094 70 1144 86
rect 1180 191 1246 196
rect 1180 157 1196 191
rect 1230 157 1246 191
rect 1180 116 1246 157
rect 1180 82 1196 116
rect 1230 82 1246 116
rect 1180 17 1246 82
rect 1280 176 1282 210
rect 1316 176 1332 210
rect 1280 120 1332 176
rect 1280 86 1282 120
rect 1316 86 1332 120
rect 1280 70 1332 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a21boi_4
flabel pwell s 0 0 1536 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 1536 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 1536 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 1536 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 1279 316 1313 350 0 FreeSans 340 0 0 0 B1_N
port 3 nsew
flabel corelocali s 1375 316 1409 350 0 FreeSans 340 0 0 0 B1_N
port 3 nsew
flabel corelocali s 1471 316 1505 350 0 FreeSans 340 0 0 0 B1_N
port 3 nsew
flabel corelocali s 799 242 833 276 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 895 242 929 276 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 1536 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 4097934
string GDS_START 4084966
<< end >>
