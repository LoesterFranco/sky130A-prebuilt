magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 552 561
rect 134 381 200 527
rect 305 265 351 491
rect 387 357 532 491
rect 19 153 87 265
rect 121 199 249 265
rect 285 199 351 265
rect 387 199 447 323
rect 17 17 85 119
rect 121 53 171 199
rect 489 163 532 357
rect 236 125 532 163
rect 236 53 273 125
rect 309 17 375 91
rect 411 53 456 125
rect 0 -17 552 17
<< obsli1 >>
rect 50 345 100 491
rect 234 345 271 491
rect 50 305 271 345
<< metal1 >>
rect 0 496 552 592
rect 0 -48 552 48
<< labels >>
rlabel locali s 121 199 249 265 6 A1
port 1 nsew signal input
rlabel locali s 121 53 171 199 6 A1
port 1 nsew signal input
rlabel locali s 19 153 87 265 6 A2
port 2 nsew signal input
rlabel locali s 305 265 351 491 6 B1
port 3 nsew signal input
rlabel locali s 285 199 351 265 6 B1
port 3 nsew signal input
rlabel locali s 387 199 447 323 6 C1
port 4 nsew signal input
rlabel locali s 489 163 532 357 6 Y
port 5 nsew signal output
rlabel locali s 411 53 456 125 6 Y
port 5 nsew signal output
rlabel locali s 387 357 532 491 6 Y
port 5 nsew signal output
rlabel locali s 236 125 532 163 6 Y
port 5 nsew signal output
rlabel locali s 236 53 273 125 6 Y
port 5 nsew signal output
rlabel locali s 309 17 375 91 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 17 17 85 119 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 552 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 552 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 134 381 200 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 552 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 552 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 552 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3955922
string GDS_START 3949274
<< end >>
