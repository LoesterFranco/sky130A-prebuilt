magic
tech sky130A
magscale 1 2
timestamp 1601050039
<< nwell >>
rect -38 261 1326 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 96 47 126 177
rect 180 47 210 177
rect 264 47 294 177
rect 348 47 378 177
rect 536 47 566 177
rect 620 47 650 177
rect 704 47 734 177
rect 788 47 818 177
rect 888 47 918 177
rect 972 47 1002 177
rect 1056 47 1086 177
rect 1140 47 1170 177
<< pmoshvt >>
rect 96 297 126 497
rect 180 297 210 497
rect 264 297 294 497
rect 348 297 378 497
rect 536 297 566 497
rect 620 297 650 497
rect 704 297 734 497
rect 788 297 818 497
rect 888 297 918 497
rect 972 297 1002 497
rect 1056 297 1086 497
rect 1140 297 1170 497
<< ndiff >>
rect 40 95 96 177
rect 40 61 52 95
rect 86 61 96 95
rect 40 47 96 61
rect 126 163 180 177
rect 126 129 136 163
rect 170 129 180 163
rect 126 95 180 129
rect 126 61 136 95
rect 170 61 180 95
rect 126 47 180 61
rect 210 95 264 177
rect 210 61 220 95
rect 254 61 264 95
rect 210 47 264 61
rect 294 163 348 177
rect 294 129 304 163
rect 338 129 348 163
rect 294 95 348 129
rect 294 61 304 95
rect 338 61 348 95
rect 294 47 348 61
rect 378 95 536 177
rect 378 61 388 95
rect 422 61 492 95
rect 526 61 536 95
rect 378 47 536 61
rect 566 95 620 177
rect 566 61 576 95
rect 610 61 620 95
rect 566 47 620 61
rect 650 163 704 177
rect 650 129 660 163
rect 694 129 704 163
rect 650 47 704 129
rect 734 95 788 177
rect 734 61 744 95
rect 778 61 788 95
rect 734 47 788 61
rect 818 95 888 177
rect 818 61 837 95
rect 871 61 888 95
rect 818 47 888 61
rect 918 95 972 177
rect 918 61 928 95
rect 962 61 972 95
rect 918 47 972 61
rect 1002 163 1056 177
rect 1002 129 1012 163
rect 1046 129 1056 163
rect 1002 47 1056 129
rect 1086 163 1140 177
rect 1086 129 1096 163
rect 1130 129 1140 163
rect 1086 95 1140 129
rect 1086 61 1096 95
rect 1130 61 1140 95
rect 1086 47 1140 61
rect 1170 163 1222 177
rect 1170 129 1180 163
rect 1214 129 1222 163
rect 1170 95 1222 129
rect 1170 61 1180 95
rect 1214 61 1222 95
rect 1170 47 1222 61
<< pdiff >>
rect 40 483 96 497
rect 40 449 52 483
rect 86 449 96 483
rect 40 415 96 449
rect 40 381 52 415
rect 86 381 96 415
rect 40 297 96 381
rect 126 477 180 497
rect 126 443 136 477
rect 170 443 180 477
rect 126 409 180 443
rect 126 375 136 409
rect 170 375 180 409
rect 126 341 180 375
rect 126 307 136 341
rect 170 307 180 341
rect 126 297 180 307
rect 210 483 264 497
rect 210 449 220 483
rect 254 449 264 483
rect 210 415 264 449
rect 210 381 220 415
rect 254 381 264 415
rect 210 297 264 381
rect 294 477 348 497
rect 294 443 304 477
rect 338 443 348 477
rect 294 409 348 443
rect 294 375 304 409
rect 338 375 348 409
rect 294 341 348 375
rect 294 307 304 341
rect 338 307 348 341
rect 294 297 348 307
rect 378 477 430 497
rect 378 443 388 477
rect 422 443 430 477
rect 378 297 430 443
rect 484 477 536 497
rect 484 443 492 477
rect 526 443 536 477
rect 484 297 536 443
rect 566 409 620 497
rect 566 375 576 409
rect 610 375 620 409
rect 566 297 620 375
rect 650 477 704 497
rect 650 443 660 477
rect 694 443 704 477
rect 650 297 704 443
rect 734 409 788 497
rect 734 375 744 409
rect 778 375 788 409
rect 734 297 788 375
rect 818 477 888 497
rect 818 443 835 477
rect 869 443 888 477
rect 818 409 888 443
rect 818 375 835 409
rect 869 375 888 409
rect 818 297 888 375
rect 918 477 972 497
rect 918 443 928 477
rect 962 443 972 477
rect 918 297 972 443
rect 1002 477 1056 497
rect 1002 443 1012 477
rect 1046 443 1056 477
rect 1002 409 1056 443
rect 1002 375 1012 409
rect 1046 375 1056 409
rect 1002 297 1056 375
rect 1086 477 1140 497
rect 1086 443 1096 477
rect 1130 443 1140 477
rect 1086 297 1140 443
rect 1170 477 1227 497
rect 1170 443 1181 477
rect 1215 443 1227 477
rect 1170 409 1227 443
rect 1170 375 1181 409
rect 1215 375 1227 409
rect 1170 341 1227 375
rect 1170 307 1181 341
rect 1215 307 1227 341
rect 1170 297 1227 307
<< ndiffc >>
rect 52 61 86 95
rect 136 129 170 163
rect 136 61 170 95
rect 220 61 254 95
rect 304 129 338 163
rect 304 61 338 95
rect 388 61 422 95
rect 492 61 526 95
rect 576 61 610 95
rect 660 129 694 163
rect 744 61 778 95
rect 837 61 871 95
rect 928 61 962 95
rect 1012 129 1046 163
rect 1096 129 1130 163
rect 1096 61 1130 95
rect 1180 129 1214 163
rect 1180 61 1214 95
<< pdiffc >>
rect 52 449 86 483
rect 52 381 86 415
rect 136 443 170 477
rect 136 375 170 409
rect 136 307 170 341
rect 220 449 254 483
rect 220 381 254 415
rect 304 443 338 477
rect 304 375 338 409
rect 304 307 338 341
rect 388 443 422 477
rect 492 443 526 477
rect 576 375 610 409
rect 660 443 694 477
rect 744 375 778 409
rect 835 443 869 477
rect 835 375 869 409
rect 928 443 962 477
rect 1012 443 1046 477
rect 1012 375 1046 409
rect 1096 443 1130 477
rect 1181 443 1215 477
rect 1181 375 1215 409
rect 1181 307 1215 341
<< poly >>
rect 96 497 126 523
rect 180 497 210 523
rect 264 497 294 523
rect 348 497 378 523
rect 536 497 566 523
rect 620 497 650 523
rect 704 497 734 523
rect 788 497 818 523
rect 888 497 918 523
rect 972 497 1002 523
rect 1056 497 1086 523
rect 1140 497 1170 523
rect 96 265 126 297
rect 180 265 210 297
rect 264 265 294 297
rect 348 265 378 297
rect 536 265 566 297
rect 620 265 650 297
rect 704 265 734 297
rect 788 265 818 297
rect 888 265 918 297
rect 972 265 1002 297
rect 1056 265 1086 297
rect 1140 265 1170 297
rect 96 249 378 265
rect 96 215 124 249
rect 158 215 192 249
rect 226 215 260 249
rect 294 215 328 249
rect 362 215 378 249
rect 96 199 378 215
rect 524 249 578 265
rect 524 215 534 249
rect 568 215 578 249
rect 524 199 578 215
rect 620 249 734 265
rect 620 215 660 249
rect 694 215 734 249
rect 620 199 734 215
rect 776 249 830 265
rect 776 215 786 249
rect 820 215 830 249
rect 776 199 830 215
rect 876 249 930 265
rect 876 215 886 249
rect 920 215 930 249
rect 876 199 930 215
rect 972 249 1086 265
rect 972 215 1012 249
rect 1046 215 1086 249
rect 972 199 1086 215
rect 1128 249 1182 265
rect 1128 215 1138 249
rect 1172 215 1182 249
rect 1128 199 1182 215
rect 96 177 126 199
rect 180 177 210 199
rect 264 177 294 199
rect 348 177 378 199
rect 536 177 566 199
rect 620 177 650 199
rect 704 177 734 199
rect 788 177 818 199
rect 888 177 918 199
rect 972 177 1002 199
rect 1056 177 1086 199
rect 1140 177 1170 199
rect 96 21 126 47
rect 180 21 210 47
rect 264 21 294 47
rect 348 21 378 47
rect 536 21 566 47
rect 620 21 650 47
rect 704 21 734 47
rect 788 21 818 47
rect 888 21 918 47
rect 972 21 1002 47
rect 1056 21 1086 47
rect 1140 21 1170 47
<< polycont >>
rect 124 215 158 249
rect 192 215 226 249
rect 260 215 294 249
rect 328 215 362 249
rect 534 215 568 249
rect 660 215 694 249
rect 786 215 820 249
rect 886 215 920 249
rect 1012 215 1046 249
rect 1138 215 1172 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 44 483 94 527
rect 44 449 52 483
rect 86 449 94 483
rect 44 415 94 449
rect 44 381 52 415
rect 86 381 94 415
rect 44 365 94 381
rect 128 477 178 493
rect 128 443 136 477
rect 170 443 178 477
rect 128 409 178 443
rect 128 375 136 409
rect 170 375 178 409
rect 128 341 178 375
rect 212 483 262 527
rect 212 449 220 483
rect 254 449 262 483
rect 212 415 262 449
rect 212 381 220 415
rect 254 381 262 415
rect 212 359 262 381
rect 296 477 346 493
rect 296 443 304 477
rect 338 443 346 477
rect 296 409 346 443
rect 380 477 430 527
rect 380 443 388 477
rect 422 443 430 477
rect 380 425 430 443
rect 484 477 886 493
rect 484 443 492 477
rect 526 459 660 477
rect 526 443 534 459
rect 484 425 534 443
rect 652 443 660 459
rect 694 459 835 477
rect 694 443 702 459
rect 652 425 702 443
rect 820 443 835 459
rect 869 443 886 477
rect 296 375 304 409
rect 338 375 346 409
rect 568 409 618 425
rect 568 391 576 409
rect 128 323 136 341
rect 17 307 136 323
rect 170 323 178 341
rect 296 341 346 375
rect 296 323 304 341
rect 170 307 304 323
rect 338 307 346 341
rect 17 289 346 307
rect 380 375 576 391
rect 610 391 618 409
rect 736 409 786 425
rect 736 391 744 409
rect 610 375 744 391
rect 778 375 786 409
rect 380 357 786 375
rect 820 409 886 443
rect 920 477 970 527
rect 920 443 928 477
rect 962 443 970 477
rect 920 425 970 443
rect 1004 477 1054 493
rect 1004 443 1012 477
rect 1046 443 1054 477
rect 820 375 835 409
rect 869 391 886 409
rect 1004 409 1054 443
rect 1088 477 1138 527
rect 1088 443 1096 477
rect 1130 443 1138 477
rect 1088 425 1138 443
rect 1181 477 1222 493
rect 1215 443 1222 477
rect 1004 391 1012 409
rect 869 375 1012 391
rect 1046 391 1054 409
rect 1181 409 1222 443
rect 1046 375 1181 391
rect 1215 375 1222 409
rect 820 357 1222 375
rect 17 181 74 289
rect 380 255 446 357
rect 1181 341 1222 357
rect 108 249 446 255
rect 108 215 124 249
rect 158 215 192 249
rect 226 215 260 249
rect 294 215 328 249
rect 362 215 446 249
rect 484 289 836 323
rect 484 249 591 289
rect 484 215 534 249
rect 568 215 591 249
rect 625 249 736 255
rect 625 215 660 249
rect 694 215 736 249
rect 770 249 836 289
rect 770 215 786 249
rect 820 215 836 249
rect 870 289 1147 323
rect 1215 307 1222 341
rect 1181 291 1222 307
rect 870 249 936 289
rect 1113 255 1147 289
rect 870 215 886 249
rect 920 215 936 249
rect 980 249 1079 255
rect 980 215 1012 249
rect 1046 215 1079 249
rect 1113 249 1271 255
rect 1113 215 1138 249
rect 1172 215 1271 249
rect 388 181 446 215
rect 17 163 354 181
rect 17 145 136 163
rect 120 129 136 145
rect 170 145 304 163
rect 170 129 186 145
rect 52 95 86 111
rect 52 17 86 61
rect 120 95 186 129
rect 288 129 304 145
rect 338 129 354 163
rect 388 163 1062 181
rect 388 147 660 163
rect 634 129 660 147
rect 694 147 1012 163
rect 694 129 721 147
rect 987 129 1012 147
rect 1046 129 1062 163
rect 1096 163 1146 179
rect 1130 129 1146 163
rect 120 61 136 95
rect 170 61 186 95
rect 120 53 186 61
rect 220 95 254 111
rect 220 17 254 61
rect 288 95 354 129
rect 288 61 304 95
rect 338 61 354 95
rect 288 51 354 61
rect 388 95 526 111
rect 837 95 871 111
rect 1096 95 1146 129
rect 422 61 492 95
rect 388 17 526 61
rect 560 61 576 95
rect 610 61 744 95
rect 778 61 794 95
rect 560 51 794 61
rect 837 17 871 61
rect 912 61 928 95
rect 962 61 1096 95
rect 1130 61 1146 95
rect 912 51 1146 61
rect 1180 163 1214 179
rect 1180 95 1214 129
rect 1180 17 1214 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
flabel corelocali s 677 221 711 255 0 FreeSans 400 0 0 0 B1
port 3 nsew
flabel corelocali s 493 221 527 255 0 FreeSans 400 0 0 0 B2
port 4 nsew
flabel corelocali s 29 221 63 255 0 FreeSans 400 0 0 0 X
port 9 nsew
flabel corelocali s 1225 221 1259 255 0 FreeSans 400 180 0 0 A2
port 2 nsew
flabel corelocali s 1045 221 1079 255 0 FreeSans 400 180 0 0 A1
port 1 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
rlabel comment s 0 0 0 0 4 a22o_4
<< properties >>
string FIXED_BBOX 0 0 1288 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 4151268
string GDS_START 4141594
string path 0.000 0.000 32.200 0.000 
<< end >>
