magic
tech sky130A
magscale 1 2
timestamp 1601050058
<< locali >>
rect 119 401 153 493
rect 18 367 153 401
rect 18 177 69 367
rect 213 199 279 265
rect 325 249 359 252
rect 325 215 391 249
rect 18 143 153 177
rect 213 152 254 199
rect 325 173 359 215
rect 437 174 471 265
rect 119 51 153 143
rect 306 139 359 173
rect 393 140 471 174
rect 306 80 340 139
rect 393 83 435 140
rect 579 151 618 265
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 27 435 77 527
rect 187 367 237 527
rect 271 401 321 485
rect 363 435 429 527
rect 467 401 517 485
rect 271 367 529 401
rect 575 333 609 493
rect 111 299 609 333
rect 111 249 145 299
rect 111 215 177 249
rect 18 17 69 109
rect 203 93 237 109
rect 191 17 257 93
rect 507 101 541 299
rect 475 67 541 101
rect 492 51 541 67
rect 575 17 627 113
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 437 174 471 265 6 A1
port 1 nsew signal input
rlabel locali s 393 140 471 174 6 A1
port 1 nsew signal input
rlabel locali s 393 83 435 140 6 A1
port 1 nsew signal input
rlabel locali s 325 249 359 252 6 A2
port 2 nsew signal input
rlabel locali s 325 215 391 249 6 A2
port 2 nsew signal input
rlabel locali s 325 173 359 215 6 A2
port 2 nsew signal input
rlabel locali s 306 139 359 173 6 A2
port 2 nsew signal input
rlabel locali s 306 80 340 139 6 A2
port 2 nsew signal input
rlabel locali s 213 199 279 265 6 A3
port 3 nsew signal input
rlabel locali s 213 152 254 199 6 A3
port 3 nsew signal input
rlabel locali s 579 151 618 265 6 B1
port 4 nsew signal input
rlabel locali s 119 401 153 493 6 X
port 5 nsew signal output
rlabel locali s 119 51 153 143 6 X
port 5 nsew signal output
rlabel locali s 18 367 153 401 6 X
port 5 nsew signal output
rlabel locali s 18 177 69 367 6 X
port 5 nsew signal output
rlabel locali s 18 143 153 177 6 X
port 5 nsew signal output
rlabel metal1 s 0 -48 644 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3562758
string GDS_START 3556270
<< end >>
