magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 828 561
rect 87 297 121 527
rect 255 367 303 527
rect 56 215 237 263
rect 339 323 373 493
rect 407 367 473 527
rect 507 323 541 493
rect 575 367 641 527
rect 675 323 709 493
rect 339 289 709 323
rect 743 297 809 527
rect 442 181 709 289
rect 339 147 709 181
rect 87 17 121 113
rect 255 17 289 113
rect 339 51 373 147
rect 407 17 473 113
rect 507 51 541 147
rect 575 17 641 113
rect 675 51 709 147
rect 743 17 809 177
rect 0 -17 828 17
<< obsli1 >>
rect 155 331 221 493
rect 155 297 305 331
rect 271 249 305 297
rect 271 215 365 249
rect 271 181 305 215
rect 155 147 305 181
rect 155 51 221 147
<< metal1 >>
rect 0 496 828 592
rect 0 -48 828 48
<< labels >>
rlabel locali s 56 215 237 263 6 A
port 1 nsew signal input
rlabel locali s 675 323 709 493 6 X
port 2 nsew signal output
rlabel locali s 675 51 709 147 6 X
port 2 nsew signal output
rlabel locali s 507 323 541 493 6 X
port 2 nsew signal output
rlabel locali s 507 51 541 147 6 X
port 2 nsew signal output
rlabel locali s 442 181 709 289 6 X
port 2 nsew signal output
rlabel locali s 339 323 373 493 6 X
port 2 nsew signal output
rlabel locali s 339 289 709 323 6 X
port 2 nsew signal output
rlabel locali s 339 147 709 181 6 X
port 2 nsew signal output
rlabel locali s 339 51 373 147 6 X
port 2 nsew signal output
rlabel locali s 743 17 809 177 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 575 17 641 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 407 17 473 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 255 17 289 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 87 17 121 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 0 -17 828 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 828 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 743 297 809 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 575 367 641 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 407 367 473 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 255 367 303 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 87 297 121 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 0 527 828 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 496 828 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3048374
string GDS_START 3041396
<< end >>
