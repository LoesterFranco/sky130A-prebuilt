magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 1369 424 1435 547
rect 1549 424 1615 547
rect 889 390 1615 424
rect 25 270 349 356
rect 483 270 839 356
rect 889 236 938 390
rect 985 270 1223 356
rect 1273 270 1703 356
rect 889 226 1705 236
rect 870 202 1705 226
rect 870 193 1168 202
rect 870 154 937 193
rect 1102 119 1168 193
rect 1302 70 1368 202
rect 1639 70 1705 202
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 23 424 79 596
rect 113 458 179 649
rect 213 424 259 587
rect 293 458 359 649
rect 393 430 439 590
rect 473 464 539 649
rect 573 430 639 596
rect 673 458 739 649
rect 773 492 839 596
rect 873 526 939 649
rect 973 492 1135 586
rect 1169 526 1235 649
rect 1269 581 1705 615
rect 1269 492 1335 581
rect 773 458 1335 492
rect 393 424 639 430
rect 773 424 839 458
rect 1475 458 1515 581
rect 23 390 839 424
rect 1651 390 1705 581
rect 383 364 449 390
rect 26 202 824 236
rect 26 70 76 202
rect 112 17 178 168
rect 214 70 248 202
rect 284 17 350 168
rect 384 66 434 202
rect 470 85 531 168
rect 565 119 624 202
rect 658 85 724 168
rect 758 119 824 202
rect 987 85 1053 159
rect 1202 85 1268 168
rect 470 51 1268 85
rect 1402 17 1605 168
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
<< metal1 >>
rect 0 683 1728 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 0 617 1728 649
rect 0 17 1728 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
rect 0 -49 1728 -17
<< labels >>
rlabel locali s 985 270 1223 356 6 A1
port 1 nsew signal input
rlabel locali s 483 270 839 356 6 A2
port 2 nsew signal input
rlabel locali s 25 270 349 356 6 A3
port 3 nsew signal input
rlabel locali s 1273 270 1703 356 6 B1
port 4 nsew signal input
rlabel locali s 1639 70 1705 202 6 Y
port 5 nsew signal output
rlabel locali s 1549 424 1615 547 6 Y
port 5 nsew signal output
rlabel locali s 1369 424 1435 547 6 Y
port 5 nsew signal output
rlabel locali s 1302 70 1368 202 6 Y
port 5 nsew signal output
rlabel locali s 1102 119 1168 193 6 Y
port 5 nsew signal output
rlabel locali s 889 390 1615 424 6 Y
port 5 nsew signal output
rlabel locali s 889 236 938 390 6 Y
port 5 nsew signal output
rlabel locali s 889 226 1705 236 6 Y
port 5 nsew signal output
rlabel locali s 870 202 1705 226 6 Y
port 5 nsew signal output
rlabel locali s 870 193 1168 202 6 Y
port 5 nsew signal output
rlabel locali s 870 154 937 193 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -49 1728 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 1728 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1728 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3865218
string GDS_START 3851158
<< end >>
