magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 614 704
<< pwell >>
rect 0 0 576 49
<< scnmos >>
rect 91 136 121 264
rect 203 136 233 264
rect 298 120 328 248
rect 414 100 444 248
<< pmoshvt >>
rect 86 398 116 566
rect 196 398 226 566
rect 286 398 316 566
rect 460 368 490 592
<< ndiff >>
rect 34 210 91 264
rect 34 176 46 210
rect 80 176 91 210
rect 34 136 91 176
rect 121 136 203 264
rect 233 248 283 264
rect 233 136 298 248
rect 248 120 298 136
rect 328 230 414 248
rect 328 196 355 230
rect 389 196 414 230
rect 328 146 414 196
rect 328 120 355 146
rect 343 112 355 120
rect 389 112 414 146
rect 343 100 414 112
rect 444 220 501 248
rect 444 186 455 220
rect 489 186 501 220
rect 444 146 501 186
rect 444 112 455 146
rect 489 112 501 146
rect 444 100 501 112
<< pdiff >>
rect 334 566 460 592
rect 27 554 86 566
rect 27 520 39 554
rect 73 520 86 554
rect 27 444 86 520
rect 27 410 39 444
rect 73 410 86 444
rect 27 398 86 410
rect 116 508 196 566
rect 116 474 139 508
rect 173 474 196 508
rect 116 398 196 474
rect 226 554 286 566
rect 226 520 239 554
rect 273 520 286 554
rect 226 444 286 520
rect 226 410 239 444
rect 273 410 286 444
rect 226 398 286 410
rect 316 560 460 566
rect 316 526 341 560
rect 375 526 412 560
rect 446 526 460 560
rect 316 492 460 526
rect 316 458 330 492
rect 364 458 412 492
rect 446 458 460 492
rect 316 398 460 458
rect 407 368 460 398
rect 490 580 549 592
rect 490 546 503 580
rect 537 546 549 580
rect 490 500 549 546
rect 490 466 503 500
rect 537 466 549 500
rect 490 420 549 466
rect 490 386 503 420
rect 537 386 549 420
rect 490 368 549 386
<< ndiffc >>
rect 46 176 80 210
rect 355 196 389 230
rect 355 112 389 146
rect 455 186 489 220
rect 455 112 489 146
<< pdiffc >>
rect 39 520 73 554
rect 39 410 73 444
rect 139 474 173 508
rect 239 520 273 554
rect 239 410 273 444
rect 341 526 375 560
rect 412 526 446 560
rect 330 458 364 492
rect 412 458 446 492
rect 503 546 537 580
rect 503 466 537 500
rect 503 386 537 420
<< poly >>
rect 460 592 490 618
rect 86 566 116 592
rect 196 566 226 592
rect 286 566 316 592
rect 86 383 116 398
rect 196 383 226 398
rect 286 383 316 398
rect 83 309 119 383
rect 193 352 229 383
rect 283 356 319 383
rect 169 336 235 352
rect 83 279 121 309
rect 169 302 185 336
rect 219 302 235 336
rect 169 286 235 302
rect 283 340 363 356
rect 460 353 490 368
rect 283 306 313 340
rect 347 306 363 340
rect 457 336 493 353
rect 283 290 363 306
rect 414 320 493 336
rect 91 264 121 279
rect 203 264 233 286
rect 298 248 328 290
rect 414 286 430 320
rect 464 286 493 320
rect 414 270 493 286
rect 414 248 444 270
rect 91 114 121 136
rect 21 98 155 114
rect 203 110 233 136
rect 21 64 37 98
rect 71 64 105 98
rect 139 64 155 98
rect 298 94 328 120
rect 414 74 444 100
rect 21 48 155 64
<< polycont >>
rect 185 302 219 336
rect 313 306 347 340
rect 430 286 464 320
rect 37 64 71 98
rect 105 64 139 98
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 23 554 89 570
rect 23 520 39 554
rect 73 520 89 554
rect 23 444 89 520
rect 123 508 189 649
rect 123 474 139 508
rect 173 474 189 508
rect 123 458 189 474
rect 223 554 280 570
rect 223 520 239 554
rect 273 520 280 554
rect 23 410 39 444
rect 73 424 89 444
rect 223 444 280 520
rect 314 560 462 649
rect 314 526 341 560
rect 375 526 412 560
rect 446 526 462 560
rect 314 492 462 526
rect 314 458 330 492
rect 364 458 412 492
rect 446 458 462 492
rect 496 580 553 596
rect 496 546 503 580
rect 537 546 553 580
rect 496 500 553 546
rect 496 466 503 500
rect 537 466 553 500
rect 223 424 239 444
rect 73 410 239 424
rect 273 424 280 444
rect 273 410 448 424
rect 23 390 448 410
rect 23 210 96 390
rect 169 336 263 356
rect 169 302 185 336
rect 219 302 263 336
rect 169 236 263 302
rect 297 340 363 356
rect 297 306 313 340
rect 347 306 363 340
rect 297 290 363 306
rect 414 336 448 390
rect 496 420 553 466
rect 496 386 503 420
rect 537 386 553 420
rect 496 370 553 386
rect 414 320 480 336
rect 414 286 430 320
rect 464 286 480 320
rect 414 270 480 286
rect 519 236 553 370
rect 23 176 46 210
rect 80 176 96 210
rect 23 148 96 176
rect 339 230 405 236
rect 339 196 355 230
rect 389 196 405 230
rect 339 146 405 196
rect 217 114 263 134
rect 21 98 263 114
rect 21 64 37 98
rect 71 64 105 98
rect 139 64 263 98
rect 21 51 263 64
rect 339 112 355 146
rect 389 112 405 146
rect 339 17 405 112
rect 439 220 553 236
rect 439 186 455 220
rect 489 202 553 220
rect 489 186 505 202
rect 439 146 505 186
rect 439 112 455 146
rect 489 112 505 146
rect 439 96 505 112
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
rlabel comment s 0 0 0 0 4 and3_1
flabel pwell s 0 0 576 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 576 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 576 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 576 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 223 94 257 128 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 223 242 257 276 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 511 390 545 424 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 511 464 545 498 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 511 538 545 572 0 FreeSans 340 0 0 0 X
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 576 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3875928
string GDS_START 3869962
<< end >>
