magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 1862 704
rect 127 311 1183 332
<< pwell >>
rect 0 0 1824 49
<< scnmos >>
rect 84 79 114 227
rect 213 79 243 227
rect 357 79 387 227
rect 457 79 487 227
rect 535 79 565 227
rect 671 79 701 227
rect 757 79 787 227
rect 875 79 905 227
rect 989 79 1019 227
rect 1089 79 1119 227
rect 1175 79 1205 227
rect 1253 79 1283 227
rect 1396 79 1426 227
rect 1482 79 1512 227
rect 1624 79 1654 227
rect 1710 79 1740 227
<< pmoshvt >>
rect 86 378 116 578
rect 216 347 246 547
rect 306 347 336 547
rect 454 347 484 547
rect 538 347 568 547
rect 653 347 683 547
rect 754 378 784 578
rect 872 347 902 547
rect 962 347 992 547
rect 1064 347 1094 547
rect 1172 368 1202 568
rect 1256 368 1286 568
rect 1370 368 1400 592
rect 1479 368 1509 592
rect 1617 368 1647 592
rect 1707 368 1737 592
<< ndiff >>
rect 27 210 84 227
rect 27 176 39 210
rect 73 176 84 210
rect 27 125 84 176
rect 27 91 39 125
rect 73 91 84 125
rect 27 79 84 91
rect 114 128 213 227
rect 114 94 139 128
rect 173 94 213 128
rect 114 79 213 94
rect 243 134 357 227
rect 243 100 283 134
rect 317 100 357 134
rect 243 79 357 100
rect 387 202 457 227
rect 387 168 412 202
rect 446 168 457 202
rect 387 125 457 168
rect 387 91 412 125
rect 446 91 457 125
rect 387 79 457 91
rect 487 79 535 227
rect 565 125 671 227
rect 565 91 594 125
rect 628 91 671 125
rect 565 79 671 91
rect 701 129 757 227
rect 701 95 712 129
rect 746 95 757 129
rect 701 79 757 95
rect 787 82 875 227
rect 787 79 814 82
rect 802 48 814 79
rect 848 79 875 82
rect 905 134 989 227
rect 905 100 930 134
rect 964 100 989 134
rect 905 79 989 100
rect 1019 129 1089 227
rect 1019 95 1044 129
rect 1078 95 1089 129
rect 1019 79 1089 95
rect 1119 79 1175 227
rect 1205 79 1253 227
rect 1283 81 1396 227
rect 1283 79 1322 81
rect 848 48 860 79
rect 802 36 860 48
rect 1298 47 1322 79
rect 1356 79 1396 81
rect 1426 217 1482 227
rect 1426 183 1437 217
rect 1471 183 1482 217
rect 1426 79 1482 183
rect 1512 81 1624 227
rect 1512 79 1551 81
rect 1356 47 1381 79
rect 1298 36 1381 47
rect 1527 47 1551 79
rect 1585 79 1624 81
rect 1654 214 1710 227
rect 1654 180 1665 214
rect 1699 180 1710 214
rect 1654 125 1710 180
rect 1654 91 1665 125
rect 1699 91 1710 125
rect 1654 79 1710 91
rect 1740 215 1797 227
rect 1740 181 1751 215
rect 1785 181 1797 215
rect 1740 125 1797 181
rect 1740 91 1751 125
rect 1785 91 1797 125
rect 1740 79 1797 91
rect 1585 47 1609 79
rect 1527 36 1609 47
<< pdiff >>
rect 27 566 86 578
rect 27 532 39 566
rect 73 532 86 566
rect 27 498 86 532
rect 27 464 39 498
rect 73 464 86 498
rect 27 424 86 464
rect 27 390 35 424
rect 69 390 86 424
rect 27 378 86 390
rect 116 566 198 578
rect 116 532 145 566
rect 179 547 198 566
rect 701 547 754 578
rect 179 532 216 547
rect 116 378 216 532
rect 163 347 216 378
rect 246 535 306 547
rect 246 501 259 535
rect 293 501 306 535
rect 246 467 306 501
rect 246 433 259 467
rect 293 433 306 467
rect 246 347 306 433
rect 336 508 454 547
rect 336 474 383 508
rect 417 474 454 508
rect 336 347 454 474
rect 484 347 538 547
rect 568 508 653 547
rect 568 474 581 508
rect 615 474 653 508
rect 568 347 653 474
rect 683 514 754 547
rect 683 480 697 514
rect 731 480 754 514
rect 683 378 754 480
rect 784 566 854 578
rect 784 532 802 566
rect 836 547 854 566
rect 1311 573 1370 592
rect 1311 568 1323 573
rect 1119 547 1172 568
rect 836 532 872 547
rect 784 378 872 532
rect 683 347 736 378
rect 819 347 872 378
rect 902 505 962 547
rect 902 471 915 505
rect 949 471 962 505
rect 902 347 962 471
rect 992 535 1064 547
rect 992 501 1017 535
rect 1051 501 1064 535
rect 992 456 1064 501
rect 992 422 1017 456
rect 1051 422 1064 456
rect 992 347 1064 422
rect 1094 368 1172 547
rect 1202 368 1256 568
rect 1286 539 1323 568
rect 1357 539 1370 573
rect 1286 368 1370 539
rect 1400 414 1479 592
rect 1400 380 1422 414
rect 1456 380 1479 414
rect 1400 368 1479 380
rect 1509 580 1617 592
rect 1509 546 1541 580
rect 1575 546 1617 580
rect 1509 368 1617 546
rect 1647 580 1707 592
rect 1647 546 1660 580
rect 1694 546 1707 580
rect 1647 497 1707 546
rect 1647 463 1660 497
rect 1694 463 1707 497
rect 1647 414 1707 463
rect 1647 380 1660 414
rect 1694 380 1707 414
rect 1647 368 1707 380
rect 1737 580 1796 592
rect 1737 546 1750 580
rect 1784 546 1796 580
rect 1737 497 1796 546
rect 1737 463 1750 497
rect 1784 463 1796 497
rect 1737 414 1796 463
rect 1737 380 1750 414
rect 1784 380 1796 414
rect 1737 368 1796 380
rect 1094 347 1147 368
<< ndiffc >>
rect 39 176 73 210
rect 39 91 73 125
rect 139 94 173 128
rect 283 100 317 134
rect 412 168 446 202
rect 412 91 446 125
rect 594 91 628 125
rect 712 95 746 129
rect 814 48 848 82
rect 930 100 964 134
rect 1044 95 1078 129
rect 1322 47 1356 81
rect 1437 183 1471 217
rect 1551 47 1585 81
rect 1665 180 1699 214
rect 1665 91 1699 125
rect 1751 181 1785 215
rect 1751 91 1785 125
<< pdiffc >>
rect 39 532 73 566
rect 39 464 73 498
rect 35 390 69 424
rect 145 532 179 566
rect 259 501 293 535
rect 259 433 293 467
rect 383 474 417 508
rect 581 474 615 508
rect 697 480 731 514
rect 802 532 836 566
rect 915 471 949 505
rect 1017 501 1051 535
rect 1017 422 1051 456
rect 1323 539 1357 573
rect 1422 380 1456 414
rect 1541 546 1575 580
rect 1660 546 1694 580
rect 1660 463 1694 497
rect 1660 380 1694 414
rect 1750 546 1784 580
rect 1750 463 1784 497
rect 1750 380 1784 414
<< poly >>
rect 213 615 1205 645
rect 86 578 116 604
rect 213 562 249 615
rect 216 547 246 562
rect 306 547 336 573
rect 451 562 487 615
rect 751 593 787 615
rect 754 578 784 593
rect 1169 583 1205 615
rect 454 547 484 562
rect 538 547 568 573
rect 653 547 683 573
rect 86 363 116 378
rect 83 326 119 363
rect 872 547 902 573
rect 962 547 992 573
rect 1064 547 1094 573
rect 1172 568 1202 583
rect 1256 568 1286 594
rect 1370 592 1400 618
rect 1479 592 1509 618
rect 1617 592 1647 618
rect 1707 592 1737 618
rect 754 363 784 378
rect 216 332 246 347
rect 306 332 336 347
rect 454 332 484 347
rect 538 332 568 347
rect 653 332 683 347
rect 21 310 119 326
rect 213 315 246 332
rect 303 315 339 332
rect 21 276 37 310
rect 71 296 119 310
rect 167 299 243 315
rect 71 276 114 296
rect 21 260 114 276
rect 84 227 114 260
rect 167 265 183 299
rect 217 265 243 299
rect 167 249 243 265
rect 303 299 409 315
rect 303 265 359 299
rect 393 265 409 299
rect 303 249 409 265
rect 213 227 243 249
rect 357 227 387 249
rect 451 242 487 332
rect 457 227 487 242
rect 535 315 571 332
rect 650 315 686 332
rect 535 299 601 315
rect 535 265 551 299
rect 585 265 601 299
rect 535 249 601 265
rect 643 299 709 315
rect 643 265 659 299
rect 693 265 709 299
rect 643 249 709 265
rect 535 227 565 249
rect 671 227 701 249
rect 751 242 787 363
rect 1172 353 1202 368
rect 1256 353 1286 368
rect 1370 353 1400 368
rect 1479 353 1509 368
rect 1617 353 1647 368
rect 1707 353 1737 368
rect 872 332 902 347
rect 962 332 992 347
rect 1064 332 1094 347
rect 869 315 905 332
rect 959 315 995 332
rect 1061 315 1097 332
rect 839 299 905 315
rect 839 265 855 299
rect 889 265 905 299
rect 839 249 905 265
rect 953 299 1019 315
rect 953 265 969 299
rect 1003 265 1019 299
rect 953 249 1019 265
rect 1061 299 1127 315
rect 1061 265 1077 299
rect 1111 265 1127 299
rect 1061 249 1127 265
rect 757 227 787 242
rect 875 227 905 249
rect 989 227 1019 249
rect 1089 227 1119 249
rect 1169 242 1205 353
rect 1175 227 1205 242
rect 1253 336 1289 353
rect 1253 320 1319 336
rect 1253 286 1269 320
rect 1303 286 1319 320
rect 1253 270 1319 286
rect 1367 317 1403 353
rect 1367 301 1433 317
rect 1253 227 1283 270
rect 1367 267 1383 301
rect 1417 281 1433 301
rect 1476 281 1512 353
rect 1614 330 1650 353
rect 1417 267 1512 281
rect 1367 251 1512 267
rect 1581 314 1654 330
rect 1581 280 1597 314
rect 1631 294 1654 314
rect 1704 294 1740 353
rect 1631 280 1740 294
rect 1581 264 1740 280
rect 1396 227 1426 251
rect 1482 227 1512 251
rect 1624 227 1654 264
rect 1710 227 1740 264
rect 84 53 114 79
rect 213 53 243 79
rect 357 53 387 79
rect 457 53 487 79
rect 535 53 565 79
rect 671 53 701 79
rect 757 53 787 79
rect 875 53 905 79
rect 989 53 1019 79
rect 1089 53 1119 79
rect 1175 53 1205 79
rect 1253 53 1283 79
rect 1396 53 1426 79
rect 1482 53 1512 79
rect 1624 53 1654 79
rect 1710 53 1740 79
<< polycont >>
rect 37 276 71 310
rect 183 265 217 299
rect 359 265 393 299
rect 551 265 585 299
rect 659 265 693 299
rect 855 265 889 299
rect 969 265 1003 299
rect 1077 265 1111 299
rect 1269 286 1303 320
rect 1383 267 1417 301
rect 1597 280 1631 314
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 19 566 89 582
rect 19 532 39 566
rect 73 532 89 566
rect 123 566 202 649
rect 123 532 145 566
rect 179 532 202 566
rect 243 535 309 551
rect 19 498 89 532
rect 243 501 259 535
rect 293 501 309 535
rect 243 498 309 501
rect 19 464 39 498
rect 73 467 309 498
rect 73 464 259 467
rect 19 424 85 464
rect 243 433 259 464
rect 293 433 309 467
rect 19 390 35 424
rect 69 390 85 424
rect 121 384 167 430
rect 243 417 309 433
rect 343 508 437 524
rect 343 474 383 508
rect 417 474 437 508
rect 343 458 437 474
rect 565 508 631 649
rect 781 566 858 649
rect 565 474 581 508
rect 615 474 631 508
rect 565 458 631 474
rect 681 514 747 551
rect 781 532 802 566
rect 836 532 858 566
rect 1307 573 1373 649
rect 681 480 697 514
rect 731 498 747 514
rect 899 505 965 551
rect 899 498 915 505
rect 731 480 915 498
rect 681 471 915 480
rect 949 471 965 505
rect 681 464 965 471
rect 21 350 87 356
rect 21 316 31 350
rect 65 316 87 350
rect 21 310 87 316
rect 21 276 37 310
rect 71 276 87 310
rect 21 260 87 276
rect 133 315 167 384
rect 343 383 377 458
rect 899 455 965 464
rect 1001 535 1067 551
rect 1001 501 1017 535
rect 1051 501 1067 535
rect 1307 539 1323 573
rect 1357 539 1373 573
rect 1506 580 1610 649
rect 1506 546 1541 580
rect 1575 546 1610 580
rect 1644 580 1715 596
rect 1644 546 1660 580
rect 1694 546 1715 580
rect 1307 532 1373 539
rect 1001 498 1067 501
rect 1001 464 1610 498
rect 1001 456 1067 464
rect 675 424 839 430
rect 275 349 377 383
rect 411 421 839 424
rect 1001 422 1017 456
rect 1051 422 1067 456
rect 411 390 907 421
rect 1001 417 1067 422
rect 133 299 233 315
rect 133 265 183 299
rect 217 265 233 299
rect 133 249 233 265
rect 23 215 89 226
rect 275 218 309 349
rect 411 315 445 390
rect 675 387 907 390
rect 343 299 445 315
rect 343 265 359 299
rect 393 265 445 299
rect 343 252 445 265
rect 505 350 551 356
rect 505 316 511 350
rect 545 316 551 350
rect 505 315 551 316
rect 675 315 709 387
rect 873 383 907 387
rect 1397 414 1511 430
rect 505 299 601 315
rect 505 265 551 299
rect 585 265 601 299
rect 505 252 601 265
rect 643 299 709 315
rect 643 265 659 299
rect 693 265 709 299
rect 643 252 709 265
rect 793 350 839 353
rect 793 316 799 350
rect 833 316 839 350
rect 873 349 1127 383
rect 1397 380 1422 414
rect 1456 380 1511 414
rect 1397 364 1511 380
rect 793 315 839 316
rect 793 299 905 315
rect 793 265 855 299
rect 889 265 905 299
rect 793 252 905 265
rect 953 299 1019 315
rect 953 265 969 299
rect 1003 265 1019 299
rect 953 218 1019 265
rect 1061 299 1127 349
rect 1061 265 1077 299
rect 1111 265 1127 299
rect 1253 350 1319 356
rect 1253 320 1279 350
rect 1253 286 1269 320
rect 1313 316 1319 350
rect 1303 286 1319 316
rect 1253 270 1319 286
rect 1353 301 1433 317
rect 1061 252 1127 265
rect 1353 267 1383 301
rect 1417 267 1433 301
rect 1353 251 1433 267
rect 1353 218 1387 251
rect 23 210 241 215
rect 23 176 39 210
rect 73 181 241 210
rect 275 202 1387 218
rect 1477 217 1511 364
rect 275 184 412 202
rect 73 176 89 181
rect 23 125 89 176
rect 207 150 241 181
rect 396 168 412 184
rect 446 184 1387 202
rect 446 168 462 184
rect 1421 183 1437 217
rect 1471 183 1511 217
rect 1576 330 1610 464
rect 1644 497 1715 546
rect 1644 463 1660 497
rect 1694 463 1715 497
rect 1644 414 1715 463
rect 1644 380 1660 414
rect 1694 380 1715 414
rect 1644 364 1715 380
rect 1750 580 1800 649
rect 1784 546 1800 580
rect 1750 497 1800 546
rect 1784 463 1800 497
rect 1750 414 1800 463
rect 1784 380 1800 414
rect 1750 364 1800 380
rect 1576 314 1647 330
rect 1576 280 1597 314
rect 1631 280 1647 314
rect 1576 264 1647 280
rect 23 91 39 125
rect 73 91 89 125
rect 23 75 89 91
rect 123 128 173 147
rect 123 94 139 128
rect 123 17 173 94
rect 207 134 362 150
rect 207 100 283 134
rect 317 100 362 134
rect 207 84 362 100
rect 396 125 462 168
rect 396 91 412 125
rect 446 91 462 125
rect 396 75 462 91
rect 560 125 662 141
rect 560 91 594 125
rect 628 91 662 125
rect 560 17 662 91
rect 696 134 994 150
rect 696 129 930 134
rect 696 95 712 129
rect 746 116 930 129
rect 746 95 762 116
rect 696 75 762 95
rect 900 100 930 116
rect 964 100 994 134
rect 900 84 994 100
rect 1028 149 1094 150
rect 1576 149 1610 264
rect 1681 230 1715 364
rect 1028 129 1610 149
rect 1028 95 1044 129
rect 1078 115 1610 129
rect 1649 214 1715 230
rect 1649 180 1665 214
rect 1699 180 1715 214
rect 1649 125 1715 180
rect 1078 95 1094 115
rect 798 48 814 82
rect 848 48 864 82
rect 1028 75 1094 95
rect 1649 91 1665 125
rect 1699 91 1715 125
rect 798 17 864 48
rect 1294 47 1322 81
rect 1356 47 1385 81
rect 1294 17 1385 47
rect 1523 47 1551 81
rect 1585 47 1613 81
rect 1649 75 1715 91
rect 1751 215 1801 231
rect 1785 181 1801 215
rect 1751 125 1801 181
rect 1785 91 1801 125
rect 1523 17 1613 47
rect 1751 17 1801 91
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 31 316 65 350
rect 511 316 545 350
rect 799 316 833 350
rect 1279 320 1313 350
rect 1279 316 1303 320
rect 1303 316 1313 320
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
<< metal1 >>
rect 0 683 1824 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 0 617 1824 649
rect 19 350 77 356
rect 19 316 31 350
rect 65 347 77 350
rect 499 350 557 356
rect 499 347 511 350
rect 65 319 511 347
rect 65 316 77 319
rect 19 310 77 316
rect 499 316 511 319
rect 545 347 557 350
rect 787 350 845 356
rect 787 347 799 350
rect 545 319 799 347
rect 545 316 557 319
rect 499 310 557 316
rect 787 316 799 319
rect 833 347 845 350
rect 1267 350 1325 356
rect 1267 347 1279 350
rect 833 319 1279 347
rect 833 316 845 319
rect 787 310 845 316
rect 1267 316 1279 319
rect 1313 316 1325 350
rect 1267 310 1325 316
rect 0 17 1824 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
rect 0 -49 1824 -17
<< labels >>
rlabel comment s 0 0 0 0 4 fa_2
flabel pwell s 0 0 1824 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 0 617 1824 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel metal1 s 0 617 1824 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 1824 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 703 390 737 424 0 FreeSans 340 0 0 0 CIN
port 3 nsew
flabel corelocali s 799 390 833 424 0 FreeSans 340 0 0 0 CIN
port 3 nsew
flabel corelocali s 127 390 161 424 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 1471 390 1505 424 0 FreeSans 340 0 0 0 COUT
port 8 nsew
flabel corelocali s 1663 390 1697 424 0 FreeSans 340 0 0 0 SUM
port 9 nsew
flabel corelocali s 1663 464 1697 498 0 FreeSans 340 0 0 0 SUM
port 9 nsew
flabel corelocali s 1663 538 1697 572 0 FreeSans 340 0 0 0 SUM
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 1824 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2215502
string GDS_START 2202056
<< end >>
