magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 1574 704
rect 822 301 1173 332
<< pwell >>
rect 0 0 1536 49
<< scnmos >>
rect 89 88 119 198
rect 305 85 335 233
rect 484 149 514 233
rect 562 149 592 233
rect 685 85 715 233
rect 958 82 988 230
rect 1076 82 1106 230
rect 1277 82 1307 230
rect 1422 82 1452 230
<< pmoshvt >>
rect 86 424 116 592
rect 288 392 318 592
rect 389 392 419 476
rect 591 392 621 592
rect 698 508 728 592
rect 924 337 954 561
rect 1048 337 1078 505
rect 1302 368 1332 536
rect 1419 368 1449 592
<< ndiff >>
rect 27 160 89 198
rect 27 126 39 160
rect 73 126 89 160
rect 27 88 89 126
rect 119 160 185 198
rect 255 182 305 233
rect 119 126 139 160
rect 173 126 185 160
rect 119 88 185 126
rect 239 150 305 182
rect 239 116 251 150
rect 285 116 305 150
rect 239 85 305 116
rect 335 208 484 233
rect 335 174 351 208
rect 385 174 484 208
rect 335 149 484 174
rect 514 149 562 233
rect 592 221 685 233
rect 592 187 620 221
rect 654 187 685 221
rect 592 149 685 187
rect 335 85 385 149
rect 635 85 685 149
rect 715 153 775 233
rect 901 218 958 230
rect 901 184 913 218
rect 947 184 958 218
rect 715 119 727 153
rect 761 119 775 153
rect 715 85 775 119
rect 901 128 958 184
rect 901 94 913 128
rect 947 94 958 128
rect 901 82 958 94
rect 988 82 1076 230
rect 1106 218 1163 230
rect 1106 184 1117 218
rect 1151 184 1163 218
rect 1106 82 1163 184
rect 1217 218 1277 230
rect 1217 184 1230 218
rect 1264 184 1277 218
rect 1217 82 1277 184
rect 1307 82 1422 230
rect 1452 214 1509 230
rect 1452 180 1463 214
rect 1497 180 1509 214
rect 1452 128 1509 180
rect 1452 94 1463 128
rect 1497 94 1509 128
rect 1452 82 1509 94
rect 1003 48 1015 82
rect 1049 48 1061 82
rect 1003 36 1061 48
rect 1322 48 1347 82
rect 1381 48 1407 82
rect 1322 36 1407 48
<< pdiff >>
rect 336 625 395 637
rect 336 592 348 625
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 470 86 546
rect 27 436 39 470
rect 73 436 86 470
rect 27 424 86 436
rect 116 580 175 592
rect 116 546 129 580
rect 163 546 175 580
rect 116 470 175 546
rect 116 436 129 470
rect 163 436 175 470
rect 116 424 175 436
rect 229 580 288 592
rect 229 546 241 580
rect 275 546 288 580
rect 229 509 288 546
rect 229 475 241 509
rect 275 475 288 509
rect 229 438 288 475
rect 229 404 241 438
rect 275 404 288 438
rect 229 392 288 404
rect 318 591 348 592
rect 382 591 395 625
rect 972 619 1030 631
rect 746 603 804 615
rect 746 592 758 603
rect 318 562 395 591
rect 532 581 591 592
rect 318 476 371 562
rect 532 547 544 581
rect 578 547 591 581
rect 318 392 389 476
rect 419 451 478 476
rect 419 417 432 451
rect 466 417 478 451
rect 419 392 478 417
rect 532 392 591 547
rect 621 508 698 592
rect 728 569 758 592
rect 792 569 804 603
rect 728 508 804 569
rect 972 585 984 619
rect 1018 585 1030 619
rect 972 561 1030 585
rect 621 445 680 508
rect 621 411 634 445
rect 668 411 680 445
rect 621 392 680 411
rect 858 383 924 561
rect 858 349 873 383
rect 907 349 924 383
rect 858 337 924 349
rect 954 505 1030 561
rect 1350 536 1419 592
rect 1243 524 1302 536
rect 954 337 1048 505
rect 1078 451 1137 505
rect 1078 417 1091 451
rect 1125 417 1137 451
rect 1078 383 1137 417
rect 1078 349 1091 383
rect 1125 349 1137 383
rect 1243 490 1255 524
rect 1289 490 1302 524
rect 1243 440 1302 490
rect 1243 406 1255 440
rect 1289 406 1302 440
rect 1243 368 1302 406
rect 1332 524 1419 536
rect 1332 490 1362 524
rect 1396 490 1419 524
rect 1332 440 1419 490
rect 1332 406 1362 440
rect 1396 406 1419 440
rect 1332 368 1419 406
rect 1449 580 1508 592
rect 1449 546 1462 580
rect 1496 546 1508 580
rect 1449 497 1508 546
rect 1449 463 1462 497
rect 1496 463 1508 497
rect 1449 414 1508 463
rect 1449 380 1462 414
rect 1496 380 1508 414
rect 1449 368 1508 380
rect 1078 337 1137 349
<< ndiffc >>
rect 39 126 73 160
rect 139 126 173 160
rect 251 116 285 150
rect 351 174 385 208
rect 620 187 654 221
rect 913 184 947 218
rect 727 119 761 153
rect 913 94 947 128
rect 1117 184 1151 218
rect 1230 184 1264 218
rect 1463 180 1497 214
rect 1463 94 1497 128
rect 1015 48 1049 82
rect 1347 48 1381 82
<< pdiffc >>
rect 39 546 73 580
rect 39 436 73 470
rect 129 546 163 580
rect 129 436 163 470
rect 241 546 275 580
rect 241 475 275 509
rect 241 404 275 438
rect 348 591 382 625
rect 544 547 578 581
rect 432 417 466 451
rect 758 569 792 603
rect 984 585 1018 619
rect 634 411 668 445
rect 873 349 907 383
rect 1091 417 1125 451
rect 1091 349 1125 383
rect 1255 490 1289 524
rect 1255 406 1289 440
rect 1362 490 1396 524
rect 1362 406 1396 440
rect 1462 546 1496 580
rect 1462 463 1496 497
rect 1462 380 1496 414
<< poly >>
rect 86 592 116 618
rect 288 592 318 618
rect 86 409 116 424
rect 83 370 119 409
rect 591 592 621 618
rect 698 592 728 618
rect 389 476 419 502
rect 924 561 954 587
rect 1419 592 1449 618
rect 698 493 728 508
rect 288 377 318 392
rect 389 377 419 392
rect 591 377 621 392
rect 53 354 119 370
rect 53 320 69 354
rect 103 320 119 354
rect 53 286 119 320
rect 53 252 69 286
rect 103 252 119 286
rect 53 236 119 252
rect 89 198 119 236
rect 167 338 233 354
rect 167 304 183 338
rect 217 304 233 338
rect 167 278 233 304
rect 285 278 321 377
rect 386 356 422 377
rect 386 326 514 356
rect 588 353 624 377
rect 695 356 731 493
rect 167 270 335 278
rect 167 236 183 270
rect 217 248 335 270
rect 217 236 233 248
rect 167 220 233 236
rect 305 233 335 248
rect 484 233 514 326
rect 562 337 637 353
rect 562 303 587 337
rect 621 303 637 337
rect 695 326 771 356
rect 1302 536 1332 562
rect 1048 505 1078 531
rect 1302 353 1332 368
rect 1419 353 1449 368
rect 562 287 637 303
rect 701 305 771 326
rect 924 322 954 337
rect 1048 322 1078 337
rect 1299 336 1335 353
rect 562 233 592 287
rect 701 278 721 305
rect 685 271 721 278
rect 755 271 771 305
rect 921 275 957 322
rect 1045 300 1081 322
rect 1169 320 1235 336
rect 1169 300 1185 320
rect 1045 286 1185 300
rect 1219 286 1235 320
rect 685 248 771 271
rect 685 233 715 248
rect 813 245 988 275
rect 1045 270 1235 286
rect 1277 320 1343 336
rect 1416 330 1452 353
rect 1277 286 1293 320
rect 1327 286 1343 320
rect 1277 270 1343 286
rect 1385 314 1452 330
rect 1385 280 1401 314
rect 1435 280 1452 314
rect 89 62 119 88
rect 484 117 514 149
rect 562 123 592 149
rect 435 101 514 117
rect 305 59 335 85
rect 435 67 451 101
rect 485 67 514 101
rect 813 205 879 245
rect 958 230 988 245
rect 1076 230 1106 270
rect 1277 230 1307 270
rect 1385 264 1452 280
rect 1422 230 1452 264
rect 813 171 829 205
rect 863 171 879 205
rect 813 155 879 171
rect 435 51 514 67
rect 685 59 715 85
rect 958 56 988 82
rect 1076 56 1106 82
rect 1277 56 1307 82
rect 1422 56 1452 82
<< polycont >>
rect 69 320 103 354
rect 69 252 103 286
rect 183 304 217 338
rect 183 236 217 270
rect 587 303 621 337
rect 721 271 755 305
rect 1185 286 1219 320
rect 1293 286 1327 320
rect 1401 280 1435 314
rect 451 67 485 101
rect 829 171 863 205
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 23 580 89 649
rect 332 625 399 649
rect 23 546 39 580
rect 73 546 89 580
rect 23 470 89 546
rect 23 436 39 470
rect 73 436 89 470
rect 23 420 89 436
rect 129 580 189 596
rect 163 546 189 580
rect 129 470 189 546
rect 163 436 189 470
rect 129 420 189 436
rect 25 354 119 370
rect 25 320 69 354
rect 103 320 119 354
rect 25 286 119 320
rect 25 252 69 286
rect 103 252 119 286
rect 25 236 119 252
rect 155 354 189 420
rect 225 580 291 596
rect 332 591 348 625
rect 382 591 399 625
rect 968 619 1034 649
rect 225 546 241 580
rect 275 557 291 580
rect 433 581 594 597
rect 433 557 544 581
rect 275 547 544 557
rect 578 547 594 581
rect 628 569 758 603
rect 792 569 808 603
rect 968 585 984 619
rect 1018 585 1034 619
rect 968 569 1034 585
rect 275 546 467 547
rect 225 523 467 546
rect 225 509 291 523
rect 628 513 662 569
rect 1068 535 1305 540
rect 225 475 241 509
rect 275 475 291 509
rect 501 489 662 513
rect 225 438 291 475
rect 225 404 241 438
rect 275 404 291 438
rect 225 388 291 404
rect 416 479 662 489
rect 718 524 1305 535
rect 718 501 1255 524
rect 416 455 535 479
rect 416 451 466 455
rect 416 417 432 451
rect 569 421 634 445
rect 416 388 466 417
rect 503 411 634 421
rect 668 411 684 445
rect 503 387 603 411
rect 155 338 233 354
rect 155 304 183 338
rect 217 304 233 338
rect 155 270 233 304
rect 155 236 183 270
rect 217 236 233 270
rect 155 220 233 236
rect 267 271 469 305
rect 155 202 189 220
rect 23 160 89 202
rect 23 126 39 160
rect 73 126 89 160
rect 23 17 89 126
rect 123 160 189 202
rect 267 186 301 271
rect 123 126 139 160
rect 173 126 189 160
rect 123 84 189 126
rect 235 150 301 186
rect 235 116 251 150
rect 285 116 301 150
rect 235 81 301 116
rect 335 208 401 237
rect 335 174 351 208
rect 385 174 401 208
rect 335 17 401 174
rect 435 185 469 271
rect 503 253 537 387
rect 718 377 752 501
rect 1169 490 1255 501
rect 1289 490 1305 524
rect 637 353 752 377
rect 571 343 752 353
rect 786 451 1125 467
rect 786 433 1091 451
rect 571 337 671 343
rect 571 303 587 337
rect 621 303 671 337
rect 786 309 820 433
rect 1075 417 1091 433
rect 854 383 963 399
rect 854 349 873 383
rect 907 349 963 383
rect 854 333 963 349
rect 571 287 671 303
rect 705 305 820 309
rect 705 271 721 305
rect 755 271 820 305
rect 705 255 820 271
rect 503 221 671 253
rect 503 219 620 221
rect 603 187 620 219
rect 654 205 879 221
rect 654 187 829 205
rect 435 153 569 185
rect 813 171 829 187
rect 863 171 879 205
rect 813 155 879 171
rect 913 218 963 333
rect 947 184 963 218
rect 1075 383 1125 417
rect 1075 349 1091 383
rect 1075 234 1125 349
rect 1169 440 1305 490
rect 1169 406 1255 440
rect 1289 406 1305 440
rect 1169 390 1305 406
rect 1346 524 1412 649
rect 1346 490 1362 524
rect 1396 490 1412 524
rect 1346 440 1412 490
rect 1346 406 1362 440
rect 1396 406 1412 440
rect 1346 390 1412 406
rect 1446 580 1519 596
rect 1446 546 1462 580
rect 1496 546 1519 580
rect 1446 497 1519 546
rect 1446 463 1462 497
rect 1496 463 1519 497
rect 1446 414 1519 463
rect 1169 320 1235 390
rect 1446 380 1462 414
rect 1496 380 1519 414
rect 1446 364 1519 380
rect 1169 286 1185 320
rect 1219 286 1235 320
rect 1169 270 1235 286
rect 1273 320 1343 356
rect 1273 286 1293 320
rect 1327 286 1343 320
rect 1273 270 1343 286
rect 1379 314 1451 330
rect 1379 280 1401 314
rect 1435 280 1451 314
rect 1201 234 1235 270
rect 1379 264 1451 280
rect 1075 218 1167 234
rect 1075 184 1117 218
rect 1151 184 1167 218
rect 1201 218 1282 234
rect 1201 184 1230 218
rect 1264 184 1282 218
rect 435 151 727 153
rect 535 119 727 151
rect 761 119 779 153
rect 913 150 963 184
rect 1379 150 1413 264
rect 1485 230 1519 364
rect 913 128 1413 150
rect 435 101 501 117
rect 435 67 451 101
rect 485 85 501 101
rect 947 116 1413 128
rect 1447 214 1519 230
rect 1447 180 1463 214
rect 1497 180 1519 214
rect 1447 128 1519 180
rect 947 94 963 116
rect 913 85 963 94
rect 485 67 963 85
rect 1447 94 1463 128
rect 1497 94 1519 128
rect 435 51 963 67
rect 999 48 1015 82
rect 1049 48 1065 82
rect 999 17 1065 48
rect 1318 48 1347 82
rect 1381 48 1411 82
rect 1447 78 1519 94
rect 1318 17 1411 48
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dlxtp_1
flabel pwell s 0 0 1536 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 0 617 1536 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 0 617 1536 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 1536 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 D
port 1 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 D
port 1 nsew
flabel corelocali s 1471 390 1505 424 0 FreeSans 340 0 0 0 Q
port 7 nsew
flabel corelocali s 1471 464 1505 498 0 FreeSans 340 0 0 0 Q
port 7 nsew
flabel corelocali s 1471 538 1505 572 0 FreeSans 340 0 0 0 Q
port 7 nsew
flabel corelocali s 1279 316 1313 350 0 FreeSans 340 0 0 0 GATE
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 1536 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3059886
string GDS_START 3048266
<< end >>
