magic
tech sky130A
magscale 1 2
timestamp 1604502741
<< locali >>
rect 151 424 217 547
rect 25 390 217 424
rect 25 236 71 390
rect 121 270 263 356
rect 301 270 551 356
rect 601 236 743 310
rect 793 270 935 356
rect 970 270 1036 356
rect 25 202 500 236
rect 232 70 298 202
rect 434 195 500 202
rect 800 195 866 226
rect 434 154 866 195
rect 434 70 500 154
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 61 581 487 615
rect 61 458 111 581
rect 257 390 291 581
rect 331 424 397 547
rect 437 458 487 581
rect 525 581 771 615
rect 525 458 581 581
rect 615 424 665 547
rect 331 390 665 424
rect 705 424 771 581
rect 811 458 845 649
rect 885 424 935 596
rect 975 458 1041 649
rect 1081 424 1131 596
rect 705 390 1131 424
rect 615 364 665 390
rect 1081 364 1131 390
rect 132 17 198 168
rect 332 17 400 168
rect 902 202 1126 236
rect 902 120 936 202
rect 714 70 936 120
rect 972 17 1040 168
rect 1076 70 1126 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
rlabel locali s 793 270 935 356 6 A1
port 1 nsew signal input
rlabel locali s 970 270 1036 356 6 A2
port 2 nsew signal input
rlabel locali s 601 236 743 310 6 B1
port 3 nsew signal input
rlabel locali s 301 270 551 356 6 C1
port 4 nsew signal input
rlabel locali s 121 270 263 356 6 D1
port 5 nsew signal input
rlabel locali s 800 195 866 226 6 Y
port 6 nsew signal output
rlabel locali s 434 195 500 202 6 Y
port 6 nsew signal output
rlabel locali s 434 154 866 195 6 Y
port 6 nsew signal output
rlabel locali s 434 70 500 154 6 Y
port 6 nsew signal output
rlabel locali s 232 70 298 202 6 Y
port 6 nsew signal output
rlabel locali s 151 424 217 547 6 Y
port 6 nsew signal output
rlabel locali s 25 390 217 424 6 Y
port 6 nsew signal output
rlabel locali s 25 236 71 390 6 Y
port 6 nsew signal output
rlabel locali s 25 202 500 236 6 Y
port 6 nsew signal output
rlabel metal1 s 0 -49 1152 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 617 1152 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3862148
string GDS_START 3852556
<< end >>
