magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 1286 704
<< pwell >>
rect 0 0 1248 49
<< scnmos >>
rect 118 123 148 251
rect 236 100 266 248
rect 322 100 352 248
rect 408 100 438 248
rect 494 100 524 248
rect 592 123 622 251
rect 678 123 708 251
rect 834 123 864 251
rect 932 123 962 251
rect 1018 123 1048 251
rect 1104 123 1134 251
<< pmoshvt >>
rect 84 392 114 592
rect 187 368 217 592
rect 277 368 307 592
rect 367 368 397 592
rect 457 368 487 592
rect 651 392 681 592
rect 741 392 771 592
rect 831 392 861 592
rect 921 392 951 592
rect 1011 392 1041 592
rect 1101 392 1131 592
<< ndiff >>
rect 65 228 118 251
rect 65 194 73 228
rect 107 194 118 228
rect 65 123 118 194
rect 148 248 221 251
rect 542 248 592 251
rect 148 239 236 248
rect 148 205 175 239
rect 209 205 236 239
rect 148 146 236 205
rect 148 123 175 146
rect 163 112 175 123
rect 209 112 236 146
rect 163 100 236 112
rect 266 220 322 248
rect 266 186 277 220
rect 311 186 322 220
rect 266 146 322 186
rect 266 112 277 146
rect 311 112 322 146
rect 266 100 322 112
rect 352 149 408 248
rect 352 115 363 149
rect 397 115 408 149
rect 352 100 408 115
rect 438 220 494 248
rect 438 186 449 220
rect 483 186 494 220
rect 438 146 494 186
rect 438 112 449 146
rect 483 112 494 146
rect 438 100 494 112
rect 524 172 592 248
rect 524 138 535 172
rect 569 138 592 172
rect 524 123 592 138
rect 622 239 678 251
rect 622 205 633 239
rect 667 205 678 239
rect 622 169 678 205
rect 622 135 633 169
rect 667 135 678 169
rect 622 123 678 135
rect 708 172 834 251
rect 708 138 719 172
rect 753 138 834 172
rect 708 123 834 138
rect 864 170 932 251
rect 864 136 887 170
rect 921 136 932 170
rect 864 123 932 136
rect 962 239 1018 251
rect 962 205 973 239
rect 1007 205 1018 239
rect 962 169 1018 205
rect 962 135 973 169
rect 1007 135 1018 169
rect 962 123 1018 135
rect 1048 239 1104 251
rect 1048 205 1059 239
rect 1093 205 1104 239
rect 1048 169 1104 205
rect 1048 135 1059 169
rect 1093 135 1104 169
rect 1048 123 1104 135
rect 1134 239 1187 251
rect 1134 205 1145 239
rect 1179 205 1187 239
rect 1134 169 1187 205
rect 1134 135 1145 169
rect 1179 135 1187 169
rect 1134 123 1187 135
rect 524 100 577 123
<< pdiff >>
rect 29 580 84 592
rect 29 546 37 580
rect 71 546 84 580
rect 29 509 84 546
rect 29 475 37 509
rect 71 475 84 509
rect 29 438 84 475
rect 29 404 37 438
rect 71 404 84 438
rect 29 392 84 404
rect 114 572 187 592
rect 114 538 140 572
rect 174 538 187 572
rect 114 392 187 538
rect 132 368 187 392
rect 217 417 277 592
rect 217 383 230 417
rect 264 383 277 417
rect 217 368 277 383
rect 307 572 367 592
rect 307 538 320 572
rect 354 538 367 572
rect 307 368 367 538
rect 397 420 457 592
rect 397 386 410 420
rect 444 386 457 420
rect 397 368 457 386
rect 487 572 542 592
rect 487 538 500 572
rect 534 538 542 572
rect 487 368 542 538
rect 596 580 651 592
rect 596 546 604 580
rect 638 546 651 580
rect 596 488 651 546
rect 596 454 604 488
rect 638 454 651 488
rect 596 392 651 454
rect 681 531 741 592
rect 681 497 694 531
rect 728 497 741 531
rect 681 440 741 497
rect 681 406 694 440
rect 728 406 741 440
rect 681 392 741 406
rect 771 580 831 592
rect 771 546 784 580
rect 818 546 831 580
rect 771 509 831 546
rect 771 475 784 509
rect 818 475 831 509
rect 771 438 831 475
rect 771 404 784 438
rect 818 404 831 438
rect 771 392 831 404
rect 861 580 921 592
rect 861 546 874 580
rect 908 546 921 580
rect 861 508 921 546
rect 861 474 874 508
rect 908 474 921 508
rect 861 392 921 474
rect 951 580 1011 592
rect 951 546 964 580
rect 998 546 1011 580
rect 951 510 1011 546
rect 951 476 964 510
rect 998 476 1011 510
rect 951 440 1011 476
rect 951 406 964 440
rect 998 406 1011 440
rect 951 392 1011 406
rect 1041 580 1101 592
rect 1041 546 1054 580
rect 1088 546 1101 580
rect 1041 508 1101 546
rect 1041 474 1054 508
rect 1088 474 1101 508
rect 1041 392 1101 474
rect 1131 580 1186 592
rect 1131 546 1144 580
rect 1178 546 1186 580
rect 1131 509 1186 546
rect 1131 475 1144 509
rect 1178 475 1186 509
rect 1131 438 1186 475
rect 1131 404 1144 438
rect 1178 404 1186 438
rect 1131 392 1186 404
<< ndiffc >>
rect 73 194 107 228
rect 175 205 209 239
rect 175 112 209 146
rect 277 186 311 220
rect 277 112 311 146
rect 363 115 397 149
rect 449 186 483 220
rect 449 112 483 146
rect 535 138 569 172
rect 633 205 667 239
rect 633 135 667 169
rect 719 138 753 172
rect 887 136 921 170
rect 973 205 1007 239
rect 973 135 1007 169
rect 1059 205 1093 239
rect 1059 135 1093 169
rect 1145 205 1179 239
rect 1145 135 1179 169
<< pdiffc >>
rect 37 546 71 580
rect 37 475 71 509
rect 37 404 71 438
rect 140 538 174 572
rect 230 383 264 417
rect 320 538 354 572
rect 410 386 444 420
rect 500 538 534 572
rect 604 546 638 580
rect 604 454 638 488
rect 694 497 728 531
rect 694 406 728 440
rect 784 546 818 580
rect 784 475 818 509
rect 784 404 818 438
rect 874 546 908 580
rect 874 474 908 508
rect 964 546 998 580
rect 964 476 998 510
rect 964 406 998 440
rect 1054 546 1088 580
rect 1054 474 1088 508
rect 1144 546 1178 580
rect 1144 475 1178 509
rect 1144 404 1178 438
<< poly >>
rect 84 592 114 618
rect 187 592 217 618
rect 277 592 307 618
rect 367 592 397 618
rect 457 592 487 618
rect 651 592 681 618
rect 741 592 771 618
rect 831 592 861 618
rect 921 592 951 618
rect 1011 592 1041 618
rect 1101 592 1131 618
rect 84 377 114 392
rect 81 296 117 377
rect 651 377 681 392
rect 741 377 771 392
rect 831 377 861 392
rect 921 377 951 392
rect 1011 377 1041 392
rect 1101 377 1131 392
rect 187 353 217 368
rect 277 353 307 368
rect 367 353 397 368
rect 457 353 487 368
rect 648 356 684 377
rect 187 338 220 353
rect 190 336 220 338
rect 274 336 310 353
rect 364 336 400 353
rect 454 336 490 353
rect 592 340 684 356
rect 190 320 524 336
rect 81 266 148 296
rect 190 286 334 320
rect 368 286 402 320
rect 436 286 470 320
rect 504 286 524 320
rect 190 270 524 286
rect 118 251 148 266
rect 236 248 266 270
rect 322 248 352 270
rect 408 248 438 270
rect 494 248 524 270
rect 592 306 608 340
rect 642 320 684 340
rect 738 320 774 377
rect 642 306 774 320
rect 592 290 774 306
rect 592 251 622 290
rect 678 251 708 290
rect 828 266 864 377
rect 918 356 954 377
rect 1008 356 1044 377
rect 918 340 1044 356
rect 918 306 934 340
rect 968 320 1044 340
rect 968 306 1048 320
rect 918 290 1048 306
rect 834 251 864 266
rect 932 251 962 290
rect 1018 251 1048 290
rect 1098 266 1134 377
rect 1104 251 1134 266
rect 118 101 148 123
rect 59 85 148 101
rect 59 51 75 85
rect 109 51 148 85
rect 236 74 266 100
rect 322 74 352 100
rect 408 74 438 100
rect 494 74 524 100
rect 592 97 622 123
rect 678 97 708 123
rect 834 101 864 123
rect 787 85 864 101
rect 932 97 962 123
rect 1018 97 1048 123
rect 59 35 148 51
rect 787 51 803 85
rect 837 55 864 85
rect 1104 55 1134 123
rect 837 51 1134 55
rect 787 25 1134 51
<< polycont >>
rect 334 286 368 320
rect 402 286 436 320
rect 470 286 504 320
rect 608 306 642 340
rect 934 306 968 340
rect 75 51 109 85
rect 803 51 837 85
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 21 580 87 596
rect 21 546 37 580
rect 71 546 87 580
rect 21 509 87 546
rect 124 572 190 649
rect 124 538 140 572
rect 174 538 190 572
rect 124 522 190 538
rect 304 572 370 649
rect 304 538 320 572
rect 354 538 370 572
rect 304 522 370 538
rect 484 572 550 649
rect 484 538 500 572
rect 534 538 550 572
rect 484 522 550 538
rect 588 581 818 615
rect 588 580 654 581
rect 588 546 604 580
rect 638 546 654 580
rect 784 580 818 581
rect 21 475 37 509
rect 71 488 87 509
rect 588 488 654 546
rect 71 475 528 488
rect 21 454 528 475
rect 21 438 87 454
rect 21 404 37 438
rect 71 404 87 438
rect 21 255 87 404
rect 121 417 410 420
rect 121 383 230 417
rect 264 386 410 417
rect 444 386 460 420
rect 264 383 460 386
rect 121 370 460 383
rect 494 404 528 454
rect 588 454 604 488
rect 638 454 654 488
rect 588 438 654 454
rect 694 531 744 547
rect 728 497 744 531
rect 694 440 744 497
rect 728 406 744 440
rect 494 370 658 404
rect 121 302 284 370
rect 592 340 658 370
rect 21 228 123 255
rect 21 194 73 228
rect 107 194 123 228
rect 21 168 123 194
rect 159 239 209 255
rect 159 205 175 239
rect 159 146 209 205
rect 25 101 71 134
rect 159 112 175 146
rect 25 85 125 101
rect 25 51 75 85
rect 109 51 125 85
rect 159 17 209 112
rect 250 236 284 302
rect 318 320 551 336
rect 318 286 334 320
rect 368 286 402 320
rect 436 286 470 320
rect 504 286 551 320
rect 592 306 608 340
rect 642 306 658 340
rect 592 290 658 306
rect 318 270 551 286
rect 517 256 551 270
rect 694 256 744 406
rect 784 509 818 546
rect 784 438 818 475
rect 858 580 908 649
rect 858 546 874 580
rect 858 508 908 546
rect 858 474 874 508
rect 858 458 908 474
rect 948 580 1014 596
rect 948 546 964 580
rect 998 546 1014 580
rect 948 510 1014 546
rect 948 476 964 510
rect 998 476 1014 510
rect 948 440 1014 476
rect 1054 580 1104 649
rect 1088 546 1104 580
rect 1054 508 1104 546
rect 1088 474 1104 508
rect 1054 458 1104 474
rect 1144 580 1194 596
rect 1178 546 1194 580
rect 1144 509 1194 546
rect 1178 475 1194 509
rect 948 424 964 440
rect 818 406 964 424
rect 998 424 1014 440
rect 1144 438 1194 475
rect 998 406 1144 424
rect 818 404 1144 406
rect 1178 404 1194 438
rect 784 390 1194 404
rect 784 388 818 390
rect 1144 388 1194 390
rect 889 340 1040 356
rect 889 306 934 340
rect 968 306 1040 340
rect 889 290 1040 306
rect 517 239 1007 256
rect 250 220 483 236
rect 517 222 633 239
rect 250 186 277 220
rect 311 202 449 220
rect 250 146 311 186
rect 433 186 449 202
rect 617 205 633 222
rect 667 222 973 239
rect 667 205 683 222
rect 250 112 277 146
rect 250 96 311 112
rect 347 149 397 168
rect 347 115 363 149
rect 347 17 397 115
rect 433 146 483 186
rect 433 112 449 146
rect 433 96 483 112
rect 519 172 569 188
rect 519 138 535 172
rect 519 17 569 138
rect 617 169 683 205
rect 957 205 973 222
rect 617 135 633 169
rect 667 135 683 169
rect 617 119 683 135
rect 719 172 753 188
rect 719 17 753 138
rect 887 170 921 188
rect 787 85 853 134
rect 787 51 803 85
rect 837 51 853 85
rect 887 85 921 136
rect 957 169 1007 205
rect 957 135 973 169
rect 957 119 1007 135
rect 1043 239 1109 255
rect 1043 205 1059 239
rect 1093 205 1109 239
rect 1043 169 1109 205
rect 1043 135 1059 169
rect 1093 135 1109 169
rect 1043 85 1109 135
rect 887 51 1109 85
rect 1145 239 1195 255
rect 1179 205 1195 239
rect 1145 169 1195 205
rect 1179 135 1195 169
rect 1145 17 1195 135
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
<< metal1 >>
rect 0 683 1248 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 0 617 1248 649
rect 0 17 1248 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
rect 0 -49 1248 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a21bo_4
flabel pwell s 0 0 1248 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 0 617 1248 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 1248 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 1248 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 31 94 65 128 0 FreeSans 340 0 0 0 B1_N
port 3 nsew
flabel corelocali s 799 94 833 128 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 X
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 1248 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 4042894
string GDS_START 4032920
<< end >>
