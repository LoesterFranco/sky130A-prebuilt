magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 1786 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 89 47 119 177
rect 183 47 213 177
rect 277 47 307 177
rect 371 47 401 177
rect 455 47 485 177
rect 549 47 579 177
rect 643 47 673 177
rect 747 47 777 177
rect 955 47 985 177
rect 1049 47 1079 177
rect 1143 47 1173 177
rect 1237 47 1267 177
rect 1331 47 1361 177
rect 1425 47 1455 177
rect 1519 47 1549 177
rect 1613 47 1643 177
<< pmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 457 297 493 497
rect 551 297 587 497
rect 645 297 681 497
rect 739 297 775 497
rect 837 297 873 497
rect 931 297 967 497
rect 1025 297 1061 497
rect 1119 297 1155 497
rect 1323 297 1359 497
rect 1417 297 1453 497
rect 1511 297 1547 497
rect 1605 297 1641 497
<< ndiff >>
rect 27 101 89 177
rect 27 67 35 101
rect 69 67 89 101
rect 27 47 89 67
rect 119 93 183 177
rect 119 59 129 93
rect 163 59 183 93
rect 119 47 183 59
rect 213 101 277 177
rect 213 67 223 101
rect 257 67 277 101
rect 213 47 277 67
rect 307 93 371 177
rect 307 59 317 93
rect 351 59 371 93
rect 307 47 371 59
rect 401 101 455 177
rect 401 67 411 101
rect 445 67 455 101
rect 401 47 455 67
rect 485 93 549 177
rect 485 59 505 93
rect 539 59 549 93
rect 485 47 549 59
rect 579 161 643 177
rect 579 127 599 161
rect 633 127 643 161
rect 579 47 643 127
rect 673 93 747 177
rect 673 59 693 93
rect 727 59 747 93
rect 673 47 747 59
rect 777 161 829 177
rect 777 127 787 161
rect 821 127 829 161
rect 777 47 829 127
rect 893 161 955 177
rect 893 127 901 161
rect 935 127 955 161
rect 893 47 955 127
rect 985 93 1049 177
rect 985 59 995 93
rect 1029 59 1049 93
rect 985 47 1049 59
rect 1079 161 1143 177
rect 1079 127 1089 161
rect 1123 127 1143 161
rect 1079 47 1143 127
rect 1173 93 1237 177
rect 1173 59 1183 93
rect 1217 59 1237 93
rect 1173 47 1237 59
rect 1267 161 1331 177
rect 1267 127 1277 161
rect 1311 127 1331 161
rect 1267 47 1331 127
rect 1361 93 1425 177
rect 1361 59 1371 93
rect 1405 59 1425 93
rect 1361 47 1425 59
rect 1455 101 1519 177
rect 1455 67 1465 101
rect 1499 67 1519 101
rect 1455 47 1519 67
rect 1549 93 1613 177
rect 1549 59 1559 93
rect 1593 59 1613 93
rect 1549 47 1613 59
rect 1643 101 1707 177
rect 1643 67 1653 101
rect 1687 67 1707 101
rect 1643 47 1707 67
<< pdiff >>
rect 27 477 81 497
rect 27 443 35 477
rect 69 443 81 477
rect 27 409 81 443
rect 27 375 35 409
rect 69 375 81 409
rect 27 297 81 375
rect 117 485 175 497
rect 117 451 129 485
rect 163 451 175 485
rect 117 417 175 451
rect 117 383 129 417
rect 163 383 175 417
rect 117 297 175 383
rect 211 477 269 497
rect 211 443 223 477
rect 257 443 269 477
rect 211 409 269 443
rect 211 375 223 409
rect 257 375 269 409
rect 211 297 269 375
rect 305 485 363 497
rect 305 451 317 485
rect 351 451 363 485
rect 305 417 363 451
rect 305 383 317 417
rect 351 383 363 417
rect 305 297 363 383
rect 399 477 457 497
rect 399 443 411 477
rect 445 443 457 477
rect 399 409 457 443
rect 399 375 411 409
rect 445 375 457 409
rect 399 297 457 375
rect 493 485 551 497
rect 493 451 505 485
rect 539 451 551 485
rect 493 417 551 451
rect 493 383 505 417
rect 539 383 551 417
rect 493 297 551 383
rect 587 477 645 497
rect 587 443 599 477
rect 633 443 645 477
rect 587 409 645 443
rect 587 375 599 409
rect 633 375 645 409
rect 587 297 645 375
rect 681 485 739 497
rect 681 451 693 485
rect 727 451 739 485
rect 681 417 739 451
rect 681 383 693 417
rect 727 383 739 417
rect 681 297 739 383
rect 775 477 837 497
rect 775 443 787 477
rect 821 443 837 477
rect 775 409 837 443
rect 775 375 787 409
rect 821 375 837 409
rect 775 297 837 375
rect 873 485 931 497
rect 873 451 885 485
rect 919 451 931 485
rect 873 417 931 451
rect 873 383 885 417
rect 919 383 931 417
rect 873 297 931 383
rect 967 477 1025 497
rect 967 443 979 477
rect 1013 443 1025 477
rect 967 409 1025 443
rect 967 375 979 409
rect 1013 375 1025 409
rect 967 297 1025 375
rect 1061 485 1119 497
rect 1061 451 1073 485
rect 1107 451 1119 485
rect 1061 297 1119 451
rect 1155 477 1323 497
rect 1155 443 1167 477
rect 1201 443 1323 477
rect 1155 377 1323 443
rect 1155 343 1167 377
rect 1201 343 1323 377
rect 1155 297 1323 343
rect 1359 417 1417 497
rect 1359 383 1371 417
rect 1405 383 1417 417
rect 1359 297 1417 383
rect 1453 485 1511 497
rect 1453 451 1465 485
rect 1499 451 1511 485
rect 1453 297 1511 451
rect 1547 417 1605 497
rect 1547 383 1559 417
rect 1593 383 1605 417
rect 1547 297 1605 383
rect 1641 485 1707 497
rect 1641 451 1653 485
rect 1687 451 1707 485
rect 1641 417 1707 451
rect 1641 383 1653 417
rect 1687 383 1707 417
rect 1641 349 1707 383
rect 1641 315 1653 349
rect 1687 315 1707 349
rect 1641 297 1707 315
<< ndiffc >>
rect 35 67 69 101
rect 129 59 163 93
rect 223 67 257 101
rect 317 59 351 93
rect 411 67 445 101
rect 505 59 539 93
rect 599 127 633 161
rect 693 59 727 93
rect 787 127 821 161
rect 901 127 935 161
rect 995 59 1029 93
rect 1089 127 1123 161
rect 1183 59 1217 93
rect 1277 127 1311 161
rect 1371 59 1405 93
rect 1465 67 1499 101
rect 1559 59 1593 93
rect 1653 67 1687 101
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 129 451 163 485
rect 129 383 163 417
rect 223 443 257 477
rect 223 375 257 409
rect 317 451 351 485
rect 317 383 351 417
rect 411 443 445 477
rect 411 375 445 409
rect 505 451 539 485
rect 505 383 539 417
rect 599 443 633 477
rect 599 375 633 409
rect 693 451 727 485
rect 693 383 727 417
rect 787 443 821 477
rect 787 375 821 409
rect 885 451 919 485
rect 885 383 919 417
rect 979 443 1013 477
rect 979 375 1013 409
rect 1073 451 1107 485
rect 1167 443 1201 477
rect 1167 343 1201 377
rect 1371 383 1405 417
rect 1465 451 1499 485
rect 1559 383 1593 417
rect 1653 451 1687 485
rect 1653 383 1687 417
rect 1653 315 1687 349
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 457 497 493 523
rect 551 497 587 523
rect 645 497 681 523
rect 739 497 775 523
rect 837 497 873 523
rect 931 497 967 523
rect 1025 497 1061 523
rect 1119 497 1155 523
rect 1323 497 1359 523
rect 1417 497 1453 523
rect 1511 497 1547 523
rect 1605 497 1641 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 457 282 493 297
rect 551 282 587 297
rect 645 282 681 297
rect 739 282 775 297
rect 837 282 873 297
rect 931 282 967 297
rect 1025 282 1061 297
rect 1119 282 1155 297
rect 1323 282 1359 297
rect 1417 282 1453 297
rect 1511 282 1547 297
rect 1605 282 1641 297
rect 79 265 119 282
rect 173 265 213 282
rect 267 265 307 282
rect 361 265 401 282
rect 22 249 401 265
rect 22 215 40 249
rect 74 215 124 249
rect 158 215 198 249
rect 232 215 282 249
rect 316 215 401 249
rect 22 199 401 215
rect 89 177 119 199
rect 183 177 213 199
rect 277 177 307 199
rect 371 177 401 199
rect 455 265 495 282
rect 549 265 589 282
rect 643 265 683 282
rect 737 265 777 282
rect 455 249 777 265
rect 455 215 465 249
rect 499 215 549 249
rect 583 215 633 249
rect 667 215 717 249
rect 751 215 777 249
rect 455 199 777 215
rect 835 269 875 282
rect 929 269 969 282
rect 1023 269 1063 282
rect 1117 269 1157 282
rect 835 265 1157 269
rect 1321 265 1361 282
rect 1415 265 1455 282
rect 1509 265 1549 282
rect 1603 265 1643 282
rect 835 249 1267 265
rect 835 215 845 249
rect 879 215 929 249
rect 963 215 1013 249
rect 1047 215 1097 249
rect 1131 215 1267 249
rect 835 202 1267 215
rect 835 199 1173 202
rect 455 177 485 199
rect 549 177 579 199
rect 643 177 673 199
rect 747 177 777 199
rect 955 177 985 199
rect 1049 177 1079 199
rect 1143 177 1173 199
rect 1237 177 1267 202
rect 1309 249 1643 265
rect 1309 215 1319 249
rect 1353 215 1403 249
rect 1437 215 1487 249
rect 1521 215 1643 249
rect 1309 199 1643 215
rect 1331 177 1361 199
rect 1425 177 1455 199
rect 1519 177 1549 199
rect 1613 177 1643 199
rect 89 21 119 47
rect 183 21 213 47
rect 277 21 307 47
rect 371 21 401 47
rect 455 21 485 47
rect 549 21 579 47
rect 643 21 673 47
rect 747 21 777 47
rect 955 21 985 47
rect 1049 21 1079 47
rect 1143 21 1173 47
rect 1237 21 1267 47
rect 1331 21 1361 47
rect 1425 21 1455 47
rect 1519 21 1549 47
rect 1613 21 1643 47
<< polycont >>
rect 40 215 74 249
rect 124 215 158 249
rect 198 215 232 249
rect 282 215 316 249
rect 465 215 499 249
rect 549 215 583 249
rect 633 215 667 249
rect 717 215 751 249
rect 845 215 879 249
rect 929 215 963 249
rect 1013 215 1047 249
rect 1097 215 1131 249
rect 1319 215 1353 249
rect 1403 215 1437 249
rect 1487 215 1521 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 35 477 69 493
rect 35 409 69 443
rect 103 485 179 527
rect 103 451 129 485
rect 163 451 179 485
rect 103 417 179 451
rect 103 383 129 417
rect 163 383 179 417
rect 223 477 257 493
rect 223 409 257 443
rect 35 333 69 375
rect 291 485 367 527
rect 291 451 317 485
rect 351 451 367 485
rect 291 417 367 451
rect 291 383 317 417
rect 351 383 367 417
rect 411 477 445 493
rect 411 409 445 443
rect 223 333 257 375
rect 479 485 555 527
rect 479 451 505 485
rect 539 451 555 485
rect 479 417 555 451
rect 479 383 505 417
rect 539 383 555 417
rect 599 477 633 493
rect 599 409 633 443
rect 411 333 445 375
rect 667 485 743 527
rect 667 451 693 485
rect 727 451 743 485
rect 667 417 743 451
rect 667 383 693 417
rect 727 383 743 417
rect 787 477 821 493
rect 787 409 821 443
rect 599 333 633 375
rect 859 485 935 527
rect 859 451 885 485
rect 919 451 935 485
rect 859 417 935 451
rect 859 383 885 417
rect 919 383 935 417
rect 979 477 1013 493
rect 1047 485 1123 527
rect 1047 451 1073 485
rect 1107 451 1123 485
rect 1167 485 1201 493
rect 1167 477 1465 485
rect 979 409 1013 443
rect 787 333 821 375
rect 979 333 1013 375
rect 1201 451 1465 477
rect 1499 451 1653 485
rect 1687 451 1703 485
rect 1167 377 1201 443
rect 1653 417 1703 451
rect 1345 383 1371 417
rect 1405 383 1559 417
rect 1593 383 1617 417
rect 1167 333 1201 343
rect 35 299 1201 333
rect 24 249 377 265
rect 24 215 40 249
rect 74 215 124 249
rect 158 215 198 249
rect 232 215 282 249
rect 316 215 377 249
rect 24 199 377 215
rect 427 249 790 265
rect 427 215 465 249
rect 499 215 549 249
rect 583 215 633 249
rect 667 215 717 249
rect 751 215 790 249
rect 427 199 790 215
rect 845 249 1204 265
rect 879 215 929 249
rect 963 215 1013 249
rect 1047 215 1097 249
rect 1131 215 1204 249
rect 845 199 1204 215
rect 1254 249 1521 326
rect 1254 215 1319 249
rect 1353 215 1403 249
rect 1437 215 1487 249
rect 1254 199 1521 215
rect 1569 161 1617 383
rect 1687 383 1703 417
rect 1653 349 1703 383
rect 1687 315 1703 349
rect 1653 299 1703 315
rect 35 127 599 161
rect 633 127 787 161
rect 821 127 837 161
rect 885 127 901 161
rect 935 127 1089 161
rect 1123 127 1277 161
rect 1311 127 1687 161
rect 35 101 69 127
rect 223 101 257 127
rect 35 51 69 67
rect 103 59 129 93
rect 163 59 179 93
rect 103 17 179 59
rect 411 101 445 127
rect 223 51 257 67
rect 291 59 317 93
rect 351 59 367 93
rect 291 17 367 59
rect 1465 101 1499 127
rect 411 51 445 67
rect 479 59 505 93
rect 539 59 693 93
rect 727 59 995 93
rect 1029 59 1183 93
rect 1217 59 1233 93
rect 1345 59 1371 93
rect 1405 59 1421 93
rect 1345 17 1421 59
rect 1653 101 1687 127
rect 1465 51 1499 67
rect 1533 59 1559 93
rect 1593 59 1609 93
rect 1533 17 1609 59
rect 1653 51 1687 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
<< metal1 >>
rect 0 561 1748 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 0 496 1748 527
rect 0 17 1748 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
rect 0 -48 1748 -17
<< labels >>
flabel corelocali s 1579 153 1613 187 0 FreeSans 200 0 0 0 Y
port 9 nsew
flabel corelocali s 1579 221 1613 255 0 FreeSans 200 0 0 0 Y
port 9 nsew
flabel corelocali s 1579 289 1613 323 0 FreeSans 200 0 0 0 Y
port 9 nsew
flabel corelocali s 1579 357 1613 391 0 FreeSans 200 0 0 0 Y
port 9 nsew
flabel corelocali s 1487 289 1521 323 0 FreeSans 200 0 0 0 B1
port 4 nsew
flabel corelocali s 756 221 790 255 0 FreeSans 200 0 0 0 A2
port 2 nsew
flabel corelocali s 302 221 336 255 0 FreeSans 200 0 0 0 A3
port 3 nsew
flabel corelocali s 1134 221 1168 255 0 FreeSans 200 0 0 0 A1
port 1 nsew
flabel corelocali s 1318 289 1352 323 0 FreeSans 200 0 0 0 B1
port 4 nsew
flabel corelocali s 1411 289 1445 323 0 FreeSans 200 0 0 0 B1
port 4 nsew
flabel corelocali s 1318 221 1352 255 0 FreeSans 200 0 0 0 B1
port 4 nsew
flabel corelocali s 1411 221 1445 255 0 FreeSans 200 0 0 0 B1
port 4 nsew
flabel corelocali s 578 221 612 255 0 FreeSans 200 0 0 0 A2
port 2 nsew
flabel corelocali s 1487 221 1521 255 0 FreeSans 200 0 0 0 B1
port 4 nsew
flabel corelocali s 466 238 466 238 0 FreeSans 200 0 0 0 A2
port 2 nsew
flabel corelocali s 1043 221 1077 255 0 FreeSans 200 0 0 0 A1
port 1 nsew
flabel corelocali s 213 221 247 255 0 FreeSans 200 0 0 0 A3
port 3 nsew
flabel corelocali s 122 221 156 255 0 FreeSans 200 0 0 0 A3
port 3 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 200 0 0 0 A3
port 3 nsew
flabel corelocali s 672 221 706 255 0 FreeSans 200 0 0 0 A2
port 2 nsew
flabel corelocali s 952 221 986 255 0 FreeSans 200 0 0 0 A1
port 1 nsew
flabel corelocali s 860 221 894 255 0 FreeSans 200 0 0 0 A1
port 1 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 1748 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1415778
string GDS_START 1402186
<< end >>
