magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 375 364 463 596
rect 22 236 88 310
rect 207 236 273 310
rect 429 230 463 364
rect 307 196 463 230
rect 307 70 357 196
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 63 378 129 540
rect 185 412 251 649
rect 63 344 341 378
rect 122 202 156 344
rect 307 330 341 344
rect 307 264 395 330
rect 51 136 156 202
rect 190 17 256 202
rect 391 17 446 162
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< metal1 >>
rect 0 683 480 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 0 617 480 649
rect 0 17 480 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
rect 0 -49 480 -17
<< labels >>
rlabel locali s 207 236 273 310 6 A
port 1 nsew signal input
rlabel locali s 22 236 88 310 6 B_N
port 2 nsew signal input
rlabel locali s 429 230 463 364 6 Y
port 3 nsew signal output
rlabel locali s 375 364 463 596 6 Y
port 3 nsew signal output
rlabel locali s 307 196 463 230 6 Y
port 3 nsew signal output
rlabel locali s 307 70 357 196 6 Y
port 3 nsew signal output
rlabel metal1 s 0 -49 480 49 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 617 480 715 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 480 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1526404
string GDS_START 1521582
<< end >>
