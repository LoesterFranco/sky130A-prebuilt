magic
tech sky130A
magscale 1 2
timestamp 1599588244
<< locali >>
rect 21 252 223 354
rect 294 290 455 356
rect 769 270 839 356
rect 883 270 949 356
rect 1051 378 1117 596
rect 1251 378 1317 596
rect 1051 344 1317 378
rect 1251 210 1317 344
rect 1051 162 1317 210
rect 1051 70 1117 162
rect 1251 70 1317 162
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 37 424 103 596
rect 143 458 177 649
rect 217 581 463 615
rect 217 424 283 581
rect 37 390 283 424
rect 323 424 357 547
rect 397 458 463 581
rect 509 464 575 649
rect 720 558 786 649
rect 934 558 1000 649
rect 633 490 1017 524
rect 633 430 667 490
rect 599 424 667 430
rect 323 390 667 424
rect 37 388 103 390
rect 599 364 667 390
rect 701 390 893 456
rect 701 326 735 390
rect 498 260 735 326
rect 983 310 1017 490
rect 1151 412 1217 649
rect 1351 364 1417 649
rect 701 226 735 260
rect 983 244 1213 310
rect 23 184 667 218
rect 701 192 806 226
rect 983 224 1017 244
rect 23 70 89 184
rect 223 156 667 184
rect 123 17 189 150
rect 223 70 289 156
rect 323 17 389 122
rect 501 85 567 122
rect 601 119 667 156
rect 740 127 806 192
rect 840 190 1017 224
rect 840 85 874 190
rect 501 51 874 85
rect 908 17 1016 156
rect 1151 17 1217 128
rect 1351 17 1417 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 683 1440 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 0 617 1440 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 1440 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -49 1440 -17
<< labels >>
rlabel locali s 883 270 949 356 6 A1_N
port 1 nsew signal input
rlabel locali s 769 270 839 356 6 A2_N
port 2 nsew signal input
rlabel locali s 21 252 223 354 6 B1
port 3 nsew signal input
rlabel locali s 294 290 455 356 6 B2
port 4 nsew signal input
rlabel locali s 1251 378 1317 596 6 X
port 5 nsew signal output
rlabel locali s 1251 210 1317 344 6 X
port 5 nsew signal output
rlabel locali s 1251 70 1317 162 6 X
port 5 nsew signal output
rlabel locali s 1051 378 1117 596 6 X
port 5 nsew signal output
rlabel locali s 1051 344 1317 378 6 X
port 5 nsew signal output
rlabel locali s 1051 162 1317 210 6 X
port 5 nsew signal output
rlabel locali s 1051 70 1117 162 6 X
port 5 nsew signal output
rlabel metal1 s 0 -49 1440 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 7 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 617 1440 715 6 VPWR
port 9 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1440 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1213542
string GDS_START 1202516
<< end >>
