magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 83 47 113 177
rect 187 47 217 177
rect 271 47 301 177
rect 375 47 405 177
rect 586 47 616 177
rect 690 47 720 177
<< pmoshvt >>
rect 85 297 121 497
rect 179 297 215 497
rect 273 297 309 497
rect 367 297 403 497
rect 588 297 624 497
rect 682 297 718 497
<< ndiff >>
rect 28 163 83 177
rect 28 129 39 163
rect 73 129 83 163
rect 28 95 83 129
rect 28 61 39 95
rect 73 61 83 95
rect 28 47 83 61
rect 113 163 187 177
rect 113 129 133 163
rect 167 129 187 163
rect 113 95 187 129
rect 113 61 133 95
rect 167 61 187 95
rect 113 47 187 61
rect 217 95 271 177
rect 217 61 227 95
rect 261 61 271 95
rect 217 47 271 61
rect 301 163 375 177
rect 301 129 321 163
rect 355 129 375 163
rect 301 95 375 129
rect 301 61 321 95
rect 355 61 375 95
rect 301 47 375 61
rect 405 95 457 177
rect 405 61 415 95
rect 449 61 457 95
rect 405 47 457 61
rect 534 95 586 177
rect 534 61 542 95
rect 576 61 586 95
rect 534 47 586 61
rect 616 163 690 177
rect 616 129 636 163
rect 670 129 690 163
rect 616 95 690 129
rect 616 61 636 95
rect 670 61 690 95
rect 616 47 690 61
rect 720 95 772 177
rect 720 61 730 95
rect 764 61 772 95
rect 720 47 772 61
<< pdiff >>
rect 27 477 85 497
rect 27 443 39 477
rect 73 443 85 477
rect 27 409 85 443
rect 27 375 39 409
rect 73 375 85 409
rect 27 341 85 375
rect 27 307 39 341
rect 73 307 85 341
rect 27 297 85 307
rect 121 477 179 497
rect 121 443 133 477
rect 167 443 179 477
rect 121 409 179 443
rect 121 375 133 409
rect 167 375 179 409
rect 121 297 179 375
rect 215 477 273 497
rect 215 443 227 477
rect 261 443 273 477
rect 215 409 273 443
rect 215 375 227 409
rect 261 375 273 409
rect 215 341 273 375
rect 215 307 227 341
rect 261 307 273 341
rect 215 297 273 307
rect 309 477 367 497
rect 309 443 321 477
rect 355 443 367 477
rect 309 409 367 443
rect 309 375 321 409
rect 355 375 367 409
rect 309 297 367 375
rect 403 409 461 497
rect 403 375 415 409
rect 449 375 461 409
rect 403 341 461 375
rect 403 307 415 341
rect 449 307 461 341
rect 403 297 461 307
rect 534 477 588 497
rect 534 443 542 477
rect 576 443 588 477
rect 534 409 588 443
rect 534 375 542 409
rect 576 375 588 409
rect 534 297 588 375
rect 624 409 682 497
rect 624 375 636 409
rect 670 375 682 409
rect 624 341 682 375
rect 624 307 636 341
rect 670 307 682 341
rect 624 297 682 307
rect 718 477 772 497
rect 718 443 730 477
rect 764 443 772 477
rect 718 409 772 443
rect 718 375 730 409
rect 764 375 772 409
rect 718 297 772 375
<< ndiffc >>
rect 39 129 73 163
rect 39 61 73 95
rect 133 129 167 163
rect 133 61 167 95
rect 227 61 261 95
rect 321 129 355 163
rect 321 61 355 95
rect 415 61 449 95
rect 542 61 576 95
rect 636 129 670 163
rect 636 61 670 95
rect 730 61 764 95
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 133 443 167 477
rect 133 375 167 409
rect 227 443 261 477
rect 227 375 261 409
rect 227 307 261 341
rect 321 443 355 477
rect 321 375 355 409
rect 415 375 449 409
rect 415 307 449 341
rect 542 443 576 477
rect 542 375 576 409
rect 636 375 670 409
rect 636 307 670 341
rect 730 443 764 477
rect 730 375 764 409
<< poly >>
rect 85 497 121 523
rect 179 497 215 523
rect 273 497 309 523
rect 367 497 403 523
rect 588 497 624 523
rect 682 497 718 523
rect 85 282 121 297
rect 179 282 215 297
rect 273 282 309 297
rect 367 282 403 297
rect 588 282 624 297
rect 682 282 718 297
rect 83 265 123 282
rect 177 265 217 282
rect 83 249 217 265
rect 83 215 112 249
rect 146 215 217 249
rect 83 199 217 215
rect 83 177 113 199
rect 187 177 217 199
rect 271 265 311 282
rect 365 265 405 282
rect 271 249 405 265
rect 271 215 318 249
rect 352 215 405 249
rect 271 199 405 215
rect 271 177 301 199
rect 375 177 405 199
rect 586 265 626 282
rect 680 265 720 282
rect 586 249 720 265
rect 586 215 602 249
rect 636 215 720 249
rect 586 199 720 215
rect 586 177 616 199
rect 690 177 720 199
rect 83 21 113 47
rect 187 21 217 47
rect 271 21 301 47
rect 375 21 405 47
rect 586 21 616 47
rect 690 21 720 47
<< polycont >>
rect 112 215 146 249
rect 318 215 352 249
rect 602 215 636 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 30 477 81 493
rect 30 443 39 477
rect 73 443 81 477
rect 30 409 81 443
rect 30 375 39 409
rect 73 375 81 409
rect 30 341 81 375
rect 125 477 175 527
rect 125 443 133 477
rect 167 443 175 477
rect 125 409 175 443
rect 125 375 133 409
rect 167 375 175 409
rect 125 359 175 375
rect 219 477 269 493
rect 219 443 227 477
rect 261 443 269 477
rect 219 409 269 443
rect 219 375 227 409
rect 261 375 269 409
rect 30 307 39 341
rect 73 325 81 341
rect 219 341 269 375
rect 313 477 772 493
rect 313 443 321 477
rect 355 459 542 477
rect 355 443 363 459
rect 313 409 363 443
rect 576 459 730 477
rect 576 443 584 459
rect 313 375 321 409
rect 355 375 363 409
rect 313 359 363 375
rect 407 409 455 425
rect 407 375 415 409
rect 449 375 455 409
rect 219 325 227 341
rect 73 307 227 325
rect 261 325 269 341
rect 407 341 455 375
rect 542 409 584 443
rect 722 443 730 459
rect 764 443 772 477
rect 576 375 584 409
rect 542 359 584 375
rect 636 409 678 425
rect 670 375 678 409
rect 407 325 415 341
rect 261 307 415 325
rect 449 307 455 341
rect 636 341 678 375
rect 722 409 772 443
rect 722 375 730 409
rect 764 375 772 409
rect 722 359 772 375
rect 30 291 455 307
rect 489 257 587 325
rect 670 325 678 341
rect 670 307 799 325
rect 636 291 799 307
rect 27 249 203 257
rect 27 215 112 249
rect 146 215 203 249
rect 247 249 455 257
rect 247 215 318 249
rect 352 215 455 249
rect 489 249 662 257
rect 489 215 602 249
rect 636 215 662 249
rect 696 181 799 291
rect 18 163 73 181
rect 18 129 39 163
rect 18 95 73 129
rect 18 61 39 95
rect 18 17 73 61
rect 107 163 799 181
rect 107 129 133 163
rect 167 145 321 163
rect 167 129 183 145
rect 107 95 183 129
rect 295 129 321 145
rect 355 145 636 163
rect 355 129 371 145
rect 107 61 133 95
rect 167 61 183 95
rect 107 51 183 61
rect 227 95 261 111
rect 227 17 261 61
rect 295 95 371 129
rect 610 129 636 145
rect 670 145 799 163
rect 670 129 686 145
rect 295 61 321 95
rect 355 61 371 95
rect 295 51 371 61
rect 415 95 576 111
rect 449 61 542 95
rect 415 17 576 61
rect 610 95 686 129
rect 610 61 636 95
rect 670 61 686 95
rect 610 51 686 61
rect 730 95 788 111
rect 764 61 788 95
rect 730 17 788 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel corelocali s 493 221 527 255 0 FreeSans 400 0 0 0 C
port 3 nsew
flabel corelocali s 714 306 714 306 0 FreeSans 400 0 0 0 Y
port 8 nsew
flabel corelocali s 132 221 166 255 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 307 221 341 255 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
rlabel comment s 0 0 0 0 4 nor3_2
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2441178
string GDS_START 2434278
<< end >>
