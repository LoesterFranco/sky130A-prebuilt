magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 2208 561
rect 22 299 88 493
rect 123 333 157 493
rect 193 367 259 493
rect 295 333 329 493
rect 365 367 431 493
rect 467 333 501 493
rect 537 367 603 493
rect 639 333 673 493
rect 709 367 775 493
rect 811 333 845 493
rect 885 367 951 493
rect 1016 333 1050 493
rect 1090 367 1156 493
rect 1193 333 1227 493
rect 1263 367 1329 493
rect 1365 333 1399 493
rect 1435 367 1501 493
rect 1537 333 1571 493
rect 1607 367 1673 493
rect 1709 333 1743 493
rect 1779 367 1845 493
rect 1881 333 1915 493
rect 1951 367 2017 493
rect 2053 333 2087 493
rect 2122 367 2188 493
rect 123 291 2096 333
rect 465 283 1751 291
rect 69 179 431 255
rect 371 17 425 122
rect 465 56 510 283
rect 544 17 597 122
rect 631 56 682 283
rect 716 17 769 122
rect 803 56 851 283
rect 893 17 946 122
rect 981 56 1051 283
rect 1098 17 1151 122
rect 1185 56 1235 283
rect 1270 17 1315 122
rect 1357 56 1407 283
rect 1442 17 1495 122
rect 1529 56 1579 283
rect 1614 17 1667 122
rect 1701 56 1751 283
rect 1786 179 2142 255
rect 1786 17 1839 122
rect 0 -17 2208 17
<< metal1 >>
rect 0 496 2208 592
rect 14 428 2194 468
rect 14 416 72 428
rect 186 416 244 428
rect 366 416 424 428
rect 542 416 600 428
rect 726 416 784 428
rect 898 416 956 428
rect 1078 416 1136 428
rect 1262 416 1320 428
rect 1434 416 1492 428
rect 1614 416 1672 428
rect 1780 416 1838 428
rect 1952 416 2010 428
rect 2132 416 2190 428
rect 293 252 443 261
rect 1857 252 2007 261
rect 293 224 2007 252
rect 293 215 443 224
rect 1857 215 2007 224
rect 0 -48 2208 48
<< labels >>
rlabel locali s 69 179 431 255 6 A
port 1 nsew signal input
rlabel locali s 1786 179 2142 255 6 A
port 1 nsew signal input
rlabel metal1 s 1857 252 2007 261 6 A
port 1 nsew signal input
rlabel metal1 s 1857 215 2007 224 6 A
port 1 nsew signal input
rlabel metal1 s 293 252 443 261 6 A
port 1 nsew signal input
rlabel metal1 s 293 224 2007 252 6 A
port 1 nsew signal input
rlabel metal1 s 293 215 443 224 6 A
port 1 nsew signal input
rlabel locali s 2053 333 2087 493 6 Y
port 2 nsew signal output
rlabel locali s 1881 333 1915 493 6 Y
port 2 nsew signal output
rlabel locali s 1709 333 1743 493 6 Y
port 2 nsew signal output
rlabel locali s 1701 56 1751 283 6 Y
port 2 nsew signal output
rlabel locali s 1537 333 1571 493 6 Y
port 2 nsew signal output
rlabel locali s 1529 56 1579 283 6 Y
port 2 nsew signal output
rlabel locali s 1365 333 1399 493 6 Y
port 2 nsew signal output
rlabel locali s 1357 56 1407 283 6 Y
port 2 nsew signal output
rlabel locali s 1193 333 1227 493 6 Y
port 2 nsew signal output
rlabel locali s 1185 56 1235 283 6 Y
port 2 nsew signal output
rlabel locali s 1016 333 1050 493 6 Y
port 2 nsew signal output
rlabel locali s 981 56 1051 283 6 Y
port 2 nsew signal output
rlabel locali s 811 333 845 493 6 Y
port 2 nsew signal output
rlabel locali s 803 56 851 283 6 Y
port 2 nsew signal output
rlabel locali s 639 333 673 493 6 Y
port 2 nsew signal output
rlabel locali s 631 56 682 283 6 Y
port 2 nsew signal output
rlabel locali s 467 333 501 493 6 Y
port 2 nsew signal output
rlabel locali s 465 283 1751 291 6 Y
port 2 nsew signal output
rlabel locali s 465 56 510 283 6 Y
port 2 nsew signal output
rlabel locali s 295 333 329 493 6 Y
port 2 nsew signal output
rlabel locali s 123 333 157 493 6 Y
port 2 nsew signal output
rlabel locali s 123 291 2096 333 6 Y
port 2 nsew signal output
rlabel locali s 22 299 88 493 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 193 367 259 493 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 365 367 431 493 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 2122 367 2188 493 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 537 367 603 493 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 709 367 775 493 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 885 367 951 493 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 1090 367 1156 493 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 1263 367 1329 493 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 1435 367 1501 493 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 1607 367 1673 493 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 1779 367 1845 493 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 1951 367 2017 493 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 2132 416 2190 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 1952 416 2010 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 1780 416 1838 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 1614 416 1672 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 1434 416 1492 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 1262 416 1320 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 1078 416 1136 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 898 416 956 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 726 416 784 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 542 416 600 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 366 416 424 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 186 416 244 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 14 428 2194 468 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 14 416 72 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 1786 17 1839 122 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 1614 17 1667 122 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 1442 17 1495 122 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 1270 17 1315 122 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 1098 17 1151 122 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 893 17 946 122 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 716 17 769 122 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 544 17 597 122 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 371 17 425 122 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 2208 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 2208 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 527 2208 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 2208 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2208 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2250552
string GDS_START 2235310
<< end >>
