magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 295 333 371 425
rect 295 289 462 333
rect 18 215 172 255
rect 206 215 380 255
rect 419 181 462 289
rect 107 147 462 181
rect 107 145 371 147
rect 107 51 183 145
rect 295 51 371 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 18 333 73 493
rect 107 367 183 527
rect 227 459 475 493
rect 227 333 261 459
rect 18 291 261 333
rect 415 367 475 459
rect 18 17 73 181
rect 227 17 261 111
rect 428 17 496 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
rlabel locali s 18 215 172 255 6 A
port 1 nsew signal input
rlabel locali s 206 215 380 255 6 B
port 2 nsew signal input
rlabel locali s 419 181 462 289 6 Y
port 3 nsew signal output
rlabel locali s 295 333 371 425 6 Y
port 3 nsew signal output
rlabel locali s 295 289 462 333 6 Y
port 3 nsew signal output
rlabel locali s 295 51 371 145 6 Y
port 3 nsew signal output
rlabel locali s 107 147 462 181 6 Y
port 3 nsew signal output
rlabel locali s 107 145 371 147 6 Y
port 3 nsew signal output
rlabel locali s 107 51 183 145 6 Y
port 3 nsew signal output
rlabel metal1 s 0 -48 552 48 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 496 552 592 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 552 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2390238
string GDS_START 2385208
<< end >>
