magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 710 704
<< pwell >>
rect 0 0 672 49
<< scnmos >>
rect 84 74 114 202
rect 299 74 329 222
rect 385 74 415 222
rect 471 74 501 222
rect 558 74 588 222
<< pmoshvt >>
rect 86 368 116 568
rect 286 368 316 592
rect 376 368 406 592
rect 466 368 496 592
rect 556 368 586 592
<< ndiff >>
rect 27 190 84 202
rect 27 156 39 190
rect 73 156 84 190
rect 27 120 84 156
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 164 164 202
rect 249 196 299 222
rect 242 188 299 196
rect 114 152 167 164
rect 114 118 125 152
rect 159 118 167 152
rect 114 74 167 118
rect 242 154 254 188
rect 288 154 299 188
rect 242 120 299 154
rect 242 86 254 120
rect 288 86 299 120
rect 242 74 299 86
rect 329 182 385 222
rect 329 148 340 182
rect 374 148 385 182
rect 329 74 385 148
rect 415 210 471 222
rect 415 176 426 210
rect 460 176 471 210
rect 415 120 471 176
rect 415 86 426 120
rect 460 86 471 120
rect 415 74 471 86
rect 501 210 558 222
rect 501 176 512 210
rect 546 176 558 210
rect 501 120 558 176
rect 501 86 512 120
rect 546 86 558 120
rect 501 74 558 86
rect 588 210 645 222
rect 588 176 599 210
rect 633 176 645 210
rect 588 120 645 176
rect 588 86 599 120
rect 633 86 645 120
rect 588 74 645 86
<< pdiff >>
rect 165 570 286 592
rect 165 568 173 570
rect 27 556 86 568
rect 27 522 39 556
rect 73 522 86 556
rect 27 440 86 522
rect 27 406 39 440
rect 73 406 86 440
rect 27 368 86 406
rect 116 536 173 568
rect 207 536 286 570
rect 116 498 286 536
rect 116 464 166 498
rect 200 464 286 498
rect 116 368 286 464
rect 316 419 376 592
rect 316 385 329 419
rect 363 385 376 419
rect 316 368 376 385
rect 406 578 466 592
rect 406 544 419 578
rect 453 544 466 578
rect 406 368 466 544
rect 496 440 556 592
rect 496 406 509 440
rect 543 406 556 440
rect 496 368 556 406
rect 586 578 645 592
rect 586 544 599 578
rect 633 544 645 578
rect 586 368 645 544
<< ndiffc >>
rect 39 156 73 190
rect 39 86 73 120
rect 125 118 159 152
rect 254 154 288 188
rect 254 86 288 120
rect 340 148 374 182
rect 426 176 460 210
rect 426 86 460 120
rect 512 176 546 210
rect 512 86 546 120
rect 599 176 633 210
rect 599 86 633 120
<< pdiffc >>
rect 39 522 73 556
rect 39 406 73 440
rect 173 536 207 570
rect 166 464 200 498
rect 329 385 363 419
rect 419 544 453 578
rect 509 406 543 440
rect 599 544 633 578
<< poly >>
rect 86 568 116 594
rect 286 592 316 618
rect 376 592 406 618
rect 466 592 496 618
rect 556 592 586 618
rect 86 353 116 368
rect 286 353 316 368
rect 376 353 406 368
rect 466 353 496 368
rect 556 353 586 368
rect 83 342 116 353
rect 83 336 114 342
rect 48 320 114 336
rect 48 286 64 320
rect 98 286 114 320
rect 283 294 319 353
rect 373 294 409 353
rect 463 336 499 353
rect 553 336 589 353
rect 463 320 589 336
rect 48 270 114 286
rect 84 202 114 270
rect 161 278 415 294
rect 161 244 177 278
rect 211 264 415 278
rect 463 286 505 320
rect 539 286 589 320
rect 463 270 589 286
rect 211 244 227 264
rect 161 228 227 244
rect 299 222 329 264
rect 385 222 415 264
rect 471 222 501 270
rect 558 222 588 270
rect 84 48 114 74
rect 299 48 329 74
rect 385 48 415 74
rect 471 48 501 74
rect 558 48 588 74
<< polycont >>
rect 64 286 98 320
rect 177 244 211 278
rect 505 286 539 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 23 556 89 572
rect 23 522 39 556
rect 73 522 89 556
rect 23 440 89 522
rect 145 570 219 649
rect 145 536 173 570
rect 207 536 219 570
rect 403 578 469 649
rect 403 544 419 578
rect 453 544 469 578
rect 403 542 469 544
rect 583 578 649 649
rect 583 544 599 578
rect 633 544 649 578
rect 583 542 649 544
rect 145 498 219 536
rect 145 464 166 498
rect 200 464 219 498
rect 145 458 219 464
rect 261 474 649 508
rect 23 406 39 440
rect 73 424 89 440
rect 73 406 195 424
rect 23 390 195 406
rect 25 320 114 356
rect 25 286 64 320
rect 98 286 114 320
rect 25 270 114 286
rect 161 294 195 390
rect 161 278 227 294
rect 161 244 177 278
rect 211 244 227 278
rect 161 236 227 244
rect 23 228 227 236
rect 23 202 195 228
rect 23 190 89 202
rect 261 194 295 474
rect 329 419 509 440
rect 363 406 509 419
rect 543 406 559 440
rect 363 390 559 406
rect 363 385 455 390
rect 329 364 455 385
rect 409 278 455 364
rect 340 244 455 278
rect 489 320 555 356
rect 489 286 505 320
rect 539 286 555 320
rect 489 270 555 286
rect 23 156 39 190
rect 73 156 89 190
rect 238 188 304 194
rect 23 120 89 156
rect 23 86 39 120
rect 73 86 89 120
rect 23 70 89 86
rect 123 152 175 168
rect 123 118 125 152
rect 159 118 175 152
rect 123 17 175 118
rect 238 154 254 188
rect 288 154 304 188
rect 238 120 304 154
rect 340 182 374 244
rect 615 226 649 474
rect 512 210 546 226
rect 340 126 374 148
rect 410 176 426 210
rect 460 176 476 210
rect 238 86 254 120
rect 288 86 304 120
rect 238 85 304 86
rect 410 120 476 176
rect 410 86 426 120
rect 460 86 476 120
rect 410 85 476 86
rect 238 51 476 85
rect 512 120 546 176
rect 512 17 546 86
rect 583 210 649 226
rect 583 176 599 210
rect 633 176 649 210
rect 583 120 649 176
rect 583 86 599 120
rect 633 86 649 120
rect 583 70 649 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel comment s 0 0 0 0 4 nand2b_2
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 Y
port 7 nsew
flabel corelocali s 415 390 449 424 0 FreeSans 340 0 0 0 Y
port 7 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 672 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1656174
string GDS_START 1650326
<< end >>
