magic
tech sky130A
magscale 1 2
timestamp 1604502697
<< nwell >>
rect -38 261 1326 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 89 47 119 131
rect 183 47 213 131
rect 381 47 411 131
rect 475 47 505 131
rect 583 47 613 119
rect 688 47 718 119
rect 783 47 813 131
rect 991 47 1021 177
rect 1085 47 1115 177
rect 1179 47 1209 177
<< pmoshvt >>
rect 81 363 117 491
rect 175 363 211 491
rect 373 369 409 497
rect 467 369 503 497
rect 572 413 608 497
rect 703 413 739 497
rect 785 413 821 497
rect 983 297 1019 497
rect 1077 297 1113 497
rect 1171 297 1207 497
<< ndiff >>
rect 27 119 89 131
rect 27 85 35 119
rect 69 85 89 119
rect 27 47 89 85
rect 119 93 183 131
rect 119 59 129 93
rect 163 59 183 93
rect 119 47 183 59
rect 213 119 265 131
rect 213 85 223 119
rect 257 85 265 119
rect 213 47 265 85
rect 319 119 381 131
rect 319 85 327 119
rect 361 85 381 119
rect 319 47 381 85
rect 411 89 475 131
rect 411 55 421 89
rect 455 55 475 89
rect 411 47 475 55
rect 505 119 555 131
rect 929 133 991 177
rect 733 119 783 131
rect 505 47 583 119
rect 613 107 688 119
rect 613 73 633 107
rect 667 73 688 107
rect 613 47 688 73
rect 718 47 783 119
rect 813 106 875 131
rect 813 72 833 106
rect 867 72 875 106
rect 813 47 875 72
rect 929 99 937 133
rect 971 99 991 133
rect 929 47 991 99
rect 1021 127 1085 177
rect 1021 93 1031 127
rect 1065 93 1085 127
rect 1021 47 1085 93
rect 1115 133 1179 177
rect 1115 99 1125 133
rect 1159 99 1179 133
rect 1115 47 1179 99
rect 1209 93 1261 177
rect 1209 59 1219 93
rect 1253 59 1261 93
rect 1209 47 1261 59
<< pdiff >>
rect 27 477 81 491
rect 27 443 35 477
rect 69 443 81 477
rect 27 409 81 443
rect 27 375 35 409
rect 69 375 81 409
rect 27 363 81 375
rect 117 461 175 491
rect 117 427 129 461
rect 163 427 175 461
rect 117 363 175 427
rect 211 477 265 491
rect 211 443 223 477
rect 257 443 265 477
rect 211 409 265 443
rect 211 375 223 409
rect 257 375 265 409
rect 211 363 265 375
rect 319 483 373 497
rect 319 449 327 483
rect 361 449 373 483
rect 319 415 373 449
rect 319 381 327 415
rect 361 381 373 415
rect 319 369 373 381
rect 409 485 467 497
rect 409 451 421 485
rect 455 451 467 485
rect 409 417 467 451
rect 409 383 421 417
rect 455 383 467 417
rect 409 369 467 383
rect 503 413 572 497
rect 608 485 703 497
rect 608 451 645 485
rect 679 451 703 485
rect 608 413 703 451
rect 739 413 785 497
rect 821 477 875 497
rect 821 443 833 477
rect 867 443 875 477
rect 821 413 875 443
rect 929 471 983 497
rect 929 437 937 471
rect 971 437 983 471
rect 503 369 555 413
rect 929 368 983 437
rect 929 334 937 368
rect 971 334 983 368
rect 929 297 983 334
rect 1019 484 1077 497
rect 1019 450 1031 484
rect 1065 450 1077 484
rect 1019 364 1077 450
rect 1019 330 1031 364
rect 1065 330 1077 364
rect 1019 297 1077 330
rect 1113 475 1171 497
rect 1113 441 1125 475
rect 1159 441 1171 475
rect 1113 384 1171 441
rect 1113 350 1125 384
rect 1159 350 1171 384
rect 1113 297 1171 350
rect 1207 485 1261 497
rect 1207 451 1219 485
rect 1253 451 1261 485
rect 1207 417 1261 451
rect 1207 383 1219 417
rect 1253 383 1261 417
rect 1207 297 1261 383
<< ndiffc >>
rect 35 85 69 119
rect 129 59 163 93
rect 223 85 257 119
rect 327 85 361 119
rect 421 55 455 89
rect 633 73 667 107
rect 833 72 867 106
rect 937 99 971 133
rect 1031 93 1065 127
rect 1125 99 1159 133
rect 1219 59 1253 93
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 129 427 163 461
rect 223 443 257 477
rect 223 375 257 409
rect 327 449 361 483
rect 327 381 361 415
rect 421 451 455 485
rect 421 383 455 417
rect 645 451 679 485
rect 833 443 867 477
rect 937 437 971 471
rect 937 334 971 368
rect 1031 450 1065 484
rect 1031 330 1065 364
rect 1125 441 1159 475
rect 1125 350 1159 384
rect 1219 451 1253 485
rect 1219 383 1253 417
<< poly >>
rect 81 491 117 517
rect 175 491 211 517
rect 373 497 409 523
rect 467 497 503 523
rect 572 497 608 523
rect 703 497 739 523
rect 785 497 821 523
rect 983 497 1019 523
rect 1077 497 1113 523
rect 1171 497 1207 523
rect 572 398 608 413
rect 703 398 739 413
rect 785 398 821 413
rect 81 348 117 363
rect 175 348 211 363
rect 373 354 409 369
rect 467 354 503 369
rect 46 318 119 348
rect 46 280 76 318
rect 21 264 76 280
rect 173 274 213 348
rect 21 230 32 264
rect 66 230 76 264
rect 21 214 76 230
rect 128 264 213 274
rect 128 230 144 264
rect 178 230 213 264
rect 371 241 411 354
rect 128 220 213 230
rect 46 176 76 214
rect 46 146 119 176
rect 89 131 119 146
rect 183 131 213 220
rect 318 225 411 241
rect 318 191 328 225
rect 362 191 411 225
rect 465 219 505 354
rect 570 337 610 398
rect 701 375 741 398
rect 547 321 610 337
rect 652 365 741 375
rect 652 331 668 365
rect 702 331 741 365
rect 652 321 741 331
rect 783 373 823 398
rect 783 357 881 373
rect 783 323 837 357
rect 871 323 881 357
rect 547 287 557 321
rect 591 287 610 321
rect 547 279 610 287
rect 783 307 881 323
rect 547 271 718 279
rect 571 249 718 271
rect 318 175 411 191
rect 381 131 411 175
rect 454 203 518 219
rect 454 169 464 203
rect 498 169 518 203
rect 454 153 518 169
rect 573 191 637 207
rect 573 157 583 191
rect 617 157 637 191
rect 475 131 505 153
rect 573 141 637 157
rect 583 119 613 141
rect 688 119 718 249
rect 783 131 813 307
rect 983 282 1019 297
rect 1077 282 1113 297
rect 1171 282 1207 297
rect 981 265 1021 282
rect 1075 265 1115 282
rect 1169 265 1209 282
rect 865 249 1021 265
rect 865 215 875 249
rect 909 215 1021 249
rect 865 199 1021 215
rect 1063 249 1209 265
rect 1063 215 1073 249
rect 1107 215 1209 249
rect 1063 199 1209 215
rect 991 177 1021 199
rect 1085 177 1115 199
rect 1179 177 1209 199
rect 89 21 119 47
rect 183 21 213 47
rect 381 21 411 47
rect 475 21 505 47
rect 583 21 613 47
rect 688 21 718 47
rect 783 21 813 47
rect 991 21 1021 47
rect 1085 21 1115 47
rect 1179 21 1209 47
<< polycont >>
rect 32 230 66 264
rect 144 230 178 264
rect 328 191 362 225
rect 668 331 702 365
rect 837 323 871 357
rect 557 287 591 321
rect 464 169 498 203
rect 583 157 617 191
rect 875 215 909 249
rect 1073 215 1107 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 35 477 69 493
rect 35 409 69 443
rect 103 461 179 527
rect 103 427 129 461
rect 163 427 179 461
rect 223 477 268 493
rect 421 485 484 527
rect 257 443 268 477
rect 223 409 268 443
rect 69 375 166 393
rect 35 359 166 375
rect 17 264 66 325
rect 17 230 32 264
rect 17 197 66 230
rect 132 323 166 359
rect 132 280 166 289
rect 257 391 268 409
rect 223 357 234 375
rect 223 337 268 357
rect 311 449 327 483
rect 361 449 377 483
rect 311 415 377 449
rect 311 381 327 415
rect 361 381 377 415
rect 132 264 178 280
rect 132 230 144 264
rect 132 214 178 230
rect 132 161 166 214
rect 35 127 166 161
rect 35 119 69 127
rect 223 119 257 337
rect 311 333 377 381
rect 455 451 484 485
rect 629 451 645 485
rect 679 451 789 485
rect 421 417 484 451
rect 455 383 484 417
rect 421 367 484 383
rect 534 391 591 401
rect 568 357 591 391
rect 311 299 458 333
rect 293 225 378 265
rect 293 191 328 225
rect 362 191 378 225
rect 424 219 458 299
rect 534 321 591 357
rect 534 287 557 321
rect 534 271 591 287
rect 634 365 702 399
rect 634 331 668 365
rect 634 323 702 331
rect 634 289 635 323
rect 669 289 702 323
rect 634 283 702 289
rect 424 203 508 219
rect 634 207 668 283
rect 755 265 789 451
rect 833 477 893 527
rect 867 443 893 477
rect 833 427 893 443
rect 937 471 981 487
rect 971 437 981 471
rect 937 373 981 437
rect 837 368 981 373
rect 837 357 937 368
rect 871 334 937 357
rect 971 334 981 368
rect 871 323 981 334
rect 837 307 981 323
rect 947 265 981 307
rect 1027 484 1081 527
rect 1027 450 1031 484
rect 1065 450 1081 484
rect 1027 364 1081 450
rect 1027 330 1031 364
rect 1065 330 1081 364
rect 1027 299 1081 330
rect 1125 475 1182 491
rect 1159 441 1182 475
rect 1125 384 1182 441
rect 1159 350 1182 384
rect 1219 485 1269 527
rect 1253 451 1269 485
rect 1219 417 1269 451
rect 1253 383 1269 417
rect 1219 351 1269 383
rect 1125 299 1182 350
rect 1148 265 1182 299
rect 755 249 909 265
rect 755 233 875 249
rect 424 169 464 203
rect 498 169 508 203
rect 424 157 508 169
rect 35 69 69 85
rect 103 59 129 93
rect 163 59 179 93
rect 223 69 257 85
rect 327 153 508 157
rect 583 191 668 207
rect 617 157 668 191
rect 327 123 458 153
rect 583 141 668 157
rect 725 215 875 233
rect 725 199 909 215
rect 947 249 1107 265
rect 947 215 1073 249
rect 947 199 1107 215
rect 1148 199 1269 265
rect 327 119 361 123
rect 725 107 759 199
rect 947 165 981 199
rect 1148 165 1182 199
rect 327 69 361 85
rect 103 17 179 59
rect 395 55 421 89
rect 455 55 471 89
rect 617 73 633 107
rect 667 73 759 107
rect 807 106 883 165
rect 395 17 471 55
rect 807 72 833 106
rect 867 72 883 106
rect 937 133 981 165
rect 971 99 981 133
rect 937 83 981 99
rect 1027 127 1081 165
rect 1027 93 1031 127
rect 1065 93 1081 127
rect 807 17 883 72
rect 1027 17 1081 93
rect 1125 133 1182 165
rect 1159 99 1182 133
rect 1125 83 1182 99
rect 1219 93 1271 110
rect 1253 59 1271 93
rect 1219 17 1271 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 132 289 166 323
rect 234 375 257 391
rect 257 375 268 391
rect 234 357 268 375
rect 534 357 568 391
rect 635 289 669 323
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 222 391 280 397
rect 222 357 234 391
rect 268 388 280 391
rect 522 391 580 397
rect 522 388 534 391
rect 268 360 534 388
rect 268 357 280 360
rect 222 351 280 357
rect 522 357 534 360
rect 568 357 580 391
rect 522 351 580 357
rect 120 323 178 329
rect 120 289 132 323
rect 166 320 178 323
rect 623 323 681 329
rect 623 320 635 323
rect 166 292 635 320
rect 166 289 178 292
rect 120 283 178 289
rect 623 289 635 292
rect 669 289 681 323
rect 623 283 681 289
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
flabel corelocali s 309 221 343 255 0 FreeSans 200 0 0 0 D
port 1 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 200 0 0 0 GATE_N
port 2 nsew
flabel corelocali s 1136 357 1170 391 0 FreeSans 200 0 0 0 Q
port 7 nsew
flabel corelocali s 30 289 64 323 0 FreeSans 200 0 0 0 GATE_N
port 2 nsew
flabel corelocali s 1136 425 1170 459 0 FreeSans 200 0 0 0 Q
port 7 nsew
flabel corelocali s 1136 85 1170 119 0 FreeSans 200 0 0 0 Q
port 7 nsew
flabel corelocali s 1225 221 1259 255 0 FreeSans 200 0 0 0 Q
port 7 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew
rlabel comment s 0 0 0 0 4 dlxtn_2
<< properties >>
string FIXED_BBOX 0 0 1288 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1948698
string GDS_START 1938194
<< end >>
