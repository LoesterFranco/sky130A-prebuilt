magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 509 349 543 425
rect 697 349 731 425
rect 509 289 898 349
rect 28 215 390 255
rect 464 215 767 255
rect 819 181 898 289
rect 107 145 898 181
rect 107 51 183 145
rect 295 51 371 145
rect 483 51 559 145
rect 671 51 747 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 18 333 73 493
rect 107 367 183 527
rect 227 333 261 493
rect 295 367 355 527
rect 389 459 858 493
rect 389 333 465 459
rect 18 291 465 333
rect 577 387 653 459
rect 765 383 858 459
rect 18 17 73 181
rect 227 17 261 111
rect 415 17 449 111
rect 603 17 637 111
rect 791 17 848 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
rlabel locali s 28 215 390 255 6 A
port 1 nsew signal input
rlabel locali s 464 215 767 255 6 B
port 2 nsew signal input
rlabel locali s 819 181 898 289 6 Y
port 3 nsew signal output
rlabel locali s 697 349 731 425 6 Y
port 3 nsew signal output
rlabel locali s 671 51 747 145 6 Y
port 3 nsew signal output
rlabel locali s 509 349 543 425 6 Y
port 3 nsew signal output
rlabel locali s 509 289 898 349 6 Y
port 3 nsew signal output
rlabel locali s 483 51 559 145 6 Y
port 3 nsew signal output
rlabel locali s 295 51 371 145 6 Y
port 3 nsew signal output
rlabel locali s 107 145 898 181 6 Y
port 3 nsew signal output
rlabel locali s 107 51 183 145 6 Y
port 3 nsew signal output
rlabel metal1 s 0 -48 920 48 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 496 920 592 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 920 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2397758
string GDS_START 2390296
<< end >>
