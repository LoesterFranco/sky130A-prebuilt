magic
tech sky130A
magscale 1 2
timestamp 1601050082
<< locali >>
rect 121 364 184 596
rect 123 226 157 364
rect 123 70 178 226
rect 305 236 371 310
rect 409 236 485 310
rect 533 236 647 310
rect 681 236 747 310
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 37 364 87 649
rect 218 412 325 649
rect 359 446 425 572
rect 470 480 536 649
rect 577 446 643 572
rect 359 412 643 446
rect 677 378 745 572
rect 227 344 745 378
rect 227 326 261 344
rect 191 260 261 326
rect 23 17 89 226
rect 227 202 261 260
rect 227 168 636 202
rect 212 17 346 120
rect 570 70 636 168
rect 672 17 738 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel locali s 533 236 647 310 6 A1
port 1 nsew signal input
rlabel locali s 409 236 485 310 6 A2
port 2 nsew signal input
rlabel locali s 305 236 371 310 6 A3
port 3 nsew signal input
rlabel locali s 681 236 747 310 6 B1
port 4 nsew signal input
rlabel locali s 123 226 157 364 6 X
port 5 nsew signal output
rlabel locali s 123 70 178 226 6 X
port 5 nsew signal output
rlabel locali s 121 364 184 596 6 X
port 5 nsew signal output
rlabel metal1 s 0 -49 768 49 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 617 768 715 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3692238
string GDS_START 3685232
<< end >>
