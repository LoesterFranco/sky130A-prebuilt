magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 134 704
<< pwell >>
rect 0 0 96 49
<< locali >>
rect 0 649 31 683
rect 65 649 96 683
rect 0 -17 31 17
rect 65 -17 96 17
<< viali >>
rect 31 649 65 683
rect 31 -17 65 17
<< metal1 >>
rect 0 683 96 715
rect 0 649 31 683
rect 65 649 96 683
rect 0 617 96 649
rect 0 17 96 49
rect 0 -17 31 17
rect 65 -17 96 17
rect 0 -49 96 -17
<< labels >>
flabel pwell s 0 0 96 49 0 FreeSans 200 0 0 0 VNB
port 2 nsew
flabel nwell s 0 617 96 666 0 FreeSans 200 0 0 0 VPB
port 3 nsew
rlabel comment s 0 0 0 0 4 fill_1
flabel metal1 s 0 617 96 666 0 FreeSans 200 0 0 0 VPWR
port 4 nsew
flabel metal1 s 0 0 96 49 0 FreeSans 200 0 0 0 VGND
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 96 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2200526
string GDS_START 2199234
<< end >>
