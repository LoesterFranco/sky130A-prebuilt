magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 998 704
<< pwell >>
rect 0 0 960 49
<< scnmos >>
rect 91 74 121 222
rect 169 74 199 222
rect 283 74 313 222
rect 411 74 441 222
rect 519 74 549 222
rect 635 74 665 222
rect 747 74 777 222
<< pmoshvt >>
rect 86 392 116 592
rect 196 392 226 592
rect 286 392 316 592
rect 432 392 462 592
rect 522 392 552 592
rect 744 368 774 592
rect 834 368 864 592
<< ndiff >>
rect 34 195 91 222
rect 34 161 46 195
rect 80 161 91 195
rect 34 120 91 161
rect 34 86 46 120
rect 80 86 91 120
rect 34 74 91 86
rect 121 74 169 222
rect 199 74 283 222
rect 313 74 411 222
rect 441 210 519 222
rect 441 176 462 210
rect 496 176 519 210
rect 441 120 519 176
rect 441 86 462 120
rect 496 86 519 120
rect 441 74 519 86
rect 549 188 635 222
rect 549 154 574 188
rect 608 154 635 188
rect 549 120 635 154
rect 549 86 574 120
rect 608 86 635 120
rect 549 74 635 86
rect 665 188 747 222
rect 665 154 693 188
rect 727 154 747 188
rect 665 116 747 154
rect 665 82 693 116
rect 727 82 747 116
rect 665 74 747 82
rect 777 120 933 222
rect 777 86 793 120
rect 827 86 887 120
rect 921 86 933 120
rect 777 74 933 86
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 509 86 546
rect 27 475 39 509
rect 73 475 86 509
rect 27 438 86 475
rect 27 404 39 438
rect 73 404 86 438
rect 27 392 86 404
rect 116 582 196 592
rect 116 548 139 582
rect 173 548 196 582
rect 116 514 196 548
rect 116 480 139 514
rect 173 480 196 514
rect 116 446 196 480
rect 116 412 139 446
rect 173 412 196 446
rect 116 392 196 412
rect 226 580 286 592
rect 226 546 239 580
rect 273 546 286 580
rect 226 509 286 546
rect 226 475 239 509
rect 273 475 286 509
rect 226 438 286 475
rect 226 404 239 438
rect 273 404 286 438
rect 226 392 286 404
rect 316 580 432 592
rect 316 546 357 580
rect 391 546 432 580
rect 316 492 432 546
rect 316 458 357 492
rect 391 458 432 492
rect 316 392 432 458
rect 462 580 522 592
rect 462 546 475 580
rect 509 546 522 580
rect 462 510 522 546
rect 462 476 475 510
rect 509 476 522 510
rect 462 440 522 476
rect 462 406 475 440
rect 509 406 522 440
rect 462 392 522 406
rect 552 580 621 592
rect 552 546 575 580
rect 609 546 621 580
rect 552 510 621 546
rect 552 476 575 510
rect 609 476 621 510
rect 552 440 621 476
rect 552 406 575 440
rect 609 406 621 440
rect 552 392 621 406
rect 675 580 744 592
rect 675 546 687 580
rect 721 546 744 580
rect 675 493 744 546
rect 675 459 687 493
rect 721 459 744 493
rect 675 368 744 459
rect 774 580 834 592
rect 774 546 787 580
rect 821 546 834 580
rect 774 497 834 546
rect 774 463 787 497
rect 821 463 834 497
rect 774 414 834 463
rect 774 380 787 414
rect 821 380 834 414
rect 774 368 834 380
rect 864 580 933 592
rect 864 546 887 580
rect 921 546 933 580
rect 864 497 933 546
rect 864 463 887 497
rect 921 463 933 497
rect 864 414 933 463
rect 864 380 887 414
rect 921 380 933 414
rect 864 368 933 380
<< ndiffc >>
rect 46 161 80 195
rect 46 86 80 120
rect 462 176 496 210
rect 462 86 496 120
rect 574 154 608 188
rect 574 86 608 120
rect 693 154 727 188
rect 693 82 727 116
rect 793 86 827 120
rect 887 86 921 120
<< pdiffc >>
rect 39 546 73 580
rect 39 475 73 509
rect 39 404 73 438
rect 139 548 173 582
rect 139 480 173 514
rect 139 412 173 446
rect 239 546 273 580
rect 239 475 273 509
rect 239 404 273 438
rect 357 546 391 580
rect 357 458 391 492
rect 475 546 509 580
rect 475 476 509 510
rect 475 406 509 440
rect 575 546 609 580
rect 575 476 609 510
rect 575 406 609 440
rect 687 546 721 580
rect 687 459 721 493
rect 787 546 821 580
rect 787 463 821 497
rect 787 380 821 414
rect 887 546 921 580
rect 887 463 921 497
rect 887 380 921 414
<< poly >>
rect 86 592 116 618
rect 196 592 226 618
rect 286 592 316 618
rect 432 592 462 618
rect 522 592 552 618
rect 744 592 774 618
rect 834 592 864 618
rect 86 377 116 392
rect 196 377 226 392
rect 286 377 316 392
rect 432 377 462 392
rect 522 377 552 392
rect 83 310 119 377
rect 193 310 229 377
rect 283 310 319 377
rect 429 356 465 377
rect 519 356 555 377
rect 405 340 471 356
rect 25 294 121 310
rect 25 260 41 294
rect 75 260 121 294
rect 25 244 121 260
rect 91 222 121 244
rect 169 294 235 310
rect 169 260 185 294
rect 219 260 235 294
rect 169 244 235 260
rect 283 294 363 310
rect 283 260 313 294
rect 347 260 363 294
rect 405 306 421 340
rect 455 306 471 340
rect 405 290 471 306
rect 519 340 585 356
rect 744 353 774 368
rect 834 353 864 368
rect 519 306 535 340
rect 569 306 585 340
rect 741 310 777 353
rect 831 310 867 353
rect 519 290 585 306
rect 635 294 867 310
rect 283 244 363 260
rect 169 222 199 244
rect 283 222 313 244
rect 411 222 441 290
rect 519 222 549 290
rect 635 260 651 294
rect 685 260 719 294
rect 753 260 867 294
rect 635 244 867 260
rect 635 222 665 244
rect 747 222 777 244
rect 91 48 121 74
rect 169 48 199 74
rect 283 48 313 74
rect 411 48 441 74
rect 519 48 549 74
rect 635 48 665 74
rect 747 48 777 74
<< polycont >>
rect 41 260 75 294
rect 185 260 219 294
rect 313 260 347 294
rect 421 306 455 340
rect 535 306 569 340
rect 651 260 685 294
rect 719 260 753 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 23 580 89 596
rect 23 546 39 580
rect 73 546 89 580
rect 23 509 89 546
rect 23 475 39 509
rect 73 475 89 509
rect 23 438 89 475
rect 23 404 39 438
rect 73 404 89 438
rect 123 582 189 649
rect 123 548 139 582
rect 173 548 189 582
rect 123 514 189 548
rect 123 480 139 514
rect 173 480 189 514
rect 123 446 189 480
rect 123 412 139 446
rect 173 412 189 446
rect 223 580 289 596
rect 223 546 239 580
rect 273 546 289 580
rect 223 509 289 546
rect 223 475 239 509
rect 273 475 289 509
rect 223 438 289 475
rect 323 580 425 649
rect 323 546 357 580
rect 391 546 425 580
rect 323 492 425 546
rect 323 458 357 492
rect 391 458 425 492
rect 459 580 525 596
rect 459 546 475 580
rect 509 546 525 580
rect 459 510 525 546
rect 459 476 475 510
rect 509 476 525 510
rect 23 378 89 404
rect 223 404 239 438
rect 273 424 289 438
rect 459 440 525 476
rect 459 424 475 440
rect 273 406 475 424
rect 509 406 525 440
rect 273 404 525 406
rect 223 390 525 404
rect 559 580 625 596
rect 559 546 575 580
rect 609 546 625 580
rect 559 510 625 546
rect 559 476 575 510
rect 609 476 625 510
rect 559 440 625 476
rect 671 580 737 649
rect 671 546 687 580
rect 721 546 737 580
rect 671 493 737 546
rect 671 459 687 493
rect 721 459 737 493
rect 671 454 737 459
rect 771 580 837 596
rect 771 546 787 580
rect 821 546 837 580
rect 771 497 837 546
rect 771 463 787 497
rect 821 463 837 497
rect 559 406 575 440
rect 609 424 625 440
rect 609 406 653 424
rect 559 390 653 406
rect 223 378 289 390
rect 23 344 289 378
rect 405 340 471 356
rect 25 294 91 310
rect 25 260 41 294
rect 75 260 91 294
rect 25 236 91 260
rect 169 294 263 310
rect 169 260 185 294
rect 219 260 263 294
rect 30 195 96 202
rect 30 161 46 195
rect 80 161 96 195
rect 30 120 96 161
rect 30 86 46 120
rect 80 86 96 120
rect 169 88 263 260
rect 297 294 363 310
rect 297 260 313 294
rect 347 260 363 294
rect 405 306 421 340
rect 455 306 471 340
rect 405 290 471 306
rect 505 340 585 356
rect 505 306 535 340
rect 569 306 585 340
rect 505 290 585 306
rect 619 310 653 390
rect 771 414 837 463
rect 771 380 787 414
rect 821 380 837 414
rect 771 364 837 380
rect 871 580 937 649
rect 871 546 887 580
rect 921 546 937 580
rect 871 497 937 546
rect 871 463 887 497
rect 921 463 937 497
rect 871 414 937 463
rect 871 380 887 414
rect 921 380 937 414
rect 871 364 937 380
rect 619 294 769 310
rect 297 88 363 260
rect 619 260 651 294
rect 685 260 719 294
rect 753 260 769 294
rect 619 256 769 260
rect 446 222 769 256
rect 446 210 512 222
rect 446 176 462 210
rect 496 176 512 210
rect 803 188 837 364
rect 446 120 512 176
rect 30 17 96 86
rect 446 86 462 120
rect 496 86 512 120
rect 446 70 512 86
rect 558 154 574 188
rect 608 154 624 188
rect 558 120 624 154
rect 558 86 574 120
rect 608 86 624 120
rect 558 17 624 86
rect 677 154 693 188
rect 727 154 837 188
rect 677 116 743 154
rect 677 82 693 116
rect 727 82 743 116
rect 677 70 743 82
rect 777 86 793 120
rect 827 86 887 120
rect 921 86 937 120
rect 777 17 937 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a41o_2
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 319 94 353 128 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 319 168 353 202 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 319 242 353 276 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 223 94 257 128 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 223 168 257 202 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 223 242 257 276 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 A4
port 4 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 B1
port 5 nsew
flabel corelocali s 703 94 737 128 0 FreeSans 340 0 0 0 X
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 960 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3768320
string GDS_START 3759576
<< end >>
