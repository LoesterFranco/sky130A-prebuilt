magic
tech sky130A
magscale 1 2
timestamp 1604502710
<< nwell >>
rect -38 332 710 704
<< pwell >>
rect 0 0 672 49
<< scpmos >>
rect 82 392 118 592
rect 284 368 320 592
rect 374 368 410 592
rect 464 368 500 592
rect 554 368 590 592
<< nmoslvt >>
rect 151 94 181 222
rect 272 74 302 222
rect 368 74 398 222
rect 458 74 488 222
rect 554 74 584 222
<< ndiff >>
rect 94 210 151 222
rect 94 176 106 210
rect 140 176 151 210
rect 94 140 151 176
rect 94 106 106 140
rect 140 106 151 140
rect 94 94 151 106
rect 181 192 272 222
rect 181 158 213 192
rect 247 158 272 192
rect 181 124 272 158
rect 181 94 213 124
rect 201 90 213 94
rect 247 90 272 124
rect 201 74 272 90
rect 302 192 368 222
rect 302 158 313 192
rect 347 158 368 192
rect 302 120 368 158
rect 302 86 313 120
rect 347 86 368 120
rect 302 74 368 86
rect 398 142 458 222
rect 398 108 413 142
rect 447 108 458 142
rect 398 74 458 108
rect 488 210 554 222
rect 488 176 499 210
rect 533 176 554 210
rect 488 120 554 176
rect 488 86 499 120
rect 533 86 554 120
rect 488 74 554 86
rect 584 152 645 222
rect 584 118 599 152
rect 633 118 645 152
rect 584 74 645 118
<< pdiff >>
rect 27 580 82 592
rect 27 546 38 580
rect 72 546 82 580
rect 27 509 82 546
rect 27 475 38 509
rect 72 475 82 509
rect 27 438 82 475
rect 27 404 38 438
rect 72 404 82 438
rect 27 392 82 404
rect 118 580 174 592
rect 118 546 128 580
rect 162 546 174 580
rect 118 512 174 546
rect 118 478 128 512
rect 162 478 174 512
rect 118 444 174 478
rect 118 410 128 444
rect 162 410 174 444
rect 118 392 174 410
rect 228 580 284 592
rect 228 546 240 580
rect 274 546 284 580
rect 228 497 284 546
rect 228 463 240 497
rect 274 463 284 497
rect 228 414 284 463
rect 228 380 240 414
rect 274 380 284 414
rect 228 368 284 380
rect 320 531 374 592
rect 320 497 330 531
rect 364 497 374 531
rect 320 414 374 497
rect 320 380 330 414
rect 364 380 374 414
rect 320 368 374 380
rect 410 580 464 592
rect 410 546 420 580
rect 454 546 464 580
rect 410 504 464 546
rect 410 470 420 504
rect 454 470 464 504
rect 410 424 464 470
rect 410 390 420 424
rect 454 390 464 424
rect 410 368 464 390
rect 500 580 554 592
rect 500 546 510 580
rect 544 546 554 580
rect 500 508 554 546
rect 500 474 510 508
rect 544 474 554 508
rect 500 368 554 474
rect 590 580 645 592
rect 590 546 600 580
rect 634 546 645 580
rect 590 497 645 546
rect 590 463 600 497
rect 634 463 645 497
rect 590 414 645 463
rect 590 380 600 414
rect 634 380 645 414
rect 590 368 645 380
<< ndiffc >>
rect 106 176 140 210
rect 106 106 140 140
rect 213 158 247 192
rect 213 90 247 124
rect 313 158 347 192
rect 313 86 347 120
rect 413 108 447 142
rect 499 176 533 210
rect 499 86 533 120
rect 599 118 633 152
<< pdiffc >>
rect 38 546 72 580
rect 38 475 72 509
rect 38 404 72 438
rect 128 546 162 580
rect 128 478 162 512
rect 128 410 162 444
rect 240 546 274 580
rect 240 463 274 497
rect 240 380 274 414
rect 330 497 364 531
rect 330 380 364 414
rect 420 546 454 580
rect 420 470 454 504
rect 420 390 454 424
rect 510 546 544 580
rect 510 474 544 508
rect 600 546 634 580
rect 600 463 634 497
rect 600 380 634 414
<< poly >>
rect 82 592 118 618
rect 284 592 320 618
rect 374 592 410 618
rect 464 592 500 618
rect 554 592 590 618
rect 82 360 118 392
rect 82 344 181 360
rect 284 352 320 368
rect 82 310 122 344
rect 156 310 181 344
rect 272 322 320 352
rect 374 322 410 368
rect 464 336 500 368
rect 554 336 590 368
rect 272 310 410 322
rect 82 294 181 310
rect 151 222 181 294
rect 229 294 410 310
rect 229 260 245 294
rect 279 260 410 294
rect 229 244 410 260
rect 458 320 590 336
rect 458 286 474 320
rect 508 300 590 320
rect 508 286 584 300
rect 458 270 584 286
rect 272 222 302 244
rect 368 222 398 244
rect 458 222 488 270
rect 554 222 584 270
rect 151 68 181 94
rect 272 48 302 74
rect 368 48 398 74
rect 458 48 488 74
rect 554 48 584 74
<< polycont >>
rect 122 310 156 344
rect 245 260 279 294
rect 474 286 508 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 22 580 72 596
rect 22 546 38 580
rect 22 509 72 546
rect 22 475 38 509
rect 22 438 72 475
rect 22 404 38 438
rect 22 260 72 404
rect 112 580 178 649
rect 112 546 128 580
rect 162 546 178 580
rect 112 512 178 546
rect 112 478 128 512
rect 162 478 178 512
rect 112 444 178 478
rect 112 410 128 444
rect 162 410 178 444
rect 112 394 178 410
rect 224 581 470 615
rect 224 580 290 581
rect 224 546 240 580
rect 274 546 290 580
rect 404 580 470 581
rect 224 497 290 546
rect 224 463 240 497
rect 274 463 290 497
rect 224 414 290 463
rect 224 380 240 414
rect 274 380 290 414
rect 224 364 290 380
rect 329 531 364 547
rect 329 497 330 531
rect 329 414 364 497
rect 329 380 330 414
rect 404 546 420 580
rect 454 546 470 580
rect 404 504 470 546
rect 404 470 420 504
rect 454 470 470 504
rect 404 424 470 470
rect 510 580 560 649
rect 544 546 560 580
rect 510 508 560 546
rect 544 474 560 508
rect 510 458 560 474
rect 600 580 650 596
rect 634 546 650 580
rect 600 497 650 546
rect 634 463 650 497
rect 600 424 650 463
rect 404 390 420 424
rect 454 414 650 424
rect 454 390 600 414
rect 106 344 172 360
rect 106 310 122 344
rect 156 310 172 344
rect 106 294 172 310
rect 229 294 295 310
rect 229 260 245 294
rect 279 260 295 294
rect 22 226 295 260
rect 329 236 364 380
rect 634 380 650 414
rect 600 364 650 380
rect 409 320 551 356
rect 409 286 474 320
rect 508 286 551 320
rect 409 270 551 286
rect 601 236 647 282
rect 22 210 156 226
rect 22 176 106 210
rect 140 176 156 210
rect 329 210 647 236
rect 329 192 499 210
rect 22 140 156 176
rect 22 106 106 140
rect 140 106 156 140
rect 22 90 156 106
rect 197 158 213 192
rect 247 158 263 192
rect 197 124 263 158
rect 197 90 213 124
rect 247 90 263 124
rect 197 17 263 90
rect 297 158 313 192
rect 347 158 363 192
rect 533 202 647 210
rect 533 176 549 202
rect 297 120 363 158
rect 297 86 313 120
rect 347 86 363 120
rect 297 70 363 86
rect 397 142 463 158
rect 397 108 413 142
rect 447 108 463 142
rect 397 17 463 108
rect 499 120 549 176
rect 533 86 549 120
rect 499 70 549 86
rect 583 152 649 168
rect 583 118 599 152
rect 633 118 649 152
rect 583 17 649 118
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
rlabel comment s 0 0 0 0 4 nor2b_2
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 B_N
port 2 nsew
flabel corelocali s 607 242 641 276 0 FreeSans 340 0 0 0 Y
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 672 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1482390
string GDS_START 1476142
<< end >>
