magic
tech sky130A
magscale 1 2
timestamp 1599588244
<< locali >>
rect 87 260 167 356
rect 201 236 267 302
rect 469 404 535 596
rect 669 424 735 596
rect 955 424 1021 596
rect 1155 424 1221 596
rect 669 404 1221 424
rect 469 390 1221 404
rect 469 370 839 390
rect 1155 370 1221 390
rect 469 364 535 370
rect 793 252 839 370
rect 889 270 1077 356
rect 1273 336 1319 356
rect 1125 270 1319 336
rect 537 218 839 252
rect 537 168 571 218
rect 469 134 571 168
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 19 482 89 572
rect 130 516 196 649
rect 369 516 435 649
rect 19 448 435 482
rect 19 390 89 448
rect 19 206 53 390
rect 237 364 335 414
rect 301 236 335 364
rect 369 270 435 448
rect 569 438 635 649
rect 769 458 921 649
rect 1055 458 1121 649
rect 1255 390 1321 649
rect 625 320 759 336
rect 469 286 759 320
rect 469 236 503 286
rect 19 70 92 206
rect 301 202 503 236
rect 126 17 192 202
rect 226 70 335 202
rect 882 202 1320 236
rect 369 100 435 168
rect 605 150 836 184
rect 605 100 639 150
rect 882 124 948 202
rect 369 66 639 100
rect 673 85 739 116
rect 982 85 1048 163
rect 673 51 1048 85
rect 1084 70 1134 202
rect 1168 17 1234 163
rect 1270 70 1320 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
<< metal1 >>
rect 0 683 1344 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 0 617 1344 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 1344 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
rect 0 -49 1344 -17
<< labels >>
rlabel locali s 87 260 167 356 6 A_N
port 1 nsew signal input
rlabel locali s 201 236 267 302 6 B_N
port 2 nsew signal input
rlabel locali s 889 270 1077 356 6 C
port 3 nsew signal input
rlabel locali s 1273 336 1319 356 6 D
port 4 nsew signal input
rlabel locali s 1125 270 1319 336 6 D
port 4 nsew signal input
rlabel locali s 1155 424 1221 596 6 Y
port 5 nsew signal output
rlabel locali s 1155 370 1221 390 6 Y
port 5 nsew signal output
rlabel locali s 955 424 1021 596 6 Y
port 5 nsew signal output
rlabel locali s 793 252 839 370 6 Y
port 5 nsew signal output
rlabel locali s 669 424 735 596 6 Y
port 5 nsew signal output
rlabel locali s 669 404 1221 424 6 Y
port 5 nsew signal output
rlabel locali s 537 218 839 252 6 Y
port 5 nsew signal output
rlabel locali s 537 168 571 218 6 Y
port 5 nsew signal output
rlabel locali s 469 404 535 596 6 Y
port 5 nsew signal output
rlabel locali s 469 390 1221 404 6 Y
port 5 nsew signal output
rlabel locali s 469 370 839 390 6 Y
port 5 nsew signal output
rlabel locali s 469 364 535 370 6 Y
port 5 nsew signal output
rlabel locali s 469 134 571 168 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -49 1344 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 7 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 617 1344 715 6 VPWR
port 9 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1344 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1456894
string GDS_START 1446598
<< end >>
