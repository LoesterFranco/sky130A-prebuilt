magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 18 337 71 491
rect 18 53 85 337
rect 203 199 339 265
rect 373 199 478 265
rect 518 199 615 265
rect 661 199 717 265
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 105 383 181 527
rect 219 419 271 491
rect 305 453 417 527
rect 461 419 513 491
rect 219 373 513 419
rect 641 337 709 491
rect 121 301 709 337
rect 121 163 169 301
rect 121 125 707 163
rect 131 17 280 91
rect 439 53 504 125
rect 540 17 616 91
rect 662 53 707 125
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel locali s 373 199 478 265 6 A1
port 1 nsew signal input
rlabel locali s 203 199 339 265 6 A2
port 2 nsew signal input
rlabel locali s 518 199 615 265 6 B1
port 3 nsew signal input
rlabel locali s 661 199 717 265 6 C1
port 4 nsew signal input
rlabel locali s 18 337 71 491 6 X
port 5 nsew signal output
rlabel locali s 18 53 85 337 6 X
port 5 nsew signal output
rlabel metal1 s 0 -48 736 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 736 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1083298
string GDS_START 1076632
<< end >>
