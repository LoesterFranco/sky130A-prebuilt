magic
tech sky130A
magscale 1 2
timestamp 1601050088
<< locali >>
rect 23 424 73 596
rect 219 424 253 547
rect 383 424 449 547
rect 583 424 649 479
rect 783 424 849 479
rect 23 390 849 424
rect 23 364 73 390
rect 107 270 377 356
rect 505 336 647 356
rect 445 270 647 336
rect 697 310 849 390
rect 23 236 73 237
rect 783 236 817 310
rect 1416 236 1895 308
rect 23 202 817 236
rect 23 81 73 202
rect 211 119 245 202
rect 384 187 817 202
rect 384 119 450 187
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 113 581 1312 615
rect 113 458 179 581
rect 293 458 343 581
rect 483 513 1026 547
rect 1060 546 1312 581
rect 1346 546 1412 649
rect 483 458 549 513
rect 683 458 749 513
rect 992 512 1026 513
rect 1446 512 1512 596
rect 1546 546 1612 649
rect 1646 512 1712 596
rect 992 478 1712 512
rect 1752 444 1802 649
rect 895 410 1802 444
rect 895 368 1216 410
rect 1837 376 1891 540
rect 1927 410 1993 649
rect 1334 342 1965 376
rect 1334 334 1368 342
rect 1030 268 1368 334
rect 109 85 175 168
rect 851 200 1343 234
rect 1931 202 1965 342
rect 281 85 347 168
rect 851 153 885 200
rect 1277 184 1343 200
rect 1481 168 1765 202
rect 484 119 885 153
rect 919 150 1105 166
rect 1481 150 1547 168
rect 919 132 1547 150
rect 919 85 953 132
rect 1071 116 1547 132
rect 109 51 953 85
rect 987 17 1037 98
rect 1175 17 1241 82
rect 1379 17 1445 82
rect 1481 78 1547 116
rect 1581 17 1665 128
rect 1699 78 1765 168
rect 1799 17 1865 202
rect 1899 78 1965 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
rlabel locali s 505 336 647 356 6 A0
port 1 nsew signal input
rlabel locali s 445 270 647 336 6 A0
port 1 nsew signal input
rlabel locali s 107 270 377 356 6 A1
port 2 nsew signal input
rlabel locali s 1416 236 1895 308 6 S
port 3 nsew signal input
rlabel locali s 783 424 849 479 6 Y
port 4 nsew signal output
rlabel locali s 783 236 817 310 6 Y
port 4 nsew signal output
rlabel locali s 697 310 849 390 6 Y
port 4 nsew signal output
rlabel locali s 583 424 649 479 6 Y
port 4 nsew signal output
rlabel locali s 384 187 817 202 6 Y
port 4 nsew signal output
rlabel locali s 384 119 450 187 6 Y
port 4 nsew signal output
rlabel locali s 383 424 449 547 6 Y
port 4 nsew signal output
rlabel locali s 219 424 253 547 6 Y
port 4 nsew signal output
rlabel locali s 211 119 245 202 6 Y
port 4 nsew signal output
rlabel locali s 23 424 73 596 6 Y
port 4 nsew signal output
rlabel locali s 23 390 849 424 6 Y
port 4 nsew signal output
rlabel locali s 23 364 73 390 6 Y
port 4 nsew signal output
rlabel locali s 23 236 73 237 6 Y
port 4 nsew signal output
rlabel locali s 23 202 817 236 6 Y
port 4 nsew signal output
rlabel locali s 23 81 73 202 6 Y
port 4 nsew signal output
rlabel metal1 s 0 -49 2016 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 617 2016 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2016 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1951968
string GDS_START 1938184
<< end >>
