magic
tech sky130A
magscale 1 2
timestamp 1599588238
<< locali >>
rect 17 423 89 596
rect 17 389 569 423
rect 17 364 89 389
rect 870 368 1162 402
rect 17 202 51 364
rect 85 236 263 310
rect 307 286 647 355
rect 697 286 935 368
rect 17 85 90 202
rect 1096 270 1162 368
rect 516 85 582 116
rect 17 51 582 85
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 123 491 189 596
rect 615 593 694 649
rect 337 559 479 591
rect 842 570 911 649
rect 337 536 705 559
rect 952 536 1018 596
rect 337 525 1018 536
rect 671 502 1018 525
rect 123 468 637 491
rect 123 457 801 468
rect 603 402 801 457
rect 952 436 1018 502
rect 1052 436 1118 649
rect 1159 436 1230 572
rect 348 218 806 252
rect 128 153 194 202
rect 348 187 414 218
rect 730 200 806 218
rect 982 236 1048 334
rect 1196 236 1230 436
rect 982 202 1230 236
rect 448 166 650 184
rect 448 153 1023 166
rect 128 150 1023 153
rect 128 119 482 150
rect 616 132 1023 150
rect 947 100 1023 132
rect 628 17 694 98
rect 842 17 911 98
rect 1057 17 1123 168
rect 1159 114 1230 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
<< metal1 >>
rect 0 683 1248 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 0 617 1248 649
rect 0 17 1248 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
rect 0 -49 1248 -17
<< labels >>
rlabel locali s 85 236 263 310 6 A0
port 1 nsew signal input
rlabel locali s 307 286 647 355 6 A1
port 2 nsew signal input
rlabel locali s 1096 270 1162 368 6 S
port 3 nsew signal input
rlabel locali s 870 368 1162 402 6 S
port 3 nsew signal input
rlabel locali s 697 286 935 368 6 S
port 3 nsew signal input
rlabel locali s 516 85 582 116 6 Y
port 4 nsew signal output
rlabel locali s 17 423 89 596 6 Y
port 4 nsew signal output
rlabel locali s 17 389 569 423 6 Y
port 4 nsew signal output
rlabel locali s 17 364 89 389 6 Y
port 4 nsew signal output
rlabel locali s 17 202 51 364 6 Y
port 4 nsew signal output
rlabel locali s 17 85 90 202 6 Y
port 4 nsew signal output
rlabel locali s 17 51 582 85 6 Y
port 4 nsew signal output
rlabel metal1 s 0 -49 1248 49 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1248 715 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1248 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1615916
string GDS_START 1606070
<< end >>
