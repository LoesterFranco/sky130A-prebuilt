magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 806 704
<< pwell >>
rect 0 0 768 49
<< scnmos >>
rect 115 112 145 222
rect 222 74 252 222
rect 308 74 338 222
rect 471 74 501 222
rect 557 74 587 222
rect 651 74 681 222
<< pmoshvt >>
rect 87 368 117 536
rect 190 368 220 592
rect 280 368 310 592
rect 474 392 504 592
rect 564 392 594 592
rect 654 392 684 592
<< ndiff >>
rect 62 172 115 222
rect 62 138 70 172
rect 104 138 115 172
rect 62 112 115 138
rect 145 118 222 222
rect 145 112 177 118
rect 165 84 177 112
rect 211 84 222 118
rect 165 74 222 84
rect 252 127 308 222
rect 252 93 263 127
rect 297 93 308 127
rect 252 74 308 93
rect 338 134 471 222
rect 338 100 349 134
rect 383 100 426 134
rect 460 100 471 134
rect 338 74 471 100
rect 501 202 557 222
rect 501 168 512 202
rect 546 168 557 202
rect 501 120 557 168
rect 501 86 512 120
rect 546 86 557 120
rect 501 74 557 86
rect 587 74 651 222
rect 681 202 738 222
rect 681 168 692 202
rect 726 168 738 202
rect 681 120 738 168
rect 681 86 692 120
rect 726 86 738 120
rect 681 74 738 86
<< pdiff >>
rect 135 566 190 592
rect 135 536 143 566
rect 32 524 87 536
rect 32 490 40 524
rect 74 490 87 524
rect 32 414 87 490
rect 32 380 40 414
rect 74 380 87 414
rect 32 368 87 380
rect 117 532 143 536
rect 177 532 190 566
rect 117 368 190 532
rect 220 414 280 592
rect 220 380 233 414
rect 267 380 280 414
rect 220 368 280 380
rect 310 566 365 592
rect 310 532 323 566
rect 357 532 365 566
rect 310 368 365 532
rect 419 580 474 592
rect 419 546 427 580
rect 461 546 474 580
rect 419 462 474 546
rect 419 428 427 462
rect 461 428 474 462
rect 419 392 474 428
rect 504 580 564 592
rect 504 546 517 580
rect 551 546 564 580
rect 504 470 564 546
rect 504 436 517 470
rect 551 436 564 470
rect 504 392 564 436
rect 594 559 654 592
rect 594 525 607 559
rect 641 525 654 559
rect 594 392 654 525
rect 684 580 739 592
rect 684 546 697 580
rect 731 546 739 580
rect 684 510 739 546
rect 684 476 697 510
rect 731 476 739 510
rect 684 440 739 476
rect 684 406 697 440
rect 731 406 739 440
rect 684 392 739 406
<< ndiffc >>
rect 70 138 104 172
rect 177 84 211 118
rect 263 93 297 127
rect 349 100 383 134
rect 426 100 460 134
rect 512 168 546 202
rect 512 86 546 120
rect 692 168 726 202
rect 692 86 726 120
<< pdiffc >>
rect 40 490 74 524
rect 40 380 74 414
rect 143 532 177 566
rect 233 380 267 414
rect 323 532 357 566
rect 427 546 461 580
rect 427 428 461 462
rect 517 546 551 580
rect 517 436 551 470
rect 607 525 641 559
rect 697 546 731 580
rect 697 476 731 510
rect 697 406 731 440
<< poly >>
rect 190 592 220 618
rect 280 592 310 618
rect 474 592 504 618
rect 564 592 594 618
rect 654 592 684 618
rect 87 536 117 562
rect 474 377 504 392
rect 564 377 594 392
rect 654 377 684 392
rect 87 353 117 368
rect 190 353 220 368
rect 280 353 310 368
rect 84 310 120 353
rect 36 294 145 310
rect 36 260 52 294
rect 86 260 145 294
rect 36 244 145 260
rect 187 274 223 353
rect 277 310 313 353
rect 471 346 507 377
rect 471 318 501 346
rect 561 318 597 377
rect 651 356 687 377
rect 651 340 747 356
rect 272 294 338 310
rect 272 274 288 294
rect 187 260 288 274
rect 322 260 338 294
rect 187 244 338 260
rect 380 302 501 318
rect 380 268 396 302
rect 430 268 501 302
rect 380 252 501 268
rect 543 302 609 318
rect 543 268 559 302
rect 593 268 609 302
rect 543 252 609 268
rect 651 306 697 340
rect 731 306 747 340
rect 651 290 747 306
rect 115 222 145 244
rect 222 222 252 244
rect 308 222 338 244
rect 471 222 501 252
rect 557 222 587 252
rect 651 222 681 290
rect 115 86 145 112
rect 222 48 252 74
rect 308 48 338 74
rect 471 48 501 74
rect 557 48 587 74
rect 651 48 681 74
<< polycont >>
rect 52 260 86 294
rect 288 260 322 294
rect 396 268 430 302
rect 559 268 593 302
rect 697 306 731 340
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 127 566 193 649
rect 24 524 90 540
rect 24 490 40 524
rect 74 490 90 524
rect 127 532 143 566
rect 177 532 193 566
rect 127 516 193 532
rect 307 566 373 649
rect 307 532 323 566
rect 357 532 373 566
rect 307 516 373 532
rect 411 580 483 596
rect 411 546 427 580
rect 461 546 483 580
rect 24 482 90 490
rect 24 448 362 482
rect 24 414 90 448
rect 24 380 40 414
rect 74 380 90 414
rect 24 364 90 380
rect 25 294 102 310
rect 25 260 52 294
rect 86 260 102 294
rect 25 236 102 260
rect 136 202 170 448
rect 54 172 170 202
rect 54 138 70 172
rect 104 168 170 172
rect 204 380 233 414
rect 267 380 283 414
rect 204 364 283 380
rect 321 378 362 448
rect 411 462 483 546
rect 411 428 427 462
rect 461 428 483 462
rect 411 412 483 428
rect 517 580 551 596
rect 517 470 551 546
rect 591 559 641 649
rect 591 525 607 559
rect 591 488 641 525
rect 681 580 747 596
rect 681 546 697 580
rect 731 546 747 580
rect 681 510 747 546
rect 681 476 697 510
rect 731 476 747 510
rect 681 454 747 476
rect 551 440 747 454
rect 551 436 697 440
rect 517 420 697 436
rect 449 386 483 412
rect 681 406 697 420
rect 731 406 747 440
rect 681 390 747 406
rect 204 208 238 364
rect 321 344 415 378
rect 449 352 511 386
rect 381 318 415 344
rect 272 294 347 310
rect 272 260 288 294
rect 322 260 347 294
rect 272 244 347 260
rect 381 302 443 318
rect 381 268 396 302
rect 430 268 443 302
rect 381 252 443 268
rect 313 218 347 244
rect 477 218 511 352
rect 545 302 647 356
rect 545 268 559 302
rect 593 268 647 302
rect 681 340 747 356
rect 681 306 697 340
rect 731 306 747 340
rect 681 290 747 306
rect 545 252 647 268
rect 204 168 279 208
rect 313 202 562 218
rect 313 184 512 202
rect 104 138 120 168
rect 54 108 120 138
rect 245 150 279 168
rect 496 168 512 184
rect 546 168 562 202
rect 161 118 211 134
rect 161 84 177 118
rect 161 17 211 84
rect 245 127 313 150
rect 245 93 263 127
rect 297 93 313 127
rect 245 70 313 93
rect 347 134 462 150
rect 347 100 349 134
rect 383 100 426 134
rect 460 100 462 134
rect 347 17 462 100
rect 496 120 562 168
rect 496 86 512 120
rect 546 86 562 120
rect 496 70 562 86
rect 676 202 742 218
rect 676 168 692 202
rect 726 168 742 202
rect 676 120 742 168
rect 676 86 692 120
rect 726 86 742 120
rect 676 17 742 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a21bo_2
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 B1_N
port 3 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 223 168 257 202 0 FreeSans 340 0 0 0 X
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 768 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 4049678
string GDS_START 4042950
<< end >>
