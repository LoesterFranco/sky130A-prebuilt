magic
tech sky130A
magscale 1 2
timestamp 1604502693
<< nwell >>
rect -38 261 1694 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 415 47 445 177
rect 499 47 529 177
rect 583 47 613 177
rect 667 47 697 177
rect 855 47 885 177
rect 939 47 969 177
rect 1023 47 1053 177
rect 1107 47 1137 177
rect 1191 47 1221 177
rect 1275 47 1305 177
rect 1359 47 1389 177
rect 1454 47 1484 177
rect 1547 47 1577 177
<< pmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 415 297 445 497
rect 499 297 529 497
rect 583 297 613 497
rect 667 297 697 497
rect 855 297 885 497
rect 939 297 969 497
rect 1023 297 1053 497
rect 1107 297 1137 497
rect 1191 297 1221 497
rect 1275 297 1305 497
rect 1359 297 1389 497
rect 1454 297 1484 497
rect 1547 297 1577 497
<< ndiff >>
rect 27 97 79 177
rect 27 63 35 97
rect 69 63 79 97
rect 27 47 79 63
rect 109 165 163 177
rect 109 131 119 165
rect 153 131 163 165
rect 109 47 163 131
rect 193 97 247 177
rect 193 63 203 97
rect 237 63 247 97
rect 193 47 247 63
rect 277 165 331 177
rect 277 131 287 165
rect 321 131 331 165
rect 277 47 331 131
rect 361 97 415 177
rect 361 63 371 97
rect 405 63 415 97
rect 361 47 415 63
rect 445 165 499 177
rect 445 131 455 165
rect 489 131 499 165
rect 445 47 499 131
rect 529 97 583 177
rect 529 63 539 97
rect 573 63 583 97
rect 529 47 583 63
rect 613 165 667 177
rect 613 131 623 165
rect 657 131 667 165
rect 613 47 667 131
rect 697 97 749 177
rect 697 63 707 97
rect 741 63 749 97
rect 697 47 749 63
rect 803 93 855 177
rect 803 59 811 93
rect 845 59 855 93
rect 803 47 855 59
rect 885 101 939 177
rect 885 67 895 101
rect 929 67 939 101
rect 885 47 939 67
rect 969 93 1023 177
rect 969 59 979 93
rect 1013 59 1023 93
rect 969 47 1023 59
rect 1053 101 1107 177
rect 1053 67 1063 101
rect 1097 67 1107 101
rect 1053 47 1107 67
rect 1137 102 1191 177
rect 1137 68 1147 102
rect 1181 68 1191 102
rect 1137 47 1191 68
rect 1221 101 1275 177
rect 1221 67 1231 101
rect 1265 67 1275 101
rect 1221 47 1275 67
rect 1305 93 1359 177
rect 1305 59 1315 93
rect 1349 59 1359 93
rect 1305 47 1359 59
rect 1389 152 1454 177
rect 1389 118 1399 152
rect 1433 118 1454 152
rect 1389 47 1454 118
rect 1484 93 1547 177
rect 1484 59 1503 93
rect 1537 59 1547 93
rect 1484 47 1547 59
rect 1577 101 1629 177
rect 1577 67 1587 101
rect 1621 67 1629 101
rect 1577 47 1629 67
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 297 79 451
rect 109 349 163 497
rect 109 315 119 349
rect 153 315 163 349
rect 109 297 163 315
rect 193 485 247 497
rect 193 451 203 485
rect 237 451 247 485
rect 193 297 247 451
rect 277 349 331 497
rect 277 315 287 349
rect 321 315 331 349
rect 277 297 331 315
rect 361 485 415 497
rect 361 451 371 485
rect 405 451 415 485
rect 361 297 415 451
rect 445 417 499 497
rect 445 383 455 417
rect 489 383 499 417
rect 445 297 499 383
rect 529 485 583 497
rect 529 451 539 485
rect 573 451 583 485
rect 529 297 583 451
rect 613 417 667 497
rect 613 383 623 417
rect 657 383 667 417
rect 613 297 667 383
rect 697 485 749 497
rect 697 451 707 485
rect 741 451 749 485
rect 697 297 749 451
rect 803 485 855 497
rect 803 451 811 485
rect 845 451 855 485
rect 803 297 855 451
rect 885 349 939 497
rect 885 315 895 349
rect 929 315 939 349
rect 885 297 939 315
rect 969 485 1023 497
rect 969 451 979 485
rect 1013 451 1023 485
rect 969 297 1023 451
rect 1053 349 1107 497
rect 1053 315 1063 349
rect 1097 315 1107 349
rect 1053 297 1107 315
rect 1137 485 1191 497
rect 1137 451 1147 485
rect 1181 451 1191 485
rect 1137 297 1191 451
rect 1221 477 1275 497
rect 1221 443 1231 477
rect 1265 443 1275 477
rect 1221 409 1275 443
rect 1221 375 1231 409
rect 1265 375 1275 409
rect 1221 297 1275 375
rect 1305 485 1359 497
rect 1305 451 1315 485
rect 1349 451 1359 485
rect 1305 297 1359 451
rect 1389 477 1454 497
rect 1389 443 1399 477
rect 1433 443 1454 477
rect 1389 409 1454 443
rect 1389 375 1399 409
rect 1433 375 1454 409
rect 1389 297 1454 375
rect 1484 485 1547 497
rect 1484 451 1503 485
rect 1537 451 1547 485
rect 1484 297 1547 451
rect 1577 477 1629 497
rect 1577 443 1587 477
rect 1621 443 1629 477
rect 1577 409 1629 443
rect 1577 375 1587 409
rect 1621 375 1629 409
rect 1577 297 1629 375
<< ndiffc >>
rect 35 63 69 97
rect 119 131 153 165
rect 203 63 237 97
rect 287 131 321 165
rect 371 63 405 97
rect 455 131 489 165
rect 539 63 573 97
rect 623 131 657 165
rect 707 63 741 97
rect 811 59 845 93
rect 895 67 929 101
rect 979 59 1013 93
rect 1063 67 1097 101
rect 1147 68 1181 102
rect 1231 67 1265 101
rect 1315 59 1349 93
rect 1399 118 1433 152
rect 1503 59 1537 93
rect 1587 67 1621 101
<< pdiffc >>
rect 35 451 69 485
rect 119 315 153 349
rect 203 451 237 485
rect 287 315 321 349
rect 371 451 405 485
rect 455 383 489 417
rect 539 451 573 485
rect 623 383 657 417
rect 707 451 741 485
rect 811 451 845 485
rect 895 315 929 349
rect 979 451 1013 485
rect 1063 315 1097 349
rect 1147 451 1181 485
rect 1231 443 1265 477
rect 1231 375 1265 409
rect 1315 451 1349 485
rect 1399 443 1433 477
rect 1399 375 1433 409
rect 1503 451 1537 485
rect 1587 443 1621 477
rect 1587 375 1621 409
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 415 497 445 523
rect 499 497 529 523
rect 583 497 613 523
rect 667 497 697 523
rect 855 497 885 523
rect 939 497 969 523
rect 1023 497 1053 523
rect 1107 497 1137 523
rect 1191 497 1221 523
rect 1275 497 1305 523
rect 1359 497 1389 523
rect 1454 497 1484 523
rect 1547 497 1577 523
rect 79 265 109 297
rect 163 265 193 297
rect 247 265 277 297
rect 331 265 361 297
rect 79 249 361 265
rect 79 215 112 249
rect 146 215 180 249
rect 214 215 361 249
rect 79 199 361 215
rect 79 177 109 199
rect 163 177 193 199
rect 247 177 277 199
rect 331 177 361 199
rect 415 265 445 297
rect 499 265 529 297
rect 583 265 613 297
rect 667 265 697 297
rect 855 265 885 297
rect 939 265 969 297
rect 1023 265 1053 297
rect 1107 265 1137 297
rect 415 249 697 265
rect 415 215 431 249
rect 465 215 499 249
rect 533 215 567 249
rect 601 215 635 249
rect 669 215 697 249
rect 415 199 697 215
rect 798 249 1137 265
rect 798 215 815 249
rect 849 215 883 249
rect 917 215 951 249
rect 985 215 1019 249
rect 1053 215 1087 249
rect 1121 215 1137 249
rect 798 199 1137 215
rect 415 177 445 199
rect 499 177 529 199
rect 583 177 613 199
rect 667 177 697 199
rect 855 177 885 199
rect 939 177 969 199
rect 1023 177 1053 199
rect 1107 177 1137 199
rect 1191 265 1221 297
rect 1275 265 1305 297
rect 1359 265 1389 297
rect 1454 265 1484 297
rect 1547 265 1577 297
rect 1191 249 1484 265
rect 1191 215 1362 249
rect 1396 215 1434 249
rect 1468 215 1484 249
rect 1191 199 1484 215
rect 1526 249 1580 265
rect 1526 215 1536 249
rect 1570 215 1580 249
rect 1526 199 1580 215
rect 1191 177 1221 199
rect 1275 177 1305 199
rect 1359 177 1389 199
rect 1454 177 1484 199
rect 1547 177 1577 199
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 415 21 445 47
rect 499 21 529 47
rect 583 21 613 47
rect 667 21 697 47
rect 855 21 885 47
rect 939 21 969 47
rect 1023 21 1053 47
rect 1107 21 1137 47
rect 1191 21 1221 47
rect 1275 21 1305 47
rect 1359 21 1389 47
rect 1454 21 1484 47
rect 1547 21 1577 47
<< polycont >>
rect 112 215 146 249
rect 180 215 214 249
rect 431 215 465 249
rect 499 215 533 249
rect 567 215 601 249
rect 635 215 669 249
rect 815 215 849 249
rect 883 215 917 249
rect 951 215 985 249
rect 1019 215 1053 249
rect 1087 215 1121 249
rect 1362 215 1396 249
rect 1434 215 1468 249
rect 1536 215 1570 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 795 485 861 527
rect 19 451 35 485
rect 69 451 203 485
rect 237 451 371 485
rect 405 451 539 485
rect 573 451 707 485
rect 741 451 757 485
rect 795 451 811 485
rect 845 451 861 485
rect 963 485 1029 527
rect 963 451 979 485
rect 1013 451 1029 485
rect 1131 485 1197 527
rect 1131 451 1147 485
rect 1181 451 1197 485
rect 1231 477 1265 493
rect 19 97 64 451
rect 1299 485 1365 527
rect 1299 451 1315 485
rect 1349 451 1365 485
rect 1399 477 1433 493
rect 1231 417 1265 443
rect 1487 485 1553 527
rect 1487 451 1503 485
rect 1537 451 1553 485
rect 1587 477 1639 493
rect 1399 417 1433 443
rect 439 383 455 417
rect 489 383 623 417
rect 657 409 1433 417
rect 657 383 1231 409
rect 1265 383 1399 409
rect 1231 359 1265 375
rect 1399 359 1433 375
rect 1621 443 1639 477
rect 1587 409 1639 443
rect 1621 375 1639 409
rect 1587 359 1639 375
rect 103 315 119 349
rect 153 315 287 349
rect 321 315 895 349
rect 929 315 1063 349
rect 1097 315 1116 349
rect 1152 285 1570 319
rect 112 249 248 265
rect 146 215 180 249
rect 214 221 248 249
rect 391 249 710 265
rect 1152 258 1186 285
rect 112 199 214 215
rect 391 215 431 249
rect 465 215 499 249
rect 533 215 567 249
rect 601 215 635 249
rect 669 215 710 249
rect 769 249 1186 258
rect 1536 249 1570 285
rect 769 215 815 249
rect 849 215 883 249
rect 917 215 951 249
rect 985 215 1019 249
rect 1053 215 1087 249
rect 1121 215 1186 249
rect 1346 215 1362 249
rect 1396 215 1434 249
rect 391 199 710 215
rect 271 165 306 187
rect 103 131 119 165
rect 153 131 287 165
rect 321 131 340 153
rect 439 131 455 165
rect 489 131 623 165
rect 657 131 1097 165
rect 895 101 929 131
rect 19 63 35 97
rect 69 63 203 97
rect 237 63 371 97
rect 405 63 539 97
rect 573 63 707 97
rect 741 63 757 97
rect 795 59 811 93
rect 845 59 861 93
rect 795 17 861 59
rect 1063 101 1097 131
rect 1264 181 1290 187
rect 1264 153 1433 181
rect 1230 152 1433 153
rect 1230 143 1399 152
rect 895 51 929 67
rect 963 59 979 93
rect 1013 59 1029 93
rect 963 17 1029 59
rect 1063 51 1097 67
rect 1131 102 1196 118
rect 1131 68 1147 102
rect 1181 68 1196 102
rect 1131 17 1196 68
rect 1230 101 1265 143
rect 1468 165 1502 249
rect 1536 199 1570 215
rect 1604 165 1639 359
rect 1468 131 1639 165
rect 1230 67 1231 101
rect 1230 51 1265 67
rect 1309 93 1359 109
rect 1399 102 1433 118
rect 1587 101 1639 131
rect 1309 59 1315 93
rect 1349 59 1359 93
rect 1309 17 1359 59
rect 1487 59 1503 93
rect 1537 59 1553 93
rect 1487 17 1553 59
rect 1621 67 1639 101
rect 1587 51 1639 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 306 165 340 187
rect 306 153 321 165
rect 321 153 340 165
rect 1230 153 1264 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
<< metal1 >>
rect 0 561 1656 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 0 496 1656 527
rect 294 187 352 193
rect 294 153 306 187
rect 340 184 352 187
rect 1218 187 1276 193
rect 1218 184 1230 187
rect 340 156 1230 184
rect 340 153 352 156
rect 294 147 352 153
rect 1218 153 1230 156
rect 1264 153 1276 187
rect 1218 147 1276 153
rect 0 17 1656 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
rect 0 -48 1656 -17
<< labels >>
flabel corelocali s 1046 221 1080 255 0 FreeSans 200 0 0 0 S
port 3 nsew
flabel corelocali s 954 221 988 255 0 FreeSans 200 0 0 0 S
port 3 nsew
flabel corelocali s 862 221 896 255 0 FreeSans 200 0 0 0 S
port 3 nsew
flabel corelocali s 770 221 804 255 0 FreeSans 200 0 0 0 S
port 3 nsew
flabel corelocali s 582 221 616 255 0 FreeSans 200 0 0 0 A1
port 2 nsew
flabel corelocali s 490 221 524 255 0 FreeSans 200 0 0 0 A1
port 2 nsew
flabel corelocali s 398 221 432 255 0 FreeSans 200 0 0 0 A1
port 2 nsew
flabel corelocali s 1138 221 1172 255 0 FreeSans 200 0 0 0 S
port 3 nsew
flabel corelocali s 214 221 248 255 0 FreeSans 200 0 0 0 A0
port 1 nsew
flabel corelocali s 122 221 156 255 0 FreeSans 200 0 0 0 A0
port 1 nsew
flabel corelocali s 30 425 64 459 0 FreeSans 200 0 0 0 Y
port 8 nsew
flabel corelocali s 30 153 64 187 0 FreeSans 200 0 0 0 Y
port 8 nsew
flabel corelocali s 30 289 64 323 0 FreeSans 200 0 0 0 Y
port 8 nsew
flabel corelocali s 30 357 64 391 0 FreeSans 200 0 0 0 Y
port 8 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 200 0 0 0 Y
port 8 nsew
flabel corelocali s 674 221 708 255 0 FreeSans 200 0 0 0 A1
port 2 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
rlabel comment s 0 0 0 0 4 mux2i_4
<< properties >>
string FIXED_BBOX 0 0 1656 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1734198
string GDS_START 1722056
string path 0.000 0.000 41.400 0.000 
<< end >>
