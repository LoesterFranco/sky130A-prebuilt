magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 111 486 167 591
rect 111 420 265 486
rect 85 356 151 386
rect 25 236 151 356
rect 85 184 151 236
rect 217 136 265 420
rect 123 70 265 136
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 288 683
rect 21 420 71 649
rect 201 520 267 649
rect 23 17 89 150
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 288 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
<< metal1 >>
rect 0 683 288 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 288 683
rect 0 617 288 649
rect 0 17 288 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 288 17
rect 0 -49 288 -17
<< labels >>
rlabel locali s 85 356 151 386 6 A
port 1 nsew signal input
rlabel locali s 85 184 151 236 6 A
port 1 nsew signal input
rlabel locali s 25 236 151 356 6 A
port 1 nsew signal input
rlabel locali s 217 136 265 420 6 Y
port 2 nsew signal output
rlabel locali s 123 70 265 136 6 Y
port 2 nsew signal output
rlabel locali s 111 486 167 591 6 Y
port 2 nsew signal output
rlabel locali s 111 420 265 486 6 Y
port 2 nsew signal output
rlabel metal1 s 0 -49 288 49 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 617 288 715 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 288 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3354728
string GDS_START 3350728
<< end >>
