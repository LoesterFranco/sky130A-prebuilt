magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 2630 704
<< pwell >>
rect 0 0 2592 49
<< scnmos >>
rect 85 74 115 222
rect 267 94 297 222
rect 492 74 522 202
rect 578 74 608 202
rect 714 119 744 247
rect 846 119 876 247
rect 1057 81 1087 229
rect 1203 81 1233 209
rect 1289 81 1319 209
rect 1602 81 1632 209
rect 1702 81 1732 209
rect 1879 116 1909 264
rect 1974 136 2004 264
rect 2163 136 2193 264
rect 2278 120 2308 248
rect 2478 100 2508 248
<< pmoshvt >>
rect 88 368 118 592
rect 226 368 256 568
rect 495 418 525 586
rect 593 418 623 586
rect 700 379 730 547
rect 843 379 873 547
rect 1054 368 1084 592
rect 1167 368 1197 568
rect 1284 400 1314 568
rect 1565 400 1595 568
rect 1683 368 1713 568
rect 1824 368 1854 592
rect 2026 384 2056 552
rect 2116 384 2146 552
rect 2340 368 2370 568
rect 2476 368 2506 592
<< ndiff >>
rect 28 210 85 222
rect 28 176 40 210
rect 74 176 85 210
rect 28 120 85 176
rect 28 86 40 120
rect 74 86 85 120
rect 28 74 85 86
rect 115 152 267 222
rect 115 118 140 152
rect 174 118 267 152
rect 115 94 267 118
rect 297 180 354 222
rect 657 237 714 247
rect 657 203 669 237
rect 703 203 714 237
rect 657 202 714 203
rect 297 146 308 180
rect 342 146 354 180
rect 297 94 354 146
rect 439 173 492 202
rect 439 139 447 173
rect 481 139 492 173
rect 115 74 186 94
rect 439 74 492 139
rect 522 127 578 202
rect 522 93 533 127
rect 567 93 578 127
rect 522 74 578 93
rect 608 169 714 202
rect 608 135 669 169
rect 703 135 714 169
rect 608 119 714 135
rect 744 197 846 247
rect 744 163 755 197
rect 789 163 846 197
rect 744 119 846 163
rect 876 201 937 247
rect 876 167 891 201
rect 925 167 937 201
rect 876 119 937 167
rect 608 74 658 119
rect 997 202 1057 229
rect 997 168 1009 202
rect 1043 168 1057 202
rect 997 134 1057 168
rect 997 100 1009 134
rect 1043 100 1057 134
rect 997 81 1057 100
rect 1087 209 1137 229
rect 1829 209 1879 264
rect 1087 127 1203 209
rect 1087 93 1126 127
rect 1160 93 1203 127
rect 1087 81 1203 93
rect 1233 197 1289 209
rect 1233 163 1244 197
rect 1278 163 1289 197
rect 1233 127 1289 163
rect 1233 93 1244 127
rect 1278 93 1289 127
rect 1233 81 1289 93
rect 1319 197 1602 209
rect 1319 163 1344 197
rect 1378 163 1415 197
rect 1449 163 1486 197
rect 1520 163 1557 197
rect 1591 163 1602 197
rect 1319 129 1602 163
rect 1319 95 1344 129
rect 1378 95 1415 129
rect 1449 95 1486 129
rect 1520 95 1557 129
rect 1591 95 1602 129
rect 1319 81 1602 95
rect 1632 197 1702 209
rect 1632 163 1657 197
rect 1691 163 1702 197
rect 1632 127 1702 163
rect 1632 93 1657 127
rect 1691 93 1702 127
rect 1632 81 1702 93
rect 1732 195 1879 209
rect 1732 161 1758 195
rect 1792 161 1879 195
rect 1732 127 1879 161
rect 1732 93 1758 127
rect 1792 116 1879 127
rect 1909 252 1974 264
rect 1909 218 1927 252
rect 1961 218 1974 252
rect 1909 182 1974 218
rect 1909 148 1927 182
rect 1961 148 1974 182
rect 1909 136 1974 148
rect 2004 250 2163 264
rect 2004 216 2030 250
rect 2064 216 2118 250
rect 2152 216 2163 250
rect 2004 182 2163 216
rect 2004 148 2030 182
rect 2064 148 2118 182
rect 2152 148 2163 182
rect 2004 136 2163 148
rect 2193 248 2243 264
rect 2193 240 2278 248
rect 2193 206 2233 240
rect 2267 206 2278 240
rect 2193 166 2278 206
rect 2193 136 2233 166
rect 1909 116 1959 136
rect 1792 93 1805 116
rect 1732 81 1805 93
rect 2221 132 2233 136
rect 2267 132 2278 166
rect 2221 120 2278 132
rect 2308 146 2478 248
rect 2308 120 2402 146
rect 2373 112 2402 120
rect 2436 112 2478 146
rect 2373 100 2478 112
rect 2508 236 2565 248
rect 2508 202 2519 236
rect 2553 202 2565 236
rect 2508 149 2565 202
rect 2508 115 2519 149
rect 2553 115 2565 149
rect 2508 100 2565 115
<< pdiff >>
rect 29 580 88 592
rect 29 546 41 580
rect 75 546 88 580
rect 29 497 88 546
rect 29 463 41 497
rect 75 463 88 497
rect 29 414 88 463
rect 29 380 41 414
rect 75 380 88 414
rect 29 368 88 380
rect 118 580 177 592
rect 118 546 131 580
rect 165 568 177 580
rect 165 546 226 568
rect 118 510 226 546
rect 118 476 131 510
rect 165 476 226 510
rect 118 440 226 476
rect 118 406 131 440
rect 165 406 226 440
rect 118 368 226 406
rect 256 531 315 568
rect 256 497 269 531
rect 303 497 315 531
rect 256 414 315 497
rect 430 473 495 586
rect 430 439 447 473
rect 481 439 495 473
rect 430 418 495 439
rect 525 547 593 586
rect 525 513 546 547
rect 580 513 593 547
rect 525 462 593 513
rect 525 428 546 462
rect 580 428 593 462
rect 525 418 593 428
rect 623 547 676 586
rect 623 531 700 547
rect 623 497 653 531
rect 687 497 700 531
rect 623 425 700 497
rect 623 418 653 425
rect 256 380 269 414
rect 303 380 315 414
rect 256 368 315 380
rect 641 391 653 418
rect 687 391 700 425
rect 641 379 700 391
rect 730 503 843 547
rect 730 469 753 503
rect 787 469 843 503
rect 730 379 843 469
rect 873 531 935 547
rect 873 497 889 531
rect 923 497 935 531
rect 873 425 935 497
rect 873 391 889 425
rect 923 391 935 425
rect 873 379 935 391
rect 995 428 1054 592
rect 995 394 1007 428
rect 1041 394 1054 428
rect 995 368 1054 394
rect 1084 580 1149 592
rect 1084 546 1100 580
rect 1134 568 1149 580
rect 2164 598 2227 610
rect 1765 580 1824 592
rect 1765 568 1777 580
rect 1134 546 1167 568
rect 1084 368 1167 546
rect 1197 428 1284 568
rect 1197 394 1210 428
rect 1244 400 1284 428
rect 1314 517 1565 568
rect 1314 483 1367 517
rect 1401 483 1483 517
rect 1517 483 1565 517
rect 1314 400 1565 483
rect 1595 531 1683 568
rect 1595 497 1625 531
rect 1659 497 1683 531
rect 1595 414 1683 497
rect 1595 400 1625 414
rect 1244 394 1256 400
rect 1197 368 1256 394
rect 1613 380 1625 400
rect 1659 380 1683 414
rect 1613 368 1683 380
rect 1713 546 1777 568
rect 1811 546 1824 580
rect 1713 449 1824 546
rect 1713 415 1777 449
rect 1811 415 1824 449
rect 1713 368 1824 415
rect 1854 580 1913 592
rect 1854 546 1867 580
rect 1901 546 1913 580
rect 2164 564 2178 598
rect 2212 564 2227 598
rect 2417 580 2476 592
rect 2417 568 2429 580
rect 2164 552 2227 564
rect 1854 508 1913 546
rect 1854 474 1867 508
rect 1901 474 1913 508
rect 1854 433 1913 474
rect 1854 399 1867 433
rect 1901 399 1913 433
rect 1854 368 1913 399
rect 1967 531 2026 552
rect 1967 497 1979 531
rect 2013 497 2026 531
rect 1967 430 2026 497
rect 1967 396 1979 430
rect 2013 396 2026 430
rect 1967 384 2026 396
rect 2056 430 2116 552
rect 2056 396 2069 430
rect 2103 396 2116 430
rect 2056 384 2116 396
rect 2146 384 2227 552
rect 2281 531 2340 568
rect 2281 497 2293 531
rect 2327 497 2340 531
rect 2281 420 2340 497
rect 2281 386 2293 420
rect 2327 386 2340 420
rect 2281 368 2340 386
rect 2370 546 2429 568
rect 2463 546 2476 580
rect 2370 500 2476 546
rect 2370 466 2429 500
rect 2463 466 2476 500
rect 2370 420 2476 466
rect 2370 386 2429 420
rect 2463 386 2476 420
rect 2370 368 2476 386
rect 2506 580 2565 592
rect 2506 546 2519 580
rect 2553 546 2565 580
rect 2506 497 2565 546
rect 2506 463 2519 497
rect 2553 463 2565 497
rect 2506 414 2565 463
rect 2506 380 2519 414
rect 2553 380 2565 414
rect 2506 368 2565 380
<< ndiffc >>
rect 40 176 74 210
rect 40 86 74 120
rect 140 118 174 152
rect 669 203 703 237
rect 308 146 342 180
rect 447 139 481 173
rect 533 93 567 127
rect 669 135 703 169
rect 755 163 789 197
rect 891 167 925 201
rect 1009 168 1043 202
rect 1009 100 1043 134
rect 1126 93 1160 127
rect 1244 163 1278 197
rect 1244 93 1278 127
rect 1344 163 1378 197
rect 1415 163 1449 197
rect 1486 163 1520 197
rect 1557 163 1591 197
rect 1344 95 1378 129
rect 1415 95 1449 129
rect 1486 95 1520 129
rect 1557 95 1591 129
rect 1657 163 1691 197
rect 1657 93 1691 127
rect 1758 161 1792 195
rect 1758 93 1792 127
rect 1927 218 1961 252
rect 1927 148 1961 182
rect 2030 216 2064 250
rect 2118 216 2152 250
rect 2030 148 2064 182
rect 2118 148 2152 182
rect 2233 206 2267 240
rect 2233 132 2267 166
rect 2402 112 2436 146
rect 2519 202 2553 236
rect 2519 115 2553 149
<< pdiffc >>
rect 41 546 75 580
rect 41 463 75 497
rect 41 380 75 414
rect 131 546 165 580
rect 131 476 165 510
rect 131 406 165 440
rect 269 497 303 531
rect 447 439 481 473
rect 546 513 580 547
rect 546 428 580 462
rect 653 497 687 531
rect 269 380 303 414
rect 653 391 687 425
rect 753 469 787 503
rect 889 497 923 531
rect 889 391 923 425
rect 1007 394 1041 428
rect 1100 546 1134 580
rect 1210 394 1244 428
rect 1367 483 1401 517
rect 1483 483 1517 517
rect 1625 497 1659 531
rect 1625 380 1659 414
rect 1777 546 1811 580
rect 1777 415 1811 449
rect 1867 546 1901 580
rect 2178 564 2212 598
rect 1867 474 1901 508
rect 1867 399 1901 433
rect 1979 497 2013 531
rect 1979 396 2013 430
rect 2069 396 2103 430
rect 2293 497 2327 531
rect 2293 386 2327 420
rect 2429 546 2463 580
rect 2429 466 2463 500
rect 2429 386 2463 420
rect 2519 546 2553 580
rect 2519 463 2553 497
rect 2519 380 2553 414
<< poly >>
rect 88 592 118 618
rect 590 615 980 645
rect 226 568 256 594
rect 495 586 525 612
rect 590 601 626 615
rect 593 586 623 601
rect 700 547 730 573
rect 840 562 876 615
rect 843 547 873 562
rect 495 403 525 418
rect 88 353 118 368
rect 226 353 256 368
rect 85 336 121 353
rect 85 320 175 336
rect 85 286 125 320
rect 159 286 175 320
rect 85 270 175 286
rect 223 326 259 353
rect 492 333 528 403
rect 593 392 623 418
rect 700 364 730 379
rect 697 342 733 364
rect 843 353 873 379
rect 697 333 798 342
rect 492 326 798 333
rect 223 310 297 326
rect 223 276 239 310
rect 273 276 297 310
rect 85 222 115 270
rect 223 260 297 276
rect 267 222 297 260
rect 492 292 748 326
rect 782 292 798 326
rect 492 276 798 292
rect 950 317 980 615
rect 1054 592 1084 618
rect 1167 568 1197 594
rect 1284 568 1314 594
rect 1565 568 1595 594
rect 1683 568 1713 594
rect 1824 592 1854 618
rect 1284 385 1314 400
rect 1565 385 1595 400
rect 1281 368 1317 385
rect 1562 375 1598 385
rect 1054 353 1084 368
rect 1167 353 1197 368
rect 1051 317 1087 353
rect 1164 317 1200 353
rect 1281 352 1354 368
rect 1281 318 1304 352
rect 1338 318 1354 352
rect 950 301 1087 317
rect 950 287 991 301
rect 492 202 522 276
rect 714 247 744 276
rect 846 247 876 273
rect 952 267 991 287
rect 1025 267 1087 301
rect 952 251 1087 267
rect 1135 301 1233 317
rect 1281 302 1354 318
rect 1441 352 1598 375
rect 2026 552 2056 578
rect 2116 552 2146 578
rect 2340 568 2370 594
rect 2476 592 2506 618
rect 2026 369 2056 384
rect 2116 369 2146 384
rect 1683 353 1713 368
rect 1824 353 1854 368
rect 1441 318 1457 352
rect 1491 345 1598 352
rect 1491 318 1507 345
rect 1135 267 1151 301
rect 1185 267 1233 301
rect 1135 251 1233 267
rect 1441 284 1507 318
rect 1680 309 1716 353
rect 1821 309 1857 353
rect 2023 309 2059 369
rect 1441 254 1457 284
rect 578 202 608 228
rect 85 48 115 74
rect 267 68 297 94
rect 714 93 744 119
rect 492 48 522 74
rect 578 51 608 74
rect 846 51 876 119
rect 952 51 982 251
rect 1057 229 1087 251
rect 1203 209 1233 251
rect 1289 250 1457 254
rect 1491 250 1507 284
rect 1289 224 1507 250
rect 1549 281 1632 297
rect 1549 247 1565 281
rect 1599 247 1632 281
rect 1549 231 1632 247
rect 1680 281 1909 309
rect 1680 247 1757 281
rect 1791 279 1909 281
rect 1791 247 1807 279
rect 1879 264 1909 279
rect 1974 279 2059 309
rect 2113 352 2149 369
rect 2340 353 2370 368
rect 2476 353 2506 368
rect 2113 336 2203 352
rect 2337 336 2373 353
rect 2473 336 2509 353
rect 2113 302 2153 336
rect 2187 302 2203 336
rect 2113 286 2203 302
rect 2278 320 2373 336
rect 2278 286 2323 320
rect 2357 286 2373 320
rect 1974 264 2004 279
rect 2163 264 2193 286
rect 2278 270 2373 286
rect 2424 320 2509 336
rect 2424 286 2440 320
rect 2474 286 2509 320
rect 2424 270 2509 286
rect 1680 231 1807 247
rect 1289 209 1319 224
rect 1602 209 1632 231
rect 1702 209 1732 231
rect 2278 248 2308 270
rect 2478 248 2508 270
rect 1879 90 1909 116
rect 1974 114 2004 136
rect 1974 98 2115 114
rect 2163 110 2193 136
rect 1057 55 1087 81
rect 1203 55 1233 81
rect 1289 55 1319 81
rect 1602 55 1632 81
rect 1702 55 1732 81
rect 1974 64 1997 98
rect 2031 64 2065 98
rect 2099 64 2115 98
rect 2278 94 2308 120
rect 2478 74 2508 100
rect 578 21 982 51
rect 1974 48 2115 64
<< polycont >>
rect 125 286 159 320
rect 239 276 273 310
rect 748 292 782 326
rect 1304 318 1338 352
rect 991 267 1025 301
rect 1457 318 1491 352
rect 1151 267 1185 301
rect 1457 250 1491 284
rect 1565 247 1599 281
rect 1757 247 1791 281
rect 2153 302 2187 336
rect 2323 286 2357 320
rect 2440 286 2474 320
rect 1997 64 2031 98
rect 2065 64 2099 98
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2592 683
rect 24 580 75 596
rect 24 546 41 580
rect 24 497 75 546
rect 24 463 41 497
rect 24 414 75 463
rect 24 380 41 414
rect 115 580 165 649
rect 115 546 131 580
rect 115 510 165 546
rect 115 476 131 510
rect 115 440 165 476
rect 115 406 131 440
rect 115 390 165 406
rect 201 581 787 615
rect 24 236 75 380
rect 109 320 167 356
rect 109 286 125 320
rect 159 286 167 320
rect 109 270 167 286
rect 201 326 235 581
rect 269 531 546 547
rect 303 513 546 531
rect 580 513 596 547
rect 303 497 367 513
rect 269 414 367 497
rect 303 380 367 414
rect 269 364 367 380
rect 409 473 497 479
rect 409 439 447 473
rect 481 439 497 473
rect 409 424 497 439
rect 409 390 415 424
rect 449 414 497 424
rect 531 462 596 513
rect 531 428 546 462
rect 580 428 596 462
rect 449 390 483 414
rect 531 409 596 428
rect 409 378 483 390
rect 201 310 289 326
rect 201 276 239 310
rect 273 276 289 310
rect 201 260 289 276
rect 201 236 258 260
rect 24 210 258 236
rect 24 176 40 210
rect 74 202 258 210
rect 323 204 367 364
rect 74 176 90 202
rect 24 120 90 176
rect 24 86 40 120
rect 74 86 90 120
rect 24 70 90 86
rect 124 152 190 168
rect 124 118 140 152
rect 174 118 190 152
rect 124 17 190 118
rect 224 85 258 202
rect 295 180 367 204
rect 295 146 308 180
rect 342 146 367 180
rect 295 123 367 146
rect 433 173 483 378
rect 562 218 596 409
rect 637 531 703 547
rect 637 497 653 531
rect 687 497 703 531
rect 637 425 703 497
rect 737 503 787 581
rect 737 469 753 503
rect 737 450 787 469
rect 821 581 1009 615
rect 637 391 653 425
rect 687 410 703 425
rect 821 410 855 581
rect 687 391 855 410
rect 637 376 855 391
rect 889 531 941 547
rect 923 497 941 531
rect 889 425 941 497
rect 975 512 1009 581
rect 1081 580 1153 649
rect 1081 546 1100 580
rect 1134 546 1153 580
rect 1230 581 1743 615
rect 1230 512 1330 581
rect 975 478 1330 512
rect 923 424 941 425
rect 889 390 895 391
rect 929 390 941 424
rect 637 375 703 376
rect 889 375 941 390
rect 669 237 703 375
rect 737 326 798 342
rect 737 292 748 326
rect 782 310 798 326
rect 782 292 857 310
rect 737 276 857 292
rect 562 184 635 218
rect 433 139 447 173
rect 481 139 483 173
rect 433 123 483 139
rect 517 127 567 150
rect 517 93 533 127
rect 517 85 567 93
rect 224 51 567 85
rect 601 85 635 184
rect 669 169 703 203
rect 669 119 703 135
rect 739 197 789 225
rect 739 163 755 197
rect 739 85 789 163
rect 601 51 789 85
rect 823 85 857 276
rect 891 201 941 375
rect 991 428 1057 444
rect 991 394 1007 428
rect 1041 398 1057 428
rect 1194 428 1262 444
rect 1041 394 1160 398
rect 991 364 1160 394
rect 1194 394 1210 428
rect 1244 394 1262 428
rect 1194 364 1262 394
rect 1126 317 1160 364
rect 975 301 1041 317
rect 975 267 991 301
rect 1025 267 1041 301
rect 975 236 1041 267
rect 1126 301 1194 317
rect 1126 267 1151 301
rect 1185 267 1194 301
rect 1126 251 1194 267
rect 1126 202 1160 251
rect 925 167 941 201
rect 891 134 941 167
rect 993 168 1009 202
rect 1043 168 1160 202
rect 1228 213 1262 364
rect 1296 368 1330 478
rect 1364 517 1523 533
rect 1364 483 1367 517
rect 1401 483 1483 517
rect 1517 483 1523 517
rect 1364 467 1523 483
rect 1296 352 1346 368
rect 1296 318 1304 352
rect 1338 318 1346 352
rect 1296 302 1346 318
rect 1380 262 1414 467
rect 1228 197 1294 213
rect 993 134 1059 168
rect 993 100 1009 134
rect 1043 100 1059 134
rect 1228 163 1244 197
rect 1278 163 1294 197
rect 1228 127 1294 163
rect 993 85 1059 100
rect 823 51 1059 85
rect 1093 93 1126 127
rect 1160 93 1194 127
rect 1093 17 1194 93
rect 1228 93 1244 127
rect 1278 93 1294 127
rect 1228 77 1294 93
rect 1328 197 1414 262
rect 1448 424 1511 430
rect 1448 390 1471 424
rect 1505 390 1511 424
rect 1448 352 1511 390
rect 1448 318 1457 352
rect 1491 318 1511 352
rect 1448 284 1511 318
rect 1557 297 1591 581
rect 1625 531 1675 547
rect 1659 497 1675 531
rect 1625 414 1675 497
rect 1659 380 1675 414
rect 1625 364 1675 380
rect 1448 250 1457 284
rect 1491 250 1511 284
rect 1448 234 1511 250
rect 1549 281 1607 297
rect 1549 247 1565 281
rect 1599 247 1607 281
rect 1549 231 1607 247
rect 1641 213 1675 364
rect 1709 365 1743 581
rect 1777 580 1811 649
rect 1777 449 1811 546
rect 1777 399 1811 415
rect 1851 598 2395 615
rect 1851 581 2178 598
rect 1851 580 1945 581
rect 1851 546 1867 580
rect 1901 546 1945 580
rect 2160 564 2178 581
rect 2212 581 2395 598
rect 2212 564 2231 581
rect 2160 548 2231 564
rect 1851 508 1945 546
rect 1851 474 1867 508
rect 1901 474 1945 508
rect 1851 433 1945 474
rect 1851 399 1867 433
rect 1901 399 1945 433
rect 1709 331 1877 365
rect 1741 281 1807 297
rect 1741 247 1757 281
rect 1791 247 1807 281
rect 1741 231 1807 247
rect 1641 197 1707 213
rect 1328 163 1344 197
rect 1378 163 1415 197
rect 1449 163 1486 197
rect 1520 163 1557 197
rect 1591 163 1607 197
rect 1328 129 1607 163
rect 1328 95 1344 129
rect 1378 95 1415 129
rect 1449 95 1486 129
rect 1520 95 1557 129
rect 1591 95 1607 129
rect 1328 88 1607 95
rect 1641 163 1657 197
rect 1691 163 1707 197
rect 1641 127 1707 163
rect 1641 93 1657 127
rect 1691 93 1707 127
rect 1641 77 1707 93
rect 1741 195 1809 197
rect 1741 161 1758 195
rect 1792 161 1809 195
rect 1741 127 1809 161
rect 1741 93 1758 127
rect 1792 93 1809 127
rect 1741 17 1809 93
rect 1843 114 1877 331
rect 1911 268 1945 399
rect 1979 531 2013 547
rect 2277 531 2327 547
rect 2277 514 2293 531
rect 2013 497 2293 514
rect 1979 480 2327 497
rect 1979 430 2013 480
rect 1979 380 2013 396
rect 2053 430 2103 446
rect 2053 396 2069 430
rect 1911 252 1977 268
rect 2053 252 2103 396
rect 2137 424 2203 430
rect 2137 390 2143 424
rect 2177 390 2203 424
rect 2137 336 2203 390
rect 2137 302 2153 336
rect 2187 302 2203 336
rect 2137 286 2203 302
rect 2239 420 2327 480
rect 2239 386 2293 420
rect 2239 370 2327 386
rect 1911 218 1927 252
rect 1961 218 1977 252
rect 1911 182 1977 218
rect 1911 148 1927 182
rect 1961 148 1977 182
rect 2014 250 2183 252
rect 2239 250 2273 370
rect 2361 336 2395 581
rect 2429 580 2479 649
rect 2463 546 2479 580
rect 2429 500 2479 546
rect 2463 466 2479 500
rect 2429 420 2479 466
rect 2463 386 2479 420
rect 2429 370 2479 386
rect 2519 580 2569 596
rect 2553 546 2569 580
rect 2519 497 2569 546
rect 2553 463 2569 497
rect 2519 414 2569 463
rect 2553 380 2569 414
rect 2307 320 2395 336
rect 2307 286 2323 320
rect 2357 286 2395 320
rect 2307 270 2395 286
rect 2429 320 2485 336
rect 2429 286 2440 320
rect 2474 286 2485 320
rect 2014 216 2030 250
rect 2064 216 2118 250
rect 2152 216 2183 250
rect 2014 182 2183 216
rect 2014 148 2030 182
rect 2064 148 2118 182
rect 2152 148 2183 182
rect 1843 98 2115 114
rect 1843 64 1997 98
rect 2031 64 2065 98
rect 2099 64 2115 98
rect 2149 98 2183 148
rect 2217 244 2273 250
rect 2217 240 2283 244
rect 2217 206 2233 240
rect 2267 206 2283 240
rect 2429 236 2485 286
rect 2217 166 2283 206
rect 2217 132 2233 166
rect 2267 132 2283 166
rect 2317 202 2485 236
rect 2519 236 2569 380
rect 2553 202 2569 236
rect 2317 98 2351 202
rect 2519 168 2569 202
rect 2149 64 2351 98
rect 2385 146 2469 162
rect 2385 112 2402 146
rect 2436 112 2469 146
rect 1843 51 2115 64
rect 2385 17 2469 112
rect 2503 149 2569 168
rect 2503 115 2519 149
rect 2553 115 2569 149
rect 2503 88 2569 115
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2592 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 415 390 449 424
rect 895 391 923 424
rect 923 391 929 424
rect 895 390 929 391
rect 1471 390 1505 424
rect 2143 390 2177 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
<< metal1 >>
rect 0 683 2592 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2592 683
rect 0 617 2592 649
rect 403 424 461 430
rect 403 390 415 424
rect 449 421 461 424
rect 883 424 941 430
rect 883 421 895 424
rect 449 393 895 421
rect 449 390 461 393
rect 403 384 461 390
rect 883 390 895 393
rect 929 421 941 424
rect 1459 424 1517 430
rect 1459 421 1471 424
rect 929 393 1471 421
rect 929 390 941 393
rect 883 384 941 390
rect 1459 390 1471 393
rect 1505 421 1517 424
rect 2131 424 2189 430
rect 2131 421 2143 424
rect 1505 393 2143 421
rect 1505 390 1517 393
rect 1459 384 1517 390
rect 2131 390 2143 393
rect 2177 390 2189 424
rect 2131 384 2189 390
rect 0 17 2592 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2592 17
rect 0 -49 2592 -17
<< labels >>
rlabel comment s 0 0 0 0 4 fahcin_1
flabel pwell s 0 0 2592 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 2592 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 2592 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 2592 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 1471 94 1505 128 0 FreeSans 340 0 0 0 COUT
port 8 nsew
flabel corelocali s 1567 94 1601 128 0 FreeSans 340 0 0 0 COUT
port 8 nsew
flabel corelocali s 991 242 1025 276 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 1759 242 1793 276 0 FreeSans 340 0 0 0 CIN
port 3 nsew
flabel corelocali s 2527 94 2561 128 0 FreeSans 340 0 0 0 SUM
port 9 nsew
flabel corelocali s 2527 168 2561 202 0 FreeSans 340 0 0 0 SUM
port 9 nsew
flabel corelocali s 2527 242 2561 276 0 FreeSans 340 0 0 0 SUM
port 9 nsew
flabel corelocali s 2527 316 2561 350 0 FreeSans 340 0 0 0 SUM
port 9 nsew
flabel corelocali s 2527 390 2561 424 0 FreeSans 340 0 0 0 SUM
port 9 nsew
flabel corelocali s 2527 464 2561 498 0 FreeSans 340 0 0 0 SUM
port 9 nsew
flabel corelocali s 2527 538 2561 572 0 FreeSans 340 0 0 0 SUM
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 2592 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2313866
string GDS_START 2294912
<< end >>
