magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 368 561
rect 105 371 171 493
rect 212 394 249 487
rect 283 428 350 493
rect 212 350 345 394
rect 85 149 157 248
rect 277 165 345 350
rect 208 131 345 165
rect 111 17 166 113
rect 208 51 249 131
rect 283 17 350 97
rect 0 -17 368 17
<< obsli1 >>
rect 17 316 71 487
rect 17 282 243 316
rect 17 117 51 282
rect 193 199 243 282
rect 17 51 69 117
<< metal1 >>
rect 0 496 368 592
rect 14 428 354 468
rect 110 416 168 428
rect 287 416 345 428
rect 0 -48 368 48
<< labels >>
rlabel locali s 85 149 157 248 6 A
port 1 nsew signal input
rlabel locali s 277 165 345 350 6 X
port 2 nsew signal output
rlabel locali s 212 394 249 487 6 X
port 2 nsew signal output
rlabel locali s 212 350 345 394 6 X
port 2 nsew signal output
rlabel locali s 208 131 345 165 6 X
port 2 nsew signal output
rlabel locali s 208 51 249 131 6 X
port 2 nsew signal output
rlabel locali s 105 371 171 493 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 283 428 350 493 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 287 416 345 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 110 416 168 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 14 428 354 468 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 283 17 350 97 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 111 17 166 113 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 368 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 368 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 527 368 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 368 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 368 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2194750
string GDS_START 2189962
<< end >>
