magic
tech sky130A
magscale 1 2
timestamp 1599588232
<< locali >>
rect 85 224 163 358
rect 197 88 263 361
rect 305 88 371 358
rect 409 270 479 356
rect 582 364 655 596
rect 621 226 655 364
rect 546 70 655 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 23 463 89 649
rect 123 429 189 596
rect 223 463 341 649
rect 375 429 441 596
rect 482 460 548 649
rect 17 426 441 429
rect 17 395 548 426
rect 17 190 51 395
rect 375 392 548 395
rect 17 71 154 190
rect 514 330 548 392
rect 514 264 587 330
rect 444 17 510 206
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel locali s 85 224 163 358 6 A
port 1 nsew signal input
rlabel locali s 197 88 263 361 6 B
port 2 nsew signal input
rlabel locali s 305 88 371 358 6 C
port 3 nsew signal input
rlabel locali s 409 270 479 356 6 D
port 4 nsew signal input
rlabel locali s 621 226 655 364 6 X
port 5 nsew signal output
rlabel locali s 582 364 655 596 6 X
port 5 nsew signal output
rlabel locali s 546 70 655 226 6 X
port 5 nsew signal output
rlabel metal1 s 0 -49 672 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 7 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 617 672 715 6 VPWR
port 9 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3250218
string GDS_START 3242920
<< end >>
