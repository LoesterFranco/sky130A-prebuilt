magic
tech sky130A
magscale 1 2
timestamp 1601050056
<< nwell >>
rect -38 332 2150 704
<< pwell >>
rect 0 0 2112 49
<< scpmos >>
rect 83 392 119 592
rect 183 392 219 592
rect 290 392 326 560
rect 397 392 433 520
rect 516 418 552 546
rect 623 379 659 547
rect 951 368 987 592
rect 1185 388 1221 556
rect 1321 388 1357 556
rect 1526 410 1562 538
rect 1707 368 1743 592
rect 1797 368 1833 592
rect 1903 368 1939 592
rect 1993 368 2029 592
<< nmoslvt >>
rect 84 118 114 246
rect 218 118 248 246
rect 386 118 416 246
rect 486 162 516 246
rect 606 118 636 246
rect 724 125 754 253
rect 959 74 989 222
rect 1203 123 1233 251
rect 1339 123 1369 251
rect 1625 74 1655 158
rect 1741 74 1771 222
rect 1827 74 1857 222
rect 1913 74 1943 222
rect 1999 74 2029 222
<< ndiff >>
rect 651 246 724 253
rect 27 234 84 246
rect 27 200 39 234
rect 73 200 84 234
rect 27 164 84 200
rect 27 130 39 164
rect 73 130 84 164
rect 27 118 84 130
rect 114 118 218 246
rect 248 234 386 246
rect 248 200 291 234
rect 325 200 386 234
rect 248 118 386 200
rect 416 234 486 246
rect 416 200 427 234
rect 461 200 486 234
rect 416 164 486 200
rect 416 130 427 164
rect 461 162 486 164
rect 516 221 606 246
rect 516 187 527 221
rect 561 187 606 221
rect 516 162 606 187
rect 461 130 471 162
rect 416 118 471 130
rect 556 118 606 162
rect 636 241 724 246
rect 636 207 663 241
rect 697 207 724 241
rect 636 164 724 207
rect 636 130 663 164
rect 697 130 724 164
rect 636 125 724 130
rect 754 237 843 253
rect 754 203 799 237
rect 833 203 843 237
rect 754 125 843 203
rect 636 118 709 125
rect 129 82 203 118
rect 129 48 149 82
rect 183 48 203 82
rect 129 36 203 48
rect 903 189 959 222
rect 903 155 914 189
rect 948 155 959 189
rect 903 74 959 155
rect 989 106 1094 222
rect 1148 171 1203 251
rect 1148 137 1158 171
rect 1192 137 1203 171
rect 1148 123 1203 137
rect 1233 238 1339 251
rect 1233 204 1294 238
rect 1328 204 1339 238
rect 1233 123 1339 204
rect 1369 239 1426 251
rect 1369 205 1380 239
rect 1414 205 1426 239
rect 1369 169 1426 205
rect 1369 135 1380 169
rect 1414 135 1426 169
rect 1670 201 1741 222
rect 1670 167 1696 201
rect 1730 167 1741 201
rect 1670 158 1741 167
rect 1369 123 1426 135
rect 1524 133 1625 158
rect 989 74 1050 106
rect 1004 72 1050 74
rect 1084 72 1094 106
rect 1524 99 1580 133
rect 1614 99 1625 133
rect 1524 74 1625 99
rect 1655 120 1741 158
rect 1655 86 1682 120
rect 1716 86 1741 120
rect 1655 74 1741 86
rect 1771 201 1827 222
rect 1771 167 1782 201
rect 1816 167 1827 201
rect 1771 120 1827 167
rect 1771 86 1782 120
rect 1816 86 1827 120
rect 1771 74 1827 86
rect 1857 210 1913 222
rect 1857 176 1868 210
rect 1902 176 1913 210
rect 1857 120 1913 176
rect 1857 86 1868 120
rect 1902 86 1913 120
rect 1857 74 1913 86
rect 1943 210 1999 222
rect 1943 176 1954 210
rect 1988 176 1999 210
rect 1943 120 1999 176
rect 1943 86 1954 120
rect 1988 86 1999 120
rect 1943 74 1999 86
rect 2029 210 2085 222
rect 2029 176 2040 210
rect 2074 176 2085 210
rect 2029 120 2085 176
rect 2029 86 2040 120
rect 2074 86 2085 120
rect 2029 74 2085 86
rect 1004 60 1094 72
<< pdiff >>
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 486 83 546
rect 27 452 39 486
rect 73 452 83 486
rect 27 392 83 452
rect 119 580 183 592
rect 119 546 129 580
rect 163 546 183 580
rect 119 486 183 546
rect 119 452 129 486
rect 163 452 183 486
rect 119 392 183 452
rect 219 580 275 592
rect 219 546 229 580
rect 263 560 275 580
rect 263 546 290 560
rect 219 508 290 546
rect 219 474 229 508
rect 263 474 290 508
rect 219 438 290 474
rect 219 404 229 438
rect 263 404 290 438
rect 219 392 290 404
rect 326 547 382 560
rect 326 513 336 547
rect 370 520 382 547
rect 573 546 623 547
rect 466 520 516 546
rect 370 513 397 520
rect 326 470 397 513
rect 326 436 336 470
rect 370 436 397 470
rect 326 392 397 436
rect 433 459 516 520
rect 433 425 443 459
rect 477 425 516 459
rect 433 418 516 425
rect 552 459 623 546
rect 552 425 579 459
rect 613 425 623 459
rect 552 418 623 425
rect 433 392 489 418
rect 567 379 623 418
rect 659 535 786 547
rect 659 501 731 535
rect 765 501 786 535
rect 659 431 786 501
rect 659 397 731 431
rect 765 397 786 431
rect 659 379 786 397
rect 895 580 951 592
rect 895 546 907 580
rect 941 546 951 580
rect 895 497 951 546
rect 895 463 907 497
rect 941 463 951 497
rect 895 414 951 463
rect 895 380 907 414
rect 941 380 951 414
rect 895 368 951 380
rect 987 580 1043 592
rect 1577 584 1707 592
rect 987 546 997 580
rect 1031 546 1043 580
rect 1577 580 1663 584
rect 987 497 1043 546
rect 987 463 997 497
rect 1031 463 1043 497
rect 987 414 1043 463
rect 987 380 997 414
rect 1031 380 1043 414
rect 1097 544 1185 556
rect 1097 510 1109 544
rect 1143 510 1185 544
rect 1097 434 1185 510
rect 1097 400 1109 434
rect 1143 400 1185 434
rect 1097 388 1185 400
rect 1221 531 1321 556
rect 1221 497 1277 531
rect 1311 497 1321 531
rect 1221 434 1321 497
rect 1221 400 1277 434
rect 1311 400 1321 434
rect 1221 388 1321 400
rect 1357 531 1413 556
rect 1577 546 1589 580
rect 1623 550 1663 580
rect 1697 550 1707 584
rect 1623 546 1707 550
rect 1577 538 1707 546
rect 1357 497 1367 531
rect 1401 497 1413 531
rect 1357 440 1413 497
rect 1357 406 1367 440
rect 1401 406 1413 440
rect 1470 508 1526 538
rect 1470 474 1482 508
rect 1516 474 1526 508
rect 1470 410 1526 474
rect 1562 516 1707 538
rect 1562 497 1663 516
rect 1562 463 1589 497
rect 1623 482 1663 497
rect 1697 482 1707 516
rect 1623 463 1707 482
rect 1562 414 1707 463
rect 1562 410 1589 414
rect 1357 388 1413 406
rect 987 368 1043 380
rect 1577 380 1589 410
rect 1623 380 1707 414
rect 1577 368 1707 380
rect 1743 580 1797 592
rect 1743 546 1753 580
rect 1787 546 1797 580
rect 1743 497 1797 546
rect 1743 463 1753 497
rect 1787 463 1797 497
rect 1743 414 1797 463
rect 1743 380 1753 414
rect 1787 380 1797 414
rect 1743 368 1797 380
rect 1833 580 1903 592
rect 1833 546 1859 580
rect 1893 546 1903 580
rect 1833 497 1903 546
rect 1833 463 1859 497
rect 1893 463 1903 497
rect 1833 414 1903 463
rect 1833 380 1859 414
rect 1893 380 1903 414
rect 1833 368 1903 380
rect 1939 580 1993 592
rect 1939 546 1949 580
rect 1983 546 1993 580
rect 1939 497 1993 546
rect 1939 463 1949 497
rect 1983 463 1993 497
rect 1939 414 1993 463
rect 1939 380 1949 414
rect 1983 380 1993 414
rect 1939 368 1993 380
rect 2029 580 2085 592
rect 2029 546 2039 580
rect 2073 546 2085 580
rect 2029 497 2085 546
rect 2029 463 2039 497
rect 2073 463 2085 497
rect 2029 414 2085 463
rect 2029 380 2039 414
rect 2073 380 2085 414
rect 2029 368 2085 380
<< ndiffc >>
rect 39 200 73 234
rect 39 130 73 164
rect 291 200 325 234
rect 427 200 461 234
rect 427 130 461 164
rect 527 187 561 221
rect 663 207 697 241
rect 663 130 697 164
rect 799 203 833 237
rect 149 48 183 82
rect 914 155 948 189
rect 1158 137 1192 171
rect 1294 204 1328 238
rect 1380 205 1414 239
rect 1380 135 1414 169
rect 1696 167 1730 201
rect 1050 72 1084 106
rect 1580 99 1614 133
rect 1682 86 1716 120
rect 1782 167 1816 201
rect 1782 86 1816 120
rect 1868 176 1902 210
rect 1868 86 1902 120
rect 1954 176 1988 210
rect 1954 86 1988 120
rect 2040 176 2074 210
rect 2040 86 2074 120
<< pdiffc >>
rect 39 546 73 580
rect 39 452 73 486
rect 129 546 163 580
rect 129 452 163 486
rect 229 546 263 580
rect 229 474 263 508
rect 229 404 263 438
rect 336 513 370 547
rect 336 436 370 470
rect 443 425 477 459
rect 579 425 613 459
rect 731 501 765 535
rect 731 397 765 431
rect 907 546 941 580
rect 907 463 941 497
rect 907 380 941 414
rect 997 546 1031 580
rect 997 463 1031 497
rect 997 380 1031 414
rect 1109 510 1143 544
rect 1109 400 1143 434
rect 1277 497 1311 531
rect 1277 400 1311 434
rect 1589 546 1623 580
rect 1663 550 1697 584
rect 1367 497 1401 531
rect 1367 406 1401 440
rect 1482 474 1516 508
rect 1589 463 1623 497
rect 1663 482 1697 516
rect 1589 380 1623 414
rect 1753 546 1787 580
rect 1753 463 1787 497
rect 1753 380 1787 414
rect 1859 546 1893 580
rect 1859 463 1893 497
rect 1859 380 1893 414
rect 1949 546 1983 580
rect 1949 463 1983 497
rect 1949 380 1983 414
rect 2039 546 2073 580
rect 2039 463 2073 497
rect 2039 380 2073 414
<< poly >>
rect 83 592 119 618
rect 183 592 219 618
rect 290 615 880 645
rect 290 560 326 615
rect 516 546 552 615
rect 623 547 659 573
rect 397 520 433 546
rect 516 392 552 418
rect 83 360 119 392
rect 74 344 140 360
rect 74 310 90 344
rect 124 310 140 344
rect 183 334 219 392
rect 290 366 326 392
rect 397 350 433 392
rect 623 350 659 379
rect 74 294 140 310
rect 182 318 248 334
rect 397 331 797 350
rect 397 320 747 331
rect 84 246 114 294
rect 182 284 198 318
rect 232 284 248 318
rect 182 268 248 284
rect 218 246 248 268
rect 386 246 416 272
rect 486 246 516 320
rect 724 297 747 320
rect 781 297 797 331
rect 724 281 797 297
rect 850 310 880 615
rect 951 592 987 618
rect 1707 592 1743 618
rect 1797 592 1833 618
rect 1903 592 1939 618
rect 1993 592 2029 618
rect 1185 556 1221 582
rect 1321 556 1357 582
rect 1526 538 1562 564
rect 1526 395 1562 410
rect 951 310 987 368
rect 1185 350 1221 388
rect 1321 356 1357 388
rect 1441 365 1562 395
rect 1441 356 1471 365
rect 1155 334 1233 350
rect 850 294 1048 310
rect 606 246 636 272
rect 724 253 754 281
rect 850 280 998 294
rect 486 136 516 162
rect 84 92 114 118
rect 218 92 248 118
rect 386 51 416 118
rect 606 51 636 118
rect 724 99 754 125
rect 858 51 888 280
rect 951 260 998 280
rect 1032 260 1048 294
rect 1155 300 1171 334
rect 1205 300 1233 334
rect 1155 284 1233 300
rect 1321 340 1471 356
rect 1321 306 1371 340
rect 1405 306 1471 340
rect 1707 317 1743 368
rect 1797 317 1833 368
rect 1903 317 1939 368
rect 1993 317 2029 368
rect 1321 290 1471 306
rect 951 244 1048 260
rect 1203 251 1233 284
rect 1339 251 1369 290
rect 959 222 989 244
rect 1441 203 1471 290
rect 1570 301 2029 317
rect 1570 267 1586 301
rect 1620 267 1654 301
rect 1688 267 1722 301
rect 1756 267 2029 301
rect 1570 251 2029 267
rect 1741 222 1771 251
rect 1827 222 1857 251
rect 1913 222 1943 251
rect 1999 222 2029 251
rect 1441 173 1655 203
rect 1625 158 1655 173
rect 386 21 888 51
rect 959 48 989 74
rect 1203 97 1233 123
rect 1339 97 1369 123
rect 1625 48 1655 74
rect 1741 48 1771 74
rect 1827 48 1857 74
rect 1913 48 1943 74
rect 1999 48 2029 74
<< polycont >>
rect 90 310 124 344
rect 198 284 232 318
rect 747 297 781 331
rect 998 260 1032 294
rect 1171 300 1205 334
rect 1371 306 1405 340
rect 1586 267 1620 301
rect 1654 267 1688 301
rect 1722 267 1756 301
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 17 580 73 596
rect 17 546 39 580
rect 17 486 73 546
rect 17 452 39 486
rect 17 436 73 452
rect 113 580 179 649
rect 113 546 129 580
rect 163 546 179 580
rect 113 486 179 546
rect 113 452 129 486
rect 163 452 179 486
rect 113 436 179 452
rect 213 581 765 615
rect 213 580 279 581
rect 213 546 229 580
rect 263 546 279 580
rect 731 551 765 581
rect 907 580 941 596
rect 213 508 279 546
rect 213 474 229 508
rect 263 474 279 508
rect 213 438 279 474
rect 17 250 51 436
rect 213 404 229 438
rect 263 404 279 438
rect 320 513 336 547
rect 370 513 697 547
rect 320 470 386 513
rect 320 436 336 470
rect 370 436 386 470
rect 427 459 477 479
rect 213 402 279 404
rect 427 425 443 459
rect 85 368 325 402
rect 85 344 140 368
rect 85 310 90 344
rect 124 310 140 344
rect 85 294 140 310
rect 182 318 257 334
rect 182 284 198 318
rect 232 284 257 318
rect 17 234 89 250
rect 182 236 257 284
rect 17 200 39 234
rect 73 200 89 234
rect 17 164 89 200
rect 291 234 325 368
rect 427 318 477 425
rect 511 459 629 479
rect 511 425 579 459
rect 613 425 629 459
rect 511 424 629 425
rect 545 390 629 424
rect 511 375 629 390
rect 291 184 325 200
rect 359 284 561 318
rect 17 130 39 164
rect 73 150 89 164
rect 359 150 393 284
rect 73 130 393 150
rect 17 116 393 130
rect 427 234 477 250
rect 461 200 477 234
rect 427 164 477 200
rect 461 130 477 164
rect 511 221 561 284
rect 511 187 527 221
rect 511 158 561 187
rect 427 124 477 130
rect 595 124 629 375
rect 17 114 89 116
rect 427 90 629 124
rect 663 241 697 513
rect 731 535 865 551
rect 765 501 865 535
rect 731 431 865 501
rect 765 397 865 431
rect 731 381 865 397
rect 663 164 697 207
rect 663 85 697 130
rect 731 331 797 347
rect 731 297 747 331
rect 781 297 797 331
rect 731 287 797 297
rect 731 153 765 287
rect 831 253 865 381
rect 799 237 865 253
rect 833 203 865 237
rect 799 187 865 203
rect 907 497 941 546
rect 907 414 941 463
rect 907 226 941 380
rect 981 580 1047 649
rect 981 546 997 580
rect 1031 546 1047 580
rect 1193 581 1500 615
rect 981 497 1047 546
rect 981 463 997 497
rect 1031 463 1047 497
rect 981 414 1047 463
rect 981 380 997 414
rect 1031 380 1047 414
rect 1081 544 1159 560
rect 1081 510 1109 544
rect 1143 510 1159 544
rect 1081 434 1159 510
rect 1081 424 1109 434
rect 1081 390 1087 424
rect 1143 400 1159 434
rect 1121 390 1159 400
rect 1081 384 1159 390
rect 981 364 1047 380
rect 982 294 1048 310
rect 982 260 998 294
rect 1032 260 1048 294
rect 982 236 1048 260
rect 1087 258 1121 384
rect 1193 350 1227 581
rect 1261 531 1328 547
rect 1261 497 1277 531
rect 1311 497 1328 531
rect 1261 434 1328 497
rect 1261 400 1277 434
rect 1311 424 1328 434
rect 1261 390 1279 400
rect 1313 390 1328 424
rect 1367 531 1417 547
rect 1401 497 1417 531
rect 1367 440 1417 497
rect 1466 542 1500 581
rect 1589 584 1700 649
rect 1589 580 1663 584
rect 1623 550 1663 580
rect 1697 550 1700 584
rect 1623 546 1700 550
rect 1466 508 1550 542
rect 1466 474 1482 508
rect 1516 474 1550 508
rect 1466 458 1550 474
rect 1401 424 1417 440
rect 1401 406 1482 424
rect 1367 390 1482 406
rect 1261 384 1328 390
rect 1155 334 1227 350
rect 1155 300 1171 334
rect 1205 300 1227 334
rect 1155 292 1227 300
rect 907 189 948 226
rect 1087 224 1260 258
rect 907 155 914 189
rect 907 153 948 155
rect 731 119 948 153
rect 982 171 1192 190
rect 982 156 1158 171
rect 982 85 1016 156
rect 1142 137 1158 156
rect 125 48 149 82
rect 183 48 207 82
rect 663 51 1016 85
rect 1050 106 1100 122
rect 1084 72 1100 106
rect 125 17 207 48
rect 1050 17 1100 72
rect 1142 85 1192 137
rect 1226 153 1260 224
rect 1294 238 1328 384
rect 1362 340 1414 356
rect 1362 306 1371 340
rect 1405 306 1414 340
rect 1362 290 1414 306
rect 1294 187 1328 204
rect 1364 239 1414 255
rect 1364 205 1380 239
rect 1364 169 1414 205
rect 1364 153 1380 169
rect 1226 135 1380 153
rect 1226 119 1414 135
rect 1448 85 1482 390
rect 1142 51 1482 85
rect 1516 149 1550 458
rect 1589 516 1700 546
rect 1589 497 1663 516
rect 1623 482 1663 497
rect 1697 482 1700 516
rect 1623 466 1700 482
rect 1737 580 1825 596
rect 1737 546 1753 580
rect 1787 546 1825 580
rect 1737 497 1825 546
rect 1589 414 1623 463
rect 1737 463 1753 497
rect 1787 463 1825 497
rect 1589 364 1623 380
rect 1657 424 1703 430
rect 1657 390 1663 424
rect 1697 390 1703 424
rect 1657 317 1703 390
rect 1737 414 1825 463
rect 1737 380 1753 414
rect 1787 380 1825 414
rect 1737 364 1825 380
rect 1859 580 1893 649
rect 1859 497 1893 546
rect 1859 414 1893 463
rect 1859 364 1893 380
rect 1933 580 1999 596
rect 1933 546 1949 580
rect 1983 546 1999 580
rect 1933 497 1999 546
rect 1933 463 1949 497
rect 1983 463 1999 497
rect 1933 414 1999 463
rect 1933 380 1949 414
rect 1983 380 1999 414
rect 1584 301 1757 317
rect 1584 267 1586 301
rect 1620 267 1654 301
rect 1688 267 1722 301
rect 1756 267 1757 301
rect 1584 251 1757 267
rect 1791 294 1825 364
rect 1933 310 1999 380
rect 2039 580 2089 649
rect 2073 546 2089 580
rect 2039 497 2089 546
rect 2073 463 2089 497
rect 2039 414 2089 463
rect 2073 380 2089 414
rect 2039 364 2089 380
rect 1933 294 1988 310
rect 1791 260 1988 294
rect 1791 217 1832 260
rect 1666 201 1732 217
rect 1666 167 1696 201
rect 1730 167 1732 201
rect 1516 133 1630 149
rect 1516 99 1580 133
rect 1614 99 1630 133
rect 1516 83 1630 99
rect 1666 120 1732 167
rect 1666 86 1682 120
rect 1716 86 1732 120
rect 1666 17 1732 86
rect 1766 201 1832 217
rect 1766 167 1782 201
rect 1816 167 1832 201
rect 1766 120 1832 167
rect 1766 86 1782 120
rect 1816 86 1832 120
rect 1766 70 1832 86
rect 1868 210 1902 226
rect 1868 120 1902 176
rect 1868 17 1902 86
rect 1938 210 1988 260
rect 1938 176 1954 210
rect 1938 120 1988 176
rect 1938 86 1954 120
rect 1938 70 1988 86
rect 2024 210 2090 226
rect 2024 176 2040 210
rect 2074 176 2090 210
rect 2024 120 2090 176
rect 2024 86 2040 120
rect 2074 86 2090 120
rect 2024 17 2090 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 511 390 545 424
rect 1087 400 1109 424
rect 1109 400 1121 424
rect 1087 390 1121 400
rect 1279 400 1311 424
rect 1311 400 1313 424
rect 1279 390 1313 400
rect 1663 390 1697 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
<< metal1 >>
rect 0 683 2112 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 0 617 2112 649
rect 499 424 557 430
rect 499 390 511 424
rect 545 421 557 424
rect 1075 424 1133 430
rect 1075 421 1087 424
rect 545 393 1087 421
rect 545 390 557 393
rect 499 384 557 390
rect 1075 390 1087 393
rect 1121 390 1133 424
rect 1075 384 1133 390
rect 1267 424 1325 430
rect 1267 390 1279 424
rect 1313 421 1325 424
rect 1651 424 1709 430
rect 1651 421 1663 424
rect 1313 393 1663 421
rect 1313 390 1325 393
rect 1267 384 1325 390
rect 1651 390 1663 393
rect 1697 390 1709 424
rect 1651 384 1709 390
rect 0 17 2112 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
rect 0 -49 2112 -17
<< labels >>
flabel pwell s 0 0 2112 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 2112 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
rlabel comment s 0 0 0 0 4 xor3_4
flabel metal1 s 0 617 2112 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 2112 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 1951 316 1985 350 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 1951 390 1985 424 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 1951 464 1985 498 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 1951 538 1985 572 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 991 242 1025 276 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 1375 316 1409 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 223 242 257 276 0 FreeSans 340 0 0 0 A
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 2112 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 602122
string GDS_START 586892
<< end >>
