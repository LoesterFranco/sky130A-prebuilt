magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 710 704
<< pwell >>
rect 0 0 672 49
<< scnmos >>
rect 103 136 133 264
rect 217 136 247 264
rect 295 136 325 264
rect 411 82 441 230
rect 505 82 535 230
<< pmoshvt >>
rect 100 384 130 552
rect 214 384 244 552
rect 304 384 334 552
rect 448 368 478 592
rect 538 368 568 592
<< ndiff >>
rect 46 235 103 264
rect 46 201 58 235
rect 92 201 103 235
rect 46 136 103 201
rect 133 136 217 264
rect 247 136 295 264
rect 325 230 375 264
rect 325 222 411 230
rect 325 188 352 222
rect 386 188 411 222
rect 325 136 411 188
rect 340 128 411 136
rect 340 94 352 128
rect 386 94 411 128
rect 340 82 411 94
rect 441 218 505 230
rect 441 184 452 218
rect 486 184 505 218
rect 441 128 505 184
rect 441 94 452 128
rect 486 94 505 128
rect 441 82 505 94
rect 535 218 631 230
rect 535 184 585 218
rect 619 184 631 218
rect 535 128 631 184
rect 535 94 575 128
rect 609 94 631 128
rect 535 82 631 94
<< pdiff >>
rect 379 580 448 592
rect 379 552 391 580
rect 41 540 100 552
rect 41 506 53 540
rect 87 506 100 540
rect 41 430 100 506
rect 41 396 53 430
rect 87 396 100 430
rect 41 384 100 396
rect 130 508 214 552
rect 130 474 153 508
rect 187 474 214 508
rect 130 384 214 474
rect 244 540 304 552
rect 244 506 257 540
rect 291 506 304 540
rect 244 440 304 506
rect 244 406 257 440
rect 291 406 304 440
rect 244 384 304 406
rect 334 546 391 552
rect 425 546 448 580
rect 334 508 448 546
rect 334 474 391 508
rect 425 474 448 508
rect 334 384 448 474
rect 395 368 448 384
rect 478 580 538 592
rect 478 546 491 580
rect 525 546 538 580
rect 478 499 538 546
rect 478 465 491 499
rect 525 465 538 499
rect 478 418 538 465
rect 478 384 491 418
rect 525 384 538 418
rect 478 368 538 384
rect 568 580 641 592
rect 568 546 595 580
rect 629 546 641 580
rect 568 497 641 546
rect 568 463 595 497
rect 629 463 641 497
rect 568 414 641 463
rect 568 380 595 414
rect 629 380 641 414
rect 568 368 641 380
<< ndiffc >>
rect 58 201 92 235
rect 352 188 386 222
rect 352 94 386 128
rect 452 184 486 218
rect 452 94 486 128
rect 585 184 619 218
rect 575 94 609 128
<< pdiffc >>
rect 53 506 87 540
rect 53 396 87 430
rect 153 474 187 508
rect 257 506 291 540
rect 257 406 291 440
rect 391 546 425 580
rect 391 474 425 508
rect 491 546 525 580
rect 491 465 525 499
rect 491 384 525 418
rect 595 546 629 580
rect 595 463 629 497
rect 595 380 629 414
<< poly >>
rect 448 592 478 618
rect 538 592 568 618
rect 100 552 130 578
rect 214 552 244 578
rect 304 552 334 578
rect 100 369 130 384
rect 214 369 244 384
rect 304 369 334 384
rect 97 279 133 369
rect 211 352 247 369
rect 301 352 337 369
rect 448 353 478 368
rect 538 353 568 368
rect 181 336 247 352
rect 181 302 197 336
rect 231 302 247 336
rect 181 286 247 302
rect 103 264 133 279
rect 217 264 247 286
rect 295 336 363 352
rect 295 302 313 336
rect 347 302 363 336
rect 445 334 481 353
rect 535 334 571 353
rect 295 286 363 302
rect 411 318 571 334
rect 295 264 325 286
rect 411 284 427 318
rect 461 284 571 318
rect 411 268 571 284
rect 411 230 441 268
rect 505 230 535 268
rect 103 114 133 136
rect 25 98 159 114
rect 217 110 247 136
rect 295 110 325 136
rect 25 64 41 98
rect 75 64 109 98
rect 143 64 159 98
rect 25 48 159 64
rect 411 56 441 82
rect 505 56 535 82
<< polycont >>
rect 197 302 231 336
rect 313 302 347 336
rect 427 284 461 318
rect 41 64 75 98
rect 109 64 143 98
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 37 540 103 556
rect 37 506 53 540
rect 87 506 103 540
rect 37 430 103 506
rect 137 508 203 649
rect 375 580 441 649
rect 137 474 153 508
rect 187 474 203 508
rect 137 458 203 474
rect 241 540 307 556
rect 241 506 257 540
rect 291 506 307 540
rect 37 396 53 430
rect 87 424 103 430
rect 241 440 307 506
rect 375 546 391 580
rect 425 546 441 580
rect 375 508 441 546
rect 375 474 391 508
rect 425 474 441 508
rect 375 458 441 474
rect 475 580 545 596
rect 475 546 491 580
rect 525 546 545 580
rect 475 499 545 546
rect 475 465 491 499
rect 525 465 545 499
rect 241 424 257 440
rect 87 406 257 424
rect 291 424 307 440
rect 291 406 441 424
rect 87 396 441 406
rect 37 390 441 396
rect 37 268 103 390
rect 181 336 263 356
rect 181 302 197 336
rect 231 302 263 336
rect 37 235 108 268
rect 181 236 263 302
rect 297 336 363 356
rect 297 302 313 336
rect 347 302 363 336
rect 297 286 363 302
rect 407 334 441 390
rect 475 418 545 465
rect 475 384 491 418
rect 525 384 545 418
rect 475 368 545 384
rect 407 318 477 334
rect 407 284 427 318
rect 461 284 477 318
rect 407 268 477 284
rect 37 201 58 235
rect 92 201 108 235
rect 511 234 545 368
rect 579 580 645 649
rect 579 546 595 580
rect 629 546 645 580
rect 579 497 645 546
rect 579 463 595 497
rect 629 463 645 497
rect 579 414 645 463
rect 579 380 595 414
rect 629 380 645 414
rect 579 364 645 380
rect 37 168 108 201
rect 336 222 402 234
rect 336 188 352 222
rect 386 188 402 222
rect 25 98 263 134
rect 25 64 41 98
rect 75 64 109 98
rect 143 64 263 98
rect 25 51 263 64
rect 336 128 402 188
rect 336 94 352 128
rect 386 94 402 128
rect 336 17 402 94
rect 436 218 551 234
rect 436 184 452 218
rect 486 184 551 218
rect 436 162 551 184
rect 585 218 649 234
rect 619 184 649 218
rect 436 128 502 162
rect 585 128 649 184
rect 436 94 452 128
rect 486 94 502 128
rect 436 78 502 94
rect 536 94 575 128
rect 609 94 649 128
rect 536 17 649 94
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel comment s 0 0 0 0 4 and3_2
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 511 168 545 202 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 31 94 65 128 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 127 94 161 128 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 223 94 257 128 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 223 242 257 276 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 B
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 672 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3079460
string GDS_START 3073094
<< end >>
