magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 1050 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 89 47 119 177
rect 183 47 213 177
rect 267 47 297 177
rect 371 47 401 177
rect 587 47 617 177
rect 681 47 711 177
rect 765 47 795 177
rect 859 47 889 177
<< pmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 489 297 525 497
rect 583 297 619 497
rect 767 297 803 497
rect 861 297 897 497
<< ndiff >>
rect 27 161 89 177
rect 27 127 35 161
rect 69 127 89 161
rect 27 93 89 127
rect 27 59 35 93
rect 69 59 89 93
rect 27 47 89 59
rect 119 93 183 177
rect 119 59 129 93
rect 163 59 183 93
rect 119 47 183 59
rect 213 161 267 177
rect 213 127 223 161
rect 257 127 267 161
rect 213 93 267 127
rect 213 59 223 93
rect 257 59 267 93
rect 213 47 267 59
rect 297 161 371 177
rect 297 127 317 161
rect 351 127 371 161
rect 297 47 371 127
rect 401 93 457 177
rect 401 59 415 93
rect 449 59 457 93
rect 401 47 457 59
rect 511 93 587 177
rect 511 59 529 93
rect 563 59 587 93
rect 511 47 587 59
rect 617 161 681 177
rect 617 127 627 161
rect 661 127 681 161
rect 617 47 681 127
rect 711 161 765 177
rect 711 127 721 161
rect 755 127 765 161
rect 711 93 765 127
rect 711 59 721 93
rect 755 59 765 93
rect 711 47 765 59
rect 795 161 859 177
rect 795 127 815 161
rect 849 127 859 161
rect 795 47 859 127
rect 889 161 971 177
rect 889 127 925 161
rect 959 127 971 161
rect 889 93 971 127
rect 889 59 925 93
rect 959 59 971 93
rect 889 47 971 59
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 485 175 497
rect 117 451 129 485
rect 163 451 175 485
rect 117 417 175 451
rect 117 383 129 417
rect 163 383 175 417
rect 117 349 175 383
rect 117 315 129 349
rect 163 315 175 349
rect 117 297 175 315
rect 211 485 269 497
rect 211 451 223 485
rect 257 451 269 485
rect 211 417 269 451
rect 211 383 223 417
rect 257 383 269 417
rect 211 297 269 383
rect 305 485 363 497
rect 305 451 317 485
rect 351 451 363 485
rect 305 417 363 451
rect 305 383 317 417
rect 351 383 363 417
rect 305 349 363 383
rect 305 315 317 349
rect 351 315 363 349
rect 305 297 363 315
rect 399 485 489 497
rect 399 451 427 485
rect 461 451 489 485
rect 399 417 489 451
rect 399 383 427 417
rect 461 383 489 417
rect 399 297 489 383
rect 525 485 583 497
rect 525 451 537 485
rect 571 451 583 485
rect 525 417 583 451
rect 525 383 537 417
rect 571 383 583 417
rect 525 349 583 383
rect 525 315 537 349
rect 571 315 583 349
rect 525 297 583 315
rect 619 485 767 497
rect 619 451 675 485
rect 709 451 767 485
rect 619 417 767 451
rect 619 383 675 417
rect 709 383 767 417
rect 619 297 767 383
rect 803 485 861 497
rect 803 451 815 485
rect 849 451 861 485
rect 803 417 861 451
rect 803 383 815 417
rect 849 383 861 417
rect 803 349 861 383
rect 803 315 815 349
rect 849 315 861 349
rect 803 297 861 315
rect 897 485 983 497
rect 897 451 925 485
rect 959 451 983 485
rect 897 417 983 451
rect 897 383 925 417
rect 959 383 983 417
rect 897 349 983 383
rect 897 315 925 349
rect 959 315 983 349
rect 897 297 983 315
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 129 59 163 93
rect 223 127 257 161
rect 223 59 257 93
rect 317 127 351 161
rect 415 59 449 93
rect 529 59 563 93
rect 627 127 661 161
rect 721 127 755 161
rect 721 59 755 93
rect 815 127 849 161
rect 925 127 959 161
rect 925 59 959 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 451 163 485
rect 129 383 163 417
rect 129 315 163 349
rect 223 451 257 485
rect 223 383 257 417
rect 317 451 351 485
rect 317 383 351 417
rect 317 315 351 349
rect 427 451 461 485
rect 427 383 461 417
rect 537 451 571 485
rect 537 383 571 417
rect 537 315 571 349
rect 675 451 709 485
rect 675 383 709 417
rect 815 451 849 485
rect 815 383 849 417
rect 815 315 849 349
rect 925 451 959 485
rect 925 383 959 417
rect 925 315 959 349
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 489 497 525 523
rect 583 497 619 523
rect 767 497 803 523
rect 861 497 897 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 489 282 525 297
rect 583 282 619 297
rect 767 282 803 297
rect 861 282 897 297
rect 79 261 119 282
rect 22 259 119 261
rect 173 259 213 282
rect 22 249 213 259
rect 22 215 38 249
rect 72 215 129 249
rect 163 215 213 249
rect 22 205 213 215
rect 89 177 119 205
rect 183 177 213 205
rect 267 259 307 282
rect 361 259 401 282
rect 267 249 401 259
rect 267 215 317 249
rect 351 215 401 249
rect 267 205 401 215
rect 487 259 527 282
rect 581 259 621 282
rect 765 259 805 282
rect 859 261 899 282
rect 859 259 989 261
rect 487 249 711 259
rect 487 215 503 249
rect 537 215 621 249
rect 655 215 711 249
rect 487 205 711 215
rect 267 177 297 205
rect 371 177 401 205
rect 587 177 617 205
rect 681 177 711 205
rect 765 249 989 259
rect 765 215 939 249
rect 973 215 989 249
rect 765 205 989 215
rect 765 177 795 205
rect 859 177 889 205
rect 89 21 119 47
rect 183 21 213 47
rect 267 21 297 47
rect 371 21 401 47
rect 587 21 617 47
rect 681 21 711 47
rect 765 21 795 47
rect 859 21 889 47
<< polycont >>
rect 38 215 72 249
rect 129 215 163 249
rect 317 215 351 249
rect 503 215 537 249
rect 621 215 655 249
rect 939 215 973 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 18 485 69 527
rect 18 451 35 485
rect 18 417 69 451
rect 18 383 35 417
rect 18 349 69 383
rect 18 315 35 349
rect 18 299 69 315
rect 103 485 179 493
rect 103 451 129 485
rect 163 451 179 485
rect 103 417 179 451
rect 103 383 129 417
rect 163 383 179 417
rect 103 349 179 383
rect 223 485 257 527
rect 223 417 257 451
rect 223 367 257 383
rect 291 485 367 493
rect 291 451 317 485
rect 351 451 367 485
rect 291 417 367 451
rect 291 383 317 417
rect 351 383 367 417
rect 103 315 129 349
rect 163 333 179 349
rect 291 349 367 383
rect 411 485 477 527
rect 411 451 427 485
rect 461 451 477 485
rect 411 417 477 451
rect 411 383 427 417
rect 461 383 477 417
rect 411 367 477 383
rect 511 485 587 493
rect 511 451 537 485
rect 571 451 587 485
rect 511 417 587 451
rect 511 383 537 417
rect 571 383 587 417
rect 291 333 317 349
rect 163 315 317 333
rect 351 333 367 349
rect 511 349 587 383
rect 659 485 735 527
rect 659 451 675 485
rect 709 451 735 485
rect 659 417 735 451
rect 659 383 675 417
rect 709 383 735 417
rect 659 367 735 383
rect 789 485 865 493
rect 789 451 815 485
rect 849 451 865 485
rect 789 417 865 451
rect 789 383 815 417
rect 849 383 865 417
rect 511 333 537 349
rect 351 315 537 333
rect 571 333 587 349
rect 789 349 865 383
rect 789 333 815 349
rect 571 315 815 333
rect 849 315 865 349
rect 103 289 865 315
rect 909 485 975 527
rect 909 451 925 485
rect 959 451 975 485
rect 909 417 975 451
rect 909 383 925 417
rect 959 383 975 417
rect 909 349 975 383
rect 909 315 925 349
rect 959 315 975 349
rect 909 289 975 315
rect 22 249 179 255
rect 22 215 38 249
rect 72 215 129 249
rect 163 215 179 249
rect 213 249 370 255
rect 213 215 317 249
rect 351 215 370 249
rect 487 249 676 255
rect 487 215 503 249
rect 537 215 621 249
rect 655 215 676 249
rect 744 211 865 289
rect 923 249 989 255
rect 923 215 939 249
rect 973 215 989 249
rect 18 161 257 181
rect 18 127 35 161
rect 69 147 223 161
rect 69 127 85 147
rect 18 93 85 127
rect 197 127 223 147
rect 291 161 677 181
rect 291 127 317 161
rect 351 127 627 161
rect 661 127 677 161
rect 721 161 755 177
rect 789 161 865 211
rect 789 127 815 161
rect 849 127 865 161
rect 909 161 975 181
rect 909 127 925 161
rect 959 127 975 161
rect 18 59 35 93
rect 69 59 85 93
rect 18 51 85 59
rect 129 93 163 109
rect 129 17 163 59
rect 197 93 257 127
rect 721 93 755 127
rect 909 93 975 127
rect 197 59 223 93
rect 257 59 415 93
rect 449 59 465 93
rect 197 51 465 59
rect 503 59 529 93
rect 563 59 721 93
rect 755 59 925 93
rect 959 59 975 93
rect 503 51 975 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
flabel corelocali s 642 221 676 255 0 FreeSans 250 0 0 0 B
port 2 nsew
flabel corelocali s 540 221 574 255 0 FreeSans 250 0 0 0 B
port 2 nsew
flabel corelocali s 947 221 981 255 0 FreeSans 250 0 0 0 A
port 1 nsew
flabel corelocali s 540 289 574 323 0 FreeSans 250 0 0 0 Y
port 9 nsew
flabel corelocali s 642 289 676 323 0 FreeSans 250 0 0 0 Y
port 9 nsew
flabel corelocali s 744 221 778 255 0 FreeSans 250 0 0 0 Y
port 9 nsew
flabel corelocali s 744 289 778 323 0 FreeSans 250 0 0 0 Y
port 9 nsew
flabel corelocali s 132 221 166 255 0 FreeSans 250 0 0 0 D
port 4 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 250 0 0 0 D
port 4 nsew
flabel corelocali s 336 221 370 255 0 FreeSans 250 0 0 0 C
port 3 nsew
flabel corelocali s 234 221 268 255 0 FreeSans 250 0 0 0 C
port 3 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
rlabel comment s 0 0 0 0 4 nand4_2
<< properties >>
string FIXED_BBOX 0 0 1012 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2301954
string GDS_START 2293066
<< end >>
