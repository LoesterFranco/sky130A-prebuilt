magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 2208 561
rect 103 427 169 527
rect 19 195 89 325
rect 103 17 169 93
rect 375 449 441 527
rect 352 176 386 337
rect 748 433 782 527
rect 488 271 555 337
rect 352 175 388 176
rect 352 174 389 175
rect 352 172 390 174
rect 352 171 391 172
rect 352 170 392 171
rect 352 168 393 170
rect 352 167 394 168
rect 352 164 395 167
rect 352 162 398 164
rect 352 157 402 162
rect 613 157 647 223
rect 703 211 799 331
rect 352 150 647 157
rect 358 147 647 150
rect 361 145 647 147
rect 364 143 647 145
rect 366 141 647 143
rect 368 138 647 141
rect 372 131 647 138
rect 375 123 647 131
rect 391 17 457 89
rect 491 61 526 123
rect 749 17 789 109
rect 1177 367 1211 527
rect 1553 427 1614 527
rect 1768 325 1802 527
rect 1135 17 1209 117
rect 1840 308 1906 493
rect 1840 301 1922 308
rect 1871 286 1922 301
rect 1878 165 1922 286
rect 1540 17 1614 123
rect 1836 158 1922 165
rect 2042 299 2103 527
rect 2137 289 2188 465
rect 1836 145 1912 158
rect 1768 17 1802 139
rect 1836 61 1906 145
rect 2037 17 2103 161
rect 2146 159 2188 289
rect 2137 53 2188 159
rect 0 -17 2208 17
<< obsli1 >>
rect 35 393 69 493
rect 35 391 169 393
rect 35 359 129 391
rect 123 357 129 359
rect 163 357 169 391
rect 123 194 169 357
rect 123 161 162 194
rect 35 127 162 161
rect 203 187 237 493
rect 35 69 69 127
rect 203 69 237 153
rect 284 415 341 489
rect 535 449 714 483
rect 284 372 646 415
rect 284 117 318 372
rect 420 225 454 372
rect 612 337 646 372
rect 680 399 714 449
rect 833 414 890 488
rect 929 438 1143 472
rect 833 399 867 414
rect 680 365 867 399
rect 987 391 1075 402
rect 612 271 651 337
rect 420 191 489 225
rect 833 177 867 365
rect 681 143 867 177
rect 284 51 341 117
rect 681 89 715 143
rect 560 55 715 89
rect 833 107 867 143
rect 901 207 949 381
rect 987 357 1033 391
rect 1067 357 1075 391
rect 987 331 1075 357
rect 1109 315 1143 438
rect 1245 427 1295 493
rect 1340 433 1517 467
rect 1109 297 1211 315
rect 1051 263 1211 297
rect 901 187 1017 207
rect 901 153 949 187
rect 983 153 1017 187
rect 901 141 1017 153
rect 1051 107 1085 263
rect 1177 249 1211 263
rect 1119 213 1153 219
rect 1245 213 1279 427
rect 1313 391 1351 393
rect 1313 357 1315 391
rect 1349 357 1351 391
rect 1313 249 1351 357
rect 1385 315 1449 381
rect 1119 153 1279 213
rect 1385 207 1423 315
rect 1483 281 1517 433
rect 1676 381 1734 491
rect 1551 315 1734 381
rect 833 73 903 107
rect 937 73 1085 107
rect 1245 107 1279 153
rect 1313 187 1423 207
rect 1313 153 1317 187
rect 1351 153 1423 187
rect 1313 141 1423 153
rect 1457 265 1517 281
rect 1697 265 1734 315
rect 1940 337 2006 485
rect 1457 199 1663 265
rect 1697 199 1844 265
rect 1457 107 1491 199
rect 1697 165 1734 199
rect 1245 73 1337 107
rect 1383 73 1491 107
rect 1668 60 1734 165
rect 1956 265 2006 337
rect 1956 199 2112 265
rect 1956 124 1990 199
rect 1940 69 1990 124
<< obsli1c >>
rect 129 357 163 391
rect 203 153 237 187
rect 1033 357 1067 391
rect 949 153 983 187
rect 1315 357 1349 391
rect 1317 153 1351 187
<< metal1 >>
rect 0 496 2208 592
rect 0 -48 2208 48
<< obsm1 >>
rect 117 391 175 397
rect 117 357 129 391
rect 163 388 175 391
rect 1021 391 1079 397
rect 1021 388 1033 391
rect 163 360 1033 388
rect 163 357 175 360
rect 117 351 175 357
rect 1021 357 1033 360
rect 1067 388 1079 391
rect 1303 391 1361 397
rect 1303 388 1315 391
rect 1067 360 1315 388
rect 1067 357 1079 360
rect 1021 351 1079 357
rect 1303 357 1315 360
rect 1349 357 1361 391
rect 1303 351 1361 357
rect 191 187 249 193
rect 191 153 203 187
rect 237 184 249 187
rect 937 187 995 193
rect 937 184 949 187
rect 237 156 949 184
rect 237 153 249 156
rect 191 147 249 153
rect 937 153 949 156
rect 983 184 995 187
rect 1305 187 1363 193
rect 1305 184 1317 187
rect 983 156 1317 184
rect 983 153 995 156
rect 937 147 995 153
rect 1305 153 1317 156
rect 1351 153 1363 187
rect 1305 147 1363 153
<< labels >>
rlabel locali s 488 271 555 337 6 D
port 1 nsew signal input
rlabel locali s 1878 165 1922 286 6 Q
port 2 nsew signal output
rlabel locali s 1871 286 1922 301 6 Q
port 2 nsew signal output
rlabel locali s 1840 308 1906 493 6 Q
port 2 nsew signal output
rlabel locali s 1840 301 1922 308 6 Q
port 2 nsew signal output
rlabel locali s 1836 158 1922 165 6 Q
port 2 nsew signal output
rlabel locali s 1836 145 1912 158 6 Q
port 2 nsew signal output
rlabel locali s 1836 61 1906 145 6 Q
port 2 nsew signal output
rlabel locali s 2146 159 2188 289 6 Q_N
port 3 nsew signal output
rlabel locali s 2137 289 2188 465 6 Q_N
port 3 nsew signal output
rlabel locali s 2137 53 2188 159 6 Q_N
port 3 nsew signal output
rlabel locali s 703 211 799 331 6 SCD
port 4 nsew signal input
rlabel locali s 613 157 647 223 6 SCE
port 5 nsew signal input
rlabel locali s 491 61 526 123 6 SCE
port 5 nsew signal input
rlabel locali s 375 123 647 131 6 SCE
port 5 nsew signal input
rlabel locali s 372 131 647 138 6 SCE
port 5 nsew signal input
rlabel locali s 368 138 647 141 6 SCE
port 5 nsew signal input
rlabel locali s 366 141 647 143 6 SCE
port 5 nsew signal input
rlabel locali s 364 143 647 145 6 SCE
port 5 nsew signal input
rlabel locali s 361 145 647 147 6 SCE
port 5 nsew signal input
rlabel locali s 358 147 647 150 6 SCE
port 5 nsew signal input
rlabel locali s 352 176 386 337 6 SCE
port 5 nsew signal input
rlabel locali s 352 175 388 176 6 SCE
port 5 nsew signal input
rlabel locali s 352 174 389 175 6 SCE
port 5 nsew signal input
rlabel locali s 352 172 390 174 6 SCE
port 5 nsew signal input
rlabel locali s 352 171 391 172 6 SCE
port 5 nsew signal input
rlabel locali s 352 170 392 171 6 SCE
port 5 nsew signal input
rlabel locali s 352 168 393 170 6 SCE
port 5 nsew signal input
rlabel locali s 352 167 394 168 6 SCE
port 5 nsew signal input
rlabel locali s 352 164 395 167 6 SCE
port 5 nsew signal input
rlabel locali s 352 162 398 164 6 SCE
port 5 nsew signal input
rlabel locali s 352 157 402 162 6 SCE
port 5 nsew signal input
rlabel locali s 352 150 647 157 6 SCE
port 5 nsew signal input
rlabel locali s 19 195 89 325 6 CLK
port 6 nsew clock input
rlabel locali s 2037 17 2103 161 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1768 17 1802 139 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1540 17 1614 123 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1135 17 1209 117 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 749 17 789 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 391 17 457 89 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 103 17 169 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 2208 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 2208 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 2042 299 2103 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1768 325 1802 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1553 427 1614 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1177 367 1211 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 748 433 782 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 375 449 441 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 103 427 169 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 2208 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 2208 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2208 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 343100
string GDS_START 326098
<< end >>
