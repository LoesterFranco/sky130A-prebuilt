magic
tech sky130A
magscale 1 2
timestamp 1604502711
<< locali >>
rect 27 148 67 326
rect 305 84 349 349
rect 392 84 455 339
rect 489 129 555 323
rect 668 349 709 493
rect 668 307 811 349
rect 685 165 811 307
rect 652 128 811 165
rect 652 51 709 128
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 35 400 69 493
rect 103 439 169 527
rect 203 417 237 493
rect 311 451 445 527
rect 488 417 522 493
rect 568 439 634 527
rect 35 366 161 400
rect 127 265 161 366
rect 203 393 522 417
rect 203 383 633 393
rect 203 332 263 383
rect 488 359 633 383
rect 127 199 195 265
rect 127 117 161 199
rect 229 117 263 332
rect 19 17 85 93
rect 119 51 161 117
rect 219 51 263 117
rect 599 265 633 359
rect 743 383 810 527
rect 599 199 651 265
rect 552 17 618 93
rect 743 17 810 93
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
rlabel locali s 27 148 67 326 6 A_N
port 1 nsew signal input
rlabel locali s 305 84 349 349 6 B
port 2 nsew signal input
rlabel locali s 392 84 455 339 6 C
port 3 nsew signal input
rlabel locali s 489 129 555 323 6 D
port 4 nsew signal input
rlabel locali s 685 165 811 307 6 X
port 5 nsew signal output
rlabel locali s 668 349 709 493 6 X
port 5 nsew signal output
rlabel locali s 668 307 811 349 6 X
port 5 nsew signal output
rlabel locali s 652 128 811 165 6 X
port 5 nsew signal output
rlabel locali s 652 51 709 128 6 X
port 5 nsew signal output
rlabel metal1 s 0 -48 828 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 828 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3851210
string GDS_START 3842998
<< end >>
