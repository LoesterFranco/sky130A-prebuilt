magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 18 215 85 391
rect 513 391 563 493
rect 701 391 751 493
rect 513 357 751 391
rect 616 323 751 357
rect 616 289 898 323
rect 346 215 494 255
rect 821 181 898 289
rect 495 147 898 181
rect 495 58 571 147
rect 683 58 759 147
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 18 425 69 527
rect 129 265 163 493
rect 208 323 312 493
rect 413 367 469 527
rect 607 427 657 527
rect 795 359 845 527
rect 208 299 572 323
rect 268 289 572 299
rect 129 199 234 265
rect 129 181 179 199
rect 22 147 179 181
rect 268 181 312 289
rect 538 249 572 289
rect 538 215 760 249
rect 268 147 369 181
rect 22 53 84 147
rect 128 17 259 113
rect 293 61 369 147
rect 426 17 461 181
rect 615 17 649 110
rect 803 17 837 110
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
rlabel locali s 346 215 494 255 6 A
port 1 nsew signal input
rlabel locali s 18 215 85 391 6 B_N
port 2 nsew signal input
rlabel locali s 821 181 898 289 6 X
port 3 nsew signal output
rlabel locali s 701 391 751 493 6 X
port 3 nsew signal output
rlabel locali s 683 58 759 147 6 X
port 3 nsew signal output
rlabel locali s 616 323 751 357 6 X
port 3 nsew signal output
rlabel locali s 616 289 898 323 6 X
port 3 nsew signal output
rlabel locali s 513 391 563 493 6 X
port 3 nsew signal output
rlabel locali s 513 357 751 391 6 X
port 3 nsew signal output
rlabel locali s 495 147 898 181 6 X
port 3 nsew signal output
rlabel locali s 495 58 571 147 6 X
port 3 nsew signal output
rlabel metal1 s 0 -48 920 48 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 496 920 592 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 920 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 661866
string GDS_START 654706
<< end >>
