magic
tech sky130A
magscale 1 2
timestamp 1601050039
<< nwell >>
rect -38 261 2062 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 519 47 549 177
rect 603 47 633 177
rect 687 47 717 177
rect 771 47 801 177
rect 855 47 885 177
rect 939 47 969 177
rect 1023 47 1053 177
rect 1107 47 1137 177
rect 1295 47 1325 177
rect 1379 47 1409 177
rect 1463 47 1493 177
rect 1547 47 1577 177
rect 1631 47 1661 177
rect 1715 47 1745 177
rect 1799 47 1829 177
rect 1883 47 1913 177
<< pmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 519 297 549 497
rect 603 297 633 497
rect 687 297 717 497
rect 771 297 801 497
rect 855 297 885 497
rect 939 297 969 497
rect 1023 297 1053 497
rect 1107 297 1137 497
rect 1295 297 1325 497
rect 1379 297 1409 497
rect 1463 297 1493 497
rect 1547 297 1577 497
rect 1631 297 1661 497
rect 1715 297 1745 497
rect 1799 297 1829 497
rect 1883 297 1913 497
<< ndiff >>
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 161 163 177
rect 109 127 119 161
rect 153 127 163 161
rect 109 47 163 127
rect 193 93 247 177
rect 193 59 203 93
rect 237 59 247 93
rect 193 47 247 59
rect 277 161 331 177
rect 277 127 287 161
rect 321 127 331 161
rect 277 47 331 127
rect 361 93 413 177
rect 361 59 371 93
rect 405 59 413 93
rect 361 47 413 59
rect 467 161 519 177
rect 467 127 475 161
rect 509 127 519 161
rect 467 93 519 127
rect 467 59 475 93
rect 509 59 519 93
rect 467 47 519 59
rect 549 93 603 177
rect 549 59 559 93
rect 593 59 603 93
rect 549 47 603 59
rect 633 161 687 177
rect 633 127 643 161
rect 677 127 687 161
rect 633 93 687 127
rect 633 59 643 93
rect 677 59 687 93
rect 633 47 687 59
rect 717 93 771 177
rect 717 59 727 93
rect 761 59 771 93
rect 717 47 771 59
rect 801 161 855 177
rect 801 127 811 161
rect 845 127 855 161
rect 801 93 855 127
rect 801 59 811 93
rect 845 59 855 93
rect 801 47 855 59
rect 885 93 939 177
rect 885 59 895 93
rect 929 59 939 93
rect 885 47 939 59
rect 969 161 1023 177
rect 969 127 979 161
rect 1013 127 1023 161
rect 969 93 1023 127
rect 969 59 979 93
rect 1013 59 1023 93
rect 969 47 1023 59
rect 1053 93 1107 177
rect 1053 59 1063 93
rect 1097 59 1107 93
rect 1053 47 1107 59
rect 1137 161 1189 177
rect 1137 127 1147 161
rect 1181 127 1189 161
rect 1137 93 1189 127
rect 1137 59 1147 93
rect 1181 59 1189 93
rect 1137 47 1189 59
rect 1243 161 1295 177
rect 1243 127 1251 161
rect 1285 127 1295 161
rect 1243 93 1295 127
rect 1243 59 1251 93
rect 1285 59 1295 93
rect 1243 47 1295 59
rect 1325 93 1379 177
rect 1325 59 1335 93
rect 1369 59 1379 93
rect 1325 47 1379 59
rect 1409 161 1463 177
rect 1409 127 1419 161
rect 1453 127 1463 161
rect 1409 93 1463 127
rect 1409 59 1419 93
rect 1453 59 1463 93
rect 1409 47 1463 59
rect 1493 93 1547 177
rect 1493 59 1503 93
rect 1537 59 1547 93
rect 1493 47 1547 59
rect 1577 161 1631 177
rect 1577 127 1587 161
rect 1621 127 1631 161
rect 1577 93 1631 127
rect 1577 59 1587 93
rect 1621 59 1631 93
rect 1577 47 1631 59
rect 1661 93 1715 177
rect 1661 59 1671 93
rect 1705 59 1715 93
rect 1661 47 1715 59
rect 1745 161 1799 177
rect 1745 127 1755 161
rect 1789 127 1799 161
rect 1745 93 1799 127
rect 1745 59 1755 93
rect 1789 59 1799 93
rect 1745 47 1799 59
rect 1829 93 1883 177
rect 1829 59 1839 93
rect 1873 59 1883 93
rect 1829 47 1883 59
rect 1913 161 1969 177
rect 1913 127 1923 161
rect 1957 127 1969 161
rect 1913 93 1969 127
rect 1913 59 1923 93
rect 1957 59 1969 93
rect 1913 47 1969 59
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 485 163 497
rect 109 451 119 485
rect 153 451 163 485
rect 109 417 163 451
rect 109 383 119 417
rect 153 383 163 417
rect 109 349 163 383
rect 109 315 119 349
rect 153 315 163 349
rect 109 297 163 315
rect 193 485 247 497
rect 193 451 203 485
rect 237 451 247 485
rect 193 417 247 451
rect 193 383 203 417
rect 237 383 247 417
rect 193 297 247 383
rect 277 485 331 497
rect 277 451 287 485
rect 321 451 331 485
rect 277 417 331 451
rect 277 383 287 417
rect 321 383 331 417
rect 277 349 331 383
rect 277 315 287 349
rect 321 315 331 349
rect 277 297 331 315
rect 361 485 413 497
rect 361 451 371 485
rect 405 451 413 485
rect 361 417 413 451
rect 361 383 371 417
rect 405 383 413 417
rect 361 297 413 383
rect 467 475 519 497
rect 467 441 475 475
rect 509 441 519 475
rect 467 407 519 441
rect 467 373 475 407
rect 509 373 519 407
rect 467 297 519 373
rect 549 417 603 497
rect 549 383 559 417
rect 593 383 603 417
rect 549 349 603 383
rect 549 315 559 349
rect 593 315 603 349
rect 549 297 603 315
rect 633 475 687 497
rect 633 441 643 475
rect 677 441 687 475
rect 633 407 687 441
rect 633 373 643 407
rect 677 373 687 407
rect 633 297 687 373
rect 717 417 771 497
rect 717 383 727 417
rect 761 383 771 417
rect 717 349 771 383
rect 717 315 727 349
rect 761 315 771 349
rect 717 297 771 315
rect 801 475 855 497
rect 801 441 811 475
rect 845 441 855 475
rect 801 407 855 441
rect 801 373 811 407
rect 845 373 855 407
rect 801 339 855 373
rect 801 305 811 339
rect 845 305 855 339
rect 801 297 855 305
rect 885 475 939 497
rect 885 441 895 475
rect 929 441 939 475
rect 885 407 939 441
rect 885 373 895 407
rect 929 373 939 407
rect 885 297 939 373
rect 969 417 1023 497
rect 969 383 979 417
rect 1013 383 1023 417
rect 969 349 1023 383
rect 969 315 979 349
rect 1013 315 1023 349
rect 969 297 1023 315
rect 1053 475 1107 497
rect 1053 441 1063 475
rect 1097 441 1107 475
rect 1053 407 1107 441
rect 1053 373 1063 407
rect 1097 373 1107 407
rect 1053 297 1107 373
rect 1137 417 1189 497
rect 1137 383 1147 417
rect 1181 383 1189 417
rect 1137 349 1189 383
rect 1137 315 1147 349
rect 1181 315 1189 349
rect 1137 297 1189 315
rect 1243 417 1295 497
rect 1243 383 1251 417
rect 1285 383 1295 417
rect 1243 349 1295 383
rect 1243 315 1251 349
rect 1285 315 1295 349
rect 1243 297 1295 315
rect 1325 475 1379 497
rect 1325 441 1335 475
rect 1369 441 1379 475
rect 1325 407 1379 441
rect 1325 373 1335 407
rect 1369 373 1379 407
rect 1325 297 1379 373
rect 1409 417 1463 497
rect 1409 383 1419 417
rect 1453 383 1463 417
rect 1409 349 1463 383
rect 1409 315 1419 349
rect 1453 315 1463 349
rect 1409 297 1463 315
rect 1493 475 1547 497
rect 1493 441 1503 475
rect 1537 441 1547 475
rect 1493 407 1547 441
rect 1493 373 1503 407
rect 1537 373 1547 407
rect 1493 297 1547 373
rect 1577 485 1631 497
rect 1577 451 1587 485
rect 1621 451 1631 485
rect 1577 417 1631 451
rect 1577 383 1587 417
rect 1621 383 1631 417
rect 1577 349 1631 383
rect 1577 315 1587 349
rect 1621 315 1631 349
rect 1577 297 1631 315
rect 1661 485 1715 497
rect 1661 451 1671 485
rect 1705 451 1715 485
rect 1661 417 1715 451
rect 1661 383 1671 417
rect 1705 383 1715 417
rect 1661 297 1715 383
rect 1745 485 1799 497
rect 1745 451 1755 485
rect 1789 451 1799 485
rect 1745 417 1799 451
rect 1745 383 1755 417
rect 1789 383 1799 417
rect 1745 349 1799 383
rect 1745 315 1755 349
rect 1789 315 1799 349
rect 1745 297 1799 315
rect 1829 485 1883 497
rect 1829 451 1839 485
rect 1873 451 1883 485
rect 1829 417 1883 451
rect 1829 383 1839 417
rect 1873 383 1883 417
rect 1829 297 1883 383
rect 1913 485 1969 497
rect 1913 451 1923 485
rect 1957 451 1969 485
rect 1913 417 1969 451
rect 1913 383 1923 417
rect 1957 383 1969 417
rect 1913 349 1969 383
rect 1913 315 1923 349
rect 1957 315 1969 349
rect 1913 297 1969 315
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 119 127 153 161
rect 203 59 237 93
rect 287 127 321 161
rect 371 59 405 93
rect 475 127 509 161
rect 475 59 509 93
rect 559 59 593 93
rect 643 127 677 161
rect 643 59 677 93
rect 727 59 761 93
rect 811 127 845 161
rect 811 59 845 93
rect 895 59 929 93
rect 979 127 1013 161
rect 979 59 1013 93
rect 1063 59 1097 93
rect 1147 127 1181 161
rect 1147 59 1181 93
rect 1251 127 1285 161
rect 1251 59 1285 93
rect 1335 59 1369 93
rect 1419 127 1453 161
rect 1419 59 1453 93
rect 1503 59 1537 93
rect 1587 127 1621 161
rect 1587 59 1621 93
rect 1671 59 1705 93
rect 1755 127 1789 161
rect 1755 59 1789 93
rect 1839 59 1873 93
rect 1923 127 1957 161
rect 1923 59 1957 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 119 451 153 485
rect 119 383 153 417
rect 119 315 153 349
rect 203 451 237 485
rect 203 383 237 417
rect 287 451 321 485
rect 287 383 321 417
rect 287 315 321 349
rect 371 451 405 485
rect 371 383 405 417
rect 475 441 509 475
rect 475 373 509 407
rect 559 383 593 417
rect 559 315 593 349
rect 643 441 677 475
rect 643 373 677 407
rect 727 383 761 417
rect 727 315 761 349
rect 811 441 845 475
rect 811 373 845 407
rect 811 305 845 339
rect 895 441 929 475
rect 895 373 929 407
rect 979 383 1013 417
rect 979 315 1013 349
rect 1063 441 1097 475
rect 1063 373 1097 407
rect 1147 383 1181 417
rect 1147 315 1181 349
rect 1251 383 1285 417
rect 1251 315 1285 349
rect 1335 441 1369 475
rect 1335 373 1369 407
rect 1419 383 1453 417
rect 1419 315 1453 349
rect 1503 441 1537 475
rect 1503 373 1537 407
rect 1587 451 1621 485
rect 1587 383 1621 417
rect 1587 315 1621 349
rect 1671 451 1705 485
rect 1671 383 1705 417
rect 1755 451 1789 485
rect 1755 383 1789 417
rect 1755 315 1789 349
rect 1839 451 1873 485
rect 1839 383 1873 417
rect 1923 451 1957 485
rect 1923 383 1957 417
rect 1923 315 1957 349
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 519 497 549 523
rect 603 497 633 523
rect 687 497 717 523
rect 771 497 801 523
rect 855 497 885 523
rect 939 497 969 523
rect 1023 497 1053 523
rect 1107 497 1137 523
rect 1295 497 1325 523
rect 1379 497 1409 523
rect 1463 497 1493 523
rect 1547 497 1577 523
rect 1631 497 1661 523
rect 1715 497 1745 523
rect 1799 497 1829 523
rect 1883 497 1913 523
rect 79 261 109 297
rect 21 259 109 261
rect 163 259 193 297
rect 247 259 277 297
rect 331 259 361 297
rect 519 265 549 297
rect 21 249 361 259
rect 21 215 38 249
rect 72 215 119 249
rect 153 215 203 249
rect 237 215 287 249
rect 321 215 361 249
rect 21 205 361 215
rect 21 203 109 205
rect 79 177 109 203
rect 163 177 193 205
rect 247 177 277 205
rect 331 177 361 205
rect 470 259 549 265
rect 603 259 633 297
rect 687 259 717 297
rect 771 259 801 297
rect 470 249 801 259
rect 470 215 486 249
rect 520 215 560 249
rect 594 215 643 249
rect 677 215 727 249
rect 761 215 801 249
rect 470 205 801 215
rect 470 199 549 205
rect 519 177 549 199
rect 603 177 633 205
rect 687 177 717 205
rect 771 177 801 205
rect 855 259 885 297
rect 939 259 969 297
rect 1023 259 1053 297
rect 1107 259 1137 297
rect 1295 259 1325 297
rect 1379 259 1409 297
rect 1463 259 1493 297
rect 1547 259 1577 297
rect 1631 259 1661 297
rect 1715 259 1745 297
rect 1799 259 1829 297
rect 1883 259 1913 297
rect 855 249 1203 259
rect 855 215 895 249
rect 929 215 978 249
rect 1012 215 1063 249
rect 1097 215 1146 249
rect 1180 215 1203 249
rect 855 205 1203 215
rect 1273 249 1588 259
rect 1273 215 1289 249
rect 1323 215 1377 249
rect 1411 215 1457 249
rect 1491 215 1538 249
rect 1572 215 1588 249
rect 1273 205 1588 215
rect 1631 249 1940 259
rect 1631 215 1647 249
rect 1681 215 1726 249
rect 1760 215 1802 249
rect 1836 215 1890 249
rect 1924 215 1940 249
rect 1631 205 1940 215
rect 855 177 885 205
rect 939 177 969 205
rect 1023 177 1053 205
rect 1107 177 1137 205
rect 1295 177 1325 205
rect 1379 177 1409 205
rect 1463 177 1493 205
rect 1547 177 1577 205
rect 1631 177 1661 205
rect 1715 177 1745 205
rect 1799 177 1829 205
rect 1883 177 1913 205
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 519 21 549 47
rect 603 21 633 47
rect 687 21 717 47
rect 771 21 801 47
rect 855 21 885 47
rect 939 21 969 47
rect 1023 21 1053 47
rect 1107 21 1137 47
rect 1295 21 1325 47
rect 1379 21 1409 47
rect 1463 21 1493 47
rect 1547 21 1577 47
rect 1631 21 1661 47
rect 1715 21 1745 47
rect 1799 21 1829 47
rect 1883 21 1913 47
<< polycont >>
rect 38 215 72 249
rect 119 215 153 249
rect 203 215 237 249
rect 287 215 321 249
rect 486 215 520 249
rect 560 215 594 249
rect 643 215 677 249
rect 727 215 761 249
rect 895 215 929 249
rect 978 215 1012 249
rect 1063 215 1097 249
rect 1146 215 1180 249
rect 1289 215 1323 249
rect 1377 215 1411 249
rect 1457 215 1491 249
rect 1538 215 1572 249
rect 1647 215 1681 249
rect 1726 215 1760 249
rect 1802 215 1836 249
rect 1890 215 1924 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 17 485 69 527
rect 17 451 35 485
rect 17 417 69 451
rect 17 383 35 417
rect 17 349 69 383
rect 17 315 35 349
rect 17 289 69 315
rect 103 485 169 493
rect 103 451 119 485
rect 153 451 169 485
rect 103 417 169 451
rect 103 383 119 417
rect 153 383 169 417
rect 103 349 169 383
rect 203 485 237 527
rect 203 417 237 451
rect 203 367 237 383
rect 271 485 337 493
rect 271 451 287 485
rect 321 451 337 485
rect 271 417 337 451
rect 271 383 287 417
rect 321 383 337 417
rect 103 315 119 349
rect 153 323 169 349
rect 271 349 337 383
rect 371 485 421 527
rect 405 451 421 485
rect 371 417 421 451
rect 405 383 421 417
rect 371 367 421 383
rect 459 475 845 493
rect 459 441 475 475
rect 509 459 643 475
rect 459 407 509 441
rect 677 459 811 475
rect 459 373 475 407
rect 459 357 509 373
rect 543 417 609 425
rect 543 383 559 417
rect 593 383 609 417
rect 271 323 287 349
rect 153 315 287 323
rect 321 323 337 349
rect 543 349 609 383
rect 643 407 677 441
rect 643 357 677 373
rect 711 417 777 425
rect 711 383 727 417
rect 761 383 777 417
rect 543 323 559 349
rect 321 315 559 323
rect 593 323 609 349
rect 711 349 777 383
rect 711 323 727 349
rect 593 315 727 323
rect 761 315 777 349
rect 103 289 777 315
rect 811 407 845 441
rect 811 339 845 373
rect 879 475 1537 493
rect 879 441 895 475
rect 929 459 1063 475
rect 879 407 929 441
rect 1097 459 1335 475
rect 879 373 895 407
rect 879 357 929 373
rect 963 417 1029 425
rect 963 383 979 417
rect 1013 383 1029 417
rect 963 349 1029 383
rect 1063 407 1097 441
rect 1369 459 1503 475
rect 1063 357 1097 373
rect 1131 417 1197 425
rect 1131 383 1147 417
rect 1181 383 1197 417
rect 963 323 979 349
rect 845 315 979 323
rect 1013 323 1029 349
rect 1131 349 1197 383
rect 1131 323 1147 349
rect 1013 315 1147 323
rect 1181 315 1197 349
rect 845 305 1197 315
rect 811 289 1197 305
rect 1235 417 1301 425
rect 1235 383 1251 417
rect 1285 383 1301 417
rect 1235 349 1301 383
rect 1335 407 1369 441
rect 1335 357 1369 373
rect 1403 417 1469 425
rect 1403 383 1419 417
rect 1453 383 1469 417
rect 1235 315 1251 349
rect 1285 323 1301 349
rect 1403 349 1469 383
rect 1503 407 1537 441
rect 1503 357 1537 373
rect 1571 485 1637 493
rect 1571 451 1587 485
rect 1621 451 1637 485
rect 1571 417 1637 451
rect 1571 383 1587 417
rect 1621 383 1637 417
rect 1403 323 1419 349
rect 1285 315 1419 323
rect 1453 323 1469 349
rect 1571 349 1637 383
rect 1671 485 1705 527
rect 1671 417 1705 451
rect 1671 367 1705 383
rect 1739 485 1805 493
rect 1739 451 1755 485
rect 1789 451 1805 485
rect 1739 417 1805 451
rect 1739 383 1755 417
rect 1789 383 1805 417
rect 1571 323 1587 349
rect 1453 315 1587 323
rect 1621 323 1637 349
rect 1739 349 1805 383
rect 1839 485 1873 527
rect 1839 417 1873 451
rect 1839 367 1873 383
rect 1907 485 1973 493
rect 1907 451 1923 485
rect 1957 451 1973 485
rect 1907 417 1973 451
rect 1907 383 1923 417
rect 1957 383 1973 417
rect 1739 323 1755 349
rect 1621 315 1755 323
rect 1789 323 1805 349
rect 1907 349 1973 383
rect 1907 323 1923 349
rect 1789 315 1923 323
rect 1957 315 1973 349
rect 1235 289 1973 315
rect 21 249 340 255
rect 21 215 38 249
rect 72 215 119 249
rect 153 215 203 249
rect 237 215 287 249
rect 321 215 340 249
rect 374 181 432 289
rect 470 249 804 255
rect 470 215 486 249
rect 520 215 560 249
rect 594 215 643 249
rect 677 215 727 249
rect 761 215 804 249
rect 862 249 1196 255
rect 862 215 895 249
rect 929 215 978 249
rect 1012 215 1063 249
rect 1097 215 1146 249
rect 1180 215 1196 249
rect 1234 249 1588 255
rect 1234 215 1289 249
rect 1323 215 1377 249
rect 1411 215 1457 249
rect 1491 215 1538 249
rect 1572 215 1588 249
rect 1631 249 2007 255
rect 1631 215 1647 249
rect 1681 215 1726 249
rect 1760 215 1802 249
rect 1836 215 1890 249
rect 1924 215 2007 249
rect 17 161 69 181
rect 17 127 35 161
rect 103 161 432 181
rect 103 127 119 161
rect 153 127 287 161
rect 321 127 432 161
rect 470 161 1973 181
rect 470 127 475 161
rect 509 147 643 161
rect 509 127 525 147
rect 17 93 69 127
rect 470 93 525 127
rect 627 127 643 147
rect 677 147 811 161
rect 677 127 693 147
rect 17 59 35 93
rect 69 59 203 93
rect 237 59 371 93
rect 405 59 475 93
rect 509 59 525 93
rect 17 51 525 59
rect 559 93 593 109
rect 559 17 593 59
rect 627 93 693 127
rect 795 127 811 147
rect 845 147 979 161
rect 845 127 861 147
rect 627 59 643 93
rect 677 59 693 93
rect 627 51 693 59
rect 727 93 761 109
rect 727 17 761 59
rect 795 93 861 127
rect 963 127 979 147
rect 1013 147 1147 161
rect 1013 127 1029 147
rect 795 59 811 93
rect 845 59 861 93
rect 795 51 861 59
rect 895 93 929 109
rect 895 17 929 59
rect 963 93 1029 127
rect 1131 127 1147 147
rect 1181 147 1251 161
rect 1181 127 1197 147
rect 963 59 979 93
rect 1013 59 1029 93
rect 963 51 1029 59
rect 1063 93 1097 109
rect 1063 17 1097 59
rect 1131 93 1197 127
rect 1131 59 1147 93
rect 1181 59 1197 93
rect 1131 51 1197 59
rect 1235 127 1251 147
rect 1285 147 1419 161
rect 1285 127 1301 147
rect 1235 93 1301 127
rect 1403 127 1419 147
rect 1453 147 1587 161
rect 1453 127 1469 147
rect 1235 59 1251 93
rect 1285 59 1301 93
rect 1235 52 1301 59
rect 1335 93 1369 109
rect 1335 17 1369 59
rect 1403 93 1469 127
rect 1571 127 1587 147
rect 1621 147 1755 161
rect 1621 127 1637 147
rect 1403 59 1419 93
rect 1453 59 1469 93
rect 1403 52 1469 59
rect 1503 93 1537 109
rect 1503 17 1537 59
rect 1571 93 1637 127
rect 1739 127 1755 147
rect 1789 147 1923 161
rect 1789 127 1805 147
rect 1571 59 1587 93
rect 1621 59 1637 93
rect 1571 52 1637 59
rect 1671 93 1705 109
rect 1671 17 1705 59
rect 1739 93 1805 127
rect 1907 127 1923 147
rect 1957 127 1973 161
rect 1739 59 1755 93
rect 1789 59 1805 93
rect 1739 52 1805 59
rect 1839 93 1873 109
rect 1839 17 1873 59
rect 1907 93 1973 127
rect 1907 59 1923 93
rect 1957 59 1973 93
rect 1907 52 1973 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
<< metal1 >>
rect 0 561 2024 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 0 496 2024 527
rect 0 17 2024 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
rect 0 -48 2024 -17
<< labels >>
flabel corelocali s 1970 221 2004 255 0 FreeSans 250 0 0 0 A1
port 1 nsew
flabel corelocali s 1878 221 1912 255 0 FreeSans 250 0 0 0 A1
port 1 nsew
flabel corelocali s 1786 221 1820 255 0 FreeSans 250 0 0 0 A1
port 1 nsew
flabel corelocali s 1694 221 1728 255 0 FreeSans 250 0 0 0 A1
port 1 nsew
flabel corelocali s 1510 221 1544 255 0 FreeSans 250 0 0 0 A2
port 2 nsew
flabel corelocali s 1418 221 1452 255 0 FreeSans 250 0 0 0 A2
port 2 nsew
flabel corelocali s 1326 221 1360 255 0 FreeSans 250 0 0 0 A2
port 2 nsew
flabel corelocali s 1234 221 1268 255 0 FreeSans 250 0 0 0 A2
port 2 nsew
flabel corelocali s 1138 221 1172 255 0 FreeSans 250 0 0 0 A3
port 3 nsew
flabel corelocali s 1046 221 1080 255 0 FreeSans 250 0 0 0 A3
port 3 nsew
flabel corelocali s 954 221 988 255 0 FreeSans 250 0 0 0 A3
port 3 nsew
flabel corelocali s 862 221 896 255 0 FreeSans 250 0 0 0 A3
port 3 nsew
flabel corelocali s 770 221 804 255 0 FreeSans 250 0 0 0 A4
port 4 nsew
flabel corelocali s 678 221 712 255 0 FreeSans 250 0 0 0 A4
port 4 nsew
flabel corelocali s 586 221 620 255 0 FreeSans 250 0 0 0 A4
port 4 nsew
flabel corelocali s 494 221 528 255 0 FreeSans 250 0 0 0 A4
port 4 nsew
flabel corelocali s 398 153 432 187 0 FreeSans 250 0 0 0 Y
port 10 nsew
flabel corelocali s 398 221 432 255 0 FreeSans 250 0 0 0 Y
port 10 nsew
flabel corelocali s 398 289 432 323 0 FreeSans 250 0 0 0 Y
port 10 nsew
flabel corelocali s 306 289 340 323 0 FreeSans 250 0 0 0 Y
port 10 nsew
flabel corelocali s 214 289 248 323 0 FreeSans 250 0 0 0 Y
port 10 nsew
flabel corelocali s 122 289 156 323 0 FreeSans 250 0 0 0 Y
port 10 nsew
flabel corelocali s 306 221 340 255 0 FreeSans 250 0 0 0 B1
port 5 nsew
flabel corelocali s 214 221 248 255 0 FreeSans 250 0 0 0 B1
port 5 nsew
flabel corelocali s 122 221 156 255 0 FreeSans 250 0 0 0 B1
port 5 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 250 0 0 0 B1
port 5 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew
rlabel comment s 0 0 0 0 4 o41ai_4
<< properties >>
string FIXED_BBOX 0 0 2024 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 990850
string GDS_START 972792
string path 0.000 0.000 10.120 0.000 
<< end >>
