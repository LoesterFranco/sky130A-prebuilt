magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 28 -17 62 17
<< scnmos >>
rect 94 47 124 177
rect 210 47 240 177
rect 304 47 334 177
rect 388 47 418 177
rect 504 47 534 177
rect 598 47 628 177
rect 692 47 722 177
rect 796 47 826 177
<< pmoshvt >>
rect 86 297 122 497
rect 202 297 238 497
rect 296 297 332 497
rect 390 297 426 497
rect 506 297 542 497
rect 600 297 636 497
rect 694 297 730 497
rect 788 297 824 497
<< ndiff >>
rect 32 101 94 177
rect 32 67 40 101
rect 74 67 94 101
rect 32 47 94 67
rect 124 115 210 177
rect 124 81 150 115
rect 184 81 210 115
rect 124 47 210 81
rect 240 97 304 177
rect 240 63 250 97
rect 284 63 304 97
rect 240 47 304 63
rect 334 115 388 177
rect 334 81 344 115
rect 378 81 388 115
rect 334 47 388 81
rect 418 97 504 177
rect 418 63 458 97
rect 492 63 504 97
rect 418 47 504 63
rect 534 114 598 177
rect 534 80 554 114
rect 588 80 598 114
rect 534 47 598 80
rect 628 95 692 177
rect 628 61 648 95
rect 682 61 692 95
rect 628 47 692 61
rect 722 163 796 177
rect 722 129 742 163
rect 776 129 796 163
rect 722 95 796 129
rect 722 61 742 95
rect 776 61 796 95
rect 722 47 796 61
rect 826 95 881 177
rect 826 61 836 95
rect 870 61 881 95
rect 826 47 881 61
<< pdiff >>
rect 32 485 86 497
rect 32 451 40 485
rect 74 451 86 485
rect 32 417 86 451
rect 32 383 40 417
rect 74 383 86 417
rect 32 349 86 383
rect 32 315 40 349
rect 74 315 86 349
rect 32 297 86 315
rect 122 297 202 497
rect 238 297 296 497
rect 332 297 390 497
rect 426 477 506 497
rect 426 443 449 477
rect 483 443 506 477
rect 426 409 506 443
rect 426 375 449 409
rect 483 375 506 409
rect 426 297 506 375
rect 542 477 600 497
rect 542 443 554 477
rect 588 443 600 477
rect 542 409 600 443
rect 542 375 554 409
rect 588 375 600 409
rect 542 341 600 375
rect 542 307 554 341
rect 588 307 600 341
rect 542 297 600 307
rect 636 477 694 497
rect 636 443 648 477
rect 682 443 694 477
rect 636 409 694 443
rect 636 375 648 409
rect 682 375 694 409
rect 636 297 694 375
rect 730 477 788 497
rect 730 443 742 477
rect 776 443 788 477
rect 730 409 788 443
rect 730 375 742 409
rect 776 375 788 409
rect 730 341 788 375
rect 730 307 742 341
rect 776 307 788 341
rect 730 297 788 307
rect 824 477 880 497
rect 824 443 836 477
rect 870 443 880 477
rect 824 409 880 443
rect 824 375 836 409
rect 870 375 880 409
rect 824 297 880 375
<< ndiffc >>
rect 40 67 74 101
rect 150 81 184 115
rect 250 63 284 97
rect 344 81 378 115
rect 458 63 492 97
rect 554 80 588 114
rect 648 61 682 95
rect 742 129 776 163
rect 742 61 776 95
rect 836 61 870 95
<< pdiffc >>
rect 40 451 74 485
rect 40 383 74 417
rect 40 315 74 349
rect 449 443 483 477
rect 449 375 483 409
rect 554 443 588 477
rect 554 375 588 409
rect 554 307 588 341
rect 648 443 682 477
rect 648 375 682 409
rect 742 443 776 477
rect 742 375 776 409
rect 742 307 776 341
rect 836 443 870 477
rect 836 375 870 409
<< poly >>
rect 86 497 122 523
rect 202 497 238 523
rect 296 497 332 523
rect 390 497 426 523
rect 506 497 542 523
rect 600 497 636 523
rect 694 497 730 523
rect 788 497 824 523
rect 86 282 122 297
rect 202 282 238 297
rect 296 282 332 297
rect 390 282 426 297
rect 506 282 542 297
rect 600 282 636 297
rect 694 282 730 297
rect 788 282 824 297
rect 84 265 124 282
rect 200 265 240 282
rect 294 265 334 282
rect 388 265 428 282
rect 504 265 544 282
rect 598 265 638 282
rect 692 265 732 282
rect 786 265 826 282
rect 30 249 124 265
rect 30 215 40 249
rect 74 215 124 249
rect 30 199 124 215
rect 176 249 240 265
rect 176 215 186 249
rect 220 215 240 249
rect 176 199 240 215
rect 282 249 346 265
rect 282 215 292 249
rect 326 215 346 249
rect 282 199 346 215
rect 388 249 452 265
rect 388 215 398 249
rect 432 215 452 249
rect 388 199 452 215
rect 504 249 826 265
rect 504 215 514 249
rect 548 215 592 249
rect 626 215 670 249
rect 704 215 748 249
rect 782 215 826 249
rect 504 199 826 215
rect 94 177 124 199
rect 210 177 240 199
rect 304 177 334 199
rect 388 177 418 199
rect 504 177 534 199
rect 598 177 628 199
rect 692 177 722 199
rect 796 177 826 199
rect 94 21 124 47
rect 210 21 240 47
rect 304 21 334 47
rect 388 21 418 47
rect 504 21 534 47
rect 598 21 628 47
rect 692 21 722 47
rect 796 21 826 47
<< polycont >>
rect 40 215 74 249
rect 186 215 220 249
rect 292 215 326 249
rect 398 215 432 249
rect 514 215 548 249
rect 592 215 626 249
rect 670 215 704 249
rect 748 215 782 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 23 485 90 490
rect 23 451 40 485
rect 74 451 90 485
rect 441 477 491 527
rect 23 417 90 451
rect 23 383 40 417
rect 74 383 90 417
rect 23 349 90 383
rect 23 315 40 349
rect 74 333 90 349
rect 74 315 152 333
rect 23 299 152 315
rect 17 249 74 265
rect 17 215 40 249
rect 17 151 74 215
rect 108 165 152 299
rect 186 324 266 475
rect 300 357 374 475
rect 441 443 449 477
rect 483 443 491 477
rect 441 409 491 443
rect 441 375 449 409
rect 483 375 491 409
rect 441 359 491 375
rect 546 477 596 493
rect 546 443 554 477
rect 588 443 596 477
rect 546 409 596 443
rect 546 375 554 409
rect 588 375 596 409
rect 186 249 220 324
rect 300 290 352 357
rect 546 341 596 375
rect 640 477 690 527
rect 640 443 648 477
rect 682 443 690 477
rect 640 409 690 443
rect 640 375 648 409
rect 682 375 690 409
rect 640 359 690 375
rect 734 477 784 493
rect 734 443 742 477
rect 776 443 784 477
rect 734 409 784 443
rect 734 375 742 409
rect 776 375 784 409
rect 186 199 220 215
rect 276 249 352 290
rect 276 215 292 249
rect 326 215 352 249
rect 276 199 352 215
rect 388 289 495 323
rect 546 307 554 341
rect 588 325 596 341
rect 734 341 784 375
rect 828 477 878 527
rect 828 443 836 477
rect 870 443 878 477
rect 828 409 878 443
rect 828 375 836 409
rect 870 375 878 409
rect 828 359 878 375
rect 734 325 742 341
rect 588 307 742 325
rect 776 325 784 341
rect 776 307 897 325
rect 546 291 897 307
rect 388 249 442 289
rect 388 215 398 249
rect 432 215 442 249
rect 388 199 442 215
rect 476 215 514 249
rect 548 215 592 249
rect 626 215 670 249
rect 704 215 748 249
rect 782 215 798 249
rect 476 165 510 215
rect 842 181 897 291
rect 108 131 510 165
rect 554 163 897 181
rect 554 145 742 163
rect 24 101 74 117
rect 24 67 40 101
rect 24 17 74 67
rect 150 115 184 131
rect 344 115 378 131
rect 150 61 184 81
rect 224 63 250 97
rect 284 63 300 97
rect 224 17 300 63
rect 554 114 604 145
rect 344 61 378 81
rect 432 63 458 97
rect 492 63 508 97
rect 432 17 508 63
rect 588 80 604 114
rect 716 129 742 145
rect 776 145 897 163
rect 776 129 792 145
rect 554 51 604 80
rect 648 95 682 111
rect 648 17 682 61
rect 716 95 792 129
rect 716 61 742 95
rect 776 61 792 95
rect 716 51 792 61
rect 836 95 870 111
rect 836 17 870 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel corelocali s 334 425 368 459 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel corelocali s 334 357 368 391 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel corelocali s 222 357 266 391 0 FreeSans 400 0 0 0 C
port 3 nsew
flabel corelocali s 436 289 470 323 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 222 425 266 459 0 FreeSans 400 0 0 0 C
port 3 nsew
flabel corelocali s 28 221 62 255 0 FreeSans 400 0 0 0 D
port 4 nsew
flabel corelocali s 844 153 878 187 0 FreeSans 400 0 0 0 X
port 9 nsew
flabel pwell s 28 -17 62 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 28 527 62 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 28 527 62 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
flabel metal1 s 28 -17 62 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
rlabel comment s 0 0 0 0 4 or4_4
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 513022
string GDS_START 505360
<< end >>
