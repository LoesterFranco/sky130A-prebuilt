magic
tech sky130A
magscale 1 2
timestamp 1601050082
<< locali >>
rect 123 424 189 547
rect 303 424 369 547
rect 503 424 569 547
rect 703 424 769 547
rect 123 390 1270 424
rect 25 270 359 356
rect 409 270 839 356
rect 889 270 1161 356
rect 480 226 1030 236
rect 1236 226 1270 390
rect 1347 270 1703 356
rect 1753 270 2087 356
rect 480 202 1270 226
rect 480 176 732 202
rect 480 119 546 176
rect 964 154 1270 202
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 23 581 869 615
rect 23 390 89 581
rect 229 458 263 581
rect 403 458 469 581
rect 603 458 669 581
rect 803 492 869 581
rect 921 526 987 649
rect 1021 492 1087 596
rect 1121 526 1187 649
rect 1221 492 1287 596
rect 1321 526 1387 649
rect 1421 492 1487 596
rect 803 458 1487 492
rect 1521 458 1587 649
rect 1421 424 1487 458
rect 1621 424 1687 596
rect 1721 458 1787 649
rect 1821 424 1887 596
rect 1921 458 1987 649
rect 2022 424 2088 596
rect 1421 390 2088 424
rect 23 202 444 236
rect 23 70 89 202
rect 123 17 189 168
rect 225 70 259 202
rect 295 17 361 168
rect 410 85 444 202
rect 580 85 646 142
rect 752 85 818 142
rect 410 51 818 85
rect 864 120 930 168
rect 1308 202 1987 236
rect 1308 170 1547 202
rect 1308 154 1374 170
rect 1567 120 1633 136
rect 864 70 1633 120
rect 1679 17 1745 168
rect 1781 70 1815 202
rect 1851 17 1917 168
rect 1953 70 1987 202
rect 2023 17 2089 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
<< metal1 >>
rect 0 683 2112 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 0 617 2112 649
rect 0 17 2112 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
rect 0 -49 2112 -17
<< labels >>
rlabel locali s 889 270 1161 356 6 A1
port 1 nsew signal input
rlabel locali s 1347 270 1703 356 6 A2
port 2 nsew signal input
rlabel locali s 1753 270 2087 356 6 A3
port 3 nsew signal input
rlabel locali s 409 270 839 356 6 B1
port 4 nsew signal input
rlabel locali s 25 270 359 356 6 B2
port 5 nsew signal input
rlabel locali s 1236 226 1270 390 6 Y
port 6 nsew signal output
rlabel locali s 964 154 1270 202 6 Y
port 6 nsew signal output
rlabel locali s 703 424 769 547 6 Y
port 6 nsew signal output
rlabel locali s 503 424 569 547 6 Y
port 6 nsew signal output
rlabel locali s 480 226 1030 236 6 Y
port 6 nsew signal output
rlabel locali s 480 202 1270 226 6 Y
port 6 nsew signal output
rlabel locali s 480 176 732 202 6 Y
port 6 nsew signal output
rlabel locali s 480 119 546 176 6 Y
port 6 nsew signal output
rlabel locali s 303 424 369 547 6 Y
port 6 nsew signal output
rlabel locali s 123 424 189 547 6 Y
port 6 nsew signal output
rlabel locali s 123 390 1270 424 6 Y
port 6 nsew signal output
rlabel metal1 s 0 -49 2112 49 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 617 2112 715 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2112 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3833182
string GDS_START 3815966
<< end >>
