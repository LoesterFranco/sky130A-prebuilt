magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 920 561
rect 115 359 165 527
rect 22 215 193 257
rect 227 215 528 257
rect 563 181 613 425
rect 843 308 893 527
rect 806 215 903 257
rect 18 17 73 181
rect 107 145 621 181
rect 107 51 173 145
rect 207 17 241 111
rect 275 51 341 145
rect 375 17 521 111
rect 555 51 621 145
rect 655 17 696 179
rect 843 17 901 165
rect 0 -17 920 17
<< obsli1 >>
rect 18 325 81 493
rect 199 325 249 493
rect 283 459 696 493
rect 283 359 333 459
rect 367 325 417 425
rect 18 291 417 325
rect 475 291 529 459
rect 647 291 696 459
rect 738 291 809 374
rect 738 257 772 291
rect 647 215 772 257
rect 738 181 772 215
rect 738 76 809 181
<< metal1 >>
rect 0 496 920 592
rect 0 -48 920 48
<< labels >>
rlabel locali s 22 215 193 257 6 A
port 1 nsew signal input
rlabel locali s 227 215 528 257 6 B
port 2 nsew signal input
rlabel locali s 806 215 903 257 6 C_N
port 3 nsew signal input
rlabel locali s 563 181 613 425 6 Y
port 4 nsew signal output
rlabel locali s 555 51 621 145 6 Y
port 4 nsew signal output
rlabel locali s 275 51 341 145 6 Y
port 4 nsew signal output
rlabel locali s 107 145 621 181 6 Y
port 4 nsew signal output
rlabel locali s 107 51 173 145 6 Y
port 4 nsew signal output
rlabel locali s 843 17 901 165 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 655 17 696 179 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 375 17 521 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 207 17 241 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 18 17 73 181 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 920 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 920 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 843 308 893 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 115 359 165 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 920 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 920 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 920 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1127922
string GDS_START 1120106
<< end >>
