magic
tech sky130A
magscale 1 2
timestamp 1604502729
<< locali >>
rect 25 200 103 436
rect 409 328 455 356
rect 359 262 455 328
rect 2207 394 2273 596
rect 2482 394 2548 596
rect 2207 360 2548 394
rect 2482 356 2548 360
rect 2482 322 2663 356
rect 2515 254 2663 322
rect 2515 226 2565 254
rect 2319 176 2565 226
rect 2319 73 2382 176
rect 2515 70 2565 176
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2688 683
rect 22 504 72 649
rect 112 504 178 596
rect 218 530 268 649
rect 401 536 467 649
rect 137 496 178 504
rect 606 502 672 551
rect 302 496 672 502
rect 137 468 672 496
rect 712 514 762 551
rect 880 548 946 649
rect 983 514 1036 551
rect 1166 549 1233 649
rect 712 480 1036 514
rect 137 462 336 468
rect 137 166 171 462
rect 606 446 672 468
rect 205 424 257 428
rect 205 390 223 424
rect 205 226 257 390
rect 291 362 361 428
rect 491 378 569 434
rect 606 412 759 446
rect 291 228 325 362
rect 491 344 691 378
rect 489 228 535 310
rect 291 194 535 228
rect 33 132 171 166
rect 33 74 99 132
rect 213 17 247 166
rect 291 70 375 194
rect 569 160 603 344
rect 638 312 691 344
rect 725 278 759 412
rect 409 17 475 160
rect 509 100 603 160
rect 637 244 759 278
rect 637 134 687 244
rect 793 210 827 480
rect 949 459 1036 480
rect 1079 481 1391 515
rect 1425 495 1682 561
rect 721 176 827 210
rect 861 210 914 421
rect 949 300 983 459
rect 1079 458 1145 481
rect 1017 390 1087 424
rect 1121 390 1127 424
rect 1017 334 1127 390
rect 1231 388 1323 447
rect 949 244 1197 300
rect 1231 210 1265 388
rect 1357 318 1391 481
rect 1299 252 1391 318
rect 861 176 1398 210
rect 721 134 787 176
rect 1147 144 1398 176
rect 1432 169 1466 495
rect 1548 269 1614 461
rect 1648 341 1682 495
rect 1716 489 1782 649
rect 1816 489 1896 581
rect 1930 489 1980 649
rect 1753 424 1828 455
rect 1753 390 1759 424
rect 1793 390 1828 424
rect 1753 384 1828 390
rect 1862 409 1896 489
rect 1862 375 1989 409
rect 1648 307 1921 341
rect 1869 275 1921 307
rect 1509 203 1655 269
rect 1689 241 1755 273
rect 1955 241 1989 375
rect 2023 326 2073 581
rect 2107 405 2173 649
rect 2307 428 2448 649
rect 2582 390 2648 649
rect 2023 292 2448 326
rect 1689 207 1989 241
rect 2112 260 2448 292
rect 861 108 1113 142
rect 1432 119 1587 169
rect 861 100 895 108
rect 509 66 895 100
rect 1079 85 1113 108
rect 1621 85 1655 203
rect 979 17 1045 74
rect 1079 51 1655 85
rect 1725 17 1791 169
rect 1900 77 1966 207
rect 2023 17 2078 226
rect 2112 70 2178 260
rect 2224 17 2282 226
rect 2416 17 2481 142
rect 2601 17 2667 220
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2688 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 223 390 257 424
rect 1087 390 1121 424
rect 1759 390 1793 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
<< metal1 >>
rect 0 683 2688 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2688 683
rect 0 617 2688 649
rect 211 424 269 430
rect 211 390 223 424
rect 257 421 269 424
rect 1075 424 1133 430
rect 1075 421 1087 424
rect 257 393 1087 421
rect 257 390 269 393
rect 211 384 269 390
rect 1075 390 1087 393
rect 1121 421 1133 424
rect 1747 424 1805 430
rect 1747 421 1759 424
rect 1121 393 1759 421
rect 1121 390 1133 393
rect 1075 384 1133 390
rect 1747 390 1759 393
rect 1793 390 1805 424
rect 1747 384 1805 390
rect 0 17 2688 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2688 17
rect 0 -49 2688 -17
<< labels >>
rlabel locali s 25 200 103 436 6 D
port 1 nsew signal input
rlabel locali s 2515 254 2663 322 6 Q
port 2 nsew signal output
rlabel locali s 2515 226 2565 254 6 Q
port 2 nsew signal output
rlabel locali s 2515 70 2565 176 6 Q
port 2 nsew signal output
rlabel locali s 2482 394 2548 596 6 Q
port 2 nsew signal output
rlabel locali s 2482 356 2548 360 6 Q
port 2 nsew signal output
rlabel locali s 2482 322 2663 356 6 Q
port 2 nsew signal output
rlabel locali s 2319 176 2565 226 6 Q
port 2 nsew signal output
rlabel locali s 2319 73 2382 176 6 Q
port 2 nsew signal output
rlabel locali s 2207 394 2273 596 6 Q
port 2 nsew signal output
rlabel locali s 2207 360 2548 394 6 Q
port 2 nsew signal output
rlabel metal1 s 1747 421 1805 430 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 1747 384 1805 393 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 1075 421 1133 430 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 1075 384 1133 393 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 211 421 269 430 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 211 393 1805 421 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 211 384 269 393 6 RESET_B
port 3 nsew signal input
rlabel locali s 409 328 455 356 6 CLK
port 4 nsew clock input
rlabel locali s 359 262 455 328 6 CLK
port 4 nsew clock input
rlabel metal1 s 0 -49 2688 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 617 2688 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2688 666
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 2926364
string GDS_START 2907590
<< end >>
