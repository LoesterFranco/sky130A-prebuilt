magic
tech sky130A
magscale 1 2
timestamp 1601050088
<< locali >>
rect 17 364 91 596
rect 17 226 51 364
rect 17 70 89 226
rect 193 238 263 310
rect 301 238 367 310
rect 409 238 475 310
rect 509 238 601 310
rect 658 242 743 310
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 125 412 203 649
rect 241 446 307 572
rect 360 480 426 649
rect 479 581 745 615
rect 479 446 545 581
rect 241 412 545 446
rect 579 378 645 547
rect 125 344 645 378
rect 679 364 745 581
rect 125 326 159 344
rect 85 260 159 326
rect 125 204 159 260
rect 125 170 576 204
rect 130 17 210 136
rect 440 86 576 170
rect 674 17 740 208
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel locali s 409 238 475 310 6 A1
port 1 nsew signal input
rlabel locali s 301 238 367 310 6 A2
port 2 nsew signal input
rlabel locali s 193 238 263 310 6 A3
port 3 nsew signal input
rlabel locali s 509 238 601 310 6 B1
port 4 nsew signal input
rlabel locali s 658 242 743 310 6 B2
port 5 nsew signal input
rlabel locali s 17 364 91 596 6 X
port 6 nsew signal output
rlabel locali s 17 226 51 364 6 X
port 6 nsew signal output
rlabel locali s 17 70 89 226 6 X
port 6 nsew signal output
rlabel metal1 s 0 -49 768 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 617 768 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3749166
string GDS_START 3742320
<< end >>
