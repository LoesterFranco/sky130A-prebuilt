magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 125 323 175 493
rect 313 391 363 493
rect 313 323 465 391
rect 869 357 1713 401
rect 869 323 913 357
rect 125 289 913 323
rect 947 289 1279 323
rect 18 215 380 255
rect 424 173 465 289
rect 947 255 985 289
rect 512 215 985 255
rect 1019 199 1167 255
rect 1203 215 1279 289
rect 1313 289 1864 323
rect 1313 215 1389 289
rect 1801 255 1864 289
rect 1425 215 1747 255
rect 1801 215 2027 255
rect 107 129 465 173
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 31 297 81 527
rect 219 365 269 527
rect 407 425 561 527
rect 605 391 655 493
rect 699 425 749 527
rect 793 453 1227 493
rect 793 391 835 453
rect 1271 435 1321 527
rect 1355 453 1799 493
rect 605 357 835 391
rect 1757 391 1799 453
rect 1843 425 1893 527
rect 1937 391 1987 493
rect 1757 357 1987 391
rect 23 95 73 179
rect 1937 289 1987 357
rect 2031 289 2081 527
rect 1203 164 2089 181
rect 503 147 2089 164
rect 503 129 1337 147
rect 23 51 1227 95
rect 1271 51 1337 129
rect 1449 145 1713 147
rect 1381 17 1415 111
rect 1449 51 1525 145
rect 1569 17 1603 111
rect 1637 51 1713 145
rect 1825 145 2089 147
rect 1757 17 1791 111
rect 1825 51 1901 145
rect 1945 17 1979 111
rect 2013 51 2089 145
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
<< metal1 >>
rect 0 561 2116 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 0 496 2116 527
rect 0 17 2116 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
rect 0 -48 2116 -17
<< labels >>
rlabel locali s 1801 255 1864 289 6 A1
port 1 nsew signal input
rlabel locali s 1801 215 2027 255 6 A1
port 1 nsew signal input
rlabel locali s 1313 289 1864 323 6 A1
port 1 nsew signal input
rlabel locali s 1313 215 1389 289 6 A1
port 1 nsew signal input
rlabel locali s 1425 215 1747 255 6 A2
port 2 nsew signal input
rlabel locali s 1203 215 1279 289 6 B1
port 3 nsew signal input
rlabel locali s 947 289 1279 323 6 B1
port 3 nsew signal input
rlabel locali s 947 255 985 289 6 B1
port 3 nsew signal input
rlabel locali s 512 215 985 255 6 B1
port 3 nsew signal input
rlabel locali s 1019 199 1167 255 6 B2
port 4 nsew signal input
rlabel locali s 18 215 380 255 6 C1
port 5 nsew signal input
rlabel locali s 869 357 1713 401 6 Y
port 6 nsew signal output
rlabel locali s 869 323 913 357 6 Y
port 6 nsew signal output
rlabel locali s 424 173 465 289 6 Y
port 6 nsew signal output
rlabel locali s 313 391 363 493 6 Y
port 6 nsew signal output
rlabel locali s 313 323 465 391 6 Y
port 6 nsew signal output
rlabel locali s 125 323 175 493 6 Y
port 6 nsew signal output
rlabel locali s 125 289 913 323 6 Y
port 6 nsew signal output
rlabel locali s 107 129 465 173 6 Y
port 6 nsew signal output
rlabel metal1 s 0 -48 2116 48 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 496 2116 592 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2116 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 905952
string GDS_START 891882
<< end >>
