magic
tech sky130A
magscale 1 2
timestamp 1604502710
<< nwell >>
rect -38 332 998 704
<< pwell >>
rect 0 0 960 49
<< scpmos >>
rect 84 368 120 592
rect 184 368 220 592
rect 274 368 310 592
rect 364 368 400 592
rect 566 368 602 592
rect 656 368 692 592
rect 746 368 782 592
rect 836 368 872 592
<< nmoslvt >>
rect 84 74 114 222
rect 190 74 220 222
rect 284 74 314 222
rect 384 74 414 222
rect 566 74 596 222
rect 660 74 690 222
rect 746 74 776 222
rect 846 74 876 222
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 169 190 222
rect 114 135 139 169
rect 173 135 190 169
rect 114 74 190 135
rect 220 152 284 222
rect 220 118 239 152
rect 273 118 284 152
rect 220 74 284 118
rect 314 169 384 222
rect 314 135 339 169
rect 373 135 384 169
rect 314 74 384 135
rect 414 210 566 222
rect 414 176 521 210
rect 555 176 566 210
rect 414 152 566 176
rect 414 118 425 152
rect 459 120 566 152
rect 459 118 521 120
rect 414 86 521 118
rect 555 86 566 120
rect 414 74 566 86
rect 596 142 660 222
rect 596 108 607 142
rect 641 108 660 142
rect 596 74 660 108
rect 690 210 746 222
rect 690 176 701 210
rect 735 176 746 210
rect 690 120 746 176
rect 690 86 701 120
rect 735 86 746 120
rect 690 74 746 86
rect 776 152 846 222
rect 776 118 801 152
rect 835 118 846 152
rect 776 74 846 118
rect 876 210 933 222
rect 876 176 887 210
rect 921 176 933 210
rect 876 120 933 176
rect 876 86 887 120
rect 921 86 933 120
rect 876 74 933 86
<< pdiff >>
rect 28 580 84 592
rect 28 546 40 580
rect 74 546 84 580
rect 28 510 84 546
rect 28 476 40 510
rect 74 476 84 510
rect 28 440 84 476
rect 28 406 40 440
rect 74 406 84 440
rect 28 368 84 406
rect 120 580 184 592
rect 120 546 130 580
rect 164 546 184 580
rect 120 508 184 546
rect 120 474 130 508
rect 164 474 184 508
rect 120 368 184 474
rect 220 580 274 592
rect 220 546 230 580
rect 264 546 274 580
rect 220 510 274 546
rect 220 476 230 510
rect 264 476 274 510
rect 220 440 274 476
rect 220 406 230 440
rect 264 406 274 440
rect 220 368 274 406
rect 310 531 364 592
rect 310 497 320 531
rect 354 497 364 531
rect 310 440 364 497
rect 310 406 320 440
rect 354 406 364 440
rect 310 368 364 406
rect 400 580 456 592
rect 400 546 410 580
rect 444 546 456 580
rect 400 492 456 546
rect 400 458 410 492
rect 444 458 456 492
rect 400 368 456 458
rect 510 580 566 592
rect 510 546 522 580
rect 556 546 566 580
rect 510 478 566 546
rect 510 444 522 478
rect 556 444 566 478
rect 510 368 566 444
rect 602 531 656 592
rect 602 497 612 531
rect 646 497 656 531
rect 602 414 656 497
rect 602 380 612 414
rect 646 380 656 414
rect 602 368 656 380
rect 692 580 746 592
rect 692 546 702 580
rect 736 546 746 580
rect 692 510 746 546
rect 692 476 702 510
rect 736 476 746 510
rect 692 440 746 476
rect 692 406 702 440
rect 736 406 746 440
rect 692 368 746 406
rect 782 580 836 592
rect 782 546 792 580
rect 826 546 836 580
rect 782 508 836 546
rect 782 474 792 508
rect 826 474 836 508
rect 782 368 836 474
rect 872 580 928 592
rect 872 546 882 580
rect 916 546 928 580
rect 872 510 928 546
rect 872 476 882 510
rect 916 476 928 510
rect 872 440 928 476
rect 872 406 882 440
rect 916 406 928 440
rect 872 368 928 406
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 139 135 173 169
rect 239 118 273 152
rect 339 135 373 169
rect 521 176 555 210
rect 425 118 459 152
rect 521 86 555 120
rect 607 108 641 142
rect 701 176 735 210
rect 701 86 735 120
rect 801 118 835 152
rect 887 176 921 210
rect 887 86 921 120
<< pdiffc >>
rect 40 546 74 580
rect 40 476 74 510
rect 40 406 74 440
rect 130 546 164 580
rect 130 474 164 508
rect 230 546 264 580
rect 230 476 264 510
rect 230 406 264 440
rect 320 497 354 531
rect 320 406 354 440
rect 410 546 444 580
rect 410 458 444 492
rect 522 546 556 580
rect 522 444 556 478
rect 612 497 646 531
rect 612 380 646 414
rect 702 546 736 580
rect 702 476 736 510
rect 702 406 736 440
rect 792 546 826 580
rect 792 474 826 508
rect 882 546 916 580
rect 882 476 916 510
rect 882 406 916 440
<< poly >>
rect 84 592 120 618
rect 184 592 220 618
rect 274 592 310 618
rect 364 592 400 618
rect 566 592 602 618
rect 656 592 692 618
rect 746 592 782 618
rect 836 592 872 618
rect 84 336 120 368
rect 184 336 220 368
rect 84 320 220 336
rect 84 286 100 320
rect 134 286 168 320
rect 202 286 220 320
rect 84 270 220 286
rect 274 336 310 368
rect 364 336 400 368
rect 274 320 400 336
rect 566 326 602 368
rect 656 326 692 368
rect 274 286 313 320
rect 347 300 400 320
rect 533 310 692 326
rect 347 286 414 300
rect 274 270 414 286
rect 84 222 114 270
rect 190 222 220 270
rect 284 222 314 270
rect 384 222 414 270
rect 533 276 549 310
rect 583 276 617 310
rect 651 276 692 310
rect 533 260 692 276
rect 746 336 782 368
rect 836 336 872 368
rect 746 320 916 336
rect 746 286 798 320
rect 832 286 866 320
rect 900 286 916 320
rect 746 270 916 286
rect 566 222 596 260
rect 660 222 690 260
rect 746 222 776 270
rect 846 222 876 270
rect 84 48 114 74
rect 190 48 220 74
rect 284 48 314 74
rect 384 48 414 74
rect 566 48 596 74
rect 660 48 690 74
rect 746 48 776 74
rect 846 48 876 74
<< polycont >>
rect 100 286 134 320
rect 168 286 202 320
rect 313 286 347 320
rect 549 276 583 310
rect 617 276 651 310
rect 798 286 832 320
rect 866 286 900 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 24 580 74 596
rect 24 546 40 580
rect 24 510 74 546
rect 24 476 40 510
rect 24 440 74 476
rect 114 580 180 649
rect 114 546 130 580
rect 164 546 180 580
rect 114 508 180 546
rect 114 474 130 508
rect 164 474 180 508
rect 114 458 180 474
rect 214 581 460 615
rect 214 580 280 581
rect 214 546 230 580
rect 264 546 280 580
rect 394 580 460 581
rect 214 510 280 546
rect 214 476 230 510
rect 264 476 280 510
rect 24 406 40 440
rect 214 440 280 476
rect 214 424 230 440
rect 74 406 230 424
rect 264 406 280 440
rect 24 390 280 406
rect 314 531 360 547
rect 314 497 320 531
rect 354 497 360 531
rect 314 440 360 497
rect 394 546 410 580
rect 444 546 460 580
rect 394 492 460 546
rect 394 458 410 492
rect 444 458 460 492
rect 506 581 736 615
rect 506 580 572 581
rect 506 546 522 580
rect 556 546 572 580
rect 702 580 736 581
rect 506 478 572 546
rect 314 406 320 440
rect 354 424 360 440
rect 506 444 522 478
rect 556 444 572 478
rect 506 428 572 444
rect 612 531 662 547
rect 646 497 662 531
rect 354 406 455 424
rect 314 394 455 406
rect 612 414 662 497
rect 314 390 612 394
rect 409 380 612 390
rect 646 380 662 414
rect 702 510 736 546
rect 702 440 736 476
rect 776 580 826 649
rect 776 546 792 580
rect 776 508 826 546
rect 776 474 792 508
rect 776 458 826 474
rect 866 580 932 596
rect 866 546 882 580
rect 916 546 932 580
rect 866 510 932 546
rect 866 476 882 510
rect 916 476 932 510
rect 866 440 932 476
rect 866 424 882 440
rect 736 406 882 424
rect 916 406 932 440
rect 702 390 932 406
rect 409 360 662 380
rect 25 320 263 356
rect 25 286 100 320
rect 134 286 168 320
rect 202 286 263 320
rect 25 270 263 286
rect 297 320 363 356
rect 297 286 313 320
rect 347 286 363 320
rect 297 270 363 286
rect 409 236 455 360
rect 697 326 743 356
rect 533 310 743 326
rect 533 276 549 310
rect 583 276 617 310
rect 651 278 743 310
rect 782 320 935 356
rect 782 286 798 320
rect 832 286 866 320
rect 900 286 935 320
rect 651 276 667 278
rect 533 260 667 276
rect 782 270 935 286
rect 23 210 89 226
rect 23 176 39 210
rect 73 176 89 210
rect 23 120 89 176
rect 23 86 39 120
rect 73 86 89 120
rect 123 202 455 236
rect 701 226 937 236
rect 491 210 937 226
rect 123 169 189 202
rect 123 135 139 169
rect 173 135 189 169
rect 323 169 389 202
rect 123 119 189 135
rect 223 152 289 168
rect 23 85 89 86
rect 223 118 239 152
rect 273 118 289 152
rect 323 135 339 169
rect 373 135 389 169
rect 491 176 521 210
rect 555 192 701 210
rect 555 176 557 192
rect 491 168 557 176
rect 323 119 389 135
rect 423 152 557 168
rect 735 202 887 210
rect 735 176 751 202
rect 223 85 289 118
rect 423 118 425 152
rect 459 120 557 152
rect 459 118 521 120
rect 423 86 521 118
rect 555 86 557 120
rect 423 85 557 86
rect 23 51 557 85
rect 591 142 657 158
rect 591 108 607 142
rect 641 108 657 142
rect 591 17 657 108
rect 701 120 751 176
rect 921 176 937 210
rect 735 86 751 120
rect 701 70 751 86
rect 785 152 851 168
rect 785 118 801 152
rect 835 118 851 152
rect 785 17 851 118
rect 887 120 937 176
rect 921 86 937 120
rect 887 70 937 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
rlabel comment s 0 0 0 0 4 o22ai_2
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 415 242 449 276 0 FreeSans 340 0 0 0 Y
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 960 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1259526
string GDS_START 1251096
<< end >>
