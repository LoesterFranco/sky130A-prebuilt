magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 119 367 173 527
rect 307 367 361 527
rect 495 367 549 527
rect 683 367 737 527
rect 871 367 925 527
rect 1059 297 1119 527
rect 28 215 248 255
rect 123 17 179 113
rect 301 17 361 113
rect 495 17 549 113
rect 683 17 737 113
rect 871 17 925 113
rect 1059 17 1109 177
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< obsli1 >>
rect 19 323 85 493
rect 207 323 273 493
rect 395 323 461 493
rect 583 323 649 493
rect 771 323 837 493
rect 959 323 1025 493
rect 19 289 319 323
rect 395 289 1025 323
rect 284 249 319 289
rect 858 255 1025 289
rect 284 215 809 249
rect 858 221 912 255
rect 946 221 984 255
rect 1018 221 1025 255
rect 284 181 319 215
rect 858 181 1025 221
rect 29 147 319 181
rect 395 147 1025 181
rect 29 51 89 147
rect 213 51 267 147
rect 395 51 461 147
rect 583 51 649 147
rect 771 51 837 147
rect 959 51 1025 147
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 912 221 946 255
rect 984 221 1018 255
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< via1 >>
rect 710 223 740 253
rect 774 223 804 253
<< obsm1 >>
rect 693 261 821 264
rect 693 255 1030 261
rect 693 253 912 255
rect 693 223 710 253
rect 740 223 774 253
rect 804 223 912 253
rect 693 221 912 223
rect 946 221 984 255
rect 1018 221 1030 255
rect 693 215 1030 221
rect 693 212 821 215
<< via2 >>
rect 697 253 737 258
rect 777 253 817 258
rect 697 223 710 253
rect 710 223 737 253
rect 777 223 804 253
rect 804 223 817 253
rect 697 218 737 223
rect 777 218 817 223
<< obsm2 >>
rect 689 258 825 275
rect 689 218 697 258
rect 737 253 777 258
rect 740 223 774 253
rect 737 218 777 223
rect 817 218 825 258
rect 689 201 825 218
<< obsm3 >>
rect 679 258 835 271
rect 679 218 697 258
rect 737 218 777 258
rect 817 218 835 258
rect 679 205 835 218
<< via3 >>
rect 697 218 737 258
rect 777 218 817 258
<< obsm4 >>
rect 274 334 830 372
rect 274 174 312 334
rect 472 174 632 334
rect 792 258 830 334
rect 817 218 830 258
rect 792 174 830 218
rect 274 136 830 174
<< via4 >>
rect 312 174 472 334
rect 632 258 792 334
rect 632 218 697 258
rect 697 218 737 258
rect 737 218 777 258
rect 777 218 792 258
rect 632 174 792 218
<< metal5 >>
rect 250 112 854 432
<< labels >>
rlabel locali s 28 215 248 255 6 A
port 1 nsew signal input
rlabel via4 s 632 174 792 334 6 X
port 2 nsew signal output
rlabel via4 s 312 174 472 334 6 X
port 2 nsew signal output
rlabel metal5 s 250 112 854 432 6 X
port 2 nsew signal output
rlabel metal1 s 0 -48 1196 48 8 VGND
port 3 nsew ground input
rlabel locali s 1059 17 1109 177 6 VGND
port 3 nsew ground input
rlabel locali s 871 17 925 113 6 VGND
port 3 nsew ground input
rlabel locali s 683 17 737 113 6 VGND
port 3 nsew ground input
rlabel locali s 495 17 549 113 6 VGND
port 3 nsew ground input
rlabel locali s 301 17 361 113 6 VGND
port 3 nsew ground input
rlabel locali s 123 17 179 113 6 VGND
port 3 nsew ground input
rlabel locali s 0 -17 1196 17 8 VGND
port 3 nsew ground input
rlabel metal1 s 0 496 1196 592 6 VPWR
port 4 nsew power input
rlabel locali s 1059 297 1119 527 6 VPWR
port 4 nsew power input
rlabel locali s 871 367 925 527 6 VPWR
port 4 nsew power input
rlabel locali s 683 367 737 527 6 VPWR
port 4 nsew power input
rlabel locali s 495 367 549 527 6 VPWR
port 4 nsew power input
rlabel locali s 307 367 361 527 6 VPWR
port 4 nsew power input
rlabel locali s 119 367 173 527 6 VPWR
port 4 nsew power input
rlabel locali s 0 527 1196 561 6 VPWR
port 4 nsew power input
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 156830
string GDS_START 146306
<< end >>
