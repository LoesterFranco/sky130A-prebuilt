magic
tech sky130A
magscale 1 2
timestamp 1601050082
<< locali >>
rect 340 405 416 471
rect 25 236 100 310
rect 382 356 416 405
rect 382 225 454 356
rect 1533 406 1614 596
rect 1580 226 1614 406
rect 1528 70 1614 226
rect 1832 364 1903 596
rect 1869 226 1903 364
rect 1828 70 1903 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 22 378 72 596
rect 112 412 162 649
rect 202 543 268 596
rect 311 577 377 649
rect 748 585 826 649
rect 860 581 1198 615
rect 411 551 658 577
rect 860 560 1030 581
rect 860 551 894 560
rect 411 543 894 551
rect 202 509 445 543
rect 624 517 894 543
rect 22 344 168 378
rect 202 363 287 509
rect 556 483 590 509
rect 450 409 522 475
rect 134 310 168 344
rect 23 180 89 202
rect 134 180 218 310
rect 253 297 348 363
rect 253 214 319 297
rect 488 248 522 409
rect 556 449 856 483
rect 556 316 590 449
rect 624 350 731 415
rect 556 282 663 316
rect 488 214 577 248
rect 23 146 509 180
rect 23 70 89 146
rect 125 17 201 112
rect 371 17 441 112
rect 475 85 509 146
rect 543 119 577 214
rect 613 119 663 282
rect 697 150 731 350
rect 804 326 856 449
rect 928 405 962 523
rect 890 371 962 405
rect 890 274 924 371
rect 996 337 1030 560
rect 765 237 924 274
rect 958 271 1030 337
rect 1064 423 1114 547
rect 1064 276 1098 423
rect 1164 389 1198 581
rect 1233 478 1299 649
rect 1342 444 1408 572
rect 1132 323 1198 389
rect 1246 372 1408 444
rect 1448 406 1498 649
rect 1246 338 1546 372
rect 1246 310 1312 338
rect 1360 276 1426 304
rect 1064 242 1426 276
rect 765 203 980 237
rect 1064 224 1118 242
rect 1360 238 1426 242
rect 1460 270 1546 338
rect 914 184 980 203
rect 1025 158 1118 224
rect 697 124 930 150
rect 697 116 1143 124
rect 697 85 731 116
rect 475 51 731 85
rect 796 17 862 82
rect 896 58 1143 116
rect 1216 17 1282 208
rect 1460 204 1494 270
rect 1328 170 1494 204
rect 1328 88 1394 170
rect 1428 17 1494 136
rect 1656 326 1691 540
rect 1731 364 1797 649
rect 1656 260 1835 326
rect 1656 125 1706 260
rect 1742 17 1792 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
<< metal1 >>
rect 0 683 1920 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 0 617 1920 649
rect 0 17 1920 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
rect 0 -49 1920 -17
<< labels >>
rlabel locali s 382 356 416 405 6 D
port 1 nsew signal input
rlabel locali s 382 225 454 356 6 D
port 1 nsew signal input
rlabel locali s 340 405 416 471 6 D
port 1 nsew signal input
rlabel locali s 1580 226 1614 406 6 Q
port 2 nsew signal output
rlabel locali s 1533 406 1614 596 6 Q
port 2 nsew signal output
rlabel locali s 1528 70 1614 226 6 Q
port 2 nsew signal output
rlabel locali s 1869 226 1903 364 6 Q_N
port 3 nsew signal output
rlabel locali s 1832 364 1903 596 6 Q_N
port 3 nsew signal output
rlabel locali s 1828 70 1903 226 6 Q_N
port 3 nsew signal output
rlabel locali s 25 236 100 310 6 CLK
port 4 nsew clock input
rlabel metal1 s 0 -49 1920 49 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1920 715 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1920 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2696264
string GDS_START 2681298
<< end >>
