magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 18 195 88 325
rect 291 333 356 490
rect 291 123 395 333
rect 1913 325 1971 493
rect 2101 325 2151 493
rect 1913 291 2281 325
rect 2199 181 2281 291
rect 1895 147 2281 181
rect 1895 51 1971 147
rect 2083 51 2159 147
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2300 561
rect 18 393 69 493
rect 103 427 179 527
rect 18 359 178 393
rect 132 161 178 359
rect 18 127 178 161
rect 18 69 69 127
rect 103 17 179 93
rect 223 69 257 493
rect 390 435 440 527
rect 484 427 534 493
rect 587 427 733 493
rect 484 401 518 427
rect 429 367 518 401
rect 429 95 463 367
rect 552 315 655 393
rect 507 153 587 277
rect 621 197 655 315
rect 699 271 733 427
rect 767 407 801 475
rect 858 441 924 527
rect 968 407 1002 475
rect 1061 435 1145 527
rect 767 373 1002 407
rect 1189 401 1223 493
rect 1270 425 1494 493
rect 1528 435 1578 527
rect 1101 367 1223 401
rect 1101 339 1135 367
rect 805 305 1135 339
rect 1294 333 1406 391
rect 699 237 1057 271
rect 621 153 702 197
rect 736 95 770 237
rect 835 187 989 203
rect 1023 201 1057 237
rect 835 153 857 187
rect 891 153 929 187
rect 963 153 989 187
rect 1101 167 1135 305
rect 329 17 395 89
rect 429 61 538 95
rect 589 61 770 95
rect 965 17 1031 109
rect 1073 89 1135 167
rect 1183 331 1406 333
rect 1450 349 1494 425
rect 1622 417 1656 475
rect 1692 451 1768 527
rect 1622 383 1792 417
rect 1183 299 1338 331
rect 1450 315 1724 349
rect 1183 141 1225 299
rect 1450 297 1494 315
rect 1259 141 1349 265
rect 1393 263 1494 297
rect 1393 107 1427 263
rect 1561 250 1679 281
rect 1758 259 1792 383
rect 1827 315 1861 527
rect 2015 359 2049 527
rect 2203 359 2237 527
rect 1471 173 1525 229
rect 1561 216 1574 250
rect 1608 216 1679 250
rect 1561 207 1679 216
rect 1631 187 1679 207
rect 1471 139 1587 173
rect 1073 55 1153 89
rect 1207 51 1427 107
rect 1471 17 1519 105
rect 1553 93 1587 139
rect 1631 153 1633 187
rect 1667 153 1679 187
rect 1631 127 1679 153
rect 1723 257 1792 259
rect 1723 215 2159 257
rect 1723 164 1788 215
rect 1723 93 1787 164
rect 1553 59 1787 93
rect 1827 17 1861 179
rect 2015 17 2049 111
rect 2203 17 2237 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2300 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 857 153 891 187
rect 929 153 963 187
rect 1574 216 1608 250
rect 1633 153 1667 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
<< metal1 >>
rect 0 561 2300 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2300 561
rect 0 496 2300 527
rect 1562 250 1679 256
rect 1562 216 1574 250
rect 1608 216 1679 250
rect 835 187 985 193
rect 835 153 857 187
rect 891 153 929 187
rect 963 184 985 187
rect 1562 187 1679 216
rect 1562 184 1633 187
rect 963 156 1633 184
rect 963 153 985 156
rect 835 147 985 153
rect 1621 153 1633 156
rect 1667 153 1679 187
rect 1621 147 1679 153
rect 0 17 2300 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2300 17
rect 0 -48 2300 -17
<< obsm1 >>
rect 201 388 269 397
rect 609 388 667 397
rect 1293 388 1361 397
rect 201 360 1361 388
rect 201 351 269 360
rect 609 351 667 360
rect 1293 351 1361 360
rect 120 252 178 261
rect 507 252 565 261
rect 1293 252 1361 261
rect 120 224 1361 252
rect 120 215 178 224
rect 507 215 565 224
rect 1293 215 1361 224
<< labels >>
rlabel locali s 18 195 88 325 6 CLK
port 1 nsew signal input
rlabel locali s 291 333 356 490 6 D
port 2 nsew signal input
rlabel locali s 291 123 395 333 6 D
port 2 nsew signal input
rlabel locali s 2199 181 2281 291 6 Q
port 3 nsew signal output
rlabel locali s 2101 325 2151 493 6 Q
port 3 nsew signal output
rlabel locali s 2083 51 2159 147 6 Q
port 3 nsew signal output
rlabel locali s 1913 325 1971 493 6 Q
port 3 nsew signal output
rlabel locali s 1913 291 2281 325 6 Q
port 3 nsew signal output
rlabel locali s 1895 147 2281 181 6 Q
port 3 nsew signal output
rlabel locali s 1895 51 1971 147 6 Q
port 3 nsew signal output
rlabel metal1 s 1621 147 1679 156 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 1562 184 1679 256 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 835 184 985 193 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 835 156 1679 184 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 835 147 985 156 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 0 -48 2300 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 2300 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2300 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1877270
string GDS_START 1860492
<< end >>
