magic
tech sky130A
magscale 1 2
timestamp 1599588232
<< locali >>
rect 23 364 89 596
rect 23 188 71 364
rect 297 290 363 356
rect 405 290 471 356
rect 23 58 224 188
rect 505 88 579 310
rect 627 236 743 310
rect 777 236 843 310
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 129 364 179 649
rect 229 390 327 596
rect 361 424 427 596
rect 461 458 527 649
rect 567 424 633 596
rect 361 390 633 424
rect 667 412 733 649
rect 229 310 263 390
rect 567 378 633 390
rect 771 378 837 596
rect 115 256 263 310
rect 567 344 837 378
rect 115 222 424 256
rect 258 17 324 188
rect 358 70 424 222
rect 766 17 832 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel locali s 405 290 471 356 6 A1
port 1 nsew signal input
rlabel locali s 505 88 579 310 6 A2
port 2 nsew signal input
rlabel locali s 627 236 743 310 6 A3
port 3 nsew signal input
rlabel locali s 777 236 843 310 6 A4
port 4 nsew signal input
rlabel locali s 297 290 363 356 6 B1
port 5 nsew signal input
rlabel locali s 23 364 89 596 6 X
port 6 nsew signal output
rlabel locali s 23 188 71 364 6 X
port 6 nsew signal output
rlabel locali s 23 58 224 188 6 X
port 6 nsew signal output
rlabel metal1 s 0 -49 864 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 8 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 9 nsew power bidirectional
rlabel metal1 s 0 617 864 715 6 VPWR
port 10 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3901140
string GDS_START 3893096
<< end >>
