magic
tech sky130A
magscale 1 2
timestamp 1604502711
<< locali >>
rect 17 305 69 493
rect 17 162 52 305
rect 182 199 248 323
rect 282 199 340 275
rect 17 51 69 162
rect 520 271 616 331
rect 564 153 616 271
rect 656 153 708 331
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 103 447 169 527
rect 398 474 449 493
rect 221 440 449 474
rect 483 451 549 485
rect 221 395 255 440
rect 103 361 255 395
rect 398 413 449 440
rect 103 265 137 361
rect 308 343 342 381
rect 398 379 480 413
rect 86 199 137 265
rect 308 309 412 343
rect 378 165 412 309
rect 236 131 412 165
rect 446 174 480 379
rect 515 401 549 451
rect 583 435 633 527
rect 667 401 703 493
rect 515 367 703 401
rect 446 140 516 174
rect 103 17 189 106
rect 236 51 270 131
rect 304 17 448 97
rect 482 51 516 140
rect 631 17 711 119
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel locali s 182 199 248 323 6 A1_N
port 1 nsew signal input
rlabel locali s 282 199 340 275 6 A2_N
port 2 nsew signal input
rlabel locali s 656 153 708 331 6 B1
port 3 nsew signal input
rlabel locali s 564 153 616 271 6 B2
port 4 nsew signal input
rlabel locali s 520 271 616 331 6 B2
port 4 nsew signal input
rlabel locali s 17 305 69 493 6 X
port 5 nsew signal output
rlabel locali s 17 162 52 305 6 X
port 5 nsew signal output
rlabel locali s 17 51 69 162 6 X
port 5 nsew signal output
rlabel metal1 s 0 -48 736 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 736 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3455764
string GDS_START 3448596
<< end >>
