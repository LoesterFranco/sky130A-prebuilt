magic
tech sky130A
magscale 1 2
timestamp 1599588201
<< nwell >>
rect -38 261 1510 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 415 47 445 177
rect 499 47 529 177
rect 687 47 717 177
rect 771 47 801 177
rect 855 47 885 177
rect 939 47 969 177
rect 1023 47 1053 177
rect 1107 47 1137 177
rect 1191 47 1221 177
rect 1275 47 1305 177
<< pmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 415 297 445 497
rect 499 297 529 497
rect 687 297 717 497
rect 771 297 801 497
rect 855 297 885 497
rect 939 297 969 497
rect 1023 297 1053 497
rect 1107 297 1137 497
rect 1191 297 1221 497
rect 1275 297 1305 497
<< ndiff >>
rect 27 163 79 177
rect 27 129 35 163
rect 69 129 79 163
rect 27 95 79 129
rect 27 61 35 95
rect 69 61 79 95
rect 27 47 79 61
rect 109 163 163 177
rect 109 129 119 163
rect 153 129 163 163
rect 109 47 163 129
rect 193 163 247 177
rect 193 129 203 163
rect 237 129 247 163
rect 193 95 247 129
rect 193 61 203 95
rect 237 61 247 95
rect 193 47 247 61
rect 277 163 331 177
rect 277 129 287 163
rect 321 129 331 163
rect 277 47 331 129
rect 361 95 415 177
rect 361 61 371 95
rect 405 61 415 95
rect 361 47 415 61
rect 445 163 499 177
rect 445 129 455 163
rect 489 129 499 163
rect 445 47 499 129
rect 529 93 581 177
rect 529 59 539 93
rect 573 59 581 93
rect 529 47 581 59
rect 635 93 687 177
rect 635 59 643 93
rect 677 59 687 93
rect 635 47 687 59
rect 717 169 771 177
rect 717 135 727 169
rect 761 135 771 169
rect 717 101 771 135
rect 717 67 727 101
rect 761 67 771 101
rect 717 47 771 67
rect 801 95 855 177
rect 801 61 811 95
rect 845 61 855 95
rect 801 47 855 61
rect 885 163 939 177
rect 885 129 895 163
rect 929 129 939 163
rect 885 95 939 129
rect 885 61 895 95
rect 929 61 939 95
rect 885 47 939 61
rect 969 163 1023 177
rect 969 129 979 163
rect 1013 129 1023 163
rect 969 95 1023 129
rect 969 61 979 95
rect 1013 61 1023 95
rect 969 47 1023 61
rect 1053 163 1107 177
rect 1053 129 1063 163
rect 1097 129 1107 163
rect 1053 95 1107 129
rect 1053 61 1063 95
rect 1097 61 1107 95
rect 1053 47 1107 61
rect 1137 95 1191 177
rect 1137 61 1147 95
rect 1181 61 1191 95
rect 1137 47 1191 61
rect 1221 163 1275 177
rect 1221 129 1231 163
rect 1265 129 1275 163
rect 1221 95 1275 129
rect 1221 61 1231 95
rect 1265 61 1275 95
rect 1221 47 1275 61
rect 1305 95 1357 177
rect 1305 61 1315 95
rect 1349 61 1357 95
rect 1305 47 1357 61
<< pdiff >>
rect 27 483 79 497
rect 27 449 35 483
rect 69 449 79 483
rect 27 415 79 449
rect 27 381 35 415
rect 69 381 79 415
rect 27 347 79 381
rect 27 313 35 347
rect 69 313 79 347
rect 27 297 79 313
rect 109 477 163 497
rect 109 443 119 477
rect 153 443 163 477
rect 109 409 163 443
rect 109 375 119 409
rect 153 375 163 409
rect 109 341 163 375
rect 109 307 119 341
rect 153 307 163 341
rect 109 297 163 307
rect 193 477 247 497
rect 193 443 203 477
rect 237 443 247 477
rect 193 297 247 443
rect 277 477 331 497
rect 277 443 287 477
rect 321 443 331 477
rect 277 297 331 443
rect 361 409 415 497
rect 361 375 371 409
rect 405 375 415 409
rect 361 297 415 375
rect 445 477 499 497
rect 445 443 455 477
rect 489 443 499 477
rect 445 297 499 443
rect 529 477 687 497
rect 529 443 541 477
rect 575 443 643 477
rect 677 443 687 477
rect 529 297 687 443
rect 717 477 771 497
rect 717 443 727 477
rect 761 443 771 477
rect 717 297 771 443
rect 801 409 855 497
rect 801 375 811 409
rect 845 375 855 409
rect 801 297 855 375
rect 885 477 939 497
rect 885 443 895 477
rect 929 443 939 477
rect 885 297 939 443
rect 969 477 1023 497
rect 969 443 979 477
rect 1013 443 1023 477
rect 969 297 1023 443
rect 1053 477 1107 497
rect 1053 443 1063 477
rect 1097 443 1107 477
rect 1053 409 1107 443
rect 1053 375 1063 409
rect 1097 375 1107 409
rect 1053 297 1107 375
rect 1137 477 1191 497
rect 1137 443 1147 477
rect 1181 443 1191 477
rect 1137 297 1191 443
rect 1221 477 1275 497
rect 1221 443 1231 477
rect 1265 443 1275 477
rect 1221 409 1275 443
rect 1221 375 1231 409
rect 1265 375 1275 409
rect 1221 341 1275 375
rect 1221 307 1231 341
rect 1265 307 1275 341
rect 1221 297 1275 307
rect 1305 477 1357 497
rect 1305 443 1315 477
rect 1349 443 1357 477
rect 1305 409 1357 443
rect 1305 375 1315 409
rect 1349 375 1357 409
rect 1305 297 1357 375
<< ndiffc >>
rect 35 129 69 163
rect 35 61 69 95
rect 119 129 153 163
rect 203 129 237 163
rect 203 61 237 95
rect 287 129 321 163
rect 371 61 405 95
rect 455 129 489 163
rect 539 59 573 93
rect 643 59 677 93
rect 727 135 761 169
rect 727 67 761 101
rect 811 61 845 95
rect 895 129 929 163
rect 895 61 929 95
rect 979 129 1013 163
rect 979 61 1013 95
rect 1063 129 1097 163
rect 1063 61 1097 95
rect 1147 61 1181 95
rect 1231 129 1265 163
rect 1231 61 1265 95
rect 1315 61 1349 95
<< pdiffc >>
rect 35 449 69 483
rect 35 381 69 415
rect 35 313 69 347
rect 119 443 153 477
rect 119 375 153 409
rect 119 307 153 341
rect 203 443 237 477
rect 287 443 321 477
rect 371 375 405 409
rect 455 443 489 477
rect 541 443 575 477
rect 643 443 677 477
rect 727 443 761 477
rect 811 375 845 409
rect 895 443 929 477
rect 979 443 1013 477
rect 1063 443 1097 477
rect 1063 375 1097 409
rect 1147 443 1181 477
rect 1231 443 1265 477
rect 1231 375 1265 409
rect 1231 307 1265 341
rect 1315 443 1349 477
rect 1315 375 1349 409
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 415 497 445 523
rect 499 497 529 523
rect 687 497 717 523
rect 771 497 801 523
rect 855 497 885 523
rect 939 497 969 523
rect 1023 497 1053 523
rect 1107 497 1137 523
rect 1191 497 1221 523
rect 1275 497 1305 523
rect 79 265 109 297
rect 163 265 193 297
rect 247 265 277 297
rect 331 265 361 297
rect 415 265 445 297
rect 499 265 529 297
rect 687 265 717 297
rect 22 249 193 265
rect 22 215 38 249
rect 72 215 193 249
rect 22 199 193 215
rect 235 249 289 265
rect 235 215 245 249
rect 279 215 289 249
rect 235 199 289 215
rect 331 249 445 265
rect 331 215 371 249
rect 405 215 445 249
rect 331 199 445 215
rect 489 249 543 265
rect 489 215 499 249
rect 533 215 543 249
rect 489 199 543 215
rect 661 249 717 265
rect 661 215 671 249
rect 705 215 717 249
rect 661 199 717 215
rect 79 177 109 199
rect 163 177 193 199
rect 247 177 277 199
rect 331 177 361 199
rect 415 177 445 199
rect 499 177 529 199
rect 687 177 717 199
rect 771 265 801 297
rect 855 265 885 297
rect 939 265 969 297
rect 1023 265 1053 297
rect 1107 265 1137 297
rect 1191 265 1221 297
rect 1275 265 1305 297
rect 771 249 885 265
rect 771 215 811 249
rect 845 215 885 249
rect 771 199 885 215
rect 927 249 981 265
rect 927 215 937 249
rect 971 215 981 249
rect 927 199 981 215
rect 1023 249 1305 265
rect 1023 215 1063 249
rect 1097 215 1141 249
rect 1175 215 1231 249
rect 1265 215 1305 249
rect 1023 199 1305 215
rect 771 177 801 199
rect 855 177 885 199
rect 939 177 969 199
rect 1023 177 1053 199
rect 1107 177 1137 199
rect 1191 177 1221 199
rect 1275 177 1305 199
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 415 21 445 47
rect 499 21 529 47
rect 687 21 717 47
rect 771 21 801 47
rect 855 21 885 47
rect 939 21 969 47
rect 1023 21 1053 47
rect 1107 21 1137 47
rect 1191 21 1221 47
rect 1275 21 1305 47
<< polycont >>
rect 38 215 72 249
rect 245 215 279 249
rect 371 215 405 249
rect 499 215 533 249
rect 671 215 705 249
rect 811 215 845 249
rect 937 215 971 249
rect 1063 215 1097 249
rect 1141 215 1175 249
rect 1231 215 1265 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 29 483 79 527
rect 29 449 35 483
rect 69 449 79 483
rect 29 415 79 449
rect 29 381 35 415
rect 69 381 79 415
rect 29 347 79 381
rect 29 313 35 347
rect 69 313 79 347
rect 29 291 79 313
rect 113 477 163 493
rect 113 443 119 477
rect 153 443 163 477
rect 113 409 163 443
rect 197 477 247 527
rect 197 443 203 477
rect 237 443 247 477
rect 197 425 247 443
rect 281 477 499 493
rect 281 443 287 477
rect 321 459 455 477
rect 321 443 331 459
rect 281 425 331 443
rect 449 443 455 459
rect 489 443 499 477
rect 449 425 499 443
rect 533 477 685 527
rect 533 443 541 477
rect 575 443 643 477
rect 677 443 685 477
rect 533 425 685 443
rect 719 477 937 493
rect 719 443 727 477
rect 761 459 895 477
rect 761 443 769 459
rect 719 425 769 443
rect 887 443 895 459
rect 929 443 937 477
rect 887 425 937 443
rect 971 477 1021 527
rect 971 443 979 477
rect 1013 443 1021 477
rect 971 425 1021 443
rect 1063 477 1105 493
rect 1097 443 1105 477
rect 113 375 119 409
rect 153 391 163 409
rect 365 409 415 425
rect 365 391 371 409
rect 153 375 371 391
rect 405 391 415 409
rect 803 409 853 425
rect 803 391 811 409
rect 405 375 811 391
rect 845 391 853 409
rect 1063 409 1105 443
rect 1139 477 1189 527
rect 1139 443 1147 477
rect 1181 443 1189 477
rect 1139 425 1189 443
rect 1223 477 1273 493
rect 1223 443 1231 477
rect 1265 443 1273 477
rect 845 375 1029 391
rect 113 357 1029 375
rect 1097 391 1105 409
rect 1223 409 1273 443
rect 1097 375 1180 391
rect 1063 357 1180 375
rect 113 341 169 357
rect 113 307 119 341
rect 153 307 169 341
rect 995 323 1029 357
rect 1146 323 1180 357
rect 1223 375 1231 409
rect 1265 375 1273 409
rect 1223 341 1273 375
rect 1307 477 1357 527
rect 1307 443 1315 477
rect 1349 443 1357 477
rect 1307 409 1357 443
rect 1307 375 1315 409
rect 1349 375 1357 409
rect 1307 359 1357 375
rect 1223 323 1231 341
rect 113 289 169 307
rect 18 249 88 255
rect 18 215 38 249
rect 72 215 88 249
rect 17 163 69 179
rect 122 173 169 289
rect 205 289 549 323
rect 205 249 304 289
rect 205 215 245 249
rect 279 215 304 249
rect 338 249 449 255
rect 338 215 371 249
rect 405 215 449 249
rect 483 249 549 289
rect 483 215 499 249
rect 533 215 549 249
rect 601 289 955 323
rect 995 289 1075 323
rect 1146 307 1231 323
rect 1265 323 1273 341
rect 1265 307 1384 323
rect 1146 289 1384 307
rect 601 249 721 289
rect 905 255 955 289
rect 1041 255 1075 289
rect 601 215 671 249
rect 705 215 721 249
rect 755 249 871 255
rect 755 215 811 249
rect 845 215 871 249
rect 905 249 1007 255
rect 905 215 937 249
rect 971 215 1007 249
rect 1041 249 1281 255
rect 1041 215 1063 249
rect 1097 215 1141 249
rect 1175 215 1231 249
rect 1265 215 1281 249
rect 1315 181 1384 289
rect 17 129 35 163
rect 103 163 169 173
rect 103 129 119 163
rect 153 129 169 163
rect 203 163 237 181
rect 271 169 945 181
rect 271 163 727 169
rect 271 129 287 163
rect 321 129 455 163
rect 489 143 727 163
rect 489 129 507 143
rect 711 135 727 143
rect 761 163 945 169
rect 761 145 895 163
rect 761 135 777 145
rect 17 95 69 129
rect 203 95 237 129
rect 17 61 35 95
rect 69 61 203 95
rect 237 61 371 95
rect 405 93 591 95
rect 405 61 539 93
rect 17 59 539 61
rect 573 59 591 93
rect 17 51 591 59
rect 629 93 677 109
rect 629 59 643 93
rect 629 17 677 59
rect 711 101 777 135
rect 879 129 895 145
rect 929 129 945 163
rect 711 67 727 101
rect 761 67 777 101
rect 711 51 777 67
rect 811 95 845 111
rect 811 17 845 61
rect 879 95 945 129
rect 879 61 895 95
rect 929 61 945 95
rect 879 51 945 61
rect 979 163 1013 181
rect 979 95 1013 129
rect 979 17 1013 61
rect 1047 163 1384 181
rect 1047 129 1063 163
rect 1097 145 1231 163
rect 1097 129 1113 145
rect 1047 95 1113 129
rect 1215 129 1231 145
rect 1265 147 1384 163
rect 1265 129 1281 147
rect 1047 61 1063 95
rect 1097 61 1113 95
rect 1047 51 1113 61
rect 1147 95 1181 111
rect 1147 17 1181 61
rect 1215 95 1281 129
rect 1215 61 1231 95
rect 1265 61 1281 95
rect 1215 51 1281 61
rect 1315 95 1366 113
rect 1349 61 1366 95
rect 1315 17 1366 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< labels >>
flabel corelocali s 30 221 64 255 0 FreeSans 400 0 0 0 C1
port 5 nsew
flabel corelocali s 952 221 986 255 0 FreeSans 400 180 0 0 A1
port 1 nsew
flabel corelocali s 768 221 802 255 0 FreeSans 400 180 0 0 A2
port 2 nsew
flabel corelocali s 214 221 248 255 0 FreeSans 400 0 0 0 B1
port 3 nsew
flabel corelocali s 398 221 432 255 0 FreeSans 400 0 0 0 B2
port 4 nsew
flabel corelocali s 1320 289 1354 323 0 FreeSans 400 0 0 0 X
port 10 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew
rlabel comment s 0 0 0 0 4 o221a_4
<< properties >>
string FIXED_BBOX 0 0 1472 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1438068
string GDS_START 1427258
string path 0.000 0.000 7.360 0.000 
<< end >>
