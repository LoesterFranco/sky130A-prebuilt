magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 1326 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 101 47 131 177
rect 179 47 209 177
rect 263 47 293 177
rect 349 47 379 177
rect 465 47 495 177
rect 549 47 579 177
rect 653 47 683 177
rect 737 47 767 177
rect 841 47 871 177
rect 925 47 955 177
rect 1029 47 1059 177
rect 1113 47 1143 177
<< pmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 457 297 493 497
rect 551 297 587 497
rect 645 297 681 497
rect 739 297 775 497
rect 833 297 869 497
rect 927 297 963 497
rect 1021 297 1057 497
rect 1115 297 1151 497
<< ndiff >>
rect 27 161 101 177
rect 27 127 35 161
rect 69 127 101 161
rect 27 93 101 127
rect 27 59 35 93
rect 69 59 101 93
rect 27 47 101 59
rect 131 47 179 177
rect 209 161 263 177
rect 209 127 219 161
rect 253 127 263 161
rect 209 93 263 127
rect 209 59 219 93
rect 253 59 263 93
rect 209 47 263 59
rect 293 47 349 177
rect 379 89 465 177
rect 379 55 404 89
rect 438 55 465 89
rect 379 47 465 55
rect 495 129 549 177
rect 495 95 505 129
rect 539 95 549 129
rect 495 47 549 95
rect 579 105 653 177
rect 579 71 599 105
rect 633 71 653 105
rect 579 47 653 71
rect 683 169 737 177
rect 683 135 693 169
rect 727 135 737 169
rect 683 101 737 135
rect 683 67 693 101
rect 727 67 737 101
rect 683 47 737 67
rect 767 105 841 177
rect 767 71 787 105
rect 821 71 841 105
rect 767 47 841 71
rect 871 169 925 177
rect 871 135 881 169
rect 915 135 925 169
rect 871 101 925 135
rect 871 67 881 101
rect 915 67 925 101
rect 871 47 925 67
rect 955 105 1029 177
rect 955 71 975 105
rect 1009 71 1029 105
rect 955 47 1029 71
rect 1059 169 1113 177
rect 1059 135 1069 169
rect 1103 135 1113 169
rect 1059 101 1113 135
rect 1059 67 1069 101
rect 1103 67 1113 101
rect 1059 47 1113 67
rect 1143 105 1209 177
rect 1143 71 1163 105
rect 1197 71 1209 105
rect 1143 47 1209 71
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 297 81 383
rect 117 477 175 497
rect 117 443 129 477
rect 163 443 175 477
rect 117 409 175 443
rect 117 375 129 409
rect 163 375 175 409
rect 117 297 175 375
rect 211 485 269 497
rect 211 451 223 485
rect 257 451 269 485
rect 211 297 269 451
rect 305 477 363 497
rect 305 443 317 477
rect 351 443 363 477
rect 305 409 363 443
rect 305 375 317 409
rect 351 375 363 409
rect 305 297 363 375
rect 399 466 457 497
rect 399 432 411 466
rect 445 432 457 466
rect 399 297 457 432
rect 493 477 551 497
rect 493 443 505 477
rect 539 443 551 477
rect 493 409 551 443
rect 493 375 505 409
rect 539 375 551 409
rect 493 341 551 375
rect 493 307 505 341
rect 539 307 551 341
rect 493 297 551 307
rect 587 489 645 497
rect 587 455 599 489
rect 633 455 645 489
rect 587 395 645 455
rect 587 361 599 395
rect 633 361 645 395
rect 587 297 645 361
rect 681 477 739 497
rect 681 443 693 477
rect 727 443 739 477
rect 681 409 739 443
rect 681 375 693 409
rect 727 375 739 409
rect 681 341 739 375
rect 681 307 693 341
rect 727 307 739 341
rect 681 297 739 307
rect 775 489 833 497
rect 775 455 787 489
rect 821 455 833 489
rect 775 395 833 455
rect 775 361 787 395
rect 821 361 833 395
rect 775 297 833 361
rect 869 477 927 497
rect 869 443 881 477
rect 915 443 927 477
rect 869 409 927 443
rect 869 375 881 409
rect 915 375 927 409
rect 869 341 927 375
rect 869 307 881 341
rect 915 307 927 341
rect 869 297 927 307
rect 963 489 1021 497
rect 963 455 975 489
rect 1009 455 1021 489
rect 963 395 1021 455
rect 963 361 975 395
rect 1009 361 1021 395
rect 963 297 1021 361
rect 1057 477 1115 497
rect 1057 443 1069 477
rect 1103 443 1115 477
rect 1057 409 1115 443
rect 1057 375 1069 409
rect 1103 375 1115 409
rect 1057 341 1115 375
rect 1057 307 1069 341
rect 1103 307 1115 341
rect 1057 297 1115 307
rect 1151 489 1209 497
rect 1151 455 1163 489
rect 1197 455 1209 489
rect 1151 395 1209 455
rect 1151 361 1163 395
rect 1197 361 1209 395
rect 1151 297 1209 361
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 219 127 253 161
rect 219 59 253 93
rect 404 55 438 89
rect 505 95 539 129
rect 599 71 633 105
rect 693 135 727 169
rect 693 67 727 101
rect 787 71 821 105
rect 881 135 915 169
rect 881 67 915 101
rect 975 71 1009 105
rect 1069 135 1103 169
rect 1069 67 1103 101
rect 1163 71 1197 105
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 129 443 163 477
rect 129 375 163 409
rect 223 451 257 485
rect 317 443 351 477
rect 317 375 351 409
rect 411 432 445 466
rect 505 443 539 477
rect 505 375 539 409
rect 505 307 539 341
rect 599 455 633 489
rect 599 361 633 395
rect 693 443 727 477
rect 693 375 727 409
rect 693 307 727 341
rect 787 455 821 489
rect 787 361 821 395
rect 881 443 915 477
rect 881 375 915 409
rect 881 307 915 341
rect 975 455 1009 489
rect 975 361 1009 395
rect 1069 443 1103 477
rect 1069 375 1103 409
rect 1069 307 1103 341
rect 1163 455 1197 489
rect 1163 361 1197 395
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 457 497 493 523
rect 551 497 587 523
rect 645 497 681 523
rect 739 497 775 523
rect 833 497 869 523
rect 927 497 963 523
rect 1021 497 1057 523
rect 1115 497 1151 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 457 282 493 297
rect 551 282 587 297
rect 645 282 681 297
rect 739 282 775 297
rect 833 282 869 297
rect 927 282 963 297
rect 1021 282 1057 297
rect 1115 282 1151 297
rect 79 265 119 282
rect 173 265 213 282
rect 267 265 307 282
rect 361 265 401 282
rect 455 265 495 282
rect 549 265 589 282
rect 643 265 683 282
rect 737 265 777 282
rect 831 265 871 282
rect 925 265 965 282
rect 1019 265 1059 282
rect 1113 265 1153 282
rect 65 249 131 265
rect 65 215 81 249
rect 115 215 131 249
rect 65 199 131 215
rect 173 249 307 265
rect 173 215 189 249
rect 223 215 257 249
rect 291 215 307 249
rect 173 199 307 215
rect 349 249 409 265
rect 349 215 359 249
rect 393 215 409 249
rect 349 199 409 215
rect 455 249 1153 265
rect 455 215 471 249
rect 505 215 539 249
rect 573 215 607 249
rect 641 215 675 249
rect 709 215 743 249
rect 777 215 811 249
rect 845 215 879 249
rect 913 215 947 249
rect 981 215 1015 249
rect 1049 215 1153 249
rect 455 199 1153 215
rect 101 177 131 199
rect 179 177 209 199
rect 263 177 293 199
rect 349 177 379 199
rect 465 177 495 199
rect 549 177 579 199
rect 653 177 683 199
rect 737 177 767 199
rect 841 177 871 199
rect 925 177 955 199
rect 1029 177 1059 199
rect 1113 177 1143 199
rect 101 21 131 47
rect 179 21 209 47
rect 263 21 293 47
rect 349 21 379 47
rect 465 21 495 47
rect 549 21 579 47
rect 653 21 683 47
rect 737 21 767 47
rect 841 21 871 47
rect 925 21 955 47
rect 1029 21 1059 47
rect 1113 21 1143 47
<< polycont >>
rect 81 215 115 249
rect 189 215 223 249
rect 257 215 291 249
rect 359 215 393 249
rect 471 215 505 249
rect 539 215 573 249
rect 607 215 641 249
rect 675 215 709 249
rect 743 215 777 249
rect 811 215 845 249
rect 879 215 913 249
rect 947 215 981 249
rect 1015 215 1049 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 19 485 79 527
rect 19 451 35 485
rect 69 451 79 485
rect 19 417 79 451
rect 19 383 35 417
rect 69 383 79 417
rect 19 361 79 383
rect 113 477 173 493
rect 113 443 129 477
rect 163 443 173 477
rect 113 409 173 443
rect 207 485 273 527
rect 207 451 223 485
rect 257 451 273 485
rect 207 429 273 451
rect 307 477 361 493
rect 307 443 317 477
rect 351 443 361 477
rect 113 375 129 409
rect 163 395 173 409
rect 307 409 361 443
rect 395 466 461 527
rect 395 432 411 466
rect 445 432 461 466
rect 495 477 549 493
rect 495 443 505 477
rect 539 443 549 477
rect 307 395 317 409
rect 163 375 317 395
rect 351 395 361 409
rect 495 409 549 443
rect 351 375 461 395
rect 113 361 461 375
rect 87 293 377 327
rect 87 265 123 293
rect 17 249 123 265
rect 341 265 377 293
rect 17 215 81 249
rect 115 215 123 249
rect 17 199 123 215
rect 173 249 307 259
rect 173 215 189 249
rect 223 215 257 249
rect 291 215 307 249
rect 173 199 307 215
rect 341 249 393 265
rect 341 215 359 249
rect 341 199 393 215
rect 427 253 461 361
rect 495 375 505 409
rect 539 375 549 409
rect 495 341 549 375
rect 583 489 649 527
rect 583 455 599 489
rect 633 455 649 489
rect 583 395 649 455
rect 583 361 599 395
rect 633 361 649 395
rect 583 357 649 361
rect 683 477 737 493
rect 683 443 693 477
rect 727 443 737 477
rect 683 409 737 443
rect 683 375 693 409
rect 727 375 737 409
rect 495 307 505 341
rect 539 323 549 341
rect 683 341 737 375
rect 771 489 837 527
rect 771 455 787 489
rect 821 455 837 489
rect 771 395 837 455
rect 771 361 787 395
rect 821 361 837 395
rect 771 357 837 361
rect 871 477 925 493
rect 871 443 881 477
rect 915 443 925 477
rect 871 409 925 443
rect 871 375 881 409
rect 915 375 925 409
rect 683 323 693 341
rect 539 307 693 323
rect 727 323 737 341
rect 871 341 925 375
rect 959 489 1025 527
rect 959 455 975 489
rect 1009 455 1025 489
rect 959 395 1025 455
rect 959 361 975 395
rect 1009 361 1025 395
rect 959 357 1025 361
rect 1059 477 1113 493
rect 1059 443 1069 477
rect 1103 443 1113 477
rect 1059 409 1113 443
rect 1059 375 1069 409
rect 1103 375 1113 409
rect 871 323 881 341
rect 727 307 881 323
rect 915 323 925 341
rect 1059 341 1113 375
rect 1147 489 1213 527
rect 1147 455 1163 489
rect 1197 455 1213 489
rect 1147 395 1213 455
rect 1147 361 1163 395
rect 1197 361 1213 395
rect 1147 357 1213 361
rect 1059 323 1069 341
rect 915 307 1069 323
rect 1103 323 1113 341
rect 1103 307 1183 323
rect 495 289 1183 307
rect 427 249 1065 253
rect 427 215 471 249
rect 505 215 539 249
rect 573 215 607 249
rect 641 215 675 249
rect 709 215 743 249
rect 777 215 811 249
rect 845 215 879 249
rect 913 215 947 249
rect 981 215 1015 249
rect 1049 215 1065 249
rect 427 211 1065 215
rect 427 165 461 211
rect 1099 177 1183 289
rect 19 161 85 165
rect 19 127 35 161
rect 69 127 85 161
rect 19 93 85 127
rect 19 59 35 93
rect 69 59 85 93
rect 19 17 85 59
rect 203 161 461 165
rect 203 127 219 161
rect 253 131 461 161
rect 495 169 1183 177
rect 495 143 693 169
rect 253 127 269 131
rect 203 93 269 127
rect 495 129 549 143
rect 203 59 219 93
rect 253 59 269 93
rect 203 51 269 59
rect 388 89 454 97
rect 388 55 404 89
rect 438 55 454 89
rect 388 17 454 55
rect 495 95 505 129
rect 539 95 549 129
rect 683 135 693 143
rect 727 143 881 169
rect 727 135 737 143
rect 495 51 549 95
rect 583 105 649 109
rect 583 71 599 105
rect 633 71 649 105
rect 583 17 649 71
rect 683 101 737 135
rect 871 135 881 143
rect 915 143 1069 169
rect 915 135 925 143
rect 683 67 693 101
rect 727 67 737 101
rect 683 51 737 67
rect 771 105 837 109
rect 771 71 787 105
rect 821 71 837 105
rect 771 17 837 71
rect 871 101 925 135
rect 1059 135 1069 143
rect 1103 143 1183 169
rect 1103 135 1113 143
rect 871 67 881 101
rect 915 67 925 101
rect 871 51 925 67
rect 959 105 1025 109
rect 959 71 975 105
rect 1009 71 1025 105
rect 959 17 1025 71
rect 1059 101 1113 135
rect 1059 67 1069 101
rect 1103 67 1113 101
rect 1059 51 1113 67
rect 1147 105 1213 109
rect 1147 71 1163 105
rect 1197 71 1213 105
rect 1147 17 1213 71
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
flabel corelocali s 1133 221 1167 255 0 FreeSans 340 0 0 0 X
port 7 nsew
flabel corelocali s 29 221 63 255 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 213 221 247 255 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew
rlabel comment s 0 0 0 0 4 and2_8
<< properties >>
string FIXED_BBOX 0 0 1288 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3346668
string GDS_START 3336998
<< end >>
