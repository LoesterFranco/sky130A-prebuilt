magic
tech sky130A
magscale 1 2
timestamp 1599588238
<< locali >>
rect 501 424 551 547
rect 691 424 757 596
rect 501 404 757 424
rect 871 404 937 596
rect 501 390 937 404
rect 501 364 567 390
rect 723 370 937 390
rect 25 270 263 356
rect 313 270 455 356
rect 533 236 567 364
rect 601 270 689 356
rect 737 270 939 336
rect 873 236 939 270
rect 533 202 836 236
rect 770 122 836 202
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 24 424 74 596
rect 114 458 164 649
rect 204 424 270 596
rect 310 581 657 615
rect 310 458 344 581
rect 384 424 450 547
rect 24 390 450 424
rect 591 458 657 581
rect 797 438 831 649
rect 23 202 489 236
rect 23 70 89 202
rect 123 17 189 165
rect 223 70 289 202
rect 423 168 489 202
rect 323 17 389 165
rect 423 134 734 168
rect 423 70 489 134
rect 525 17 648 100
rect 684 85 734 134
rect 870 85 936 202
rect 684 51 936 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
rlabel locali s 25 270 263 356 6 A1
port 1 nsew signal input
rlabel locali s 313 270 455 356 6 A2
port 2 nsew signal input
rlabel locali s 601 270 689 356 6 A3
port 3 nsew signal input
rlabel locali s 873 236 939 270 6 B1
port 4 nsew signal input
rlabel locali s 737 270 939 336 6 B1
port 4 nsew signal input
rlabel locali s 871 404 937 596 6 Y
port 5 nsew signal output
rlabel locali s 770 122 836 202 6 Y
port 5 nsew signal output
rlabel locali s 723 370 937 390 6 Y
port 5 nsew signal output
rlabel locali s 691 424 757 596 6 Y
port 5 nsew signal output
rlabel locali s 533 236 567 364 6 Y
port 5 nsew signal output
rlabel locali s 533 202 836 236 6 Y
port 5 nsew signal output
rlabel locali s 501 424 551 547 6 Y
port 5 nsew signal output
rlabel locali s 501 404 757 424 6 Y
port 5 nsew signal output
rlabel locali s 501 390 937 404 6 Y
port 5 nsew signal output
rlabel locali s 501 364 567 390 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -49 960 49 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 617 960 715 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 823470
string GDS_START 814690
<< end >>
