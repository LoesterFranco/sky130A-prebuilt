magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 101 270 167 356
rect 759 364 847 596
rect 269 244 337 310
rect 303 196 337 244
rect 377 236 455 310
rect 491 196 557 310
rect 303 162 557 196
rect 813 226 847 364
rect 773 70 847 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 23 446 89 540
rect 130 480 196 649
rect 230 581 625 615
rect 230 446 264 581
rect 23 412 264 446
rect 23 390 89 412
rect 23 226 57 390
rect 413 378 479 547
rect 201 344 479 378
rect 23 108 89 226
rect 125 136 167 226
rect 201 204 235 344
rect 591 330 625 581
rect 659 364 725 649
rect 201 170 269 204
rect 125 17 201 136
rect 235 128 269 170
rect 591 264 671 330
rect 705 260 779 326
rect 705 230 739 260
rect 591 196 739 230
rect 591 128 625 196
rect 235 78 625 128
rect 659 17 725 162
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel locali s 377 236 455 310 6 A0
port 1 nsew signal input
rlabel locali s 491 196 557 310 6 A1
port 2 nsew signal input
rlabel locali s 303 196 337 244 6 A1
port 2 nsew signal input
rlabel locali s 303 162 557 196 6 A1
port 2 nsew signal input
rlabel locali s 269 244 337 310 6 A1
port 2 nsew signal input
rlabel locali s 101 270 167 356 6 S
port 3 nsew signal input
rlabel locali s 813 226 847 364 6 X
port 4 nsew signal output
rlabel locali s 773 70 847 226 6 X
port 4 nsew signal output
rlabel locali s 759 364 847 596 6 X
port 4 nsew signal output
rlabel metal1 s 0 -49 864 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 617 864 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1903020
string GDS_START 1896158
<< end >>
