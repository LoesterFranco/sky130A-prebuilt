magic
tech sky130A
magscale 1 2
timestamp 1604502697
<< nwell >>
rect -38 261 1326 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 123 47 153 177
rect 209 47 239 177
rect 305 47 335 177
rect 401 47 431 177
rect 497 47 527 177
rect 709 47 739 177
rect 803 47 833 177
rect 905 47 935 177
rect 981 47 1011 177
rect 1085 47 1115 177
rect 1169 47 1199 177
<< pmoshvt >>
rect 115 297 151 497
rect 211 297 247 497
rect 307 297 343 497
rect 403 297 439 497
rect 499 297 535 497
rect 701 297 737 497
rect 795 297 831 497
rect 889 297 925 497
rect 983 297 1019 497
rect 1077 297 1113 497
rect 1171 297 1207 497
<< ndiff >>
rect 36 157 123 177
rect 36 123 52 157
rect 86 123 123 157
rect 36 89 123 123
rect 36 55 52 89
rect 86 55 123 89
rect 36 47 123 55
rect 153 89 209 177
rect 153 55 164 89
rect 198 55 209 89
rect 153 47 209 55
rect 239 157 305 177
rect 239 123 260 157
rect 294 123 305 157
rect 239 47 305 123
rect 335 89 401 177
rect 335 55 356 89
rect 390 55 401 89
rect 335 47 401 55
rect 431 157 497 177
rect 431 123 452 157
rect 486 123 497 157
rect 431 47 497 123
rect 527 89 709 177
rect 527 55 570 89
rect 604 55 651 89
rect 685 55 709 89
rect 527 47 709 55
rect 739 169 803 177
rect 739 135 749 169
rect 783 135 803 169
rect 739 101 803 135
rect 739 67 749 101
rect 783 67 803 101
rect 739 47 803 67
rect 833 89 905 177
rect 833 55 851 89
rect 885 55 905 89
rect 833 47 905 55
rect 935 47 981 177
rect 1011 131 1085 177
rect 1011 97 1031 131
rect 1065 97 1085 131
rect 1011 47 1085 97
rect 1115 47 1169 177
rect 1199 161 1261 177
rect 1199 127 1219 161
rect 1253 127 1261 161
rect 1199 93 1261 127
rect 1199 59 1219 93
rect 1253 59 1261 93
rect 1199 47 1261 59
<< pdiff >>
rect 60 477 115 497
rect 60 443 68 477
rect 102 443 115 477
rect 60 409 115 443
rect 60 375 68 409
rect 102 375 115 409
rect 60 297 115 375
rect 151 489 211 497
rect 151 455 164 489
rect 198 455 211 489
rect 151 297 211 455
rect 247 353 307 497
rect 247 319 260 353
rect 294 319 307 353
rect 247 297 307 319
rect 343 489 403 497
rect 343 455 356 489
rect 390 455 403 489
rect 343 297 403 455
rect 439 353 499 497
rect 439 319 452 353
rect 486 319 499 353
rect 439 297 499 319
rect 535 489 593 497
rect 535 455 547 489
rect 581 455 593 489
rect 535 297 593 455
rect 647 459 701 497
rect 647 425 655 459
rect 689 425 701 459
rect 647 389 701 425
rect 647 355 655 389
rect 689 355 701 389
rect 647 297 701 355
rect 737 341 795 497
rect 737 307 749 341
rect 783 307 795 341
rect 737 297 795 307
rect 831 428 889 497
rect 831 394 843 428
rect 877 394 889 428
rect 831 339 889 394
rect 831 305 843 339
rect 877 305 889 339
rect 831 297 889 305
rect 925 489 983 497
rect 925 455 937 489
rect 971 455 983 489
rect 925 297 983 455
rect 1019 421 1077 497
rect 1019 387 1031 421
rect 1065 387 1077 421
rect 1019 297 1077 387
rect 1113 489 1171 497
rect 1113 455 1125 489
rect 1159 455 1171 489
rect 1113 297 1171 455
rect 1207 419 1261 497
rect 1207 385 1219 419
rect 1253 385 1261 419
rect 1207 343 1261 385
rect 1207 309 1219 343
rect 1253 309 1261 343
rect 1207 297 1261 309
<< ndiffc >>
rect 52 123 86 157
rect 52 55 86 89
rect 164 55 198 89
rect 260 123 294 157
rect 356 55 390 89
rect 452 123 486 157
rect 570 55 604 89
rect 651 55 685 89
rect 749 135 783 169
rect 749 67 783 101
rect 851 55 885 89
rect 1031 97 1065 131
rect 1219 127 1253 161
rect 1219 59 1253 93
<< pdiffc >>
rect 68 443 102 477
rect 68 375 102 409
rect 164 455 198 489
rect 260 319 294 353
rect 356 455 390 489
rect 452 319 486 353
rect 547 455 581 489
rect 655 425 689 459
rect 655 355 689 389
rect 749 307 783 341
rect 843 394 877 428
rect 843 305 877 339
rect 937 455 971 489
rect 1031 387 1065 421
rect 1125 455 1159 489
rect 1219 385 1253 419
rect 1219 309 1253 343
<< poly >>
rect 115 497 151 523
rect 211 497 247 523
rect 307 497 343 523
rect 403 497 439 523
rect 499 497 535 523
rect 701 497 737 523
rect 795 497 831 523
rect 889 497 925 523
rect 983 497 1019 523
rect 1077 497 1113 523
rect 1171 497 1207 523
rect 115 282 151 297
rect 211 282 247 297
rect 307 282 343 297
rect 403 282 439 297
rect 499 282 535 297
rect 701 282 737 297
rect 795 282 831 297
rect 889 282 925 297
rect 983 282 1019 297
rect 1077 282 1113 297
rect 1171 282 1207 297
rect 113 265 153 282
rect 209 265 249 282
rect 305 265 345 282
rect 401 265 441 282
rect 497 265 537 282
rect 699 265 739 282
rect 793 265 833 282
rect 887 265 927 282
rect 981 265 1021 282
rect 1075 265 1115 282
rect 100 249 164 265
rect 100 215 110 249
rect 144 215 164 249
rect 100 199 164 215
rect 209 249 560 265
rect 209 215 360 249
rect 394 215 428 249
rect 462 215 506 249
rect 540 215 560 249
rect 209 199 560 215
rect 661 249 833 265
rect 661 215 671 249
rect 705 215 833 249
rect 661 199 833 215
rect 875 249 939 265
rect 875 215 885 249
rect 919 215 939 249
rect 875 199 939 215
rect 981 249 1115 265
rect 981 215 1025 249
rect 1059 215 1115 249
rect 981 199 1115 215
rect 123 177 153 199
rect 209 177 239 199
rect 305 177 335 199
rect 401 177 431 199
rect 497 177 527 199
rect 709 177 739 199
rect 803 177 833 199
rect 905 177 935 199
rect 981 177 1011 199
rect 1085 177 1115 199
rect 1169 265 1209 282
rect 1169 249 1233 265
rect 1169 215 1179 249
rect 1213 215 1233 249
rect 1169 199 1233 215
rect 1169 177 1199 199
rect 123 21 153 47
rect 209 21 239 47
rect 305 21 335 47
rect 401 21 431 47
rect 497 21 527 47
rect 709 21 739 47
rect 803 21 833 47
rect 905 21 935 47
rect 981 21 1011 47
rect 1085 21 1115 47
rect 1169 21 1199 47
<< polycont >>
rect 110 215 144 249
rect 360 215 394 249
rect 428 215 462 249
rect 506 215 540 249
rect 671 215 705 249
rect 885 215 919 249
rect 1025 215 1059 249
rect 1179 215 1213 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 21 477 104 493
rect 21 443 68 477
rect 102 443 104 477
rect 138 489 214 527
rect 138 455 164 489
rect 198 455 214 489
rect 330 489 406 527
rect 330 455 356 489
rect 390 455 406 489
rect 521 489 598 527
rect 521 455 547 489
rect 581 455 598 489
rect 911 489 987 527
rect 655 459 877 476
rect 21 421 104 443
rect 689 442 877 459
rect 911 455 937 489
rect 971 455 987 489
rect 1099 489 1175 527
rect 1099 455 1125 489
rect 1159 455 1175 489
rect 21 409 618 421
rect 21 375 68 409
rect 102 387 618 409
rect 102 375 107 387
rect 21 359 107 375
rect 21 168 60 359
rect 94 249 170 325
rect 94 215 110 249
rect 144 215 170 249
rect 94 202 170 215
rect 210 319 260 353
rect 294 319 452 353
rect 486 319 516 353
rect 21 157 102 168
rect 21 123 52 157
rect 86 123 102 157
rect 210 157 308 319
rect 584 305 618 387
rect 655 389 689 425
rect 841 428 877 442
rect 841 394 843 428
rect 877 394 1031 421
rect 841 387 1031 394
rect 1065 419 1269 421
rect 1065 387 1219 419
rect 655 339 689 355
rect 749 341 783 361
rect 584 271 705 305
rect 342 249 550 265
rect 342 215 360 249
rect 394 215 428 249
rect 462 215 506 249
rect 540 237 550 249
rect 643 249 705 271
rect 540 215 606 237
rect 342 199 606 215
rect 643 215 671 249
rect 643 199 705 215
rect 572 157 606 199
rect 749 169 783 307
rect 841 339 877 387
rect 1218 385 1219 387
rect 1253 385 1269 419
rect 841 305 843 339
rect 841 289 877 305
rect 913 319 1172 353
rect 913 255 958 319
rect 869 249 958 255
rect 869 215 885 249
rect 919 215 958 249
rect 869 202 958 215
rect 992 249 1075 272
rect 992 215 1025 249
rect 1059 215 1075 249
rect 992 202 1075 215
rect 1126 258 1172 319
rect 1218 343 1269 385
rect 1218 309 1219 343
rect 1253 309 1269 343
rect 1218 292 1269 309
rect 1126 249 1244 258
rect 1126 215 1179 249
rect 1213 215 1244 249
rect 1126 211 1244 215
rect 210 123 260 157
rect 294 123 452 157
rect 486 123 502 157
rect 572 135 749 157
rect 783 135 1077 168
rect 572 134 1077 135
rect 572 123 783 134
rect 21 89 102 123
rect 749 101 783 123
rect 21 55 52 89
rect 86 55 102 89
rect 21 51 102 55
rect 136 55 164 89
rect 198 55 214 89
rect 136 17 214 55
rect 330 55 356 89
rect 390 55 406 89
rect 330 17 406 55
rect 547 55 570 89
rect 604 55 651 89
rect 685 55 701 89
rect 547 17 701 55
rect 1021 131 1077 134
rect 1021 97 1031 131
rect 1065 97 1077 131
rect 749 51 783 67
rect 835 55 851 89
rect 885 55 901 89
rect 1021 81 1077 97
rect 1213 161 1269 177
rect 1213 127 1219 161
rect 1253 127 1269 161
rect 1213 93 1269 127
rect 835 17 901 55
rect 1213 59 1219 93
rect 1253 59 1269 93
rect 1213 17 1269 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
flabel corelocali s 115 221 159 255 0 FreeSans 340 0 0 0 B1_N
port 3 nsew
flabel corelocali s 1185 240 1185 240 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 1040 221 1074 255 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 223 289 267 323 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 1288 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1150338
string GDS_START 1141668
<< end >>
