magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 89 93 119 177
rect 287 47 317 177
rect 403 47 433 177
rect 497 47 527 177
rect 581 47 611 177
rect 697 47 727 177
rect 791 47 821 177
rect 885 47 915 177
rect 989 47 1019 177
<< pmoshvt >>
rect 81 413 117 497
rect 279 297 315 497
rect 395 297 431 497
rect 489 297 525 497
rect 583 297 619 497
rect 699 297 735 497
rect 793 297 829 497
rect 887 297 923 497
rect 981 297 1017 497
<< ndiff >>
rect 27 149 89 177
rect 27 115 35 149
rect 69 115 89 149
rect 27 93 89 115
rect 119 165 171 177
rect 119 131 129 165
rect 163 131 171 165
rect 119 120 171 131
rect 119 93 169 120
rect 227 104 287 177
rect 225 93 287 104
rect 225 59 233 93
rect 267 59 287 93
rect 225 47 287 59
rect 317 115 403 177
rect 317 81 343 115
rect 377 81 403 115
rect 317 47 403 81
rect 433 97 497 177
rect 433 63 443 97
rect 477 63 497 97
rect 433 47 497 63
rect 527 115 581 177
rect 527 81 537 115
rect 571 81 581 115
rect 527 47 581 81
rect 611 97 697 177
rect 611 63 651 97
rect 685 63 697 97
rect 611 47 697 63
rect 727 114 791 177
rect 727 80 747 114
rect 781 80 791 114
rect 727 47 791 80
rect 821 95 885 177
rect 821 61 841 95
rect 875 61 885 95
rect 821 47 885 61
rect 915 163 989 177
rect 915 129 935 163
rect 969 129 989 163
rect 915 95 989 129
rect 915 61 935 95
rect 969 61 989 95
rect 915 47 989 61
rect 1019 95 1074 177
rect 1019 61 1029 95
rect 1063 61 1074 95
rect 1019 47 1074 61
<< pdiff >>
rect 27 477 81 497
rect 27 443 35 477
rect 69 443 81 477
rect 27 413 81 443
rect 117 472 171 497
rect 117 438 129 472
rect 163 438 171 472
rect 117 413 171 438
rect 225 485 279 497
rect 225 451 233 485
rect 267 451 279 485
rect 225 417 279 451
rect 225 383 233 417
rect 267 383 279 417
rect 225 349 279 383
rect 225 315 233 349
rect 267 315 279 349
rect 225 297 279 315
rect 315 297 395 497
rect 431 297 489 497
rect 525 297 583 497
rect 619 477 699 497
rect 619 443 642 477
rect 676 443 699 477
rect 619 409 699 443
rect 619 375 642 409
rect 676 375 699 409
rect 619 297 699 375
rect 735 477 793 497
rect 735 443 747 477
rect 781 443 793 477
rect 735 409 793 443
rect 735 375 747 409
rect 781 375 793 409
rect 735 341 793 375
rect 735 307 747 341
rect 781 307 793 341
rect 735 297 793 307
rect 829 477 887 497
rect 829 443 841 477
rect 875 443 887 477
rect 829 409 887 443
rect 829 375 841 409
rect 875 375 887 409
rect 829 297 887 375
rect 923 477 981 497
rect 923 443 935 477
rect 969 443 981 477
rect 923 409 981 443
rect 923 375 935 409
rect 969 375 981 409
rect 923 341 981 375
rect 923 307 935 341
rect 969 307 981 341
rect 923 297 981 307
rect 1017 477 1071 497
rect 1017 443 1029 477
rect 1063 443 1071 477
rect 1017 409 1071 443
rect 1017 375 1029 409
rect 1063 375 1071 409
rect 1017 297 1071 375
<< ndiffc >>
rect 35 115 69 149
rect 129 131 163 165
rect 233 59 267 93
rect 343 81 377 115
rect 443 63 477 97
rect 537 81 571 115
rect 651 63 685 97
rect 747 80 781 114
rect 841 61 875 95
rect 935 129 969 163
rect 935 61 969 95
rect 1029 61 1063 95
<< pdiffc >>
rect 35 443 69 477
rect 129 438 163 472
rect 233 451 267 485
rect 233 383 267 417
rect 233 315 267 349
rect 642 443 676 477
rect 642 375 676 409
rect 747 443 781 477
rect 747 375 781 409
rect 747 307 781 341
rect 841 443 875 477
rect 841 375 875 409
rect 935 443 969 477
rect 935 375 969 409
rect 935 307 969 341
rect 1029 443 1063 477
rect 1029 375 1063 409
<< poly >>
rect 81 497 117 523
rect 279 497 315 523
rect 395 497 431 523
rect 489 497 525 523
rect 583 497 619 523
rect 699 497 735 523
rect 793 497 829 523
rect 887 497 923 523
rect 981 497 1017 523
rect 81 398 117 413
rect 79 265 119 398
rect 279 282 315 297
rect 395 282 431 297
rect 489 282 525 297
rect 583 282 619 297
rect 699 282 735 297
rect 793 282 829 297
rect 887 282 923 297
rect 981 282 1017 297
rect 277 265 317 282
rect 393 265 433 282
rect 487 265 527 282
rect 581 265 621 282
rect 697 265 737 282
rect 791 265 831 282
rect 885 265 925 282
rect 979 265 1019 282
rect 45 249 123 265
rect 45 215 55 249
rect 89 215 123 249
rect 45 199 123 215
rect 209 249 317 265
rect 209 215 219 249
rect 253 215 317 249
rect 209 199 317 215
rect 369 249 433 265
rect 369 215 379 249
rect 413 215 433 249
rect 369 199 433 215
rect 475 249 539 265
rect 475 215 491 249
rect 525 215 539 249
rect 475 199 539 215
rect 581 249 645 265
rect 581 215 591 249
rect 625 215 645 249
rect 581 199 645 215
rect 697 249 1019 265
rect 697 215 707 249
rect 741 215 785 249
rect 819 215 863 249
rect 897 215 941 249
rect 975 215 1019 249
rect 697 199 1019 215
rect 89 177 119 199
rect 287 177 317 199
rect 403 177 433 199
rect 497 177 527 199
rect 581 177 611 199
rect 697 177 727 199
rect 791 177 821 199
rect 885 177 915 199
rect 989 177 1019 199
rect 89 67 119 93
rect 287 21 317 47
rect 403 21 433 47
rect 497 21 527 47
rect 581 21 611 47
rect 697 21 727 47
rect 791 21 821 47
rect 885 21 915 47
rect 989 21 1019 47
<< polycont >>
rect 55 215 89 249
rect 219 215 253 249
rect 379 215 413 249
rect 491 215 525 249
rect 591 215 625 249
rect 707 215 741 249
rect 785 215 819 249
rect 863 215 897 249
rect 941 215 975 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 17 477 73 527
rect 17 443 35 477
rect 69 443 73 477
rect 17 427 73 443
rect 129 472 167 491
rect 163 438 167 472
rect 21 249 89 391
rect 21 215 55 249
rect 21 199 89 215
rect 129 265 167 438
rect 217 485 283 490
rect 217 451 233 485
rect 267 451 283 485
rect 634 477 684 527
rect 217 417 283 451
rect 217 383 233 417
rect 267 383 283 417
rect 217 349 283 383
rect 217 315 233 349
rect 267 315 345 349
rect 129 249 253 265
rect 129 215 219 249
rect 129 199 253 215
rect 129 165 167 199
rect 17 149 69 165
rect 17 115 35 149
rect 17 17 69 115
rect 163 131 167 165
rect 301 165 345 315
rect 379 249 437 475
rect 413 215 437 249
rect 379 199 437 215
rect 475 249 541 475
rect 634 443 642 477
rect 676 443 684 477
rect 634 409 684 443
rect 634 375 642 409
rect 676 375 684 409
rect 634 359 684 375
rect 739 477 789 493
rect 739 443 747 477
rect 781 443 789 477
rect 739 409 789 443
rect 739 375 747 409
rect 781 375 789 409
rect 739 341 789 375
rect 833 477 883 527
rect 833 443 841 477
rect 875 443 883 477
rect 833 409 883 443
rect 833 375 841 409
rect 875 375 883 409
rect 833 359 883 375
rect 927 477 977 493
rect 927 443 935 477
rect 969 443 977 477
rect 927 409 977 443
rect 927 375 935 409
rect 969 375 977 409
rect 475 215 491 249
rect 525 215 541 249
rect 475 199 541 215
rect 575 289 688 323
rect 739 307 747 341
rect 781 325 789 341
rect 927 341 977 375
rect 1021 477 1071 527
rect 1021 443 1029 477
rect 1063 443 1071 477
rect 1021 409 1071 443
rect 1021 375 1029 409
rect 1063 375 1071 409
rect 1021 359 1071 375
rect 927 325 935 341
rect 781 307 935 325
rect 969 325 977 341
rect 969 307 1083 325
rect 739 291 1083 307
rect 575 249 635 289
rect 575 215 591 249
rect 625 215 635 249
rect 575 199 635 215
rect 669 215 707 249
rect 741 215 785 249
rect 819 215 863 249
rect 897 215 941 249
rect 975 215 991 249
rect 669 165 703 215
rect 1035 181 1083 291
rect 301 131 703 165
rect 747 163 1083 181
rect 747 145 935 163
rect 129 87 167 131
rect 217 93 267 117
rect 217 59 233 93
rect 343 115 377 131
rect 537 115 571 131
rect 343 61 377 81
rect 417 63 443 97
rect 477 63 493 97
rect 217 17 267 59
rect 417 17 493 63
rect 747 114 797 145
rect 537 61 571 81
rect 625 63 651 97
rect 685 63 701 97
rect 625 17 701 63
rect 781 80 797 114
rect 909 129 935 145
rect 969 145 1083 163
rect 969 129 985 145
rect 747 51 797 80
rect 841 95 875 111
rect 841 17 875 61
rect 909 95 985 129
rect 909 61 935 95
rect 969 61 985 95
rect 909 51 985 61
rect 1029 95 1063 111
rect 1029 17 1063 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
flabel corelocali s 29 221 63 255 0 FreeSans 400 0 0 0 D_N
port 4 nsew
flabel corelocali s 492 425 526 459 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel corelocali s 492 357 526 391 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel corelocali s 399 357 433 391 0 FreeSans 400 0 0 0 C
port 3 nsew
flabel corelocali s 598 306 598 306 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 399 425 433 459 0 FreeSans 400 0 0 0 C
port 3 nsew
flabel corelocali s 1039 153 1073 187 0 FreeSans 400 0 0 0 X
port 9 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
rlabel comment s 0 0 0 0 4 or4b_4
<< properties >>
string FIXED_BBOX 0 0 1104 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 536002
string GDS_START 527266
<< end >>
