magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 1478 704
<< pwell >>
rect 0 0 1440 49
<< scnmos >>
rect 225 74 255 222
rect 311 74 341 222
rect 397 74 427 222
rect 483 74 513 222
rect 581 94 611 222
rect 667 94 697 222
rect 765 108 795 236
rect 860 123 890 251
rect 1034 123 1064 251
rect 1120 123 1150 251
rect 1206 123 1236 251
rect 1292 123 1322 251
<< pmoshvt >>
rect 108 368 138 592
rect 198 368 228 592
rect 288 368 318 592
rect 378 368 408 592
rect 572 392 602 592
rect 672 392 702 592
rect 762 392 792 592
rect 857 392 887 592
rect 948 392 978 592
rect 1109 392 1139 592
rect 1199 392 1229 592
rect 1289 392 1319 592
<< ndiff >>
rect 810 236 860 251
rect 715 222 765 236
rect 172 210 225 222
rect 172 176 180 210
rect 214 176 225 210
rect 172 120 225 176
rect 172 86 180 120
rect 214 86 225 120
rect 172 74 225 86
rect 255 210 311 222
rect 255 176 266 210
rect 300 176 311 210
rect 255 120 311 176
rect 255 86 266 120
rect 300 86 311 120
rect 255 74 311 86
rect 341 122 397 222
rect 341 88 352 122
rect 386 88 397 122
rect 341 74 397 88
rect 427 166 483 222
rect 427 132 438 166
rect 472 132 483 166
rect 427 74 483 132
rect 513 188 581 222
rect 513 154 524 188
rect 558 154 581 188
rect 513 120 581 154
rect 513 86 524 120
rect 558 94 581 120
rect 611 210 667 222
rect 611 176 622 210
rect 656 176 667 210
rect 611 140 667 176
rect 611 106 622 140
rect 656 106 667 140
rect 611 94 667 106
rect 697 140 765 222
rect 697 106 708 140
rect 742 108 765 140
rect 795 196 860 236
rect 795 162 811 196
rect 845 162 860 196
rect 795 123 860 162
rect 890 170 1034 251
rect 890 136 901 170
rect 935 136 1034 170
rect 890 123 1034 136
rect 1064 169 1120 251
rect 1064 135 1075 169
rect 1109 135 1120 169
rect 1064 123 1120 135
rect 1150 238 1206 251
rect 1150 204 1161 238
rect 1195 204 1206 238
rect 1150 123 1206 204
rect 1236 239 1292 251
rect 1236 205 1247 239
rect 1281 205 1292 239
rect 1236 169 1292 205
rect 1236 135 1247 169
rect 1281 135 1292 169
rect 1236 123 1292 135
rect 1322 239 1375 251
rect 1322 205 1333 239
rect 1367 205 1375 239
rect 1322 169 1375 205
rect 1322 135 1333 169
rect 1367 135 1375 169
rect 1322 123 1375 135
rect 795 108 845 123
rect 742 106 750 108
rect 697 94 750 106
rect 558 86 566 94
rect 513 74 566 86
<< pdiff >>
rect 53 580 108 592
rect 53 546 61 580
rect 95 546 108 580
rect 53 497 108 546
rect 53 463 61 497
rect 95 463 108 497
rect 53 414 108 463
rect 53 380 61 414
rect 95 380 108 414
rect 53 368 108 380
rect 138 580 198 592
rect 138 546 151 580
rect 185 546 198 580
rect 138 497 198 546
rect 138 463 151 497
rect 185 463 198 497
rect 138 414 198 463
rect 138 380 151 414
rect 185 380 198 414
rect 138 368 198 380
rect 228 580 288 592
rect 228 546 241 580
rect 275 546 288 580
rect 228 462 288 546
rect 228 428 241 462
rect 275 428 288 462
rect 228 368 288 428
rect 318 580 378 592
rect 318 546 331 580
rect 365 546 378 580
rect 318 497 378 546
rect 318 463 331 497
rect 365 463 378 497
rect 318 414 378 463
rect 318 380 331 414
rect 365 380 378 414
rect 318 368 378 380
rect 408 580 463 592
rect 408 546 421 580
rect 455 546 463 580
rect 408 497 463 546
rect 408 463 421 497
rect 455 463 463 497
rect 408 414 463 463
rect 408 380 421 414
rect 455 380 463 414
rect 517 530 572 592
rect 517 496 525 530
rect 559 496 572 530
rect 517 392 572 496
rect 602 582 672 592
rect 602 548 625 582
rect 659 548 672 582
rect 602 392 672 548
rect 702 446 762 592
rect 702 412 715 446
rect 749 412 762 446
rect 702 392 762 412
rect 792 582 857 592
rect 792 548 807 582
rect 841 548 857 582
rect 792 392 857 548
rect 887 582 948 592
rect 887 548 900 582
rect 934 548 948 582
rect 887 514 948 548
rect 887 480 900 514
rect 934 480 948 514
rect 887 446 948 480
rect 887 412 900 446
rect 934 412 948 446
rect 887 392 948 412
rect 978 582 1109 592
rect 978 548 992 582
rect 1026 548 1061 582
rect 1095 548 1109 582
rect 978 514 1109 548
rect 978 480 992 514
rect 1026 480 1061 514
rect 1095 480 1109 514
rect 978 392 1109 480
rect 1139 580 1199 592
rect 1139 546 1152 580
rect 1186 546 1199 580
rect 1139 510 1199 546
rect 1139 476 1152 510
rect 1186 476 1199 510
rect 1139 440 1199 476
rect 1139 406 1152 440
rect 1186 406 1199 440
rect 1139 392 1199 406
rect 1229 580 1289 592
rect 1229 546 1242 580
rect 1276 546 1289 580
rect 1229 492 1289 546
rect 1229 458 1242 492
rect 1276 458 1289 492
rect 1229 392 1289 458
rect 1319 580 1374 592
rect 1319 546 1332 580
rect 1366 546 1374 580
rect 1319 509 1374 546
rect 1319 475 1332 509
rect 1366 475 1374 509
rect 1319 438 1374 475
rect 1319 404 1332 438
rect 1366 404 1374 438
rect 1319 392 1374 404
rect 408 368 463 380
<< ndiffc >>
rect 180 176 214 210
rect 180 86 214 120
rect 266 176 300 210
rect 266 86 300 120
rect 352 88 386 122
rect 438 132 472 166
rect 524 154 558 188
rect 524 86 558 120
rect 622 176 656 210
rect 622 106 656 140
rect 708 106 742 140
rect 811 162 845 196
rect 901 136 935 170
rect 1075 135 1109 169
rect 1161 204 1195 238
rect 1247 205 1281 239
rect 1247 135 1281 169
rect 1333 205 1367 239
rect 1333 135 1367 169
<< pdiffc >>
rect 61 546 95 580
rect 61 463 95 497
rect 61 380 95 414
rect 151 546 185 580
rect 151 463 185 497
rect 151 380 185 414
rect 241 546 275 580
rect 241 428 275 462
rect 331 546 365 580
rect 331 463 365 497
rect 331 380 365 414
rect 421 546 455 580
rect 421 463 455 497
rect 421 380 455 414
rect 525 496 559 530
rect 625 548 659 582
rect 715 412 749 446
rect 807 548 841 582
rect 900 548 934 582
rect 900 480 934 514
rect 900 412 934 446
rect 992 548 1026 582
rect 1061 548 1095 582
rect 992 480 1026 514
rect 1061 480 1095 514
rect 1152 546 1186 580
rect 1152 476 1186 510
rect 1152 406 1186 440
rect 1242 546 1276 580
rect 1242 458 1276 492
rect 1332 546 1366 580
rect 1332 475 1366 509
rect 1332 404 1366 438
<< poly >>
rect 108 592 138 618
rect 198 592 228 618
rect 288 592 318 618
rect 378 592 408 618
rect 572 592 602 618
rect 672 592 702 618
rect 762 592 792 618
rect 857 592 887 618
rect 948 592 978 618
rect 1109 592 1139 618
rect 1199 592 1229 618
rect 1289 592 1319 618
rect 572 377 602 392
rect 672 377 702 392
rect 762 377 792 392
rect 857 377 887 392
rect 948 377 978 392
rect 1109 377 1139 392
rect 1199 377 1229 392
rect 1289 377 1319 392
rect 108 353 138 368
rect 198 353 228 368
rect 288 353 318 368
rect 378 353 408 368
rect 569 360 605 377
rect 105 310 141 353
rect 195 310 231 353
rect 285 310 321 353
rect 375 310 411 353
rect 555 344 621 360
rect 555 310 571 344
rect 605 310 621 344
rect 669 324 705 377
rect 759 324 795 377
rect 854 360 890 377
rect 105 294 459 310
rect 555 294 621 310
rect 667 308 795 324
rect 105 280 409 294
rect 225 222 255 280
rect 311 260 409 280
rect 443 274 459 294
rect 443 260 513 274
rect 311 244 513 260
rect 311 222 341 244
rect 397 222 427 244
rect 483 222 513 244
rect 581 222 611 294
rect 667 274 706 308
rect 740 274 795 308
rect 837 344 903 360
rect 837 310 853 344
rect 887 310 903 344
rect 837 294 903 310
rect 945 296 981 377
rect 1106 356 1142 377
rect 1196 356 1232 377
rect 1106 340 1236 356
rect 1106 306 1122 340
rect 1156 306 1236 340
rect 667 258 795 274
rect 667 222 697 258
rect 765 236 795 258
rect 860 251 890 294
rect 945 266 1064 296
rect 1106 290 1236 306
rect 1034 251 1064 266
rect 1120 251 1150 290
rect 1206 251 1236 290
rect 1286 277 1322 377
rect 1292 251 1322 277
rect 225 48 255 74
rect 311 48 341 74
rect 397 48 427 74
rect 483 48 513 74
rect 581 68 611 94
rect 667 68 697 94
rect 765 82 795 108
rect 860 97 890 123
rect 1034 101 1064 123
rect 998 85 1064 101
rect 1120 97 1150 123
rect 1206 97 1236 123
rect 998 51 1014 85
rect 1048 55 1064 85
rect 1292 55 1322 123
rect 1048 51 1322 55
rect 998 25 1322 51
<< polycont >>
rect 571 310 605 344
rect 409 260 443 294
rect 706 274 740 308
rect 853 310 887 344
rect 1122 306 1156 340
rect 1014 51 1048 85
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 45 580 95 649
rect 45 546 61 580
rect 45 497 95 546
rect 45 463 61 497
rect 45 414 95 463
rect 45 380 61 414
rect 45 364 95 380
rect 135 580 185 596
rect 135 546 151 580
rect 135 497 185 546
rect 135 463 151 497
rect 135 414 185 463
rect 135 380 151 414
rect 225 580 275 649
rect 225 546 241 580
rect 225 462 275 546
rect 225 428 241 462
rect 225 412 275 428
rect 315 580 381 596
rect 315 546 331 580
rect 365 546 381 580
rect 315 497 381 546
rect 315 463 331 497
rect 365 463 381 497
rect 315 414 381 463
rect 135 378 185 380
rect 315 380 331 414
rect 365 380 381 414
rect 315 378 381 380
rect 135 344 381 378
rect 421 580 455 649
rect 609 582 860 598
rect 421 497 455 546
rect 509 530 575 556
rect 609 548 625 582
rect 659 548 807 582
rect 841 548 860 582
rect 900 582 942 598
rect 934 548 942 582
rect 509 496 525 530
rect 559 514 575 530
rect 900 514 942 548
rect 559 496 900 514
rect 509 480 900 496
rect 934 480 942 514
rect 976 582 1111 649
rect 976 548 992 582
rect 1026 548 1061 582
rect 1095 548 1111 582
rect 976 514 1111 548
rect 976 480 992 514
rect 1026 480 1061 514
rect 1095 480 1111 514
rect 1145 580 1192 596
rect 1145 546 1152 580
rect 1186 546 1192 580
rect 1145 510 1192 546
rect 421 414 455 463
rect 884 446 942 480
rect 1145 476 1152 510
rect 1186 476 1192 510
rect 1145 446 1192 476
rect 1226 580 1292 649
rect 1226 546 1242 580
rect 1276 546 1292 580
rect 1226 492 1292 546
rect 1226 458 1242 492
rect 1276 458 1292 492
rect 1326 580 1382 596
rect 1326 546 1332 580
rect 1366 546 1382 580
rect 1326 509 1382 546
rect 1326 475 1332 509
rect 1366 475 1382 509
rect 421 364 455 380
rect 489 412 715 446
rect 749 412 765 446
rect 135 282 185 344
rect 489 310 523 412
rect 799 378 839 430
rect 884 412 900 446
rect 934 440 1192 446
rect 934 412 1152 440
rect 1136 406 1152 412
rect 1186 424 1192 440
rect 1326 438 1382 475
rect 1326 424 1332 438
rect 1186 406 1332 424
rect 1136 404 1332 406
rect 1366 404 1382 438
rect 1136 390 1382 404
rect 1316 388 1382 390
rect 393 294 523 310
rect 557 344 903 378
rect 557 310 571 344
rect 605 310 621 344
rect 793 310 853 344
rect 887 310 903 344
rect 557 294 621 310
rect 690 308 756 310
rect 135 248 359 282
rect 266 210 359 248
rect 393 260 409 294
rect 443 260 523 294
rect 690 274 706 308
rect 740 274 756 308
rect 793 294 903 310
rect 985 340 1223 356
rect 985 306 1122 340
rect 1156 306 1223 340
rect 985 290 1223 306
rect 393 226 656 260
rect 690 242 756 274
rect 164 176 180 210
rect 214 176 230 210
rect 164 120 230 176
rect 164 86 180 120
rect 214 86 230 120
rect 164 17 230 86
rect 300 192 359 210
rect 608 210 656 226
rect 300 176 474 192
rect 266 166 474 176
rect 266 158 438 166
rect 266 120 300 158
rect 436 132 438 158
rect 472 132 474 166
rect 266 70 300 86
rect 336 122 402 124
rect 336 88 352 122
rect 386 88 402 122
rect 436 109 474 132
rect 508 188 574 192
rect 508 154 524 188
rect 558 154 574 188
rect 508 120 574 154
rect 336 17 402 88
rect 508 86 524 120
rect 558 86 574 120
rect 608 176 622 210
rect 792 238 1211 256
rect 792 222 1161 238
rect 792 208 849 222
rect 656 196 849 208
rect 1145 204 1161 222
rect 1195 204 1211 238
rect 1145 203 1211 204
rect 1247 239 1281 255
rect 656 176 811 196
rect 608 174 811 176
rect 608 140 656 174
rect 792 162 811 174
rect 845 162 849 196
rect 608 106 622 140
rect 608 90 656 106
rect 692 106 708 140
rect 742 106 758 140
rect 792 119 849 162
rect 885 170 951 188
rect 885 136 901 170
rect 935 136 951 170
rect 1247 169 1281 205
rect 508 17 574 86
rect 692 17 758 106
rect 885 17 951 136
rect 1059 135 1075 169
rect 1109 135 1247 169
rect 985 101 1025 134
rect 1247 119 1281 135
rect 1317 239 1383 255
rect 1317 205 1333 239
rect 1367 205 1383 239
rect 1317 169 1383 205
rect 1317 135 1333 169
rect 1367 135 1383 169
rect 985 85 1064 101
rect 985 51 1014 85
rect 1048 51 1064 85
rect 1317 17 1383 135
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 683 1440 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 0 617 1440 649
rect 0 17 1440 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -49 1440 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a211o_4
flabel pwell s 0 0 1440 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 1440 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 1440 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 1440 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 319 168 353 202 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 319 242 353 276 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 703 242 737 276 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 799 390 833 424 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 991 94 1025 128 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 1183 316 1217 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 1440 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3950722
string GDS_START 3939174
<< end >>
