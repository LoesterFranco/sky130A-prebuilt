magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 552 561
rect 105 445 171 527
rect 21 195 67 333
rect 209 269 275 491
rect 381 381 447 527
rect 209 209 316 269
rect 185 17 231 173
rect 267 159 316 209
rect 352 199 431 269
rect 470 199 528 269
rect 267 53 353 159
rect 389 75 431 199
rect 465 17 531 163
rect 0 -17 552 17
<< obsli1 >>
rect 19 409 71 487
rect 19 369 171 409
rect 103 233 171 369
rect 309 345 347 491
rect 483 345 517 491
rect 309 305 517 345
rect 103 143 149 233
rect 73 53 149 143
<< metal1 >>
rect 0 496 552 592
rect 0 -48 552 48
<< labels >>
rlabel locali s 389 75 431 199 6 A1
port 1 nsew signal input
rlabel locali s 352 199 431 269 6 A1
port 1 nsew signal input
rlabel locali s 470 199 528 269 6 A2
port 2 nsew signal input
rlabel locali s 21 195 67 333 6 B1_N
port 3 nsew signal input
rlabel locali s 267 159 316 209 6 Y
port 4 nsew signal output
rlabel locali s 267 53 353 159 6 Y
port 4 nsew signal output
rlabel locali s 209 269 275 491 6 Y
port 4 nsew signal output
rlabel locali s 209 209 316 269 6 Y
port 4 nsew signal output
rlabel locali s 465 17 531 163 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 185 17 231 173 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 552 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 552 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 381 381 447 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 105 445 171 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 552 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 552 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 552 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 4009346
string GDS_START 4003110
<< end >>
