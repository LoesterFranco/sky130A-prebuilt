magic
tech sky130A
magscale 1 2
timestamp 1604502710
<< nwell >>
rect -38 332 1094 704
<< pwell >>
rect 0 0 1056 49
<< scpmos >>
rect 83 368 119 592
rect 173 368 209 592
rect 263 368 299 592
rect 353 368 389 592
rect 443 368 479 592
rect 533 368 569 592
rect 623 368 659 592
rect 723 368 759 592
rect 840 403 876 571
rect 930 403 966 571
<< nmoslvt >>
rect 387 74 417 222
rect 473 74 503 222
rect 687 74 717 222
rect 773 74 803 222
rect 859 74 889 222
<< ndiff >>
rect 314 84 387 222
rect 314 50 326 84
rect 360 74 387 84
rect 417 152 473 222
rect 417 118 428 152
rect 462 118 473 152
rect 417 74 473 118
rect 503 84 687 222
rect 503 74 530 84
rect 360 50 372 74
rect 314 38 372 50
rect 518 50 530 74
rect 564 50 626 84
rect 660 74 687 84
rect 717 152 773 222
rect 717 118 728 152
rect 762 118 773 152
rect 717 74 773 118
rect 803 152 859 222
rect 803 118 814 152
rect 848 118 859 152
rect 803 74 859 118
rect 889 186 1029 222
rect 889 152 900 186
rect 934 152 983 186
rect 1017 152 1029 186
rect 889 118 1029 152
rect 889 84 900 118
rect 934 84 983 118
rect 1017 84 1029 118
rect 889 74 1029 84
rect 660 50 672 74
rect 518 38 672 50
<< pdiff >>
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 500 83 546
rect 27 466 39 500
rect 73 466 83 500
rect 27 420 83 466
rect 27 386 39 420
rect 73 386 83 420
rect 27 368 83 386
rect 119 580 173 592
rect 119 546 129 580
rect 163 546 173 580
rect 119 507 173 546
rect 119 473 129 507
rect 163 473 173 507
rect 119 434 173 473
rect 119 400 129 434
rect 163 400 173 434
rect 119 368 173 400
rect 209 580 263 592
rect 209 546 219 580
rect 253 546 263 580
rect 209 502 263 546
rect 209 468 219 502
rect 253 468 263 502
rect 209 368 263 468
rect 299 580 353 592
rect 299 546 309 580
rect 343 546 353 580
rect 299 507 353 546
rect 299 473 309 507
rect 343 473 353 507
rect 299 434 353 473
rect 299 400 309 434
rect 343 400 353 434
rect 299 368 353 400
rect 389 531 443 592
rect 389 497 399 531
rect 433 497 443 531
rect 389 420 443 497
rect 389 386 399 420
rect 433 386 443 420
rect 389 368 443 386
rect 479 582 533 592
rect 479 548 489 582
rect 523 548 533 582
rect 479 514 533 548
rect 479 480 489 514
rect 523 480 533 514
rect 479 368 533 480
rect 569 531 623 592
rect 569 497 579 531
rect 613 497 623 531
rect 569 446 623 497
rect 569 412 579 446
rect 613 412 623 446
rect 569 368 623 412
rect 659 582 723 592
rect 659 548 679 582
rect 713 548 723 582
rect 659 514 723 548
rect 659 480 679 514
rect 713 480 723 514
rect 659 446 723 480
rect 659 412 679 446
rect 713 412 723 446
rect 659 368 723 412
rect 759 582 825 592
rect 759 548 779 582
rect 813 571 825 582
rect 813 548 840 571
rect 759 514 840 548
rect 759 480 779 514
rect 813 480 840 514
rect 759 446 840 480
rect 759 412 779 446
rect 813 412 840 446
rect 759 403 840 412
rect 876 559 930 571
rect 876 525 886 559
rect 920 525 930 559
rect 876 449 930 525
rect 876 415 886 449
rect 920 415 930 449
rect 876 403 930 415
rect 966 559 1022 571
rect 966 525 976 559
rect 1010 525 1022 559
rect 966 449 1022 525
rect 966 415 976 449
rect 1010 415 1022 449
rect 966 403 1022 415
rect 759 368 825 403
<< ndiffc >>
rect 326 50 360 84
rect 428 118 462 152
rect 530 50 564 84
rect 626 50 660 84
rect 728 118 762 152
rect 814 118 848 152
rect 900 152 934 186
rect 983 152 1017 186
rect 900 84 934 118
rect 983 84 1017 118
<< pdiffc >>
rect 39 546 73 580
rect 39 466 73 500
rect 39 386 73 420
rect 129 546 163 580
rect 129 473 163 507
rect 129 400 163 434
rect 219 546 253 580
rect 219 468 253 502
rect 309 546 343 580
rect 309 473 343 507
rect 309 400 343 434
rect 399 497 433 531
rect 399 386 433 420
rect 489 548 523 582
rect 489 480 523 514
rect 579 497 613 531
rect 579 412 613 446
rect 679 548 713 582
rect 679 480 713 514
rect 679 412 713 446
rect 779 548 813 582
rect 779 480 813 514
rect 779 412 813 446
rect 886 525 920 559
rect 886 415 920 449
rect 976 525 1010 559
rect 976 415 1010 449
<< poly >>
rect 83 592 119 618
rect 173 592 209 618
rect 263 592 299 618
rect 353 592 389 618
rect 443 592 479 618
rect 533 592 569 618
rect 623 592 659 618
rect 723 592 759 618
rect 840 571 876 597
rect 930 571 966 597
rect 840 388 876 403
rect 930 388 966 403
rect 83 268 119 368
rect 173 268 209 368
rect 263 268 299 368
rect 353 353 389 368
rect 443 353 479 368
rect 533 353 569 368
rect 623 353 659 368
rect 353 323 659 353
rect 83 252 299 268
rect 83 238 174 252
rect 89 218 174 238
rect 208 218 242 252
rect 276 218 299 252
rect 387 320 645 323
rect 387 286 459 320
rect 493 286 527 320
rect 561 286 595 320
rect 629 286 645 320
rect 387 245 645 286
rect 723 310 759 368
rect 840 358 1012 388
rect 859 349 1012 358
rect 859 315 962 349
rect 996 315 1012 349
rect 723 294 803 310
rect 723 274 745 294
rect 687 260 745 274
rect 779 260 803 294
rect 387 222 417 245
rect 473 222 503 245
rect 687 244 803 260
rect 687 222 717 244
rect 773 222 803 244
rect 859 299 1012 315
rect 859 222 889 299
rect 89 202 299 218
rect 387 48 417 74
rect 473 48 503 74
rect 687 48 717 74
rect 773 48 803 74
rect 859 48 889 74
<< polycont >>
rect 174 218 208 252
rect 242 218 276 252
rect 459 286 493 320
rect 527 286 561 320
rect 595 286 629 320
rect 962 315 996 349
rect 745 260 779 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 23 580 73 649
rect 23 546 39 580
rect 23 500 73 546
rect 23 466 39 500
rect 23 420 73 466
rect 23 386 39 420
rect 23 370 73 386
rect 113 580 179 596
rect 113 546 129 580
rect 163 546 179 580
rect 113 507 179 546
rect 113 473 129 507
rect 163 473 179 507
rect 113 434 179 473
rect 219 580 253 649
rect 219 502 253 546
rect 219 452 253 468
rect 293 582 729 615
rect 293 581 489 582
rect 293 580 343 581
rect 293 546 309 580
rect 473 548 489 581
rect 523 581 679 582
rect 523 548 539 581
rect 293 507 343 546
rect 293 473 309 507
rect 113 400 129 434
rect 163 418 179 434
rect 293 434 343 473
rect 293 418 309 434
rect 163 400 309 418
rect 113 384 343 400
rect 377 531 433 547
rect 377 497 399 531
rect 377 446 433 497
rect 473 514 539 548
rect 663 548 679 581
rect 713 548 729 582
rect 473 480 489 514
rect 523 480 539 514
rect 579 531 629 547
rect 613 497 629 531
rect 579 446 629 497
rect 377 420 579 446
rect 377 386 399 420
rect 433 412 579 420
rect 613 412 629 446
rect 663 514 729 548
rect 663 480 679 514
rect 713 480 729 514
rect 663 446 729 480
rect 663 412 679 446
rect 713 412 729 446
rect 763 582 829 649
rect 763 548 779 582
rect 813 548 829 582
rect 763 514 829 548
rect 763 480 779 514
rect 813 480 829 514
rect 763 446 829 480
rect 763 412 779 446
rect 813 412 829 446
rect 870 559 936 575
rect 870 525 886 559
rect 920 525 936 559
rect 870 449 936 525
rect 870 415 886 449
rect 920 415 936 449
rect 377 370 433 386
rect 870 399 936 415
rect 976 559 1026 649
rect 1010 525 1026 559
rect 976 449 1026 525
rect 1010 415 1026 449
rect 976 399 1026 415
rect 870 378 916 399
rect 377 350 411 370
rect 107 336 411 350
rect 611 344 916 378
rect 611 336 645 344
rect 37 316 411 336
rect 445 320 645 336
rect 37 302 141 316
rect 37 282 71 302
rect 445 286 459 320
rect 493 286 527 320
rect 561 286 595 320
rect 629 286 645 320
rect 25 168 71 282
rect 217 268 359 282
rect 445 270 645 286
rect 729 294 795 310
rect 158 252 359 268
rect 158 218 174 252
rect 208 218 242 252
rect 276 236 359 252
rect 729 260 745 294
rect 779 260 795 294
rect 729 236 795 260
rect 276 218 795 236
rect 158 202 795 218
rect 882 202 916 344
rect 950 349 1031 365
rect 950 315 962 349
rect 996 315 1031 349
rect 950 236 1031 315
rect 882 186 1033 202
rect 25 152 762 168
rect 25 134 428 152
rect 412 118 428 134
rect 462 134 728 152
rect 462 118 478 134
rect 412 106 478 118
rect 712 118 728 134
rect 712 102 762 118
rect 798 152 848 168
rect 798 118 814 152
rect 310 84 376 100
rect 310 50 326 84
rect 360 50 376 84
rect 310 17 376 50
rect 514 84 676 100
rect 514 50 530 84
rect 564 50 626 84
rect 660 50 676 84
rect 514 17 676 50
rect 798 17 848 118
rect 882 152 900 186
rect 934 152 983 186
rect 1017 152 1033 186
rect 882 118 1033 152
rect 882 84 900 118
rect 934 84 983 118
rect 1017 84 1033 118
rect 882 69 1033 84
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 683 1056 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 0 617 1056 649
rect 0 17 1056 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -49 1056 -17
<< labels >>
flabel pwell s 0 0 1056 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 0 617 1056 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
rlabel comment s 0 0 0 0 4 nor2b_4
flabel metal1 s 0 617 1056 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 1056 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 223 242 257 276 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 319 242 353 276 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 991 242 1025 276 0 FreeSans 340 0 0 0 B_N
port 2 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 B_N
port 2 nsew
flabel corelocali s 31 168 65 202 0 FreeSans 340 0 0 0 Y
port 7 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 Y
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 1056 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1546732
string GDS_START 1538454
<< end >>
