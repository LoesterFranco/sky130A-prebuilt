magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 125 333 176 493
rect 317 333 368 490
rect 515 333 560 493
rect 701 333 752 490
rect 893 333 941 490
rect 1091 333 1166 490
rect 1315 333 1365 490
rect 1507 333 1557 490
rect 1699 333 1749 490
rect 1891 333 1941 490
rect 2083 333 2131 490
rect 2275 333 2326 490
rect 125 291 2326 333
rect 515 283 1941 291
rect 69 221 335 255
rect 369 221 437 255
rect 69 179 471 221
rect 515 56 560 283
rect 701 56 752 283
rect 893 56 941 283
rect 1091 56 1161 283
rect 1315 56 1365 283
rect 1507 56 1557 283
rect 1699 56 1749 283
rect 1891 56 1941 283
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2484 561
rect 28 299 81 527
rect 220 367 272 527
rect 413 367 464 527
rect 604 367 656 527
rect 797 367 848 527
rect 993 367 1044 527
rect 1218 424 1270 527
rect 1218 367 1269 424
rect 1411 367 1462 527
rect 1603 367 1654 527
rect 1795 367 1846 527
rect 1987 367 2038 527
rect 2179 367 2230 527
rect 2370 367 2422 527
rect 411 17 465 122
rect 604 17 657 122
rect 796 17 849 122
rect 993 17 1046 122
rect 1218 17 1271 122
rect 1410 17 1455 122
rect 1602 17 1655 122
rect 1794 17 1847 122
rect 1986 221 2079 255
rect 2113 221 2181 255
rect 2215 221 2382 255
rect 1986 179 2382 221
rect 1986 17 2039 122
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2484 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 335 221 369 255
rect 437 221 471 255
rect 2079 221 2113 255
rect 2181 221 2215 255
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
<< metal1 >>
rect 0 561 2484 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2484 561
rect 0 496 2484 527
rect 0 17 2484 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2484 17
rect 0 -48 2484 -17
<< obsm1 >>
rect 323 255 483 261
rect 323 221 335 255
rect 369 221 437 255
rect 471 252 483 255
rect 2057 255 2227 261
rect 2057 252 2079 255
rect 471 224 2079 252
rect 471 221 483 224
rect 323 215 483 221
rect 2057 221 2079 224
rect 2113 221 2181 255
rect 2215 221 2227 255
rect 2057 215 2227 221
<< labels >>
rlabel locali s 69 179 471 255 6 A
port 1 nsew signal input
rlabel locali s 2275 333 2326 490 6 Y
port 2 nsew signal output
rlabel locali s 2083 333 2131 490 6 Y
port 2 nsew signal output
rlabel locali s 1891 333 1941 490 6 Y
port 2 nsew signal output
rlabel locali s 1891 56 1941 283 6 Y
port 2 nsew signal output
rlabel locali s 1699 333 1749 490 6 Y
port 2 nsew signal output
rlabel locali s 1699 56 1749 283 6 Y
port 2 nsew signal output
rlabel locali s 1507 333 1557 490 6 Y
port 2 nsew signal output
rlabel locali s 1507 56 1557 283 6 Y
port 2 nsew signal output
rlabel locali s 1315 333 1365 490 6 Y
port 2 nsew signal output
rlabel locali s 1315 56 1365 283 6 Y
port 2 nsew signal output
rlabel locali s 1091 333 1166 490 6 Y
port 2 nsew signal output
rlabel locali s 1091 56 1161 283 6 Y
port 2 nsew signal output
rlabel locali s 893 333 941 490 6 Y
port 2 nsew signal output
rlabel locali s 893 56 941 283 6 Y
port 2 nsew signal output
rlabel locali s 701 333 752 490 6 Y
port 2 nsew signal output
rlabel locali s 701 56 752 283 6 Y
port 2 nsew signal output
rlabel locali s 515 333 560 493 6 Y
port 2 nsew signal output
rlabel locali s 515 283 1941 291 6 Y
port 2 nsew signal output
rlabel locali s 515 56 560 283 6 Y
port 2 nsew signal output
rlabel locali s 317 333 368 490 6 Y
port 2 nsew signal output
rlabel locali s 125 333 176 493 6 Y
port 2 nsew signal output
rlabel locali s 125 291 2326 333 6 Y
port 2 nsew signal output
rlabel metal1 s 0 -48 2484 48 8 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 496 2484 592 6 VPWR
port 4 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2484 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1797500
string GDS_START 1783280
<< end >>
