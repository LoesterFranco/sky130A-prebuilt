magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 2024 561
rect 126 367 176 527
rect 294 435 344 527
rect 462 435 512 527
rect 630 435 680 527
rect 904 435 954 527
rect 1072 435 1122 527
rect 1592 409 1650 493
rect 1232 357 1650 409
rect 1684 367 1734 527
rect 1592 333 1650 357
rect 1768 333 1818 493
rect 1852 367 1902 527
rect 1936 333 2007 493
rect 337 289 1146 323
rect 1592 289 2007 333
rect 337 255 371 289
rect 1112 255 1146 289
rect 98 215 371 255
rect 435 215 1078 255
rect 1112 215 1486 255
rect 1963 181 2007 289
rect 470 17 504 111
rect 638 17 672 111
rect 807 17 862 181
rect 996 17 1030 111
rect 1164 17 1198 111
rect 1332 17 1366 111
rect 1500 17 1554 111
rect 1676 129 2007 181
rect 0 -17 2024 17
<< obsli1 >>
rect 17 323 92 493
rect 210 401 260 493
rect 378 401 428 493
rect 546 401 596 493
rect 714 401 764 493
rect 210 357 764 401
rect 807 401 870 493
rect 988 401 1038 493
rect 1156 443 1550 493
rect 1156 401 1198 443
rect 807 357 1198 401
rect 210 323 260 357
rect 17 289 213 323
rect 247 289 260 323
rect 1180 289 1225 323
rect 1259 289 1554 323
rect 17 181 64 289
rect 1520 255 1554 289
rect 1520 215 1929 255
rect 17 129 352 181
rect 386 145 772 181
rect 386 95 436 145
rect 34 51 436 95
rect 538 51 604 145
rect 706 51 772 145
rect 896 147 1642 181
rect 896 145 1486 147
rect 896 51 962 145
rect 1064 51 1130 145
rect 1232 51 1298 145
rect 1400 51 1466 145
rect 1592 95 1642 147
rect 1592 61 1994 95
<< obsli1c >>
rect 213 289 247 323
rect 1225 289 1259 323
<< metal1 >>
rect 0 496 2024 592
rect 0 -48 2024 48
<< obsm1 >>
rect 201 323 259 329
rect 201 289 213 323
rect 247 320 259 323
rect 1213 323 1271 329
rect 1213 320 1225 323
rect 247 292 1225 320
rect 247 289 259 292
rect 201 283 259 289
rect 1213 289 1225 292
rect 1259 289 1271 323
rect 1213 283 1271 289
<< labels >>
rlabel locali s 435 215 1078 255 6 A
port 1 nsew signal input
rlabel locali s 1112 255 1146 289 6 B
port 2 nsew signal input
rlabel locali s 1112 215 1486 255 6 B
port 2 nsew signal input
rlabel locali s 337 289 1146 323 6 B
port 2 nsew signal input
rlabel locali s 337 255 371 289 6 B
port 2 nsew signal input
rlabel locali s 98 215 371 255 6 B
port 2 nsew signal input
rlabel locali s 1963 181 2007 289 6 Y
port 3 nsew signal output
rlabel locali s 1936 333 2007 493 6 Y
port 3 nsew signal output
rlabel locali s 1768 333 1818 493 6 Y
port 3 nsew signal output
rlabel locali s 1676 129 2007 181 6 Y
port 3 nsew signal output
rlabel locali s 1592 409 1650 493 6 Y
port 3 nsew signal output
rlabel locali s 1592 333 1650 357 6 Y
port 3 nsew signal output
rlabel locali s 1592 289 2007 333 6 Y
port 3 nsew signal output
rlabel locali s 1232 357 1650 409 6 Y
port 3 nsew signal output
rlabel locali s 1500 17 1554 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 1332 17 1366 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 1164 17 1198 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 996 17 1030 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 807 17 862 181 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 638 17 672 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 470 17 504 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 2024 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 2024 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 1852 367 1902 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 1684 367 1734 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 1072 435 1122 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 904 435 954 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 630 435 680 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 462 435 512 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 294 435 344 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 126 367 176 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 2024 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 2024 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2024 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 618256
string GDS_START 604216
<< end >>
