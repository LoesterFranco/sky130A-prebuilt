magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1196 561
rect 115 359 165 527
rect 283 359 333 527
rect 703 393 753 425
rect 871 393 921 425
rect 703 391 921 393
rect 1123 391 1179 493
rect 703 357 1179 391
rect 703 289 1033 323
rect 703 257 737 289
rect 18 215 365 257
rect 419 215 737 257
rect 999 257 1033 289
rect 771 215 953 255
rect 999 215 1083 257
rect 1121 181 1179 357
rect 18 17 73 181
rect 107 145 1179 181
rect 107 51 173 145
rect 207 17 241 111
rect 275 51 341 145
rect 375 17 409 111
rect 443 51 509 145
rect 543 17 577 111
rect 611 51 677 145
rect 711 17 745 111
rect 779 51 845 145
rect 879 17 913 111
rect 947 51 1013 145
rect 1047 17 1081 111
rect 1121 51 1179 145
rect 0 -17 1196 17
<< obsli1 >>
rect 30 325 81 493
rect 199 325 249 493
rect 367 459 585 493
rect 367 425 489 459
rect 523 425 585 459
rect 367 417 585 425
rect 367 325 417 417
rect 30 291 417 325
rect 451 325 501 383
rect 535 359 585 417
rect 619 459 1005 493
rect 619 325 669 459
rect 787 427 837 459
rect 955 427 1005 459
rect 1039 459 1089 493
rect 1039 425 1041 459
rect 1075 425 1089 459
rect 451 291 669 325
<< obsli1c >>
rect 489 425 523 459
rect 1041 425 1075 459
<< metal1 >>
rect 0 496 1196 592
rect 0 -48 1196 48
<< obsm1 >>
rect 477 459 536 467
rect 477 425 489 459
rect 523 456 536 459
rect 1029 459 1088 467
rect 1029 456 1041 459
rect 523 428 1041 456
rect 523 425 536 428
rect 477 413 536 425
rect 1029 425 1041 428
rect 1075 425 1088 459
rect 1029 413 1088 425
<< labels >>
rlabel locali s 18 215 365 257 6 A
port 1 nsew signal input
rlabel locali s 999 257 1033 289 6 B
port 2 nsew signal input
rlabel locali s 999 215 1083 257 6 B
port 2 nsew signal input
rlabel locali s 703 289 1033 323 6 B
port 2 nsew signal input
rlabel locali s 703 257 737 289 6 B
port 2 nsew signal input
rlabel locali s 419 215 737 257 6 B
port 2 nsew signal input
rlabel locali s 771 215 953 255 6 C
port 3 nsew signal input
rlabel locali s 1123 391 1179 493 6 Y
port 4 nsew signal output
rlabel locali s 1121 181 1179 357 6 Y
port 4 nsew signal output
rlabel locali s 1121 51 1179 145 6 Y
port 4 nsew signal output
rlabel locali s 947 51 1013 145 6 Y
port 4 nsew signal output
rlabel locali s 871 393 921 425 6 Y
port 4 nsew signal output
rlabel locali s 779 51 845 145 6 Y
port 4 nsew signal output
rlabel locali s 703 393 753 425 6 Y
port 4 nsew signal output
rlabel locali s 703 391 921 393 6 Y
port 4 nsew signal output
rlabel locali s 703 357 1179 391 6 Y
port 4 nsew signal output
rlabel locali s 611 51 677 145 6 Y
port 4 nsew signal output
rlabel locali s 443 51 509 145 6 Y
port 4 nsew signal output
rlabel locali s 275 51 341 145 6 Y
port 4 nsew signal output
rlabel locali s 107 145 1179 181 6 Y
port 4 nsew signal output
rlabel locali s 107 51 173 145 6 Y
port 4 nsew signal output
rlabel locali s 1047 17 1081 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 879 17 913 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 711 17 745 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 543 17 577 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 375 17 409 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 207 17 241 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 18 17 73 181 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 1196 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1196 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 283 359 333 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 115 359 165 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 1196 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 1196 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1988588
string GDS_START 1979272
<< end >>
