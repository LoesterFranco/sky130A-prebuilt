magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 17 425 275 483
rect 121 265 169 323
rect 468 299 523 493
rect 17 199 86 265
rect 121 199 298 265
rect 489 152 523 299
rect 468 83 523 152
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 21 357 275 391
rect 319 367 375 527
rect 21 299 86 357
rect 241 333 275 357
rect 241 299 395 333
rect 361 165 395 299
rect 20 131 395 165
rect 20 61 71 131
rect 105 17 181 97
rect 225 61 259 131
rect 293 17 379 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
rlabel locali s 121 265 169 323 6 A
port 1 nsew signal input
rlabel locali s 121 199 298 265 6 A
port 1 nsew signal input
rlabel locali s 17 425 275 483 6 B
port 2 nsew signal input
rlabel locali s 17 199 86 265 6 C
port 3 nsew signal input
rlabel locali s 489 152 523 299 6 X
port 4 nsew signal output
rlabel locali s 468 299 523 493 6 X
port 4 nsew signal output
rlabel locali s 468 83 523 152 6 X
port 4 nsew signal output
rlabel metal1 s 0 -48 552 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 552 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 552 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 458900
string GDS_START 453638
<< end >>
