magic
tech sky130A
magscale 1 2
timestamp 1604502697
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 89 47 119 131
rect 186 47 216 177
rect 280 47 310 177
rect 374 47 404 177
rect 478 47 508 177
rect 572 47 602 177
rect 656 47 686 177
rect 762 47 792 177
<< pmoshvt >>
rect 81 360 117 444
rect 188 297 224 497
rect 282 297 318 497
rect 376 297 412 497
rect 470 297 506 497
rect 564 297 600 497
rect 658 297 694 497
rect 764 297 800 497
<< ndiff >>
rect 134 131 186 177
rect 27 108 89 131
rect 27 74 35 108
rect 69 74 89 108
rect 27 47 89 74
rect 119 97 186 131
rect 119 63 134 97
rect 168 63 186 97
rect 119 47 186 63
rect 216 164 280 177
rect 216 130 236 164
rect 270 130 280 164
rect 216 96 280 130
rect 216 62 236 96
rect 270 62 280 96
rect 216 47 280 62
rect 310 97 374 177
rect 310 63 330 97
rect 364 63 374 97
rect 310 47 374 63
rect 404 101 478 177
rect 404 67 414 101
rect 448 67 478 101
rect 404 47 478 67
rect 508 97 572 177
rect 508 63 518 97
rect 552 63 572 97
rect 508 47 572 63
rect 602 165 656 177
rect 602 131 612 165
rect 646 131 656 165
rect 602 47 656 131
rect 686 97 762 177
rect 686 63 706 97
rect 740 63 762 97
rect 686 47 762 63
rect 792 165 854 177
rect 792 131 812 165
rect 846 131 854 165
rect 792 47 854 131
<< pdiff >>
rect 134 476 188 497
rect 134 444 142 476
rect 27 412 81 444
rect 27 378 35 412
rect 69 378 81 412
rect 27 360 81 378
rect 117 442 142 444
rect 176 442 188 476
rect 117 360 188 442
rect 134 297 188 360
rect 224 340 282 497
rect 224 306 236 340
rect 270 306 282 340
rect 224 297 282 306
rect 318 476 376 497
rect 318 442 330 476
rect 364 442 376 476
rect 318 297 376 442
rect 412 340 470 497
rect 412 306 424 340
rect 458 306 470 340
rect 412 297 470 306
rect 506 476 564 497
rect 506 442 518 476
rect 552 442 564 476
rect 506 297 564 442
rect 600 297 658 497
rect 694 297 764 497
rect 800 476 854 497
rect 800 442 812 476
rect 846 442 854 476
rect 800 297 854 442
<< ndiffc >>
rect 35 74 69 108
rect 134 63 168 97
rect 236 130 270 164
rect 236 62 270 96
rect 330 63 364 97
rect 414 67 448 101
rect 518 63 552 97
rect 612 131 646 165
rect 706 63 740 97
rect 812 131 846 165
<< pdiffc >>
rect 35 378 69 412
rect 142 442 176 476
rect 236 306 270 340
rect 330 442 364 476
rect 424 306 458 340
rect 518 442 552 476
rect 812 442 846 476
<< poly >>
rect 188 497 224 523
rect 282 497 318 523
rect 376 497 412 523
rect 470 497 506 523
rect 564 497 600 523
rect 658 497 694 523
rect 764 497 800 523
rect 81 444 117 470
rect 81 345 117 360
rect 79 265 119 345
rect 188 282 224 297
rect 282 282 318 297
rect 376 282 412 297
rect 470 282 506 297
rect 564 282 600 297
rect 658 282 694 297
rect 764 282 800 297
rect 22 249 119 265
rect 22 215 35 249
rect 69 215 119 249
rect 22 199 119 215
rect 89 131 119 199
rect 186 265 226 282
rect 280 265 320 282
rect 374 265 414 282
rect 468 265 508 282
rect 562 265 602 282
rect 656 265 696 282
rect 762 265 802 282
rect 186 249 508 265
rect 186 215 308 249
rect 342 215 386 249
rect 420 215 464 249
rect 498 215 508 249
rect 186 199 508 215
rect 550 249 614 265
rect 550 215 560 249
rect 594 215 614 249
rect 550 199 614 215
rect 656 249 720 265
rect 656 215 666 249
rect 700 215 720 249
rect 656 199 720 215
rect 762 249 826 265
rect 762 215 772 249
rect 806 215 826 249
rect 762 199 826 215
rect 186 177 216 199
rect 280 177 310 199
rect 374 177 404 199
rect 478 177 508 199
rect 572 177 602 199
rect 656 177 686 199
rect 762 177 792 199
rect 89 21 119 47
rect 186 21 216 47
rect 280 21 310 47
rect 374 21 404 47
rect 478 21 508 47
rect 572 21 602 47
rect 656 21 686 47
rect 762 21 792 47
<< polycont >>
rect 35 215 69 249
rect 308 215 342 249
rect 386 215 420 249
rect 464 215 498 249
rect 560 215 594 249
rect 666 215 700 249
rect 772 215 806 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 120 476 192 527
rect 17 412 69 444
rect 120 442 142 476
rect 176 442 192 476
rect 304 476 380 527
rect 304 442 330 476
rect 364 442 380 476
rect 491 476 569 527
rect 491 442 518 476
rect 552 442 569 476
rect 774 476 891 485
rect 774 442 812 476
rect 846 442 891 476
rect 17 378 35 412
rect 69 378 806 408
rect 17 374 806 378
rect 17 362 163 374
rect 17 249 85 328
rect 17 215 35 249
rect 69 215 85 249
rect 129 181 163 362
rect 17 147 163 181
rect 202 306 236 340
rect 270 306 424 340
rect 458 306 484 340
rect 202 283 484 306
rect 202 181 254 283
rect 560 249 622 340
rect 288 215 308 249
rect 342 215 386 249
rect 420 215 464 249
rect 498 215 523 249
rect 202 164 448 181
rect 17 108 69 147
rect 202 130 236 164
rect 270 147 448 164
rect 270 130 286 147
rect 17 74 35 108
rect 17 58 69 74
rect 134 97 168 113
rect 134 17 168 63
rect 202 96 286 130
rect 202 62 236 96
rect 270 62 286 96
rect 202 57 286 62
rect 330 97 364 113
rect 330 17 364 63
rect 401 101 448 147
rect 489 165 523 215
rect 594 215 622 249
rect 560 199 622 215
rect 666 249 714 340
rect 700 215 714 249
rect 666 199 714 215
rect 772 249 806 374
rect 772 199 806 215
rect 850 165 891 442
rect 489 131 612 165
rect 646 131 812 165
rect 846 131 891 165
rect 401 67 414 101
rect 401 51 448 67
rect 492 63 518 97
rect 552 63 568 97
rect 492 17 568 63
rect 680 63 706 97
rect 740 63 768 97
rect 680 17 768 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel corelocali s 579 289 613 323 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 672 221 706 255 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 400 0 0 0 C_N
port 3 nsew
flabel corelocali s 438 289 472 323 0 FreeSans 200 180 0 0 X
port 8 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
rlabel comment s 0 0 0 0 4 or3b_4
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 491918
string GDS_START 485228
<< end >>
