magic
tech sky130A
magscale 1 2
timestamp 1601050088
<< locali >>
rect 85 302 219 360
rect 935 458 1031 582
rect 935 244 985 458
rect 1978 370 2279 420
rect 2192 252 2279 370
rect 2192 236 2357 252
rect 2095 202 2357 236
rect 2684 404 2750 596
rect 2884 404 2951 596
rect 2684 370 2951 404
rect 2527 270 2596 356
rect 2899 236 2949 370
rect 2711 202 2949 236
rect 2711 96 2761 202
rect 2899 96 2949 202
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3072 683
rect 17 394 73 596
rect 113 394 163 649
rect 203 560 269 596
rect 315 594 383 649
rect 633 560 699 592
rect 203 526 699 560
rect 203 394 269 526
rect 17 268 51 394
rect 267 268 333 330
rect 17 234 333 268
rect 17 70 73 234
rect 367 200 401 526
rect 846 492 901 534
rect 435 458 901 492
rect 435 358 501 458
rect 109 17 159 200
rect 195 192 401 200
rect 195 158 427 192
rect 195 70 261 158
rect 307 17 359 124
rect 393 85 427 158
rect 461 125 495 358
rect 541 356 592 424
rect 675 387 806 424
rect 846 387 901 458
rect 541 310 641 356
rect 675 276 709 387
rect 531 242 709 276
rect 743 310 833 353
rect 531 125 597 242
rect 631 85 683 208
rect 743 126 777 310
rect 867 262 901 387
rect 813 209 901 262
rect 1065 458 1131 649
rect 1171 424 1205 596
rect 1019 390 1205 424
rect 1239 581 1743 615
rect 1823 590 1937 649
rect 2085 590 2151 649
rect 2299 590 2425 649
rect 1239 430 1273 581
rect 1307 498 1357 547
rect 1398 545 1575 581
rect 1709 556 1743 581
rect 2459 556 2543 572
rect 1307 464 1507 498
rect 1239 396 1297 430
rect 1019 184 1053 390
rect 1087 275 1127 356
rect 1177 310 1229 356
rect 1087 218 1161 275
rect 1019 175 1081 184
rect 1195 175 1229 310
rect 1263 243 1297 396
rect 1331 281 1415 430
rect 1473 257 1507 464
rect 1541 330 1575 545
rect 1609 488 1675 547
rect 1709 522 2543 556
rect 1609 454 2425 488
rect 1609 419 1675 454
rect 1716 380 1843 420
rect 1809 355 1843 380
rect 1541 296 1775 330
rect 1641 264 1775 296
rect 1809 310 1895 355
rect 1263 209 1439 243
rect 1373 203 1439 209
rect 1473 221 1537 257
rect 1473 187 1775 221
rect 1809 187 1843 310
rect 1956 270 2142 336
rect 1956 236 1990 270
rect 1877 202 1990 236
rect 811 141 1081 175
rect 393 51 683 85
rect 811 51 877 141
rect 917 17 983 107
rect 1019 85 1081 141
rect 1175 119 1241 175
rect 1275 153 1341 169
rect 1741 153 1775 187
rect 1877 153 1911 202
rect 2391 168 2425 454
rect 2459 390 2543 522
rect 2584 390 2650 649
rect 2784 438 2850 649
rect 2459 236 2493 390
rect 2643 270 2865 336
rect 2459 202 2571 236
rect 2643 168 2677 270
rect 2990 364 3040 649
rect 1275 119 1707 153
rect 1741 119 1911 153
rect 1945 134 2677 168
rect 1673 85 1707 119
rect 1945 85 1979 134
rect 1019 51 1639 85
rect 1673 51 1979 85
rect 2013 17 2063 100
rect 2193 17 2259 100
rect 2393 17 2459 100
rect 2607 17 2675 100
rect 2797 17 2863 168
rect 2983 17 3049 252
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3072 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
<< metal1 >>
rect 0 683 3072 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3072 683
rect 0 617 3072 649
rect 0 17 3072 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3072 17
rect 0 -49 3072 -17
<< obsm1 >>
rect 691 421 749 430
rect 1363 421 1421 430
rect 691 393 1421 421
rect 691 384 749 393
rect 1363 384 1421 393
rect 595 347 653 356
rect 787 347 845 356
rect 1075 347 1133 356
rect 595 319 1133 347
rect 595 310 653 319
rect 787 310 845 319
rect 1075 310 1133 319
rect 1171 347 1229 356
rect 1843 347 1901 356
rect 1171 319 1901 347
rect 1171 310 1229 319
rect 1843 310 1901 319
<< labels >>
rlabel locali s 85 302 219 360 6 A
port 1 nsew signal input
rlabel locali s 935 458 1031 582 6 B
port 2 nsew signal input
rlabel locali s 935 244 985 458 6 B
port 2 nsew signal input
rlabel locali s 2527 270 2596 356 6 CI
port 3 nsew signal input
rlabel locali s 2192 252 2279 370 6 COUT
port 4 nsew signal output
rlabel locali s 2192 236 2357 252 6 COUT
port 4 nsew signal output
rlabel locali s 2095 202 2357 236 6 COUT
port 4 nsew signal output
rlabel locali s 1978 370 2279 420 6 COUT
port 4 nsew signal output
rlabel locali s 2899 236 2949 370 6 SUM
port 5 nsew signal output
rlabel locali s 2899 96 2949 202 6 SUM
port 5 nsew signal output
rlabel locali s 2884 404 2951 596 6 SUM
port 5 nsew signal output
rlabel locali s 2711 202 2949 236 6 SUM
port 5 nsew signal output
rlabel locali s 2711 96 2761 202 6 SUM
port 5 nsew signal output
rlabel locali s 2684 404 2750 596 6 SUM
port 5 nsew signal output
rlabel locali s 2684 370 2951 404 6 SUM
port 5 nsew signal output
rlabel metal1 s 0 -49 3072 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 3072 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 3072 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 2505984
string GDS_START 2484460
<< end >>
