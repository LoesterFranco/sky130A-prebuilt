magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 736 561
rect 17 299 85 493
rect 119 299 153 527
rect 207 367 257 527
rect 512 367 578 527
rect 17 177 52 299
rect 260 215 344 255
rect 378 215 444 255
rect 478 215 544 255
rect 17 51 85 177
rect 119 17 169 177
rect 307 17 352 109
rect 649 215 719 265
rect 0 -17 736 17
<< obsli1 >>
rect 386 333 452 493
rect 612 333 678 493
rect 191 299 678 333
rect 191 249 225 299
rect 86 215 225 249
rect 207 147 452 181
rect 207 51 273 147
rect 386 51 452 147
rect 578 173 612 299
rect 578 51 678 173
<< metal1 >>
rect 0 496 736 592
rect 0 -48 736 48
<< labels >>
rlabel locali s 260 215 344 255 6 A1
port 1 nsew signal input
rlabel locali s 378 215 444 255 6 A2
port 2 nsew signal input
rlabel locali s 478 215 544 255 6 B1
port 3 nsew signal input
rlabel locali s 649 215 719 265 6 C1
port 4 nsew signal input
rlabel locali s 17 299 85 493 6 X
port 5 nsew signal output
rlabel locali s 17 177 52 299 6 X
port 5 nsew signal output
rlabel locali s 17 51 85 177 6 X
port 5 nsew signal output
rlabel locali s 307 17 352 109 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 119 17 169 177 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 736 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 736 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 512 367 578 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 207 367 257 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 119 299 153 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 736 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 736 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1285988
string GDS_START 1279204
<< end >>
