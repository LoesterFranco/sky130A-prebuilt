magic
tech sky130A
magscale 1 2
timestamp 1599588232
<< locali >>
rect 85 314 217 360
rect 85 280 459 314
rect 277 88 359 246
rect 393 180 459 280
rect 561 190 641 324
rect 743 236 839 310
rect 2970 282 3021 596
rect 3373 364 3445 596
rect 2970 70 3047 282
rect 3411 226 3445 364
rect 3377 70 3445 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3391 683
rect 3425 649 3487 683
rect 3521 649 3552 683
rect 17 428 93 596
rect 127 462 193 649
rect 301 496 391 596
rect 499 530 569 649
rect 705 530 844 649
rect 878 581 1248 615
rect 301 462 777 496
rect 878 494 944 581
rect 17 394 421 428
rect 17 246 51 394
rect 355 362 421 394
rect 17 180 229 246
rect 17 70 89 180
rect 123 17 204 136
rect 493 146 527 462
rect 743 460 777 462
rect 978 460 1074 547
rect 615 392 709 428
rect 743 426 1074 460
rect 1108 459 1180 547
rect 615 358 944 392
rect 675 202 709 358
rect 878 270 944 358
rect 393 112 527 146
rect 393 80 470 112
rect 568 17 634 156
rect 675 68 730 202
rect 766 17 832 202
rect 866 85 932 202
rect 978 169 1012 426
rect 1046 258 1112 392
rect 978 119 1044 169
rect 1078 85 1112 258
rect 1146 160 1180 459
rect 1214 467 1248 581
rect 1282 501 1397 649
rect 1431 581 1633 615
rect 1431 467 1465 581
rect 1214 433 1465 467
rect 1499 459 1565 547
rect 1214 194 1261 433
rect 1499 399 1533 459
rect 1599 444 1633 581
rect 1667 478 1733 649
rect 1785 460 1851 596
rect 1885 494 1935 649
rect 1975 581 2221 615
rect 1975 460 2025 581
rect 1599 410 1713 444
rect 1785 426 2025 460
rect 1975 420 2025 426
rect 2065 442 2115 540
rect 2155 476 2221 581
rect 2273 577 2548 611
rect 2273 477 2324 577
rect 2364 462 2444 543
rect 2482 504 2548 577
rect 2588 504 2622 649
rect 2662 462 2728 596
rect 2774 496 2863 582
rect 2364 442 2795 462
rect 2065 428 2795 442
rect 1327 347 1533 399
rect 1567 350 1645 376
rect 1601 316 1645 350
rect 1295 279 1533 313
rect 1567 310 1645 316
rect 1295 160 1329 279
rect 1471 276 1533 279
rect 1679 303 1713 410
rect 2065 408 2478 428
rect 1747 374 1813 392
rect 1747 340 2410 374
rect 1747 337 1813 340
rect 2076 303 2278 306
rect 1363 208 1429 245
rect 1471 242 1610 276
rect 1679 269 2278 303
rect 1576 235 1610 242
rect 2076 240 2278 269
rect 1363 174 1542 208
rect 1576 180 1772 235
rect 1806 201 2042 235
rect 1146 94 1329 160
rect 866 51 1112 85
rect 1363 17 1430 140
rect 1476 70 1542 174
rect 1640 17 1706 136
rect 1806 70 1856 201
rect 1890 17 1956 167
rect 1992 85 2042 201
rect 2076 172 2310 206
rect 2344 180 2410 340
rect 2076 119 2142 172
rect 2276 146 2310 172
rect 2444 146 2478 408
rect 2513 226 2579 392
rect 2617 350 2687 394
rect 2617 316 2623 350
rect 2657 316 2687 350
rect 2617 260 2687 316
rect 2729 260 2795 428
rect 2829 226 2863 496
rect 2897 364 2931 649
rect 2513 192 2863 226
rect 3061 364 3127 649
rect 3173 326 3239 572
rect 3283 364 3333 649
rect 3479 364 3529 649
rect 2176 85 2242 138
rect 1992 51 2242 85
rect 2276 80 2478 146
rect 2652 17 2718 158
rect 2754 70 2820 192
rect 2870 17 2936 158
rect 3173 260 3377 326
rect 3081 17 3131 226
rect 3173 90 3244 260
rect 3291 17 3341 226
rect 3479 17 3529 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3552 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 3199 649 3233 683
rect 3295 649 3329 683
rect 3391 649 3425 683
rect 3487 649 3521 683
rect 1567 316 1601 350
rect 2623 316 2657 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
<< metal1 >>
rect 0 683 3552 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3391 683
rect 3425 649 3487 683
rect 3521 649 3552 683
rect 0 617 3552 649
rect 0 616 50 617
rect 1555 350 1613 356
rect 1555 316 1567 350
rect 1601 347 1613 350
rect 2611 350 2669 356
rect 2611 347 2623 350
rect 1601 319 2623 347
rect 1601 316 1613 319
rect 1555 310 1613 316
rect 2611 316 2623 319
rect 2657 316 2669 350
rect 2611 310 2669 316
rect 0 49 50 50
rect 0 17 3552 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3552 17
rect 0 -49 3552 -17
<< labels >>
rlabel locali s 277 88 359 246 6 D
port 1 nsew signal input
rlabel locali s 3411 226 3445 364 6 Q
port 2 nsew signal output
rlabel locali s 3377 70 3445 226 6 Q
port 2 nsew signal output
rlabel locali s 3373 364 3445 596 6 Q
port 2 nsew signal output
rlabel locali s 2970 282 3021 596 6 Q_N
port 3 nsew signal output
rlabel locali s 2970 70 3047 282 6 Q_N
port 3 nsew signal output
rlabel locali s 561 190 641 324 6 SCD
port 4 nsew signal input
rlabel locali s 393 180 459 280 6 SCE
port 5 nsew signal input
rlabel locali s 85 314 217 360 6 SCE
port 5 nsew signal input
rlabel locali s 85 280 459 314 6 SCE
port 5 nsew signal input
rlabel metal1 s 2611 347 2669 356 6 SET_B
port 6 nsew signal input
rlabel metal1 s 2611 310 2669 319 6 SET_B
port 6 nsew signal input
rlabel metal1 s 1555 347 1613 356 6 SET_B
port 6 nsew signal input
rlabel metal1 s 1555 319 2669 347 6 SET_B
port 6 nsew signal input
rlabel metal1 s 1555 310 1613 319 6 SET_B
port 6 nsew signal input
rlabel locali s 743 236 839 310 6 CLK
port 7 nsew clock input
rlabel metal1 s 0 -49 3552 49 8 VGND
port 8 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 9 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 10 nsew power bidirectional
rlabel metal1 s 0 617 3552 715 6 VPWR
port 11 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 3552 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 151104
string GDS_START 126196
<< end >>
