magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 644 561
rect 103 437 169 527
rect 30 153 90 323
rect 302 433 439 527
rect 301 329 440 391
rect 475 316 536 473
rect 573 336 627 527
rect 19 17 85 118
rect 501 155 536 316
rect 375 17 455 116
rect 489 51 536 155
rect 573 17 627 144
rect 0 -17 644 17
<< obsli1 >>
rect 35 403 69 489
rect 35 357 171 403
rect 124 227 171 357
rect 209 295 266 484
rect 209 265 381 295
rect 209 261 467 265
rect 124 161 235 227
rect 269 189 467 261
rect 124 131 167 161
rect 119 56 167 131
rect 269 122 303 189
rect 223 83 303 122
rect 223 54 257 83
<< metal1 >>
rect 0 496 644 592
rect 0 -48 644 48
<< labels >>
rlabel locali s 30 153 90 323 6 A_N
port 1 nsew signal input
rlabel locali s 301 329 440 391 6 B
port 2 nsew signal input
rlabel locali s 501 155 536 316 6 X
port 3 nsew signal output
rlabel locali s 489 51 536 155 6 X
port 3 nsew signal output
rlabel locali s 475 316 536 473 6 X
port 3 nsew signal output
rlabel locali s 573 17 627 144 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 375 17 455 116 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 19 17 85 118 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 644 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 644 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 573 336 627 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 302 433 439 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 103 437 169 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 644 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 644 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3768912
string GDS_START 3763308
<< end >>
