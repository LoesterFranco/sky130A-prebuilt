magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 828 561
rect 22 282 73 527
rect 107 359 158 493
rect 192 447 258 527
rect 432 447 513 527
rect 22 17 73 182
rect 107 165 141 359
rect 243 215 337 255
rect 371 181 405 220
rect 107 51 174 165
rect 303 154 405 181
rect 213 17 247 150
rect 303 147 404 154
rect 303 76 347 147
rect 671 265 705 485
rect 746 363 809 527
rect 594 215 705 265
rect 740 215 809 329
rect 675 17 709 111
rect 0 -17 828 17
<< obsli1 >>
rect 567 411 637 485
rect 220 377 637 411
rect 220 323 254 377
rect 175 289 254 323
rect 288 299 492 343
rect 175 199 209 289
rect 439 271 492 299
rect 526 299 637 377
rect 439 113 473 271
rect 526 249 560 299
rect 522 215 560 249
rect 522 138 556 215
rect 381 79 473 113
rect 507 64 556 138
rect 591 145 809 181
rect 591 64 637 145
rect 743 64 809 145
<< metal1 >>
rect 0 496 828 592
rect 0 -48 828 48
<< labels >>
rlabel locali s 243 215 337 255 6 A1_N
port 1 nsew signal input
rlabel locali s 371 181 405 220 6 A2_N
port 2 nsew signal input
rlabel locali s 303 154 405 181 6 A2_N
port 2 nsew signal input
rlabel locali s 303 147 404 154 6 A2_N
port 2 nsew signal input
rlabel locali s 303 76 347 147 6 A2_N
port 2 nsew signal input
rlabel locali s 740 215 809 329 6 B1
port 3 nsew signal input
rlabel locali s 671 265 705 485 6 B2
port 4 nsew signal input
rlabel locali s 594 215 705 265 6 B2
port 4 nsew signal input
rlabel locali s 107 359 158 493 6 X
port 5 nsew signal output
rlabel locali s 107 165 141 359 6 X
port 5 nsew signal output
rlabel locali s 107 51 174 165 6 X
port 5 nsew signal output
rlabel locali s 675 17 709 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 213 17 247 150 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 22 17 73 182 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 828 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 828 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 746 363 809 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 432 447 513 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 192 447 258 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 22 282 73 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 828 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 828 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1526168
string GDS_START 1519120
<< end >>
