magic
tech sky130A
magscale 1 2
timestamp 1601050088
<< locali >>
rect 113 424 179 596
rect 315 444 365 596
rect 811 444 845 547
rect 985 444 1051 547
rect 1386 504 1452 547
rect 1369 444 1452 504
rect 315 424 1452 444
rect 1566 424 1632 547
rect 113 410 1632 424
rect 113 390 365 410
rect 1369 390 1632 410
rect 315 364 365 390
rect 25 270 281 356
rect 315 236 349 364
rect 509 342 1200 376
rect 509 270 711 342
rect 837 236 1039 308
rect 1081 270 1200 342
rect 1242 252 1315 318
rect 1369 286 1607 356
rect 1657 252 1991 356
rect 109 202 349 236
rect 109 119 175 202
rect 281 119 349 202
rect 1281 218 1691 252
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 23 390 73 649
rect 213 458 279 649
rect 405 478 471 649
rect 505 512 571 596
rect 605 546 671 649
rect 705 581 1151 615
rect 705 512 771 581
rect 505 478 771 512
rect 885 478 951 581
rect 1085 478 1151 581
rect 1185 478 1251 649
rect 1285 581 1706 615
rect 1285 546 1352 581
rect 1285 530 1335 546
rect 1492 458 1526 581
rect 1672 424 1706 581
rect 1746 458 1796 649
rect 1836 424 1902 596
rect 1672 390 1902 424
rect 1942 390 1992 649
rect 23 85 75 236
rect 209 85 247 168
rect 383 202 803 236
rect 1081 202 1147 210
rect 383 154 631 202
rect 383 85 433 154
rect 667 120 701 168
rect 737 154 1147 202
rect 1181 184 1247 218
rect 1755 184 1993 218
rect 1181 150 1805 184
rect 1181 120 1247 150
rect 23 51 433 85
rect 479 70 1247 120
rect 1281 17 1347 116
rect 1381 70 1431 150
rect 1467 17 1533 116
rect 1567 70 1617 150
rect 1653 17 1721 116
rect 1755 70 1805 150
rect 1841 17 1907 150
rect 1943 70 1993 184
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
rlabel locali s 1657 252 1991 356 6 A1
port 1 nsew signal input
rlabel locali s 1281 218 1691 252 6 A1
port 1 nsew signal input
rlabel locali s 1242 252 1315 318 6 A1
port 1 nsew signal input
rlabel locali s 1369 286 1607 356 6 A2
port 2 nsew signal input
rlabel locali s 1081 270 1200 342 6 B1
port 3 nsew signal input
rlabel locali s 509 342 1200 376 6 B1
port 3 nsew signal input
rlabel locali s 509 270 711 342 6 B1
port 3 nsew signal input
rlabel locali s 837 236 1039 308 6 B2
port 4 nsew signal input
rlabel locali s 25 270 281 356 6 C1
port 5 nsew signal input
rlabel locali s 1566 424 1632 547 6 Y
port 6 nsew signal output
rlabel locali s 1386 504 1452 547 6 Y
port 6 nsew signal output
rlabel locali s 1369 444 1452 504 6 Y
port 6 nsew signal output
rlabel locali s 1369 390 1632 410 6 Y
port 6 nsew signal output
rlabel locali s 985 444 1051 547 6 Y
port 6 nsew signal output
rlabel locali s 811 444 845 547 6 Y
port 6 nsew signal output
rlabel locali s 315 444 365 596 6 Y
port 6 nsew signal output
rlabel locali s 315 424 1452 444 6 Y
port 6 nsew signal output
rlabel locali s 315 364 365 390 6 Y
port 6 nsew signal output
rlabel locali s 315 236 349 364 6 Y
port 6 nsew signal output
rlabel locali s 281 119 349 202 6 Y
port 6 nsew signal output
rlabel locali s 113 424 179 596 6 Y
port 6 nsew signal output
rlabel locali s 113 410 1632 424 6 Y
port 6 nsew signal output
rlabel locali s 113 390 365 410 6 Y
port 6 nsew signal output
rlabel locali s 109 202 349 236 6 Y
port 6 nsew signal output
rlabel locali s 109 119 175 202 6 Y
port 6 nsew signal output
rlabel metal1 s 0 -49 2016 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 617 2016 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2016 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1195944
string GDS_START 1180470
<< end >>
