magic
tech sky130A
magscale 1 2
timestamp 1601050047
<< nwell >>
rect -38 332 902 704
<< pwell >>
rect 0 0 864 49
<< scpmos >>
rect 86 368 116 592
rect 324 392 354 592
rect 424 392 454 592
rect 540 392 570 592
rect 630 392 660 592
rect 744 392 774 592
<< nmoslvt >>
rect 219 74 249 222
rect 333 74 363 222
rect 419 74 449 222
rect 513 74 543 222
rect 627 74 657 222
rect 741 74 771 222
<< ndiff >>
rect 27 188 219 222
rect 27 154 39 188
rect 73 154 174 188
rect 208 154 219 188
rect 27 120 219 154
rect 27 86 39 120
rect 73 86 174 120
rect 208 86 219 120
rect 27 74 219 86
rect 249 188 333 222
rect 249 154 274 188
rect 308 154 333 188
rect 249 120 333 154
rect 249 86 274 120
rect 308 86 333 120
rect 249 74 333 86
rect 363 210 419 222
rect 363 176 374 210
rect 408 176 419 210
rect 363 120 419 176
rect 363 86 374 120
rect 408 86 419 120
rect 363 74 419 86
rect 449 74 513 222
rect 543 74 627 222
rect 657 74 741 222
rect 771 196 828 222
rect 771 162 782 196
rect 816 162 828 196
rect 771 120 828 162
rect 771 86 782 120
rect 816 86 828 120
rect 771 74 828 86
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 497 86 546
rect 27 463 39 497
rect 73 463 86 497
rect 27 414 86 463
rect 27 380 39 414
rect 73 380 86 414
rect 27 368 86 380
rect 116 580 175 592
rect 116 546 129 580
rect 163 546 175 580
rect 116 497 175 546
rect 116 463 129 497
rect 163 463 175 497
rect 116 414 175 463
rect 116 380 129 414
rect 163 380 175 414
rect 265 580 324 592
rect 265 546 277 580
rect 311 546 324 580
rect 265 510 324 546
rect 265 476 277 510
rect 311 476 324 510
rect 265 440 324 476
rect 265 406 277 440
rect 311 406 324 440
rect 265 392 324 406
rect 354 580 424 592
rect 354 546 377 580
rect 411 546 424 580
rect 354 510 424 546
rect 354 476 377 510
rect 411 476 424 510
rect 354 440 424 476
rect 354 406 377 440
rect 411 406 424 440
rect 354 392 424 406
rect 454 580 540 592
rect 454 546 477 580
rect 511 546 540 580
rect 454 508 540 546
rect 454 474 477 508
rect 511 474 540 508
rect 454 392 540 474
rect 570 580 630 592
rect 570 546 583 580
rect 617 546 630 580
rect 570 509 630 546
rect 570 475 583 509
rect 617 475 630 509
rect 570 438 630 475
rect 570 404 583 438
rect 617 404 630 438
rect 570 392 630 404
rect 660 582 744 592
rect 660 548 683 582
rect 717 548 744 582
rect 660 514 744 548
rect 660 480 683 514
rect 717 480 744 514
rect 660 446 744 480
rect 660 412 683 446
rect 717 412 744 446
rect 660 392 744 412
rect 774 580 833 592
rect 774 546 787 580
rect 821 546 833 580
rect 774 509 833 546
rect 774 475 787 509
rect 821 475 833 509
rect 774 438 833 475
rect 774 404 787 438
rect 821 404 833 438
rect 774 392 833 404
rect 116 368 175 380
<< ndiffc >>
rect 39 154 73 188
rect 174 154 208 188
rect 39 86 73 120
rect 174 86 208 120
rect 274 154 308 188
rect 274 86 308 120
rect 374 176 408 210
rect 374 86 408 120
rect 782 162 816 196
rect 782 86 816 120
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 129 546 163 580
rect 129 463 163 497
rect 129 380 163 414
rect 277 546 311 580
rect 277 476 311 510
rect 277 406 311 440
rect 377 546 411 580
rect 377 476 411 510
rect 377 406 411 440
rect 477 546 511 580
rect 477 474 511 508
rect 583 546 617 580
rect 583 475 617 509
rect 583 404 617 438
rect 683 548 717 582
rect 683 480 717 514
rect 683 412 717 446
rect 787 546 821 580
rect 787 475 821 509
rect 787 404 821 438
<< poly >>
rect 86 592 116 618
rect 324 592 354 618
rect 424 592 454 618
rect 540 592 570 618
rect 630 592 660 618
rect 744 592 774 618
rect 324 377 354 392
rect 424 377 454 392
rect 540 377 570 392
rect 630 377 660 392
rect 744 377 774 392
rect 86 353 116 368
rect 321 356 357 377
rect 421 356 457 377
rect 83 310 119 353
rect 297 340 363 356
rect 83 294 249 310
rect 83 260 131 294
rect 165 260 199 294
rect 233 260 249 294
rect 297 306 313 340
rect 347 306 363 340
rect 297 290 363 306
rect 405 340 471 356
rect 405 306 421 340
rect 455 306 471 340
rect 537 310 573 377
rect 627 310 663 377
rect 741 310 777 377
rect 405 290 471 306
rect 513 294 579 310
rect 83 244 249 260
rect 219 222 249 244
rect 333 222 363 290
rect 419 222 449 290
rect 513 260 529 294
rect 563 260 579 294
rect 513 244 579 260
rect 627 294 693 310
rect 627 260 643 294
rect 677 260 693 294
rect 627 244 693 260
rect 741 294 843 310
rect 741 260 793 294
rect 827 260 843 294
rect 741 244 843 260
rect 513 222 543 244
rect 627 222 657 244
rect 741 222 771 244
rect 219 48 249 74
rect 333 48 363 74
rect 419 48 449 74
rect 513 48 543 74
rect 627 48 657 74
rect 741 48 771 74
<< polycont >>
rect 131 260 165 294
rect 199 260 233 294
rect 313 306 347 340
rect 421 306 455 340
rect 529 260 563 294
rect 643 260 677 294
rect 793 260 827 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 23 580 89 596
rect 23 546 39 580
rect 73 546 89 580
rect 23 497 89 546
rect 23 463 39 497
rect 73 463 89 497
rect 23 414 89 463
rect 23 380 39 414
rect 73 380 89 414
rect 23 364 89 380
rect 129 580 179 649
rect 163 546 179 580
rect 129 497 179 546
rect 163 463 179 497
rect 129 414 179 463
rect 163 380 179 414
rect 129 364 179 380
rect 229 580 327 596
rect 229 546 277 580
rect 311 546 327 580
rect 229 510 327 546
rect 229 476 277 510
rect 311 476 327 510
rect 229 440 327 476
rect 229 406 277 440
rect 311 406 327 440
rect 229 390 327 406
rect 361 580 427 596
rect 361 546 377 580
rect 411 546 427 580
rect 361 510 427 546
rect 361 476 377 510
rect 411 476 427 510
rect 361 440 427 476
rect 461 580 527 649
rect 461 546 477 580
rect 511 546 527 580
rect 461 508 527 546
rect 461 474 477 508
rect 511 474 527 508
rect 461 458 527 474
rect 567 580 633 596
rect 567 546 583 580
rect 617 546 633 580
rect 567 509 633 546
rect 567 475 583 509
rect 617 475 633 509
rect 361 406 377 440
rect 411 424 427 440
rect 567 438 633 475
rect 567 424 583 438
rect 411 406 583 424
rect 361 404 583 406
rect 617 404 633 438
rect 667 582 733 649
rect 667 548 683 582
rect 717 548 733 582
rect 667 514 733 548
rect 667 480 683 514
rect 717 480 733 514
rect 667 446 733 480
rect 667 412 683 446
rect 717 412 733 446
rect 771 580 837 596
rect 771 546 787 580
rect 821 546 837 580
rect 771 509 837 546
rect 771 475 787 509
rect 821 475 837 509
rect 771 438 837 475
rect 361 390 633 404
rect 23 188 71 364
rect 229 310 263 390
rect 567 378 633 390
rect 771 404 787 438
rect 821 404 837 438
rect 771 378 837 404
rect 115 294 263 310
rect 115 260 131 294
rect 165 260 199 294
rect 233 260 263 294
rect 297 340 363 356
rect 297 306 313 340
rect 347 306 363 340
rect 297 290 363 306
rect 405 340 471 356
rect 567 344 837 378
rect 405 306 421 340
rect 455 306 471 340
rect 405 290 471 306
rect 505 294 579 310
rect 115 256 263 260
rect 505 260 529 294
rect 563 260 579 294
rect 115 222 424 256
rect 358 210 424 222
rect 23 154 39 188
rect 73 154 174 188
rect 208 154 224 188
rect 23 120 224 154
rect 23 86 39 120
rect 73 86 174 120
rect 208 86 224 120
rect 23 58 224 86
rect 258 154 274 188
rect 308 154 324 188
rect 258 120 324 154
rect 258 86 274 120
rect 308 86 324 120
rect 258 17 324 86
rect 358 176 374 210
rect 408 176 424 210
rect 358 120 424 176
rect 358 86 374 120
rect 408 86 424 120
rect 505 88 579 260
rect 627 294 743 310
rect 627 260 643 294
rect 677 260 743 294
rect 627 236 743 260
rect 777 294 843 310
rect 777 260 793 294
rect 827 260 843 294
rect 777 236 843 260
rect 766 196 832 202
rect 766 162 782 196
rect 816 162 832 196
rect 766 120 832 162
rect 358 70 424 86
rect 766 86 782 120
rect 816 86 832 120
rect 766 17 832 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a41o_1
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 799 242 833 276 0 FreeSans 340 0 0 0 A4
port 4 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 511 94 545 128 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 511 168 545 202 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 511 242 545 276 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 703 242 737 276 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 B1
port 5 nsew
flabel corelocali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 864 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3901140
string GDS_START 3893096
<< end >>
