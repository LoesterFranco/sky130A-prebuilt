magic
tech sky130A
magscale 1 2
timestamp 1604502741
<< locali >>
rect 314 424 360 547
rect 314 394 455 424
rect 612 394 662 547
rect 314 390 662 394
rect 409 360 662 390
rect 25 270 263 356
rect 297 270 363 356
rect 409 236 455 360
rect 697 326 743 356
rect 533 278 743 326
rect 533 260 667 278
rect 782 270 935 356
rect 123 202 455 236
rect 123 119 189 202
rect 323 119 389 202
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 24 424 74 596
rect 114 458 180 649
rect 214 581 460 615
rect 214 424 280 581
rect 24 390 280 424
rect 394 458 460 581
rect 506 581 736 615
rect 506 428 572 581
rect 702 424 736 581
rect 776 458 826 649
rect 866 424 932 596
rect 702 390 932 424
rect 23 85 89 226
rect 701 226 937 236
rect 491 202 937 226
rect 223 85 289 168
rect 491 192 751 202
rect 491 168 557 192
rect 423 85 557 168
rect 23 51 557 85
rect 591 17 657 158
rect 701 70 751 192
rect 785 17 851 168
rect 887 70 937 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
rlabel locali s 782 270 935 356 6 A1
port 1 nsew signal input
rlabel locali s 697 326 743 356 6 A2
port 2 nsew signal input
rlabel locali s 533 278 743 326 6 A2
port 2 nsew signal input
rlabel locali s 533 260 667 278 6 A2
port 2 nsew signal input
rlabel locali s 25 270 263 356 6 B1
port 3 nsew signal input
rlabel locali s 297 270 363 356 6 B2
port 4 nsew signal input
rlabel locali s 612 394 662 547 6 Y
port 5 nsew signal output
rlabel locali s 409 360 662 390 6 Y
port 5 nsew signal output
rlabel locali s 409 236 455 360 6 Y
port 5 nsew signal output
rlabel locali s 323 119 389 202 6 Y
port 5 nsew signal output
rlabel locali s 314 424 360 547 6 Y
port 5 nsew signal output
rlabel locali s 314 394 455 424 6 Y
port 5 nsew signal output
rlabel locali s 314 390 662 394 6 Y
port 5 nsew signal output
rlabel locali s 123 202 455 236 6 Y
port 5 nsew signal output
rlabel locali s 123 119 189 202 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -49 960 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 960 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1259526
string GDS_START 1251096
<< end >>
