magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 19 451 837 485
rect 19 97 64 451
rect 1272 285 1730 319
rect 118 199 247 265
rect 471 199 810 265
rect 1272 258 1306 285
rect 849 215 1306 258
rect 19 63 837 97
rect 1696 199 1730 285
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 875 451 941 527
rect 1053 451 1129 527
rect 1241 451 1317 527
rect 1361 417 1395 493
rect 1429 451 1505 527
rect 1549 417 1583 493
rect 1647 451 1713 527
rect 479 383 1583 417
rect 1361 359 1395 383
rect 1549 359 1583 383
rect 1757 359 1809 493
rect 103 315 1226 349
rect 1486 215 1662 249
rect 291 165 370 187
rect 1360 181 1420 187
rect 103 131 370 165
rect 479 131 1207 165
rect 875 17 941 93
rect 985 51 1019 131
rect 1053 17 1129 93
rect 1173 51 1207 131
rect 1360 143 1583 181
rect 1241 17 1316 118
rect 1360 51 1395 143
rect 1449 17 1499 109
rect 1549 102 1583 143
rect 1618 165 1662 215
rect 1774 165 1809 359
rect 1618 131 1809 165
rect 1647 17 1713 93
rect 1757 51 1809 131
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
<< metal1 >>
rect 0 561 1840 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 0 496 1840 527
rect 0 17 1840 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
rect 0 -48 1840 -17
<< obsm1 >>
rect 324 184 382 193
rect 1338 184 1406 193
rect 324 156 1406 184
rect 324 147 382 156
rect 1338 147 1406 156
<< labels >>
rlabel locali s 118 199 247 265 6 A0
port 1 nsew signal input
rlabel locali s 471 199 810 265 6 A1
port 2 nsew signal input
rlabel locali s 1696 199 1730 285 6 S
port 3 nsew signal input
rlabel locali s 1272 285 1730 319 6 S
port 3 nsew signal input
rlabel locali s 1272 258 1306 285 6 S
port 3 nsew signal input
rlabel locali s 849 215 1306 258 6 S
port 3 nsew signal input
rlabel locali s 19 451 837 485 6 Y
port 4 nsew signal output
rlabel locali s 19 97 64 451 6 Y
port 4 nsew signal output
rlabel locali s 19 63 837 97 6 Y
port 4 nsew signal output
rlabel metal1 s 0 -48 1840 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 1840 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1840 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2187082
string GDS_START 2174124
<< end >>
