magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 1602 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 89 47 119 131
rect 173 47 203 131
rect 381 47 411 131
rect 470 47 500 131
rect 574 47 604 119
rect 678 47 708 131
rect 750 47 780 131
rect 951 47 981 177
rect 1032 47 1062 177
rect 1139 47 1169 177
rect 1223 47 1253 177
rect 1327 47 1357 177
rect 1411 47 1441 177
<< pmoshvt >>
rect 81 363 117 491
rect 175 363 211 491
rect 373 369 409 497
rect 467 369 503 497
rect 572 413 608 497
rect 666 413 702 497
rect 762 413 798 497
rect 943 297 979 497
rect 1037 297 1073 497
rect 1131 297 1167 497
rect 1225 297 1261 497
rect 1319 297 1355 497
rect 1413 297 1449 497
<< ndiff >>
rect 37 106 89 131
rect 37 72 45 106
rect 79 72 89 106
rect 37 47 89 72
rect 119 93 173 131
rect 119 59 129 93
rect 163 59 173 93
rect 119 47 173 59
rect 203 106 255 131
rect 203 72 213 106
rect 247 72 255 106
rect 203 47 255 72
rect 329 119 381 131
rect 329 85 337 119
rect 371 85 381 119
rect 329 47 381 85
rect 411 89 470 131
rect 411 55 421 89
rect 455 55 470 89
rect 411 47 470 55
rect 500 119 550 131
rect 899 165 951 177
rect 899 131 907 165
rect 941 131 951 165
rect 628 119 678 131
rect 500 47 574 119
rect 604 106 678 119
rect 604 72 624 106
rect 658 72 678 106
rect 604 47 678 72
rect 708 47 750 131
rect 780 106 832 131
rect 780 72 790 106
rect 824 72 832 106
rect 780 47 832 72
rect 899 93 951 131
rect 899 59 907 93
rect 941 59 951 93
rect 899 47 951 59
rect 981 47 1032 177
rect 1062 161 1139 177
rect 1062 127 1079 161
rect 1113 127 1139 161
rect 1062 93 1139 127
rect 1062 59 1079 93
rect 1113 59 1139 93
rect 1062 47 1139 59
rect 1169 161 1223 177
rect 1169 127 1179 161
rect 1213 127 1223 161
rect 1169 93 1223 127
rect 1169 59 1179 93
rect 1213 59 1223 93
rect 1169 47 1223 59
rect 1253 93 1327 177
rect 1253 59 1275 93
rect 1309 59 1327 93
rect 1253 47 1327 59
rect 1357 161 1411 177
rect 1357 127 1367 161
rect 1401 127 1411 161
rect 1357 93 1411 127
rect 1357 59 1367 93
rect 1401 59 1411 93
rect 1357 47 1411 59
rect 1441 161 1493 177
rect 1441 127 1451 161
rect 1485 127 1493 161
rect 1441 93 1493 127
rect 1441 59 1451 93
rect 1485 59 1493 93
rect 1441 47 1493 59
<< pdiff >>
rect 27 477 81 491
rect 27 443 35 477
rect 69 443 81 477
rect 27 409 81 443
rect 27 375 35 409
rect 69 375 81 409
rect 27 363 81 375
rect 117 461 175 491
rect 117 427 129 461
rect 163 427 175 461
rect 117 363 175 427
rect 211 477 265 491
rect 211 443 223 477
rect 257 443 265 477
rect 211 409 265 443
rect 211 375 223 409
rect 257 375 265 409
rect 211 363 265 375
rect 319 483 373 497
rect 319 449 327 483
rect 361 449 373 483
rect 319 415 373 449
rect 319 381 327 415
rect 361 381 373 415
rect 319 369 373 381
rect 409 485 467 497
rect 409 451 421 485
rect 455 451 467 485
rect 409 417 467 451
rect 409 383 421 417
rect 455 383 467 417
rect 409 369 467 383
rect 503 413 572 497
rect 608 472 666 497
rect 608 438 620 472
rect 654 438 666 472
rect 608 413 666 438
rect 702 413 762 497
rect 798 477 943 497
rect 798 443 810 477
rect 844 443 892 477
rect 926 443 943 477
rect 798 413 943 443
rect 503 369 555 413
rect 886 297 943 413
rect 979 471 1037 497
rect 979 437 991 471
rect 1025 437 1037 471
rect 979 368 1037 437
rect 979 334 991 368
rect 1025 334 1037 368
rect 979 297 1037 334
rect 1073 485 1131 497
rect 1073 451 1085 485
rect 1119 451 1131 485
rect 1073 411 1131 451
rect 1073 377 1085 411
rect 1119 377 1131 411
rect 1073 297 1131 377
rect 1167 485 1225 497
rect 1167 451 1179 485
rect 1213 451 1225 485
rect 1167 417 1225 451
rect 1167 383 1179 417
rect 1213 383 1225 417
rect 1167 349 1225 383
rect 1167 315 1179 349
rect 1213 315 1225 349
rect 1167 297 1225 315
rect 1261 485 1319 497
rect 1261 451 1273 485
rect 1307 451 1319 485
rect 1261 417 1319 451
rect 1261 383 1273 417
rect 1307 383 1319 417
rect 1261 297 1319 383
rect 1355 485 1413 497
rect 1355 451 1367 485
rect 1401 451 1413 485
rect 1355 417 1413 451
rect 1355 383 1367 417
rect 1401 383 1413 417
rect 1355 349 1413 383
rect 1355 315 1367 349
rect 1401 315 1413 349
rect 1355 297 1413 315
rect 1449 485 1503 497
rect 1449 451 1461 485
rect 1495 451 1503 485
rect 1449 417 1503 451
rect 1449 383 1461 417
rect 1495 383 1503 417
rect 1449 349 1503 383
rect 1449 315 1461 349
rect 1495 315 1503 349
rect 1449 297 1503 315
<< ndiffc >>
rect 45 72 79 106
rect 129 59 163 93
rect 213 72 247 106
rect 337 85 371 119
rect 421 55 455 89
rect 907 131 941 165
rect 624 72 658 106
rect 790 72 824 106
rect 907 59 941 93
rect 1079 127 1113 161
rect 1079 59 1113 93
rect 1179 127 1213 161
rect 1179 59 1213 93
rect 1275 59 1309 93
rect 1367 127 1401 161
rect 1367 59 1401 93
rect 1451 127 1485 161
rect 1451 59 1485 93
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 129 427 163 461
rect 223 443 257 477
rect 223 375 257 409
rect 327 449 361 483
rect 327 381 361 415
rect 421 451 455 485
rect 421 383 455 417
rect 620 438 654 472
rect 810 443 844 477
rect 892 443 926 477
rect 991 437 1025 471
rect 991 334 1025 368
rect 1085 451 1119 485
rect 1085 377 1119 411
rect 1179 451 1213 485
rect 1179 383 1213 417
rect 1179 315 1213 349
rect 1273 451 1307 485
rect 1273 383 1307 417
rect 1367 451 1401 485
rect 1367 383 1401 417
rect 1367 315 1401 349
rect 1461 451 1495 485
rect 1461 383 1495 417
rect 1461 315 1495 349
<< poly >>
rect 81 491 117 517
rect 175 491 211 517
rect 373 497 409 523
rect 467 497 503 523
rect 572 497 608 523
rect 666 497 702 523
rect 762 497 798 523
rect 943 497 979 523
rect 1037 497 1073 523
rect 1131 497 1167 523
rect 1225 497 1261 523
rect 1319 497 1355 523
rect 1413 497 1449 523
rect 572 398 608 413
rect 666 398 702 413
rect 762 398 798 413
rect 81 348 117 363
rect 175 348 211 363
rect 373 354 409 369
rect 467 354 503 369
rect 45 318 119 348
rect 173 318 213 348
rect 45 280 87 318
rect 33 264 87 280
rect 173 274 203 318
rect 33 230 43 264
rect 77 230 87 264
rect 33 214 87 230
rect 129 264 203 274
rect 371 265 411 354
rect 129 230 145 264
rect 179 230 203 264
rect 129 220 203 230
rect 45 176 87 214
rect 45 146 119 176
rect 89 131 119 146
rect 173 131 203 220
rect 293 249 411 265
rect 293 215 303 249
rect 337 215 411 249
rect 465 219 505 354
rect 570 327 610 398
rect 664 375 704 398
rect 547 305 610 327
rect 652 365 718 375
rect 652 331 668 365
rect 702 331 718 365
rect 652 321 718 331
rect 760 373 800 398
rect 760 357 852 373
rect 760 323 804 357
rect 838 323 852 357
rect 547 271 557 305
rect 591 279 610 305
rect 760 307 852 323
rect 760 285 790 307
rect 591 271 708 279
rect 547 249 708 271
rect 293 199 411 215
rect 381 131 411 199
rect 453 203 507 219
rect 453 169 463 203
rect 497 169 507 203
rect 453 153 507 169
rect 556 197 622 207
rect 556 163 572 197
rect 606 163 622 197
rect 470 131 500 153
rect 556 147 622 163
rect 574 119 604 147
rect 678 131 708 249
rect 750 255 790 285
rect 943 282 979 297
rect 1037 282 1073 297
rect 1131 282 1167 297
rect 1225 282 1261 297
rect 1319 282 1355 297
rect 1413 282 1449 297
rect 941 265 981 282
rect 1035 265 1075 282
rect 1129 265 1169 282
rect 1223 265 1263 282
rect 1317 265 1357 282
rect 1411 265 1451 282
rect 750 131 780 255
rect 832 249 981 265
rect 832 215 842 249
rect 876 235 981 249
rect 876 215 886 235
rect 832 199 886 215
rect 951 177 981 235
rect 1023 249 1077 265
rect 1023 215 1033 249
rect 1067 215 1077 249
rect 1023 199 1077 215
rect 1119 249 1451 265
rect 1119 215 1129 249
rect 1163 215 1197 249
rect 1231 215 1451 249
rect 1119 199 1451 215
rect 1032 177 1062 199
rect 1139 177 1169 199
rect 1223 177 1253 199
rect 1327 177 1357 199
rect 1411 177 1441 199
rect 89 21 119 47
rect 173 21 203 47
rect 381 21 411 47
rect 470 21 500 47
rect 574 21 604 47
rect 678 21 708 47
rect 750 21 780 47
rect 951 21 981 47
rect 1032 21 1062 47
rect 1139 21 1169 47
rect 1223 21 1253 47
rect 1327 21 1357 47
rect 1411 21 1441 47
<< polycont >>
rect 43 230 77 264
rect 145 230 179 264
rect 303 215 337 249
rect 668 331 702 365
rect 804 323 838 357
rect 557 271 591 305
rect 463 169 497 203
rect 572 163 606 197
rect 842 215 876 249
rect 1033 215 1067 249
rect 1129 215 1163 249
rect 1197 215 1231 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 17 477 79 493
rect 17 443 35 477
rect 69 443 79 477
rect 17 409 79 443
rect 113 461 179 527
rect 113 427 129 461
rect 163 427 179 461
rect 213 477 267 493
rect 213 443 223 477
rect 257 443 267 477
rect 17 375 35 409
rect 69 393 79 409
rect 213 409 267 443
rect 69 391 179 393
rect 69 375 127 391
rect 17 359 127 375
rect 121 357 127 359
rect 161 357 179 391
rect 17 264 87 325
rect 17 230 43 264
rect 77 230 87 264
rect 17 197 87 230
rect 121 264 179 357
rect 121 230 145 264
rect 121 214 179 230
rect 213 375 223 409
rect 257 375 267 409
rect 213 323 267 375
rect 213 289 219 323
rect 253 289 267 323
rect 311 483 377 493
rect 311 449 327 483
rect 361 449 377 483
rect 311 415 377 449
rect 311 381 327 415
rect 361 381 377 415
rect 311 333 377 381
rect 411 485 465 527
rect 411 451 421 485
rect 455 451 465 485
rect 804 477 941 527
rect 411 417 465 451
rect 604 472 770 477
rect 604 438 620 472
rect 654 438 770 472
rect 604 433 770 438
rect 411 383 421 417
rect 455 383 465 417
rect 411 367 465 383
rect 625 391 702 399
rect 625 357 656 391
rect 690 365 702 391
rect 311 299 423 333
rect 121 161 155 214
rect 45 127 155 161
rect 45 106 79 127
rect 213 106 247 289
rect 287 249 353 260
rect 287 215 303 249
rect 337 215 353 249
rect 287 191 353 215
rect 389 219 423 299
rect 489 323 591 337
rect 489 289 545 323
rect 579 305 591 323
rect 489 271 557 289
rect 489 253 591 271
rect 625 331 668 357
rect 625 315 702 331
rect 625 219 659 315
rect 736 265 770 433
rect 804 443 810 477
rect 844 443 892 477
rect 926 443 941 477
rect 804 427 941 443
rect 975 471 1035 487
rect 975 437 991 471
rect 1025 437 1035 471
rect 975 373 1035 437
rect 1069 485 1129 527
rect 1069 451 1085 485
rect 1119 451 1129 485
rect 1163 485 1229 493
rect 1163 451 1179 485
rect 1213 451 1229 485
rect 1069 430 1129 451
rect 1069 411 1135 430
rect 1069 377 1085 411
rect 1119 377 1135 411
rect 1069 375 1135 377
rect 1169 417 1229 451
rect 1169 383 1179 417
rect 1213 383 1229 417
rect 1169 375 1229 383
rect 804 368 1035 373
rect 804 357 991 368
rect 838 334 991 357
rect 1025 341 1035 368
rect 1179 349 1229 375
rect 1263 485 1317 527
rect 1263 451 1273 485
rect 1307 451 1317 485
rect 1263 417 1317 451
rect 1263 383 1273 417
rect 1307 383 1317 417
rect 1263 367 1317 383
rect 1351 485 1417 493
rect 1351 451 1367 485
rect 1401 451 1417 485
rect 1351 417 1417 451
rect 1351 383 1367 417
rect 1401 383 1417 417
rect 1025 334 1145 341
rect 838 323 1145 334
rect 804 307 1145 323
rect 736 249 876 265
rect 736 233 842 249
rect 389 203 507 219
rect 389 169 463 203
rect 497 169 507 203
rect 389 157 507 169
rect 45 56 79 72
rect 113 59 129 93
rect 163 59 179 93
rect 113 17 179 59
rect 213 56 247 72
rect 332 153 507 157
rect 556 197 659 219
rect 556 163 572 197
rect 606 163 659 197
rect 332 123 423 153
rect 556 147 659 163
rect 698 215 842 233
rect 698 199 876 215
rect 332 119 371 123
rect 332 85 337 119
rect 698 113 732 199
rect 910 165 944 307
rect 1111 265 1145 307
rect 1213 333 1229 349
rect 1351 349 1417 383
rect 1351 333 1367 349
rect 1213 315 1367 333
rect 1401 315 1417 349
rect 1179 299 1417 315
rect 1451 485 1502 527
rect 1451 451 1461 485
rect 1495 451 1502 485
rect 1451 417 1502 451
rect 1451 383 1461 417
rect 1495 383 1502 417
rect 1451 349 1502 383
rect 1451 315 1461 349
rect 1495 315 1502 349
rect 1451 299 1502 315
rect 1281 265 1417 299
rect 978 249 1077 265
rect 978 215 1033 249
rect 1067 215 1077 249
rect 1111 249 1247 265
rect 1111 215 1129 249
rect 1163 215 1197 249
rect 1231 215 1247 249
rect 978 199 1077 215
rect 1281 211 1453 265
rect 1281 181 1417 211
rect 891 131 907 165
rect 941 131 957 165
rect 608 106 732 113
rect 332 69 371 85
rect 405 55 421 89
rect 455 55 471 89
rect 608 72 624 106
rect 658 72 732 106
rect 608 56 732 72
rect 774 106 840 122
rect 774 72 790 106
rect 824 72 840 106
rect 405 17 471 55
rect 774 17 840 72
rect 891 93 957 131
rect 891 59 907 93
rect 941 59 957 93
rect 891 51 957 59
rect 1063 161 1129 165
rect 1063 127 1079 161
rect 1113 127 1129 161
rect 1063 93 1129 127
rect 1063 59 1079 93
rect 1113 59 1129 93
rect 1063 17 1129 59
rect 1163 161 1417 181
rect 1163 127 1179 161
rect 1213 147 1367 161
rect 1213 127 1239 147
rect 1163 93 1239 127
rect 1351 127 1367 147
rect 1401 127 1417 161
rect 1163 59 1179 93
rect 1213 59 1239 93
rect 1163 51 1239 59
rect 1275 93 1317 113
rect 1309 59 1317 93
rect 1275 17 1317 59
rect 1351 93 1417 127
rect 1351 59 1367 93
rect 1401 59 1417 93
rect 1351 51 1417 59
rect 1451 161 1493 177
rect 1485 127 1493 161
rect 1451 93 1493 127
rect 1485 59 1493 93
rect 1451 17 1493 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 127 357 161 391
rect 219 289 253 323
rect 656 365 690 391
rect 656 357 668 365
rect 668 357 690 365
rect 545 305 579 323
rect 545 289 557 305
rect 557 289 579 305
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
<< metal1 >>
rect 0 561 1564 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 0 496 1564 527
rect 115 391 173 397
rect 115 357 127 391
rect 161 388 173 391
rect 644 391 702 397
rect 644 388 656 391
rect 161 360 656 388
rect 161 357 173 360
rect 115 351 173 357
rect 644 357 656 360
rect 690 357 702 391
rect 644 351 702 357
rect 207 323 265 329
rect 207 289 219 323
rect 253 320 265 323
rect 533 323 591 329
rect 533 320 545 323
rect 253 292 545 320
rect 253 289 265 292
rect 207 283 265 289
rect 533 289 545 292
rect 579 289 591 323
rect 533 283 591 289
rect 0 17 1564 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
rect 0 -48 1564 -17
<< labels >>
flabel corelocali s 1041 221 1075 255 0 FreeSans 200 0 0 0 RESET_B
port 3 nsew
flabel corelocali s 305 221 339 255 0 FreeSans 200 0 0 0 D
port 1 nsew
flabel corelocali s 29 221 63 255 0 FreeSans 200 0 0 0 GATE_N
port 2 nsew
flabel corelocali s 1317 221 1351 255 0 FreeSans 200 0 0 0 Q
port 8 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
port 5 nsew
rlabel comment s 0 0 0 0 4 dlrtn_4
<< properties >>
string FIXED_BBOX 0 0 1564 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3577968
string GDS_START 3565504
string path 0.000 0.000 39.100 0.000 
<< end >>
