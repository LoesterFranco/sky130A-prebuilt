magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 902 704
<< pwell >>
rect 0 0 864 49
<< scnmos >>
rect 87 112 117 222
rect 190 74 220 222
rect 276 74 306 222
rect 394 94 424 222
rect 512 94 542 222
rect 641 94 671 222
rect 736 94 766 222
<< pmoshvt >>
rect 86 368 116 536
rect 193 368 223 592
rect 283 368 313 592
rect 422 392 452 592
rect 506 392 536 592
rect 608 392 638 592
rect 716 392 746 592
<< ndiff >>
rect 30 184 87 222
rect 30 150 42 184
rect 76 150 87 184
rect 30 112 87 150
rect 117 136 190 222
rect 117 112 144 136
rect 132 102 144 112
rect 178 102 190 136
rect 132 74 190 102
rect 220 210 276 222
rect 220 176 231 210
rect 265 176 276 210
rect 220 120 276 176
rect 220 86 231 120
rect 265 86 276 120
rect 220 74 276 86
rect 306 140 394 222
rect 306 106 340 140
rect 374 106 394 140
rect 306 94 394 106
rect 424 210 512 222
rect 424 176 451 210
rect 485 176 512 210
rect 424 140 512 176
rect 424 106 451 140
rect 485 106 512 140
rect 424 94 512 106
rect 542 140 641 222
rect 542 106 572 140
rect 606 106 641 140
rect 542 94 641 106
rect 671 210 736 222
rect 671 176 691 210
rect 725 176 736 210
rect 671 140 736 176
rect 671 106 691 140
rect 725 106 736 140
rect 671 94 736 106
rect 766 155 837 222
rect 766 121 791 155
rect 825 121 837 155
rect 766 94 837 121
rect 306 74 356 94
<< pdiff >>
rect 134 573 193 592
rect 134 539 146 573
rect 180 539 193 573
rect 134 536 193 539
rect 27 524 86 536
rect 27 490 39 524
rect 73 490 86 524
rect 27 440 86 490
rect 27 406 39 440
rect 73 406 86 440
rect 27 368 86 406
rect 116 368 193 536
rect 223 414 283 592
rect 223 380 236 414
rect 270 380 283 414
rect 223 368 283 380
rect 313 580 422 592
rect 313 546 350 580
rect 384 546 422 580
rect 313 392 422 546
rect 452 392 506 592
rect 536 392 608 592
rect 638 392 716 592
rect 746 580 835 592
rect 746 546 789 580
rect 823 546 835 580
rect 746 509 835 546
rect 746 475 789 509
rect 823 475 835 509
rect 746 438 835 475
rect 746 404 789 438
rect 823 404 835 438
rect 746 392 835 404
rect 313 368 366 392
<< ndiffc >>
rect 42 150 76 184
rect 144 102 178 136
rect 231 176 265 210
rect 231 86 265 120
rect 340 106 374 140
rect 451 176 485 210
rect 451 106 485 140
rect 572 106 606 140
rect 691 176 725 210
rect 691 106 725 140
rect 791 121 825 155
<< pdiffc >>
rect 146 539 180 573
rect 39 490 73 524
rect 39 406 73 440
rect 236 380 270 414
rect 350 546 384 580
rect 789 546 823 580
rect 789 475 823 509
rect 789 404 823 438
<< poly >>
rect 193 592 223 618
rect 283 592 313 618
rect 422 592 452 618
rect 506 592 536 618
rect 608 592 638 618
rect 716 592 746 618
rect 86 536 116 562
rect 422 377 452 392
rect 506 377 536 392
rect 608 377 638 392
rect 716 377 746 392
rect 86 353 116 368
rect 193 353 223 368
rect 283 353 313 368
rect 83 336 117 353
rect 44 320 117 336
rect 44 286 60 320
rect 94 286 117 320
rect 44 270 117 286
rect 87 222 117 270
rect 190 290 226 353
rect 280 326 316 353
rect 419 336 455 377
rect 503 360 539 377
rect 605 360 641 377
rect 276 310 346 326
rect 276 290 296 310
rect 190 276 296 290
rect 330 276 346 310
rect 190 260 346 276
rect 389 320 455 336
rect 389 286 405 320
rect 439 286 455 320
rect 497 344 563 360
rect 497 310 513 344
rect 547 310 563 344
rect 497 294 563 310
rect 605 344 671 360
rect 605 310 621 344
rect 655 310 671 344
rect 605 294 671 310
rect 389 270 455 286
rect 190 222 220 260
rect 276 222 306 260
rect 394 222 424 270
rect 512 222 542 294
rect 641 222 671 294
rect 713 354 749 377
rect 713 338 779 354
rect 713 304 729 338
rect 763 304 779 338
rect 713 288 779 304
rect 736 222 766 288
rect 87 86 117 112
rect 190 48 220 74
rect 276 48 306 74
rect 394 68 424 94
rect 512 68 542 94
rect 641 68 671 94
rect 736 68 766 94
<< polycont >>
rect 60 286 94 320
rect 296 276 330 310
rect 405 286 439 320
rect 513 310 547 344
rect 621 310 655 344
rect 729 304 763 338
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 130 573 196 649
rect 23 524 89 540
rect 130 539 146 573
rect 180 539 196 573
rect 310 580 425 649
rect 310 546 350 580
rect 384 546 425 580
rect 773 580 847 596
rect 130 532 196 539
rect 459 538 739 572
rect 23 490 39 524
rect 73 498 89 524
rect 459 498 493 538
rect 73 490 493 498
rect 23 464 493 490
rect 23 440 178 464
rect 23 406 39 440
rect 73 406 178 440
rect 23 390 178 406
rect 25 320 110 356
rect 25 286 60 320
rect 94 286 110 320
rect 25 270 110 286
rect 144 236 178 390
rect 26 202 178 236
rect 212 414 286 430
rect 212 380 236 414
rect 270 380 286 414
rect 212 364 286 380
rect 212 226 246 364
rect 280 310 349 326
rect 280 276 296 310
rect 330 276 349 310
rect 280 260 349 276
rect 389 320 455 430
rect 389 286 405 320
rect 439 286 455 320
rect 497 344 563 430
rect 497 310 513 344
rect 547 310 563 344
rect 497 294 563 310
rect 601 344 671 504
rect 601 310 621 344
rect 655 310 671 344
rect 601 294 671 310
rect 705 354 739 538
rect 773 546 789 580
rect 823 546 847 580
rect 773 509 847 546
rect 773 475 789 509
rect 823 475 847 509
rect 773 438 847 475
rect 773 404 789 438
rect 823 404 847 438
rect 773 388 847 404
rect 705 338 779 354
rect 705 304 729 338
rect 763 304 779 338
rect 705 288 779 304
rect 389 270 455 286
rect 315 226 349 260
rect 813 254 847 388
rect 675 226 847 254
rect 212 210 281 226
rect 26 184 92 202
rect 26 150 42 184
rect 76 150 92 184
rect 212 176 231 210
rect 265 176 281 210
rect 315 220 847 226
rect 315 210 741 220
rect 315 192 451 210
rect 26 108 92 150
rect 128 136 178 168
rect 128 102 144 136
rect 128 17 178 102
rect 212 120 281 176
rect 435 176 451 192
rect 485 192 691 210
rect 485 176 501 192
rect 212 86 231 120
rect 265 86 281 120
rect 212 70 281 86
rect 315 140 399 156
rect 315 106 340 140
rect 374 106 399 140
rect 315 17 399 106
rect 435 140 501 176
rect 675 176 691 192
rect 725 176 741 210
rect 435 106 451 140
rect 485 106 501 140
rect 435 90 501 106
rect 537 140 641 156
rect 537 106 572 140
rect 606 106 641 140
rect 537 17 641 106
rect 675 140 741 176
rect 675 106 691 140
rect 725 106 741 140
rect 675 90 741 106
rect 775 155 841 186
rect 775 121 791 155
rect 825 121 841 155
rect 775 17 841 121
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel comment s 0 0 0 0 4 or4b_2
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 415 390 449 424 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 511 390 545 424 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 607 390 641 424 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 607 464 641 498 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 D_N
port 4 nsew
flabel corelocali s 223 390 257 424 0 FreeSans 340 0 0 0 X
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 864 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1081188
string GDS_START 1073752
<< end >>
