magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1196 561
rect 103 427 169 527
rect 17 197 66 325
rect 103 17 169 93
rect 395 367 458 527
rect 296 191 362 265
rect 768 427 828 527
rect 952 299 1009 527
rect 1043 328 1093 491
rect 1127 351 1179 527
rect 1043 299 1100 328
rect 1066 265 1100 299
rect 1066 199 1179 265
rect 1066 165 1100 199
rect 379 17 445 89
rect 752 17 818 165
rect 952 17 1009 165
rect 1043 137 1100 165
rect 1043 83 1093 137
rect 1127 17 1179 110
rect 0 -17 1196 17
<< obsli1 >>
rect 35 393 69 493
rect 35 359 156 393
rect 122 323 156 359
rect 122 280 156 289
rect 203 391 248 493
rect 203 357 214 391
rect 203 337 248 357
rect 122 214 168 280
rect 122 161 156 214
rect 35 127 156 161
rect 35 69 69 127
rect 203 69 237 337
rect 295 333 361 483
rect 584 451 734 485
rect 498 391 555 401
rect 532 357 555 391
rect 295 299 432 333
rect 398 219 432 299
rect 498 271 555 357
rect 589 323 657 399
rect 589 289 590 323
rect 624 289 657 323
rect 589 283 657 289
rect 398 157 472 219
rect 589 207 623 283
rect 700 265 734 451
rect 872 373 916 487
rect 772 307 916 373
rect 882 265 916 307
rect 700 233 844 265
rect 311 153 472 157
rect 311 123 432 153
rect 547 141 623 207
rect 670 199 844 233
rect 882 199 1032 265
rect 311 69 345 123
rect 670 107 704 199
rect 882 165 916 199
rect 572 73 704 107
rect 872 83 916 165
<< obsli1c >>
rect 122 289 156 323
rect 214 357 248 391
rect 498 357 532 391
rect 590 289 624 323
<< metal1 >>
rect 0 496 1196 592
rect 0 -48 1196 48
<< obsm1 >>
rect 202 391 260 397
rect 202 357 214 391
rect 248 388 260 391
rect 486 391 544 397
rect 486 388 498 391
rect 248 360 498 388
rect 248 357 260 360
rect 202 351 260 357
rect 486 357 498 360
rect 532 357 544 391
rect 486 351 544 357
rect 110 323 168 329
rect 110 289 122 323
rect 156 320 168 323
rect 578 323 636 329
rect 578 320 590 323
rect 156 292 590 320
rect 156 289 168 292
rect 110 283 168 289
rect 578 289 590 292
rect 624 289 636 323
rect 578 283 636 289
<< labels >>
rlabel locali s 296 191 362 265 6 D
port 1 nsew signal input
rlabel locali s 1066 265 1100 299 6 Q
port 2 nsew signal output
rlabel locali s 1066 199 1179 265 6 Q
port 2 nsew signal output
rlabel locali s 1066 165 1100 199 6 Q
port 2 nsew signal output
rlabel locali s 1043 328 1093 491 6 Q
port 2 nsew signal output
rlabel locali s 1043 299 1100 328 6 Q
port 2 nsew signal output
rlabel locali s 1043 137 1100 165 6 Q
port 2 nsew signal output
rlabel locali s 1043 83 1093 137 6 Q
port 2 nsew signal output
rlabel locali s 17 197 66 325 6 GATE_N
port 3 nsew clock input
rlabel locali s 1127 17 1179 110 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 952 17 1009 165 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 752 17 818 165 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 379 17 445 89 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 103 17 169 93 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 1196 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1196 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 1127 351 1179 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 952 299 1009 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 768 427 828 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 395 367 458 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 103 427 169 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 1196 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 1196 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2784190
string GDS_START 2774118
<< end >>
