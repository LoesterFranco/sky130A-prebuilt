magic
tech sky130A
magscale 1 2
timestamp 1601050058
<< locali >>
rect 361 405 694 421
rect 809 405 1536 421
rect 361 371 1536 405
rect 193 303 726 337
rect 193 266 282 303
rect 80 215 282 266
rect 341 215 636 269
rect 670 199 726 303
rect 852 303 1400 337
rect 852 282 995 303
rect 760 199 995 282
rect 1074 215 1288 269
rect 1366 199 1400 303
rect 1434 268 1536 371
rect 1434 165 1470 268
rect 1313 131 1470 165
rect 1313 90 1347 131
rect 1056 54 1347 90
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 18 333 77 527
rect 191 455 257 527
rect 291 455 687 493
rect 111 421 155 438
rect 291 421 327 455
rect 723 439 777 527
rect 887 455 953 527
rect 1056 455 1122 527
rect 1224 455 1291 527
rect 1471 455 1537 527
rect 111 387 327 421
rect 111 372 155 387
rect 31 173 359 181
rect 31 159 626 173
rect 31 139 767 159
rect 31 125 248 139
rect 355 125 767 139
rect 801 127 1234 163
rect 31 107 71 125
rect 105 17 171 89
rect 205 85 248 125
rect 293 17 327 105
rect 721 91 767 125
rect 449 17 515 89
rect 621 17 687 89
rect 721 51 984 91
rect 1502 96 1536 119
rect 1396 62 1536 96
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
<< metal1 >>
rect 0 561 1564 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 0 496 1564 527
rect 0 17 1564 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
rect 0 -48 1564 -17
<< obsm1 >>
rect 202 116 260 125
rect 1490 116 1548 125
rect 202 88 1548 116
rect 202 79 260 88
rect 1490 79 1548 88
<< labels >>
rlabel locali s 670 199 726 303 6 A1
port 1 nsew signal input
rlabel locali s 193 303 726 337 6 A1
port 1 nsew signal input
rlabel locali s 193 266 282 303 6 A1
port 1 nsew signal input
rlabel locali s 80 215 282 266 6 A1
port 1 nsew signal input
rlabel locali s 341 215 636 269 6 A2
port 2 nsew signal input
rlabel locali s 1366 199 1400 303 6 B1
port 3 nsew signal input
rlabel locali s 852 303 1400 337 6 B1
port 3 nsew signal input
rlabel locali s 852 282 995 303 6 B1
port 3 nsew signal input
rlabel locali s 760 199 995 282 6 B1
port 3 nsew signal input
rlabel locali s 1074 215 1288 269 6 C1
port 4 nsew signal input
rlabel locali s 1434 268 1536 371 6 Y
port 5 nsew signal output
rlabel locali s 1434 165 1470 268 6 Y
port 5 nsew signal output
rlabel locali s 1313 131 1470 165 6 Y
port 5 nsew signal output
rlabel locali s 1313 90 1347 131 6 Y
port 5 nsew signal output
rlabel locali s 1056 54 1347 90 6 Y
port 5 nsew signal output
rlabel locali s 809 405 1536 421 6 Y
port 5 nsew signal output
rlabel locali s 361 405 694 421 6 Y
port 5 nsew signal output
rlabel locali s 361 371 1536 405 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -48 1564 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1564 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1564 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1308074
string GDS_START 1298054
<< end >>
