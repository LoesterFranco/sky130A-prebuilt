magic
tech sky130A
magscale 1 2
timestamp 1604502710
<< nwell >>
rect -38 332 3398 704
<< pwell >>
rect 0 0 3360 49
<< scpmos >>
rect 83 392 119 592
rect 173 392 209 592
rect 263 392 299 592
rect 363 392 399 592
rect 568 392 604 592
rect 663 392 699 592
rect 758 392 794 592
rect 848 392 884 592
rect 1050 368 1086 592
rect 1252 377 1288 577
rect 1342 377 1378 577
rect 1432 377 1468 577
rect 1522 377 1558 577
rect 1741 392 1777 592
rect 1831 392 1867 592
rect 1957 392 1993 592
rect 2047 392 2083 592
rect 2289 392 2325 592
rect 2389 392 2425 592
rect 2489 392 2525 592
rect 2589 392 2625 592
rect 2842 368 2878 592
rect 2945 368 2981 592
rect 3035 368 3071 592
rect 3135 368 3171 592
rect 3225 368 3261 592
<< nmoslvt >>
rect 84 126 114 254
rect 170 126 200 254
rect 269 126 299 254
rect 355 126 385 254
rect 585 119 615 247
rect 680 119 710 247
rect 766 119 796 247
rect 852 119 882 247
rect 1050 74 1080 222
rect 1248 121 1278 249
rect 1334 121 1364 249
rect 1420 121 1450 249
rect 1506 121 1536 249
rect 1776 74 1806 202
rect 1862 74 1892 202
rect 1948 74 1978 202
rect 2034 74 2064 202
rect 2256 74 2286 202
rect 2374 74 2404 202
rect 2544 74 2574 202
rect 2630 74 2660 202
rect 2842 74 2872 222
rect 2988 74 3018 222
rect 3074 74 3104 222
rect 3160 74 3190 222
rect 3246 74 3276 222
<< ndiff >>
rect 27 240 84 254
rect 27 206 39 240
rect 73 206 84 240
rect 27 172 84 206
rect 27 138 39 172
rect 73 138 84 172
rect 27 126 84 138
rect 114 172 170 254
rect 114 138 125 172
rect 159 138 170 172
rect 114 126 170 138
rect 200 246 269 254
rect 200 212 217 246
rect 251 212 269 246
rect 200 178 269 212
rect 200 144 217 178
rect 251 144 269 178
rect 200 126 269 144
rect 299 242 355 254
rect 299 208 310 242
rect 344 208 355 242
rect 299 126 355 208
rect 385 126 458 254
rect 400 90 458 126
rect 400 56 412 90
rect 446 56 458 90
rect 512 119 585 247
rect 615 185 680 247
rect 615 151 626 185
rect 660 151 680 185
rect 615 119 680 151
rect 710 191 766 247
rect 710 157 721 191
rect 755 157 766 191
rect 710 119 766 157
rect 796 237 852 247
rect 796 203 807 237
rect 841 203 852 237
rect 796 169 852 203
rect 796 135 807 169
rect 841 135 852 169
rect 796 119 852 135
rect 882 236 939 247
rect 882 202 893 236
rect 927 202 939 236
rect 1191 239 1248 249
rect 882 168 939 202
rect 882 134 893 168
rect 927 134 939 168
rect 882 119 939 134
rect 993 210 1050 222
rect 993 176 1005 210
rect 1039 176 1050 210
rect 993 120 1050 176
rect 512 108 570 119
rect 512 74 524 108
rect 558 74 570 108
rect 512 62 570 74
rect 400 44 458 56
rect 993 86 1005 120
rect 1039 86 1050 120
rect 993 74 1050 86
rect 1080 210 1137 222
rect 1080 176 1091 210
rect 1125 176 1137 210
rect 1080 120 1137 176
rect 1191 205 1203 239
rect 1237 205 1248 239
rect 1191 167 1248 205
rect 1191 133 1203 167
rect 1237 133 1248 167
rect 1191 121 1248 133
rect 1278 169 1334 249
rect 1278 135 1289 169
rect 1323 135 1334 169
rect 1278 121 1334 135
rect 1364 237 1420 249
rect 1364 203 1375 237
rect 1409 203 1420 237
rect 1364 169 1420 203
rect 1364 135 1375 169
rect 1409 135 1420 169
rect 1364 121 1420 135
rect 1450 237 1506 249
rect 1450 203 1461 237
rect 1495 203 1506 237
rect 1450 121 1506 203
rect 1536 169 1609 249
rect 1536 135 1563 169
rect 1597 135 1609 169
rect 1536 121 1609 135
rect 1080 86 1091 120
rect 1125 86 1137 120
rect 1080 74 1137 86
rect 1703 82 1776 202
rect 1703 48 1715 82
rect 1749 74 1776 82
rect 1806 127 1862 202
rect 1806 93 1817 127
rect 1851 93 1862 127
rect 1806 74 1862 93
rect 1892 127 1948 202
rect 1892 93 1903 127
rect 1937 93 1948 127
rect 1892 74 1948 93
rect 1978 190 2034 202
rect 1978 156 1989 190
rect 2023 156 2034 190
rect 1978 120 2034 156
rect 1978 86 1989 120
rect 2023 86 2034 120
rect 1978 74 2034 86
rect 2064 190 2121 202
rect 2064 156 2075 190
rect 2109 156 2121 190
rect 2064 120 2121 156
rect 2064 86 2075 120
rect 2109 86 2121 120
rect 2064 74 2121 86
rect 2199 179 2256 202
rect 2199 145 2211 179
rect 2245 145 2256 179
rect 2199 74 2256 145
rect 2286 85 2374 202
rect 2286 74 2313 85
rect 1749 48 1761 74
rect 2301 51 2313 74
rect 2347 74 2374 85
rect 2404 123 2544 202
rect 2404 89 2415 123
rect 2449 89 2485 123
rect 2519 89 2544 123
rect 2404 74 2544 89
rect 2574 172 2630 202
rect 2574 138 2585 172
rect 2619 138 2630 172
rect 2574 74 2630 138
rect 2660 184 2731 202
rect 2660 150 2685 184
rect 2719 150 2731 184
rect 2660 116 2731 150
rect 2660 82 2671 116
rect 2705 82 2731 116
rect 2660 74 2731 82
rect 2785 172 2842 222
rect 2785 138 2797 172
rect 2831 138 2842 172
rect 2785 74 2842 138
rect 2872 210 2988 222
rect 2872 176 2943 210
rect 2977 176 2988 210
rect 2872 120 2988 176
rect 2872 86 2943 120
rect 2977 86 2988 120
rect 2872 74 2988 86
rect 3018 210 3074 222
rect 3018 176 3029 210
rect 3063 176 3074 210
rect 3018 120 3074 176
rect 3018 86 3029 120
rect 3063 86 3074 120
rect 3018 74 3074 86
rect 3104 142 3160 222
rect 3104 108 3115 142
rect 3149 108 3160 142
rect 3104 74 3160 108
rect 3190 210 3246 222
rect 3190 176 3201 210
rect 3235 176 3246 210
rect 3190 120 3246 176
rect 3190 86 3201 120
rect 3235 86 3246 120
rect 3190 74 3246 86
rect 3276 142 3333 222
rect 3276 108 3287 142
rect 3321 108 3333 142
rect 3276 74 3333 108
rect 2347 51 2359 74
rect 1703 36 1761 48
rect 2301 39 2359 51
<< pdiff >>
rect 1668 627 1726 639
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 510 83 546
rect 27 476 39 510
rect 73 476 83 510
rect 27 440 83 476
rect 27 406 39 440
rect 73 406 83 440
rect 27 392 83 406
rect 119 580 173 592
rect 119 546 129 580
rect 163 546 173 580
rect 119 510 173 546
rect 119 476 129 510
rect 163 476 173 510
rect 119 440 173 476
rect 119 406 129 440
rect 163 406 173 440
rect 119 392 173 406
rect 209 580 263 592
rect 209 546 219 580
rect 253 546 263 580
rect 209 512 263 546
rect 209 478 219 512
rect 253 478 263 512
rect 209 392 263 478
rect 299 580 363 592
rect 299 546 319 580
rect 353 546 363 580
rect 299 512 363 546
rect 299 478 319 512
rect 353 478 363 512
rect 299 392 363 478
rect 399 580 455 592
rect 399 546 409 580
rect 443 546 455 580
rect 399 392 455 546
rect 509 580 568 592
rect 509 546 522 580
rect 556 546 568 580
rect 509 392 568 546
rect 604 531 663 592
rect 604 497 614 531
rect 648 497 663 531
rect 604 438 663 497
rect 604 404 614 438
rect 648 404 663 438
rect 604 392 663 404
rect 699 580 758 592
rect 699 546 714 580
rect 748 546 758 580
rect 699 509 758 546
rect 699 475 714 509
rect 748 475 758 509
rect 699 438 758 475
rect 699 404 714 438
rect 748 404 758 438
rect 699 392 758 404
rect 794 531 848 592
rect 794 497 804 531
rect 838 497 848 531
rect 794 438 848 497
rect 794 404 804 438
rect 838 404 848 438
rect 794 392 848 404
rect 884 580 940 592
rect 884 546 894 580
rect 928 546 940 580
rect 884 509 940 546
rect 884 475 894 509
rect 928 475 940 509
rect 884 438 940 475
rect 884 404 894 438
rect 928 404 940 438
rect 884 392 940 404
rect 994 580 1050 592
rect 994 546 1006 580
rect 1040 546 1050 580
rect 994 497 1050 546
rect 994 463 1006 497
rect 1040 463 1050 497
rect 994 414 1050 463
rect 994 380 1006 414
rect 1040 380 1050 414
rect 994 368 1050 380
rect 1086 580 1142 592
rect 1086 546 1096 580
rect 1130 546 1142 580
rect 1668 593 1680 627
rect 1714 593 1726 627
rect 1882 627 1942 639
rect 1668 592 1726 593
rect 1882 593 1895 627
rect 1929 593 1942 627
rect 1882 592 1942 593
rect 1086 497 1142 546
rect 1086 463 1096 497
rect 1130 463 1142 497
rect 1086 414 1142 463
rect 1086 380 1096 414
rect 1130 380 1142 414
rect 1086 368 1142 380
rect 1196 565 1252 577
rect 1196 531 1208 565
rect 1242 531 1252 565
rect 1196 494 1252 531
rect 1196 460 1208 494
rect 1242 460 1252 494
rect 1196 423 1252 460
rect 1196 389 1208 423
rect 1242 389 1252 423
rect 1196 377 1252 389
rect 1288 565 1342 577
rect 1288 531 1298 565
rect 1332 531 1342 565
rect 1288 480 1342 531
rect 1288 446 1298 480
rect 1332 446 1342 480
rect 1288 377 1342 446
rect 1378 531 1432 577
rect 1378 497 1388 531
rect 1422 497 1432 531
rect 1378 423 1432 497
rect 1378 389 1388 423
rect 1422 389 1432 423
rect 1378 377 1432 389
rect 1468 527 1522 577
rect 1468 493 1478 527
rect 1512 493 1522 527
rect 1468 377 1522 493
rect 1558 423 1614 577
rect 1558 389 1568 423
rect 1602 389 1614 423
rect 1668 392 1741 592
rect 1777 491 1831 592
rect 1777 457 1787 491
rect 1821 457 1831 491
rect 1777 392 1831 457
rect 1867 392 1957 592
rect 1993 580 2047 592
rect 1993 546 2003 580
rect 2037 546 2047 580
rect 1993 507 2047 546
rect 1993 473 2003 507
rect 2037 473 2047 507
rect 1993 392 2047 473
rect 2083 580 2139 592
rect 2083 546 2093 580
rect 2127 546 2139 580
rect 2083 507 2139 546
rect 2083 473 2093 507
rect 2127 473 2139 507
rect 2083 392 2139 473
rect 2233 539 2289 592
rect 2233 505 2245 539
rect 2279 505 2289 539
rect 2233 438 2289 505
rect 2233 404 2245 438
rect 2279 404 2289 438
rect 2233 392 2289 404
rect 2325 463 2389 592
rect 2325 429 2345 463
rect 2379 429 2389 463
rect 2325 392 2389 429
rect 2425 539 2489 592
rect 2425 505 2445 539
rect 2479 505 2489 539
rect 2425 440 2489 505
rect 2425 406 2445 440
rect 2479 406 2489 440
rect 2425 392 2489 406
rect 2525 582 2589 592
rect 2525 548 2545 582
rect 2579 548 2589 582
rect 2525 514 2589 548
rect 2525 480 2545 514
rect 2579 480 2589 514
rect 2525 392 2589 480
rect 2625 582 2691 592
rect 2625 548 2645 582
rect 2679 548 2691 582
rect 2625 514 2691 548
rect 2625 480 2645 514
rect 2679 480 2691 514
rect 2625 446 2691 480
rect 2625 412 2645 446
rect 2679 412 2691 446
rect 2625 392 2691 412
rect 2779 580 2842 592
rect 2779 546 2791 580
rect 2825 546 2842 580
rect 2779 497 2842 546
rect 2779 463 2791 497
rect 2825 463 2842 497
rect 2779 414 2842 463
rect 1558 377 1614 389
rect 2779 380 2791 414
rect 2825 380 2842 414
rect 2779 368 2842 380
rect 2878 580 2945 592
rect 2878 546 2891 580
rect 2925 546 2945 580
rect 2878 497 2945 546
rect 2878 463 2891 497
rect 2925 463 2945 497
rect 2878 414 2945 463
rect 2878 380 2891 414
rect 2925 380 2945 414
rect 2878 368 2945 380
rect 2981 580 3035 592
rect 2981 546 2991 580
rect 3025 546 3035 580
rect 2981 497 3035 546
rect 2981 463 2991 497
rect 3025 463 3035 497
rect 2981 414 3035 463
rect 2981 380 2991 414
rect 3025 380 3035 414
rect 2981 368 3035 380
rect 3071 580 3135 592
rect 3071 546 3081 580
rect 3115 546 3135 580
rect 3071 478 3135 546
rect 3071 444 3081 478
rect 3115 444 3135 478
rect 3071 368 3135 444
rect 3171 580 3225 592
rect 3171 546 3181 580
rect 3215 546 3225 580
rect 3171 497 3225 546
rect 3171 463 3181 497
rect 3215 463 3225 497
rect 3171 414 3225 463
rect 3171 380 3181 414
rect 3215 380 3225 414
rect 3171 368 3225 380
rect 3261 580 3327 592
rect 3261 546 3281 580
rect 3315 546 3327 580
rect 3261 478 3327 546
rect 3261 444 3281 478
rect 3315 444 3327 478
rect 3261 368 3327 444
<< ndiffc >>
rect 39 206 73 240
rect 39 138 73 172
rect 125 138 159 172
rect 217 212 251 246
rect 217 144 251 178
rect 310 208 344 242
rect 412 56 446 90
rect 626 151 660 185
rect 721 157 755 191
rect 807 203 841 237
rect 807 135 841 169
rect 893 202 927 236
rect 893 134 927 168
rect 1005 176 1039 210
rect 524 74 558 108
rect 1005 86 1039 120
rect 1091 176 1125 210
rect 1203 205 1237 239
rect 1203 133 1237 167
rect 1289 135 1323 169
rect 1375 203 1409 237
rect 1375 135 1409 169
rect 1461 203 1495 237
rect 1563 135 1597 169
rect 1091 86 1125 120
rect 1715 48 1749 82
rect 1817 93 1851 127
rect 1903 93 1937 127
rect 1989 156 2023 190
rect 1989 86 2023 120
rect 2075 156 2109 190
rect 2075 86 2109 120
rect 2211 145 2245 179
rect 2313 51 2347 85
rect 2415 89 2449 123
rect 2485 89 2519 123
rect 2585 138 2619 172
rect 2685 150 2719 184
rect 2671 82 2705 116
rect 2797 138 2831 172
rect 2943 176 2977 210
rect 2943 86 2977 120
rect 3029 176 3063 210
rect 3029 86 3063 120
rect 3115 108 3149 142
rect 3201 176 3235 210
rect 3201 86 3235 120
rect 3287 108 3321 142
<< pdiffc >>
rect 39 546 73 580
rect 39 476 73 510
rect 39 406 73 440
rect 129 546 163 580
rect 129 476 163 510
rect 129 406 163 440
rect 219 546 253 580
rect 219 478 253 512
rect 319 546 353 580
rect 319 478 353 512
rect 409 546 443 580
rect 522 546 556 580
rect 614 497 648 531
rect 614 404 648 438
rect 714 546 748 580
rect 714 475 748 509
rect 714 404 748 438
rect 804 497 838 531
rect 804 404 838 438
rect 894 546 928 580
rect 894 475 928 509
rect 894 404 928 438
rect 1006 546 1040 580
rect 1006 463 1040 497
rect 1006 380 1040 414
rect 1096 546 1130 580
rect 1680 593 1714 627
rect 1895 593 1929 627
rect 1096 463 1130 497
rect 1096 380 1130 414
rect 1208 531 1242 565
rect 1208 460 1242 494
rect 1208 389 1242 423
rect 1298 531 1332 565
rect 1298 446 1332 480
rect 1388 497 1422 531
rect 1388 389 1422 423
rect 1478 493 1512 527
rect 1568 389 1602 423
rect 1787 457 1821 491
rect 2003 546 2037 580
rect 2003 473 2037 507
rect 2093 546 2127 580
rect 2093 473 2127 507
rect 2245 505 2279 539
rect 2245 404 2279 438
rect 2345 429 2379 463
rect 2445 505 2479 539
rect 2445 406 2479 440
rect 2545 548 2579 582
rect 2545 480 2579 514
rect 2645 548 2679 582
rect 2645 480 2679 514
rect 2645 412 2679 446
rect 2791 546 2825 580
rect 2791 463 2825 497
rect 2791 380 2825 414
rect 2891 546 2925 580
rect 2891 463 2925 497
rect 2891 380 2925 414
rect 2991 546 3025 580
rect 2991 463 3025 497
rect 2991 380 3025 414
rect 3081 546 3115 580
rect 3081 444 3115 478
rect 3181 546 3215 580
rect 3181 463 3215 497
rect 3181 380 3215 414
rect 3281 546 3315 580
rect 3281 444 3315 478
<< poly >>
rect 83 592 119 618
rect 173 592 209 618
rect 263 592 299 618
rect 363 592 399 618
rect 568 592 604 618
rect 663 592 699 618
rect 758 592 794 618
rect 848 592 884 618
rect 1050 592 1086 618
rect 83 356 119 392
rect 173 356 209 392
rect 44 340 209 356
rect 44 306 60 340
rect 94 306 128 340
rect 162 306 209 340
rect 44 290 209 306
rect 263 360 299 392
rect 363 360 399 392
rect 263 344 471 360
rect 263 310 285 344
rect 319 310 353 344
rect 387 310 421 344
rect 455 310 471 344
rect 263 294 471 310
rect 84 254 114 290
rect 170 254 200 290
rect 269 254 299 294
rect 355 254 385 294
rect 568 292 604 392
rect 663 292 699 392
rect 758 336 794 392
rect 848 336 884 392
rect 1252 577 1288 603
rect 1342 577 1378 603
rect 1432 577 1468 603
rect 1522 577 1558 603
rect 1741 592 1777 618
rect 1831 592 1867 618
rect 1957 592 1993 618
rect 2047 592 2083 618
rect 2289 592 2325 618
rect 2389 592 2425 618
rect 2489 592 2525 618
rect 2589 592 2625 618
rect 2842 592 2878 618
rect 2945 592 2981 618
rect 3035 592 3071 618
rect 3135 592 3171 618
rect 3225 592 3261 618
rect 758 320 1008 336
rect 758 306 958 320
rect 568 262 615 292
rect 663 262 710 292
rect 585 247 615 262
rect 680 247 710 262
rect 766 286 958 306
rect 992 286 1008 320
rect 766 283 1008 286
rect 766 247 796 283
rect 852 247 882 283
rect 942 270 1008 283
rect 84 100 114 126
rect 170 100 200 126
rect 269 100 299 126
rect 355 100 385 126
rect 1050 237 1086 368
rect 1252 339 1288 377
rect 1342 339 1378 377
rect 1207 323 1378 339
rect 1207 289 1223 323
rect 1257 289 1291 323
rect 1325 289 1378 323
rect 1432 345 1468 377
rect 1522 345 1558 377
rect 1432 329 1661 345
rect 1432 309 1475 329
rect 1207 273 1378 289
rect 1420 295 1475 309
rect 1509 295 1543 329
rect 1577 295 1611 329
rect 1645 295 1661 329
rect 1420 279 1661 295
rect 1248 249 1278 273
rect 1334 249 1364 273
rect 1420 249 1450 279
rect 1506 249 1536 279
rect 1050 222 1080 237
rect 585 51 615 119
rect 680 51 710 119
rect 766 93 796 119
rect 852 93 882 119
rect 1248 95 1278 121
rect 1334 95 1364 121
rect 1420 95 1450 121
rect 1506 95 1536 121
rect 1050 51 1080 74
rect 1631 51 1661 279
rect 1741 318 1777 392
rect 1831 318 1867 392
rect 1957 355 1993 392
rect 2047 355 2083 392
rect 1948 339 2083 355
rect 1741 302 1892 318
rect 1741 268 1769 302
rect 1803 268 1837 302
rect 1871 268 1892 302
rect 1741 252 1892 268
rect 1776 202 1806 252
rect 1862 202 1892 252
rect 1948 305 1964 339
rect 1998 305 2032 339
rect 2066 319 2083 339
rect 2066 305 2082 319
rect 1948 289 2082 305
rect 1948 202 1978 289
rect 2052 247 2082 289
rect 2289 305 2325 392
rect 2389 305 2425 392
rect 2489 377 2525 392
rect 2589 377 2625 392
rect 2489 347 2666 377
rect 2544 344 2666 347
rect 2544 310 2616 344
rect 2650 310 2666 344
rect 2289 289 2496 305
rect 2289 269 2446 289
rect 2034 217 2082 247
rect 2256 255 2446 269
rect 2480 255 2496 289
rect 2256 239 2496 255
rect 2544 294 2666 310
rect 2708 304 2774 310
rect 2842 304 2878 368
rect 2708 294 2878 304
rect 2945 326 2981 368
rect 3035 326 3071 368
rect 3135 326 3171 368
rect 3225 326 3261 368
rect 2945 310 3276 326
rect 2945 296 3004 310
rect 2034 202 2064 217
rect 2256 202 2286 239
rect 2374 202 2404 239
rect 2544 202 2574 294
rect 2630 202 2660 294
rect 2708 260 2724 294
rect 2758 260 2878 294
rect 2708 244 2878 260
rect 2988 276 3004 296
rect 3038 276 3072 310
rect 3106 276 3140 310
rect 3174 276 3208 310
rect 3242 276 3276 310
rect 2988 260 3276 276
rect 2842 222 2872 244
rect 2988 222 3018 260
rect 3074 222 3104 260
rect 3160 222 3190 260
rect 3246 222 3276 260
rect 585 21 1661 51
rect 1776 48 1806 74
rect 1862 48 1892 74
rect 1948 48 1978 74
rect 2034 48 2064 74
rect 2256 48 2286 74
rect 2374 48 2404 74
rect 2544 48 2574 74
rect 2630 48 2660 74
rect 2842 48 2872 74
rect 2988 48 3018 74
rect 3074 48 3104 74
rect 3160 48 3190 74
rect 3246 48 3276 74
<< polycont >>
rect 60 306 94 340
rect 128 306 162 340
rect 285 310 319 344
rect 353 310 387 344
rect 421 310 455 344
rect 958 286 992 320
rect 1223 289 1257 323
rect 1291 289 1325 323
rect 1475 295 1509 329
rect 1543 295 1577 329
rect 1611 295 1645 329
rect 1769 268 1803 302
rect 1837 268 1871 302
rect 1964 305 1998 339
rect 2032 305 2066 339
rect 2616 310 2650 344
rect 2446 255 2480 289
rect 2724 260 2758 294
rect 3004 276 3038 310
rect 3072 276 3106 310
rect 3140 276 3174 310
rect 3208 276 3242 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3360 683
rect 23 580 73 649
rect 23 546 39 580
rect 23 510 73 546
rect 23 476 39 510
rect 23 440 73 476
rect 23 406 39 440
rect 23 390 73 406
rect 113 580 179 596
rect 113 546 129 580
rect 163 546 179 580
rect 113 510 179 546
rect 113 476 129 510
rect 163 476 179 510
rect 113 440 179 476
rect 219 580 269 649
rect 253 546 269 580
rect 219 512 269 546
rect 253 478 269 512
rect 219 462 269 478
rect 303 580 369 596
rect 303 546 319 580
rect 353 546 369 580
rect 303 512 369 546
rect 409 580 459 649
rect 443 546 459 580
rect 409 530 459 546
rect 505 581 944 615
rect 505 580 572 581
rect 505 546 522 580
rect 556 546 572 580
rect 698 580 764 581
rect 505 530 572 546
rect 609 531 660 547
rect 303 478 319 512
rect 353 496 369 512
rect 609 497 614 531
rect 648 497 660 531
rect 609 496 660 497
rect 353 478 660 496
rect 303 462 660 478
rect 113 406 129 440
rect 163 428 179 440
rect 598 438 660 462
rect 163 406 539 428
rect 113 394 539 406
rect 113 390 179 394
rect 25 340 178 356
rect 25 306 60 340
rect 94 306 128 340
rect 162 306 178 340
rect 25 290 178 306
rect 217 344 471 360
rect 217 310 285 344
rect 319 310 353 344
rect 387 310 421 344
rect 455 310 471 344
rect 505 354 539 394
rect 598 404 614 438
rect 648 404 660 438
rect 598 388 660 404
rect 698 546 714 580
rect 748 546 764 580
rect 875 580 944 581
rect 698 509 764 546
rect 698 475 714 509
rect 748 475 764 509
rect 698 438 764 475
rect 698 404 714 438
rect 748 404 764 438
rect 698 388 764 404
rect 804 531 838 547
rect 804 438 838 497
rect 804 354 838 404
rect 505 320 838 354
rect 875 546 894 580
rect 928 546 944 580
rect 875 509 944 546
rect 875 475 894 509
rect 928 475 944 509
rect 875 438 944 475
rect 875 404 894 438
rect 928 424 944 438
rect 875 390 895 404
rect 929 390 944 424
rect 875 384 944 390
rect 990 580 1040 596
rect 990 546 1006 580
rect 990 497 1040 546
rect 990 463 1006 497
rect 990 414 1040 463
rect 217 294 471 310
rect 505 260 841 286
rect 23 246 274 256
rect 23 240 217 246
rect 23 206 39 240
rect 73 212 217 240
rect 251 212 274 246
rect 73 206 274 212
rect 23 172 73 206
rect 209 178 274 206
rect 310 252 841 260
rect 310 242 539 252
rect 344 226 539 242
rect 791 237 841 252
rect 344 208 360 226
rect 310 192 360 208
rect 610 192 676 218
rect 23 138 39 172
rect 23 17 73 138
rect 109 138 125 172
rect 159 138 175 172
rect 109 94 175 138
rect 209 144 217 178
rect 251 144 274 178
rect 394 185 676 192
rect 394 158 626 185
rect 209 128 274 144
rect 315 124 428 158
rect 610 151 626 158
rect 660 151 676 185
rect 315 94 362 124
rect 109 55 362 94
rect 508 108 574 124
rect 610 119 676 151
rect 721 191 755 218
rect 396 56 412 90
rect 446 56 462 90
rect 396 17 462 56
rect 508 74 524 108
rect 558 85 574 108
rect 721 85 755 157
rect 791 203 807 237
rect 791 169 841 203
rect 791 135 807 169
rect 791 119 841 135
rect 875 236 909 384
rect 990 380 1006 414
rect 990 336 1040 380
rect 1080 580 1146 649
rect 1664 627 1730 649
rect 1282 581 1630 615
rect 1664 593 1680 627
rect 1714 593 1730 627
rect 1878 627 1946 649
rect 1878 593 1895 627
rect 1929 593 1946 627
rect 1080 546 1096 580
rect 1130 546 1146 580
rect 1080 497 1146 546
rect 1080 463 1096 497
rect 1130 463 1146 497
rect 1080 414 1146 463
rect 1080 380 1096 414
rect 1130 380 1146 414
rect 1080 364 1146 380
rect 1192 565 1242 581
rect 1192 531 1208 565
rect 1192 494 1242 531
rect 1192 460 1208 494
rect 1192 423 1242 460
rect 1282 565 1348 581
rect 1282 531 1298 565
rect 1332 531 1348 565
rect 1596 559 1630 581
rect 1987 580 2053 596
rect 1987 559 2003 580
rect 1282 480 1348 531
rect 1282 446 1298 480
rect 1332 446 1348 480
rect 1282 441 1348 446
rect 1388 531 1425 547
rect 1422 497 1425 531
rect 1192 389 1208 423
rect 1388 423 1425 497
rect 1462 527 1528 547
rect 1462 493 1478 527
rect 1512 493 1528 527
rect 1596 546 2003 559
rect 2037 546 2053 580
rect 1596 525 2053 546
rect 1462 491 1528 493
rect 1987 507 2053 525
rect 1462 457 1787 491
rect 1821 457 1837 491
rect 1987 473 2003 507
rect 2037 473 2053 507
rect 1987 457 2053 473
rect 2093 580 2127 649
rect 2093 507 2127 546
rect 2093 457 2127 473
rect 2161 582 2595 615
rect 2161 581 2545 582
rect 2161 423 2195 581
rect 2529 548 2545 581
rect 2579 548 2595 582
rect 1242 389 1388 407
rect 1422 389 1568 423
rect 1602 389 2195 423
rect 2229 539 2495 547
rect 2229 505 2245 539
rect 2279 513 2445 539
rect 2279 505 2295 513
rect 2229 438 2295 505
rect 2429 505 2445 513
rect 2479 505 2495 539
rect 2229 404 2245 438
rect 2279 404 2295 438
rect 1192 373 1425 389
rect 943 320 1040 336
rect 943 286 958 320
rect 992 307 1040 320
rect 1207 323 1341 339
rect 1207 307 1223 323
rect 992 289 1223 307
rect 1257 289 1291 323
rect 1325 289 1341 323
rect 992 286 1341 289
rect 943 273 1341 286
rect 943 270 1040 273
rect 875 202 893 236
rect 927 202 943 236
rect 875 168 943 202
rect 875 134 893 168
rect 927 134 943 168
rect 875 85 943 134
rect 558 74 943 85
rect 508 51 943 74
rect 989 210 1040 270
rect 1388 253 1425 373
rect 1459 329 1703 355
rect 1459 295 1475 329
rect 1509 295 1543 329
rect 1577 295 1611 329
rect 1645 295 1703 329
rect 1459 287 1703 295
rect 1753 302 1895 355
rect 1753 268 1769 302
rect 1803 268 1837 302
rect 1871 268 1895 302
rect 1945 339 2087 355
rect 1945 305 1964 339
rect 1998 305 2032 339
rect 2066 305 2087 339
rect 1945 289 2087 305
rect 1375 239 1425 253
rect 989 176 1005 210
rect 1039 176 1040 210
rect 989 120 1040 176
rect 989 86 1005 120
rect 1039 86 1040 120
rect 989 70 1040 86
rect 1075 210 1141 226
rect 1075 176 1091 210
rect 1125 176 1141 210
rect 1075 120 1141 176
rect 1075 86 1091 120
rect 1125 86 1141 120
rect 1187 205 1203 239
rect 1237 237 1425 239
rect 1237 205 1375 237
rect 1187 167 1237 205
rect 1409 203 1425 237
rect 1187 133 1203 167
rect 1187 117 1237 133
rect 1273 169 1339 171
rect 1273 135 1289 169
rect 1323 135 1339 169
rect 1075 17 1141 86
rect 1273 85 1339 135
rect 1375 169 1425 203
rect 1461 237 1665 253
rect 1753 252 1895 268
rect 1495 219 1665 237
rect 1495 203 1511 219
rect 1461 187 1511 203
rect 1631 218 1665 219
rect 1631 190 2023 218
rect 1409 153 1425 169
rect 1547 169 1597 185
rect 1631 184 1989 190
rect 1547 153 1563 169
rect 1409 135 1563 153
rect 1973 156 1989 184
rect 1375 119 1597 135
rect 1631 127 1851 150
rect 1631 116 1817 127
rect 1631 85 1665 116
rect 1273 51 1665 85
rect 1801 93 1817 116
rect 1699 48 1715 82
rect 1749 48 1765 82
rect 1801 70 1851 93
rect 1887 127 1937 150
rect 1887 93 1903 127
rect 1699 17 1765 48
rect 1887 17 1937 93
rect 1973 120 2023 156
rect 1973 86 1989 120
rect 1973 70 2023 86
rect 2059 190 2109 206
rect 2059 156 2075 190
rect 2059 120 2109 156
rect 2059 86 2075 120
rect 2059 17 2109 86
rect 2143 85 2177 389
rect 2229 206 2295 404
rect 2211 179 2295 206
rect 2329 463 2395 479
rect 2329 429 2345 463
rect 2379 429 2395 463
rect 2329 424 2395 429
rect 2329 390 2335 424
rect 2369 390 2395 424
rect 2429 446 2495 505
rect 2529 514 2595 548
rect 2529 480 2545 514
rect 2579 480 2595 514
rect 2629 582 2695 596
rect 2629 548 2645 582
rect 2679 548 2695 582
rect 2629 514 2695 548
rect 2629 480 2645 514
rect 2679 480 2695 514
rect 2629 446 2695 480
rect 2429 440 2645 446
rect 2429 406 2445 440
rect 2479 412 2645 440
rect 2679 412 2695 446
rect 2775 580 2841 596
rect 2775 546 2791 580
rect 2825 546 2841 580
rect 2775 497 2841 546
rect 2775 463 2791 497
rect 2825 463 2841 497
rect 2775 414 2841 463
rect 2479 406 2495 412
rect 2429 390 2495 406
rect 2329 221 2395 390
rect 2775 380 2791 414
rect 2825 380 2841 414
rect 2775 378 2841 380
rect 2430 289 2567 356
rect 2601 344 2841 378
rect 2875 580 2941 649
rect 2875 546 2891 580
rect 2925 546 2941 580
rect 2875 497 2941 546
rect 2875 463 2891 497
rect 2925 463 2941 497
rect 2875 414 2941 463
rect 2875 380 2891 414
rect 2925 380 2941 414
rect 2875 364 2941 380
rect 2975 580 3041 596
rect 2975 546 2991 580
rect 3025 546 3041 580
rect 2975 497 3041 546
rect 2975 463 2991 497
rect 3025 463 3041 497
rect 2975 414 3041 463
rect 3081 580 3131 649
rect 3115 546 3131 580
rect 3081 478 3131 546
rect 3115 444 3131 478
rect 3081 428 3131 444
rect 3165 580 3231 596
rect 3165 546 3181 580
rect 3215 546 3231 580
rect 3165 497 3231 546
rect 3165 463 3181 497
rect 3215 463 3231 497
rect 2975 380 2991 414
rect 3025 394 3041 414
rect 3165 414 3231 463
rect 3265 580 3331 649
rect 3265 546 3281 580
rect 3315 546 3331 580
rect 3265 478 3331 546
rect 3265 444 3281 478
rect 3315 444 3331 478
rect 3265 428 3331 444
rect 3165 394 3181 414
rect 3025 380 3181 394
rect 3215 394 3231 414
rect 3215 380 3335 394
rect 2975 360 3335 380
rect 2601 310 2616 344
rect 2650 310 2666 344
rect 2601 294 2666 310
rect 2708 294 2773 310
rect 2430 255 2446 289
rect 2480 260 2567 289
rect 2708 260 2724 294
rect 2758 260 2773 294
rect 2480 255 2773 260
rect 2533 226 2773 255
rect 2329 192 2499 221
rect 2807 192 2841 344
rect 2329 187 2635 192
rect 2245 153 2295 179
rect 2465 172 2635 187
rect 2465 158 2585 172
rect 2245 145 2431 153
rect 2211 124 2431 145
rect 2572 138 2585 158
rect 2619 138 2635 172
rect 2211 123 2535 124
rect 2211 119 2415 123
rect 2397 89 2415 119
rect 2449 89 2485 123
rect 2519 89 2535 123
rect 2572 119 2635 138
rect 2669 184 2735 192
rect 2669 150 2685 184
rect 2719 150 2735 184
rect 2397 85 2535 89
rect 2669 116 2735 150
rect 2781 172 2841 192
rect 2781 138 2797 172
rect 2831 138 2841 172
rect 2781 119 2841 138
rect 2875 310 3242 326
rect 2875 276 3004 310
rect 3038 276 3072 310
rect 3106 276 3140 310
rect 3174 276 3208 310
rect 2875 260 3242 276
rect 2669 85 2671 116
rect 2143 51 2313 85
rect 2347 51 2363 85
rect 2397 82 2671 85
rect 2705 85 2735 116
rect 2875 85 2909 260
rect 3289 226 3335 360
rect 2705 82 2909 85
rect 2397 51 2909 82
rect 2943 210 2977 226
rect 2943 120 2977 176
rect 2943 17 2977 86
rect 3013 210 3335 226
rect 3013 176 3029 210
rect 3063 192 3201 210
rect 3013 120 3063 176
rect 3185 176 3201 192
rect 3235 192 3335 210
rect 3013 86 3029 120
rect 3013 70 3063 86
rect 3099 142 3149 158
rect 3099 108 3115 142
rect 3099 17 3149 108
rect 3185 120 3235 176
rect 3185 86 3201 120
rect 3185 70 3235 86
rect 3271 142 3337 158
rect 3271 108 3287 142
rect 3321 108 3337 142
rect 3271 17 3337 108
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3360 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 3199 649 3233 683
rect 3295 649 3329 683
rect 895 404 928 424
rect 928 404 929 424
rect 895 390 929 404
rect 2335 390 2369 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
<< metal1 >>
rect 0 683 3360 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3360 683
rect 0 617 3360 649
rect 883 424 941 430
rect 883 390 895 424
rect 929 421 941 424
rect 2323 424 2381 430
rect 2323 421 2335 424
rect 929 393 2335 421
rect 929 390 941 393
rect 883 384 941 390
rect 2323 390 2335 393
rect 2369 390 2381 424
rect 2323 384 2381 390
rect 0 17 3360 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3360 17
rect 0 -49 3360 -17
<< labels >>
flabel pwell s 0 0 3360 49 0 FreeSans 200 0 0 0 VNB
port 8 nsew
flabel nbase s 0 617 3360 666 0 FreeSans 200 0 0 0 VPB
port 9 nsew
rlabel comment s 0 0 0 0 4 mux4_4
flabel metal1 s 0 617 3360 666 0 FreeSans 340 0 0 0 VPWR
port 10 nsew
flabel metal1 s 0 0 3360 49 0 FreeSans 340 0 0 0 VGND
port 7 nsew
flabel corelocali s 2527 316 2561 350 0 FreeSans 340 0 0 0 S1
port 6 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A0
port 1 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A0
port 1 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A0
port 1 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 A1
port 2 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 A1
port 2 nsew
flabel corelocali s 1759 316 1793 350 0 FreeSans 340 0 0 0 A2
port 3 nsew
flabel corelocali s 1855 316 1889 350 0 FreeSans 340 0 0 0 A2
port 3 nsew
flabel corelocali s 1951 316 1985 350 0 FreeSans 340 0 0 0 A3
port 4 nsew
flabel corelocali s 2047 316 2081 350 0 FreeSans 340 0 0 0 A3
port 4 nsew
flabel corelocali s 1471 316 1505 350 0 FreeSans 340 0 0 0 S0
port 5 nsew
flabel corelocali s 1567 316 1601 350 0 FreeSans 340 0 0 0 S0
port 5 nsew
flabel corelocali s 1663 316 1697 350 0 FreeSans 340 0 0 0 S0
port 5 nsew
flabel corelocali s 3295 242 3329 276 0 FreeSans 340 0 0 0 X
port 11 nsew
flabel corelocali s 3295 316 3329 350 0 FreeSans 340 0 0 0 X
port 11 nsew
<< properties >>
string FIXED_BBOX 0 0 3360 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1909026
string GDS_START 1884740
<< end >>
