magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 21 199 89 391
rect 379 199 437 475
rect 475 199 541 475
rect 739 325 789 493
rect 927 325 977 493
rect 575 289 688 323
rect 739 291 1083 325
rect 575 199 635 289
rect 1035 181 1083 291
rect 747 145 1083 181
rect 747 51 797 145
rect 909 51 985 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 17 427 73 527
rect 129 265 167 491
rect 217 349 283 490
rect 217 315 345 349
rect 129 199 253 265
rect 17 17 69 165
rect 129 87 167 199
rect 301 165 345 315
rect 634 359 684 527
rect 833 359 883 527
rect 1021 359 1071 527
rect 669 215 991 249
rect 669 165 703 215
rect 301 131 703 165
rect 217 17 267 117
rect 343 61 377 131
rect 417 17 493 97
rect 537 61 571 131
rect 625 17 701 97
rect 841 17 875 111
rect 1029 17 1063 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
rlabel locali s 575 289 688 323 6 A
port 1 nsew signal input
rlabel locali s 575 199 635 289 6 A
port 1 nsew signal input
rlabel locali s 475 199 541 475 6 B
port 2 nsew signal input
rlabel locali s 379 199 437 475 6 C
port 3 nsew signal input
rlabel locali s 21 199 89 391 6 D_N
port 4 nsew signal input
rlabel locali s 1035 181 1083 291 6 X
port 5 nsew signal output
rlabel locali s 927 325 977 493 6 X
port 5 nsew signal output
rlabel locali s 909 51 985 145 6 X
port 5 nsew signal output
rlabel locali s 747 145 1083 181 6 X
port 5 nsew signal output
rlabel locali s 747 51 797 145 6 X
port 5 nsew signal output
rlabel locali s 739 325 789 493 6 X
port 5 nsew signal output
rlabel locali s 739 291 1083 325 6 X
port 5 nsew signal output
rlabel metal1 s 0 -48 1104 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 1104 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1104 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 536002
string GDS_START 527266
<< end >>
