magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 91 47 121 177
rect 185 47 215 177
rect 383 47 413 177
rect 467 47 497 177
rect 571 47 601 177
rect 665 47 695 177
rect 775 47 805 177
rect 859 47 889 177
rect 963 47 993 177
rect 1057 47 1087 177
<< pmoshvt >>
rect 83 297 119 497
rect 177 297 213 497
rect 375 297 411 497
rect 469 297 505 497
rect 563 297 599 497
rect 657 297 693 497
rect 767 297 803 497
rect 861 297 897 497
rect 955 297 991 497
rect 1049 297 1085 497
<< ndiff >>
rect 27 163 91 177
rect 27 129 37 163
rect 71 129 91 163
rect 27 95 91 129
rect 27 61 37 95
rect 71 61 91 95
rect 27 47 91 61
rect 121 163 185 177
rect 121 129 131 163
rect 165 129 185 163
rect 121 95 185 129
rect 121 61 131 95
rect 165 61 185 95
rect 121 47 185 61
rect 215 95 383 177
rect 215 61 225 95
rect 259 61 329 95
rect 363 61 383 95
rect 215 47 383 61
rect 413 95 467 177
rect 413 61 423 95
rect 457 61 467 95
rect 413 47 467 61
rect 497 163 571 177
rect 497 129 517 163
rect 551 129 571 163
rect 497 47 571 129
rect 601 95 665 177
rect 601 61 611 95
rect 645 61 665 95
rect 601 47 665 61
rect 695 95 775 177
rect 695 61 714 95
rect 748 61 775 95
rect 695 47 775 61
rect 805 95 859 177
rect 805 61 815 95
rect 849 61 859 95
rect 805 47 859 61
rect 889 163 963 177
rect 889 129 909 163
rect 943 129 963 163
rect 889 47 963 129
rect 993 163 1057 177
rect 993 129 1003 163
rect 1037 129 1057 163
rect 993 95 1057 129
rect 993 61 1003 95
rect 1037 61 1057 95
rect 993 47 1057 61
rect 1087 163 1139 177
rect 1087 129 1097 163
rect 1131 129 1139 163
rect 1087 95 1139 129
rect 1087 61 1097 95
rect 1131 61 1139 95
rect 1087 47 1139 61
<< pdiff >>
rect 27 483 83 497
rect 27 449 37 483
rect 71 449 83 483
rect 27 393 83 449
rect 27 359 37 393
rect 71 359 83 393
rect 27 297 83 359
rect 119 409 177 497
rect 119 375 131 409
rect 165 375 177 409
rect 119 341 177 375
rect 119 307 131 341
rect 165 307 177 341
rect 119 297 177 307
rect 213 477 267 497
rect 213 443 225 477
rect 259 443 267 477
rect 213 349 267 443
rect 213 315 225 349
rect 259 315 267 349
rect 213 297 267 315
rect 321 477 375 497
rect 321 443 329 477
rect 363 443 375 477
rect 321 297 375 443
rect 411 409 469 497
rect 411 375 423 409
rect 457 375 469 409
rect 411 297 469 375
rect 505 477 563 497
rect 505 443 517 477
rect 551 443 563 477
rect 505 297 563 443
rect 599 409 657 497
rect 599 375 611 409
rect 645 375 657 409
rect 599 297 657 375
rect 693 477 767 497
rect 693 443 713 477
rect 747 443 767 477
rect 693 407 767 443
rect 693 373 713 407
rect 747 373 767 407
rect 693 297 767 373
rect 803 477 861 497
rect 803 443 815 477
rect 849 443 861 477
rect 803 297 861 443
rect 897 477 955 497
rect 897 443 909 477
rect 943 443 955 477
rect 897 409 955 443
rect 897 375 909 409
rect 943 375 955 409
rect 897 297 955 375
rect 991 477 1049 497
rect 991 443 1003 477
rect 1037 443 1049 477
rect 991 297 1049 443
rect 1085 477 1144 497
rect 1085 443 1098 477
rect 1132 443 1144 477
rect 1085 409 1144 443
rect 1085 375 1098 409
rect 1132 375 1144 409
rect 1085 341 1144 375
rect 1085 307 1098 341
rect 1132 307 1144 341
rect 1085 297 1144 307
<< ndiffc >>
rect 37 129 71 163
rect 37 61 71 95
rect 131 129 165 163
rect 131 61 165 95
rect 225 61 259 95
rect 329 61 363 95
rect 423 61 457 95
rect 517 129 551 163
rect 611 61 645 95
rect 714 61 748 95
rect 815 61 849 95
rect 909 129 943 163
rect 1003 129 1037 163
rect 1003 61 1037 95
rect 1097 129 1131 163
rect 1097 61 1131 95
<< pdiffc >>
rect 37 449 71 483
rect 37 359 71 393
rect 131 375 165 409
rect 131 307 165 341
rect 225 443 259 477
rect 225 315 259 349
rect 329 443 363 477
rect 423 375 457 409
rect 517 443 551 477
rect 611 375 645 409
rect 713 443 747 477
rect 713 373 747 407
rect 815 443 849 477
rect 909 443 943 477
rect 909 375 943 409
rect 1003 443 1037 477
rect 1098 443 1132 477
rect 1098 375 1132 409
rect 1098 307 1132 341
<< poly >>
rect 83 497 119 523
rect 177 497 213 523
rect 375 497 411 523
rect 469 497 505 523
rect 563 497 599 523
rect 657 497 693 523
rect 767 497 803 523
rect 861 497 897 523
rect 955 497 991 523
rect 1049 497 1085 523
rect 83 282 119 297
rect 177 282 213 297
rect 375 282 411 297
rect 469 282 505 297
rect 563 282 599 297
rect 657 282 693 297
rect 767 282 803 297
rect 861 282 897 297
rect 955 282 991 297
rect 1049 282 1085 297
rect 81 265 121 282
rect 175 265 215 282
rect 373 265 413 282
rect 467 265 507 282
rect 561 265 601 282
rect 655 265 695 282
rect 765 265 805 282
rect 859 265 899 282
rect 953 265 993 282
rect 1047 265 1087 282
rect 22 249 215 265
rect 22 215 34 249
rect 68 215 215 249
rect 22 199 215 215
rect 361 249 425 265
rect 361 215 371 249
rect 405 215 425 249
rect 361 199 425 215
rect 467 249 601 265
rect 467 215 517 249
rect 551 215 601 249
rect 467 199 601 215
rect 643 249 707 265
rect 643 215 653 249
rect 687 215 707 249
rect 643 199 707 215
rect 753 249 817 265
rect 753 215 763 249
rect 797 215 817 249
rect 753 199 817 215
rect 859 249 993 265
rect 859 215 909 249
rect 943 215 993 249
rect 859 199 993 215
rect 1035 249 1099 265
rect 1035 215 1045 249
rect 1079 215 1099 249
rect 1035 199 1099 215
rect 91 177 121 199
rect 185 177 215 199
rect 383 177 413 199
rect 467 177 497 199
rect 571 177 601 199
rect 665 177 695 199
rect 775 177 805 199
rect 859 177 889 199
rect 963 177 993 199
rect 1057 177 1087 199
rect 91 21 121 47
rect 185 21 215 47
rect 383 21 413 47
rect 467 21 497 47
rect 571 21 601 47
rect 665 21 695 47
rect 775 21 805 47
rect 859 21 889 47
rect 963 21 993 47
rect 1057 21 1087 47
<< polycont >>
rect 34 215 68 249
rect 371 215 405 249
rect 517 215 551 249
rect 653 215 687 249
rect 763 215 797 249
rect 909 215 943 249
rect 1045 215 1079 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 18 483 275 493
rect 18 449 37 483
rect 71 477 275 483
rect 71 459 225 477
rect 71 449 87 459
rect 18 393 87 449
rect 259 443 275 477
rect 18 359 37 393
rect 71 359 87 393
rect 121 409 181 425
rect 121 375 131 409
rect 165 375 181 409
rect 121 341 181 375
rect 18 249 84 323
rect 18 215 34 249
rect 68 215 84 249
rect 121 307 131 341
rect 165 307 181 341
rect 121 181 181 307
rect 225 391 275 443
rect 321 477 755 493
rect 321 443 329 477
rect 363 459 517 477
rect 363 443 371 459
rect 321 425 371 443
rect 509 443 517 459
rect 551 459 713 477
rect 551 443 559 459
rect 509 425 559 443
rect 705 443 713 459
rect 747 443 755 477
rect 415 409 465 425
rect 415 391 423 409
rect 225 375 423 391
rect 457 391 465 409
rect 603 409 653 425
rect 603 391 611 409
rect 457 375 611 391
rect 645 375 653 409
rect 225 357 653 375
rect 705 407 755 443
rect 807 477 857 527
rect 807 443 815 477
rect 849 443 857 477
rect 807 425 857 443
rect 901 477 951 493
rect 901 443 909 477
rect 943 443 951 477
rect 705 373 713 407
rect 747 391 755 407
rect 901 409 951 443
rect 995 477 1045 527
rect 995 443 1003 477
rect 1037 443 1045 477
rect 995 425 1045 443
rect 1098 477 1139 493
rect 1132 443 1139 477
rect 901 391 909 409
rect 747 375 909 391
rect 943 391 951 409
rect 1098 409 1139 443
rect 943 375 1098 391
rect 1132 375 1139 409
rect 747 373 1139 375
rect 705 357 1139 373
rect 225 349 275 357
rect 259 315 275 349
rect 1098 341 1139 357
rect 225 299 275 315
rect 346 289 713 323
rect 346 249 438 289
rect 346 215 371 249
rect 405 215 438 249
rect 472 249 603 255
rect 472 215 517 249
rect 551 215 603 249
rect 637 249 713 289
rect 637 215 653 249
rect 687 215 713 249
rect 747 289 1054 323
rect 1132 307 1139 341
rect 1098 291 1139 307
rect 747 249 813 289
rect 1020 255 1054 289
rect 747 215 763 249
rect 797 215 813 249
rect 847 249 983 255
rect 847 215 909 249
rect 943 215 983 249
rect 1020 249 1177 255
rect 1020 215 1045 249
rect 1079 215 1177 249
rect 21 163 71 179
rect 121 173 959 181
rect 21 129 37 163
rect 21 95 71 129
rect 21 61 37 95
rect 105 163 959 173
rect 105 129 131 163
rect 165 145 517 163
rect 165 129 181 145
rect 487 129 517 145
rect 551 145 909 163
rect 551 129 567 145
rect 883 129 909 145
rect 943 129 959 163
rect 1003 163 1053 181
rect 1037 129 1053 163
rect 105 95 181 129
rect 105 61 131 95
rect 165 61 181 95
rect 225 95 363 111
rect 714 95 748 111
rect 1003 95 1053 129
rect 259 61 329 95
rect 21 17 71 61
rect 225 17 363 61
rect 397 61 423 95
rect 457 61 611 95
rect 645 61 661 95
rect 397 51 661 61
rect 714 17 748 61
rect 789 61 815 95
rect 849 61 1003 95
rect 1037 61 1053 95
rect 789 51 1053 61
rect 1097 163 1131 181
rect 1097 95 1131 129
rect 1097 17 1131 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
flabel corelocali s 391 289 425 323 0 FreeSans 400 0 0 0 B2
port 4 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 400 0 0 0 C1
port 5 nsew
flabel corelocali s 1058 238 1058 238 0 FreeSans 400 180 0 0 A2
port 2 nsew
flabel corelocali s 933 238 933 238 0 FreeSans 400 180 0 0 A1
port 1 nsew
flabel corelocali s 511 238 511 238 0 FreeSans 400 0 0 0 B1
port 3 nsew
flabel corelocali s 391 221 425 255 0 FreeSans 400 0 0 0 B2
port 4 nsew
flabel corelocali s 132 221 166 255 0 FreeSans 400 0 0 0 Y
port 10 nsew
flabel corelocali s 30 289 64 323 0 FreeSans 400 0 0 0 C1
port 5 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew
rlabel comment s 0 0 0 0 4 a221oi_2
<< properties >>
string FIXED_BBOX 0 0 1196 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1231362
string GDS_START 1221708
<< end >>
