magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 1382 704
rect 356 318 766 332
<< pwell >>
rect 0 0 1344 49
<< scnmos >>
rect 84 74 114 222
rect 172 74 202 222
rect 284 74 314 222
rect 370 74 400 222
rect 484 74 514 222
rect 570 74 600 222
<< pmoshvt >>
rect 85 368 115 592
rect 175 368 205 592
rect 265 368 295 592
rect 386 368 416 592
rect 506 368 536 592
rect 628 368 658 592
rect 748 368 778 592
rect 870 368 900 592
rect 960 368 990 592
rect 1050 368 1080 592
rect 1140 368 1170 592
rect 1230 368 1260 592
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 210 172 222
rect 114 176 125 210
rect 159 176 172 210
rect 114 120 172 176
rect 114 86 125 120
rect 159 86 172 120
rect 114 74 172 86
rect 202 152 284 222
rect 202 118 225 152
rect 259 118 284 152
rect 202 74 284 118
rect 314 210 370 222
rect 314 176 325 210
rect 359 176 370 210
rect 314 120 370 176
rect 314 86 325 120
rect 359 86 370 120
rect 314 74 370 86
rect 400 127 484 222
rect 400 93 425 127
rect 459 93 484 127
rect 400 74 484 93
rect 514 202 570 222
rect 514 168 525 202
rect 559 168 570 202
rect 514 120 570 168
rect 514 86 525 120
rect 559 86 570 120
rect 514 74 570 86
rect 600 118 708 222
rect 600 84 611 118
rect 645 84 708 118
rect 600 74 708 84
rect 615 72 708 74
<< pdiff >>
rect 313 604 368 616
rect 313 592 324 604
rect 27 580 85 592
rect 27 546 38 580
rect 72 546 85 580
rect 27 497 85 546
rect 27 463 38 497
rect 72 463 85 497
rect 27 414 85 463
rect 27 380 38 414
rect 72 380 85 414
rect 27 368 85 380
rect 115 575 175 592
rect 115 541 128 575
rect 162 541 175 575
rect 115 368 175 541
rect 205 580 265 592
rect 205 546 218 580
rect 252 546 265 580
rect 205 502 265 546
rect 205 468 218 502
rect 252 468 265 502
rect 205 368 265 468
rect 295 570 324 592
rect 358 592 368 604
rect 554 604 610 616
rect 554 592 565 604
rect 358 570 386 592
rect 295 368 386 570
rect 416 400 506 592
rect 416 368 444 400
rect 434 366 444 368
rect 478 368 506 400
rect 536 570 565 592
rect 599 592 610 604
rect 796 604 852 616
rect 796 592 807 604
rect 599 570 628 592
rect 536 368 628 570
rect 658 400 748 592
rect 658 368 686 400
rect 478 366 488 368
rect 434 354 488 366
rect 676 366 686 368
rect 720 368 748 400
rect 778 570 807 592
rect 841 592 852 604
rect 841 570 870 592
rect 778 368 870 570
rect 900 526 960 592
rect 900 492 913 526
rect 947 492 960 526
rect 900 368 960 492
rect 990 577 1050 592
rect 990 543 1003 577
rect 1037 543 1050 577
rect 990 368 1050 543
rect 1080 584 1140 592
rect 1080 550 1093 584
rect 1127 550 1140 584
rect 1080 506 1140 550
rect 1080 472 1093 506
rect 1127 472 1140 506
rect 1080 368 1140 472
rect 1170 577 1230 592
rect 1170 543 1183 577
rect 1217 543 1230 577
rect 1170 368 1230 543
rect 1260 580 1317 592
rect 1260 546 1273 580
rect 1307 546 1317 580
rect 1260 497 1317 546
rect 1260 463 1273 497
rect 1307 463 1317 497
rect 1260 414 1317 463
rect 1260 380 1273 414
rect 1307 380 1317 414
rect 1260 368 1317 380
rect 720 366 730 368
rect 676 354 730 366
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 125 176 159 210
rect 125 86 159 120
rect 225 118 259 152
rect 325 176 359 210
rect 325 86 359 120
rect 425 93 459 127
rect 525 168 559 202
rect 525 86 559 120
rect 611 84 645 118
<< pdiffc >>
rect 38 546 72 580
rect 38 463 72 497
rect 38 380 72 414
rect 128 541 162 575
rect 218 546 252 580
rect 218 468 252 502
rect 324 570 358 604
rect 444 366 478 400
rect 565 570 599 604
rect 686 366 720 400
rect 807 570 841 604
rect 913 492 947 526
rect 1003 543 1037 577
rect 1093 550 1127 584
rect 1093 472 1127 506
rect 1183 543 1217 577
rect 1273 546 1307 580
rect 1273 463 1307 497
rect 1273 380 1307 414
<< poly >>
rect 85 592 115 618
rect 175 592 205 618
rect 265 592 295 618
rect 386 592 416 618
rect 506 592 536 618
rect 85 353 115 368
rect 175 353 205 368
rect 265 353 295 368
rect 386 353 416 368
rect 628 592 658 618
rect 748 592 778 618
rect 506 353 536 368
rect 628 353 658 368
rect 870 592 900 618
rect 960 592 990 618
rect 1050 592 1080 618
rect 1140 592 1170 618
rect 1230 592 1260 618
rect 748 353 778 368
rect 870 353 900 368
rect 960 353 990 368
rect 1050 353 1080 368
rect 1140 353 1170 368
rect 1230 353 1260 368
rect 82 336 118 353
rect 172 336 208 353
rect 82 320 208 336
rect 82 300 137 320
rect 84 286 137 300
rect 171 286 208 320
rect 84 270 208 286
rect 262 336 298 353
rect 383 339 419 353
rect 503 339 539 353
rect 625 339 661 353
rect 745 339 781 353
rect 262 320 328 336
rect 262 286 278 320
rect 312 286 328 320
rect 383 309 781 339
rect 84 222 114 270
rect 172 222 202 270
rect 262 267 328 286
rect 262 237 400 267
rect 284 222 314 237
rect 370 222 400 237
rect 484 222 514 309
rect 570 222 600 309
rect 84 48 114 74
rect 172 48 202 74
rect 284 48 314 74
rect 370 48 400 74
rect 484 48 514 74
rect 570 48 600 74
rect 751 134 781 309
rect 867 302 903 353
rect 957 302 993 353
rect 1047 302 1083 353
rect 1140 336 1173 353
rect 1227 336 1260 353
rect 859 286 1083 302
rect 859 252 875 286
rect 909 252 943 286
rect 977 252 1083 286
rect 859 236 1083 252
rect 1143 320 1257 336
rect 1143 286 1177 320
rect 1211 286 1257 320
rect 1143 252 1257 286
rect 1143 218 1177 252
rect 1211 218 1257 252
rect 1143 184 1257 218
rect 1143 150 1177 184
rect 1211 150 1257 184
rect 751 118 1095 134
rect 751 84 773 118
rect 807 84 841 118
rect 875 84 909 118
rect 943 84 977 118
rect 1011 84 1045 118
rect 1079 84 1095 118
rect 751 68 1095 84
rect 1143 116 1257 150
rect 1143 82 1177 116
rect 1211 82 1257 116
rect 1143 66 1257 82
<< polycont >>
rect 137 286 171 320
rect 278 286 312 320
rect 875 252 909 286
rect 943 252 977 286
rect 1177 286 1211 320
rect 1177 218 1211 252
rect 1177 150 1211 184
rect 773 84 807 118
rect 841 84 875 118
rect 909 84 943 118
rect 977 84 1011 118
rect 1045 84 1079 118
rect 1177 82 1211 116
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 22 580 72 596
rect 22 546 38 580
rect 22 502 72 546
rect 112 575 178 649
rect 308 604 1053 615
rect 112 541 128 575
rect 162 541 178 575
rect 112 536 178 541
rect 218 580 268 596
rect 252 546 268 580
rect 308 570 324 604
rect 358 570 565 604
rect 599 570 807 604
rect 841 581 1053 604
rect 841 570 857 581
rect 987 577 1053 581
rect 218 536 268 546
rect 897 536 947 547
rect 987 543 1003 577
rect 1037 543 1053 577
rect 987 540 1053 543
rect 1093 584 1127 600
rect 218 526 947 536
rect 218 502 913 526
rect 22 497 218 502
rect 22 463 38 497
rect 72 468 218 497
rect 252 468 268 502
rect 897 492 913 502
rect 1093 506 1127 550
rect 1167 577 1233 649
rect 1167 543 1183 577
rect 1217 543 1233 577
rect 1167 540 1233 543
rect 1273 580 1323 596
rect 1307 546 1323 580
rect 1273 506 1323 546
rect 947 492 1093 506
rect 897 472 1093 492
rect 1127 497 1323 506
rect 1127 472 1273 497
rect 22 414 72 463
rect 325 438 804 468
rect 1307 463 1323 497
rect 325 434 1227 438
rect 22 380 38 414
rect 22 364 72 380
rect 121 384 359 434
rect 770 404 1227 434
rect 121 320 187 384
rect 428 366 444 400
rect 478 366 686 400
rect 720 370 736 400
rect 720 366 1061 370
rect 428 350 1061 366
rect 670 336 1061 350
rect 121 286 137 320
rect 171 286 187 320
rect 121 270 187 286
rect 262 320 328 336
rect 262 286 278 320
rect 312 304 328 320
rect 312 302 551 304
rect 312 286 993 302
rect 262 270 875 286
rect 409 252 875 270
rect 909 252 943 286
rect 977 252 993 286
rect 409 236 993 252
rect 23 210 73 226
rect 23 176 39 210
rect 23 120 73 176
rect 23 86 39 120
rect 23 17 73 86
rect 109 210 375 236
rect 109 176 125 210
rect 159 202 325 210
rect 159 176 175 202
rect 109 120 175 176
rect 309 176 325 202
rect 359 202 375 210
rect 1027 202 1061 336
rect 359 176 525 202
rect 309 168 525 176
rect 559 168 1061 202
rect 1161 320 1227 404
rect 1273 414 1323 463
rect 1307 380 1323 414
rect 1273 364 1323 380
rect 1161 286 1177 320
rect 1211 286 1227 320
rect 1161 252 1227 286
rect 1161 218 1177 252
rect 1211 218 1227 252
rect 1161 184 1227 218
rect 109 86 125 120
rect 159 86 175 120
rect 109 70 175 86
rect 209 152 275 168
rect 209 118 225 152
rect 259 118 275 152
rect 209 17 275 118
rect 309 120 375 168
rect 309 86 325 120
rect 359 86 375 120
rect 309 70 375 86
rect 409 127 475 134
rect 409 93 425 127
rect 459 93 475 127
rect 409 17 475 93
rect 509 120 575 168
rect 1161 150 1177 184
rect 1211 150 1227 184
rect 509 86 525 120
rect 559 86 575 120
rect 509 70 575 86
rect 611 118 673 134
rect 645 84 673 118
rect 611 17 673 84
rect 757 118 1127 134
rect 757 84 773 118
rect 807 84 841 118
rect 875 84 909 118
rect 943 84 977 118
rect 1011 84 1045 118
rect 1079 84 1127 118
rect 757 68 1127 84
rect 1161 116 1227 150
rect 1161 82 1177 116
rect 1211 82 1227 116
rect 1161 66 1227 82
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
<< metal1 >>
rect 0 683 1344 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 0 617 1344 649
rect 0 17 1344 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
rect 0 -49 1344 -17
<< labels >>
rlabel comment s 0 0 0 0 4 nor3_4
flabel pwell s 0 0 1344 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 0 617 1344 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 1344 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 1344 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 127 390 161 424 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 223 390 257 424 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 319 390 353 424 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 415 242 449 276 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 511 242 545 276 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 799 94 833 128 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 895 94 929 128 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 991 94 1025 128 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 1087 94 1121 128 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 127 94 161 128 0 FreeSans 340 0 0 0 Y
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 1344 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1972228
string GDS_START 1962236
<< end >>
