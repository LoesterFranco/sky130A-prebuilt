magic
tech sky130A
magscale 1 2
timestamp 1604502741
<< locali >>
rect 551 364 655 596
rect 25 236 91 310
rect 407 270 473 356
rect 621 226 655 364
rect 575 70 655 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 23 386 89 596
rect 123 420 189 649
rect 260 398 326 572
rect 23 352 166 386
rect 260 364 373 398
rect 451 390 517 649
rect 132 326 166 352
rect 132 260 305 326
rect 132 202 166 260
rect 339 236 373 364
rect 507 260 587 326
rect 507 236 541 260
rect 23 136 166 202
rect 200 17 305 226
rect 339 202 541 236
rect 339 108 409 202
rect 453 17 536 168
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel locali s 407 270 473 356 6 A
port 1 nsew signal input
rlabel locali s 25 236 91 310 6 B_N
port 2 nsew signal input
rlabel locali s 621 226 655 364 6 X
port 3 nsew signal output
rlabel locali s 575 70 655 226 6 X
port 3 nsew signal output
rlabel locali s 551 364 655 596 6 X
port 3 nsew signal output
rlabel metal1 s 0 -49 672 49 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 617 672 715 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 761892
string GDS_START 756080
<< end >>
