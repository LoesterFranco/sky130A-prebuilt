magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 644 561
rect 19 299 85 527
rect 188 383 240 527
rect 390 401 446 471
rect 342 367 446 401
rect 18 195 84 265
rect 120 199 205 265
rect 239 199 291 265
rect 342 199 387 367
rect 482 333 530 467
rect 421 299 530 333
rect 19 17 85 161
rect 120 53 159 199
rect 239 132 273 199
rect 421 165 455 299
rect 489 199 537 265
rect 193 53 273 132
rect 307 131 530 165
rect 307 51 341 131
rect 381 17 447 97
rect 481 59 530 131
rect 0 -17 644 17
<< obsli1 >>
rect 120 349 154 461
rect 274 435 340 469
rect 274 349 308 435
rect 120 315 308 349
<< metal1 >>
rect 0 496 644 592
rect 0 -48 644 48
<< labels >>
rlabel locali s 239 199 291 265 6 A1
port 1 nsew signal input
rlabel locali s 239 132 273 199 6 A1
port 1 nsew signal input
rlabel locali s 193 53 273 132 6 A1
port 1 nsew signal input
rlabel locali s 120 199 205 265 6 A2
port 2 nsew signal input
rlabel locali s 120 53 159 199 6 A2
port 2 nsew signal input
rlabel locali s 18 195 84 265 6 A3
port 3 nsew signal input
rlabel locali s 390 401 446 471 6 B1
port 4 nsew signal input
rlabel locali s 342 367 446 401 6 B1
port 4 nsew signal input
rlabel locali s 342 199 387 367 6 B1
port 4 nsew signal input
rlabel locali s 489 199 537 265 6 C1
port 5 nsew signal input
rlabel locali s 482 333 530 467 6 Y
port 6 nsew signal output
rlabel locali s 481 59 530 131 6 Y
port 6 nsew signal output
rlabel locali s 421 299 530 333 6 Y
port 6 nsew signal output
rlabel locali s 421 165 455 299 6 Y
port 6 nsew signal output
rlabel locali s 307 131 530 165 6 Y
port 6 nsew signal output
rlabel locali s 307 51 341 131 6 Y
port 6 nsew signal output
rlabel locali s 381 17 447 97 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 19 17 85 161 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 644 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 644 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 188 383 240 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 19 299 85 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 644 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 644 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3601492
string GDS_START 3595338
<< end >>
