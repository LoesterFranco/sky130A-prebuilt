magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1196 561
rect 103 369 186 527
rect 396 455 462 527
rect 564 455 630 527
rect 98 153 156 335
rect 190 153 256 285
rect 379 289 1179 345
rect 1135 171 1179 289
rect 103 17 186 119
rect 469 17 535 97
rect 637 17 703 97
rect 829 123 1179 171
rect 0 -17 1196 17
<< obsli1 >>
rect 17 353 69 493
rect 220 353 271 493
rect 313 421 362 493
rect 496 421 530 493
rect 664 421 1179 493
rect 313 387 1179 421
rect 379 379 1179 387
rect 17 255 64 353
rect 17 221 30 255
rect 17 133 64 221
rect 220 319 345 353
rect 290 255 345 319
rect 290 205 762 255
rect 796 221 862 255
rect 896 221 1101 255
rect 796 205 1101 221
rect 17 56 69 133
rect 290 119 345 205
rect 220 51 345 119
rect 379 131 795 171
rect 379 51 435 131
rect 569 55 603 131
rect 737 89 795 131
rect 737 51 1147 89
<< obsli1c >>
rect 30 221 64 255
rect 862 221 896 255
<< metal1 >>
rect 0 496 1196 592
rect 0 -48 1196 48
<< obsm1 >>
rect 17 255 76 261
rect 17 221 30 255
rect 64 252 76 255
rect 850 255 908 261
rect 850 252 862 255
rect 64 224 862 252
rect 64 221 76 224
rect 17 215 76 221
rect 850 221 862 224
rect 896 221 908 255
rect 850 215 908 221
<< labels >>
rlabel locali s 98 153 156 335 6 A
port 1 nsew signal input
rlabel locali s 190 153 256 285 6 TE_B
port 2 nsew signal input
rlabel locali s 1135 171 1179 289 6 Z
port 3 nsew signal output
rlabel locali s 829 123 1179 171 6 Z
port 3 nsew signal output
rlabel locali s 379 289 1179 345 6 Z
port 3 nsew signal output
rlabel locali s 637 17 703 97 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 469 17 535 97 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 103 17 186 119 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 1196 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1196 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 564 455 630 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 396 455 462 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 103 369 186 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 1196 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 1196 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2870408
string GDS_START 2860962
<< end >>
