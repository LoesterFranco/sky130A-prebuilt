magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 113 265 165 450
rect 199 409 265 489
rect 415 409 535 493
rect 199 363 535 409
rect 199 319 265 363
rect 299 269 349 323
rect 17 199 79 265
rect 113 199 216 265
rect 284 199 349 269
rect 383 204 454 323
rect 488 165 535 363
rect 345 51 535 165
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 19 299 79 527
rect 308 455 374 527
rect 19 123 290 165
rect 19 51 80 123
rect 114 17 180 89
rect 214 51 290 123
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
rlabel locali s 17 199 79 265 6 A1
port 1 nsew signal input
rlabel locali s 113 265 165 450 6 A2
port 2 nsew signal input
rlabel locali s 113 199 216 265 6 A2
port 2 nsew signal input
rlabel locali s 299 269 349 323 6 B1
port 3 nsew signal input
rlabel locali s 284 199 349 269 6 B1
port 3 nsew signal input
rlabel locali s 383 204 454 323 6 C1
port 4 nsew signal input
rlabel locali s 488 165 535 363 6 Y
port 5 nsew signal output
rlabel locali s 415 409 535 493 6 Y
port 5 nsew signal output
rlabel locali s 345 51 535 165 6 Y
port 5 nsew signal output
rlabel locali s 199 409 265 489 6 Y
port 5 nsew signal output
rlabel locali s 199 363 535 409 6 Y
port 5 nsew signal output
rlabel locali s 199 319 265 363 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -48 552 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 552 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 552 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2589902
string GDS_START 2584602
<< end >>
