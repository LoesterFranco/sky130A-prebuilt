magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 184 47 214 131
rect 280 47 310 131
rect 376 47 406 131
rect 472 47 502 131
<< pmoshvt >>
rect 90 297 126 497
rect 186 297 222 497
rect 282 297 318 497
rect 378 297 414 497
rect 474 297 510 497
rect 570 297 606 497
<< ndiff >>
rect 108 95 184 131
rect 108 61 139 95
rect 173 61 184 95
rect 108 47 184 61
rect 214 106 280 131
rect 214 72 235 106
rect 269 72 280 106
rect 214 47 280 72
rect 310 95 376 131
rect 310 61 331 95
rect 365 61 376 95
rect 310 47 376 61
rect 406 106 472 131
rect 406 72 427 106
rect 461 72 472 106
rect 406 47 472 72
rect 502 95 591 131
rect 502 61 523 95
rect 557 61 591 95
rect 502 47 591 61
<< pdiff >>
rect 27 478 90 497
rect 27 444 43 478
rect 77 444 90 478
rect 27 410 90 444
rect 27 376 43 410
rect 77 376 90 410
rect 27 297 90 376
rect 126 471 186 497
rect 126 437 139 471
rect 173 437 186 471
rect 126 383 186 437
rect 126 349 139 383
rect 173 349 186 383
rect 126 297 186 349
rect 222 478 282 497
rect 222 444 235 478
rect 269 444 282 478
rect 222 410 282 444
rect 222 376 235 410
rect 269 376 282 410
rect 222 297 282 376
rect 318 471 378 497
rect 318 437 331 471
rect 365 437 378 471
rect 318 383 378 437
rect 318 349 331 383
rect 365 349 378 383
rect 318 297 378 349
rect 414 478 474 497
rect 414 444 427 478
rect 461 444 474 478
rect 414 410 474 444
rect 414 376 427 410
rect 461 376 474 410
rect 414 297 474 376
rect 510 471 570 497
rect 510 437 523 471
rect 557 437 570 471
rect 510 383 570 437
rect 510 349 523 383
rect 557 349 570 383
rect 510 297 570 349
rect 606 478 677 497
rect 606 444 619 478
rect 653 444 677 478
rect 606 410 677 444
rect 606 376 619 410
rect 653 376 677 410
rect 606 297 677 376
<< ndiffc >>
rect 139 61 173 95
rect 235 72 269 106
rect 331 61 365 95
rect 427 72 461 106
rect 523 61 557 95
<< pdiffc >>
rect 43 444 77 478
rect 43 376 77 410
rect 139 437 173 471
rect 139 349 173 383
rect 235 444 269 478
rect 235 376 269 410
rect 331 437 365 471
rect 331 349 365 383
rect 427 444 461 478
rect 427 376 461 410
rect 523 437 557 471
rect 523 349 557 383
rect 619 444 653 478
rect 619 376 653 410
<< poly >>
rect 90 497 126 523
rect 186 497 222 523
rect 282 497 318 523
rect 378 497 414 523
rect 474 497 510 523
rect 570 497 606 523
rect 90 282 126 297
rect 186 282 222 297
rect 282 282 318 297
rect 378 282 414 297
rect 474 282 510 297
rect 570 282 606 297
rect 88 259 128 282
rect 184 259 224 282
rect 280 259 320 282
rect 376 259 416 282
rect 472 259 512 282
rect 568 259 608 282
rect 88 249 608 259
rect 88 215 115 249
rect 149 215 193 249
rect 227 215 271 249
rect 305 215 349 249
rect 383 215 427 249
rect 461 215 495 249
rect 529 215 608 249
rect 88 205 608 215
rect 184 131 214 205
rect 280 131 310 205
rect 376 131 406 205
rect 472 131 502 205
rect 184 21 214 47
rect 280 21 310 47
rect 376 21 406 47
rect 472 21 502 47
<< polycont >>
rect 115 215 149 249
rect 193 215 227 249
rect 271 215 305 249
rect 349 215 383 249
rect 427 215 461 249
rect 495 215 529 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 17 478 86 527
rect 17 444 43 478
rect 77 444 86 478
rect 17 410 86 444
rect 17 376 43 410
rect 77 376 86 410
rect 17 360 86 376
rect 131 471 182 487
rect 131 437 139 471
rect 173 437 182 471
rect 131 383 182 437
rect 131 349 139 383
rect 173 349 182 383
rect 226 478 278 527
rect 226 444 235 478
rect 269 444 278 478
rect 226 410 278 444
rect 226 376 235 410
rect 269 376 278 410
rect 226 360 278 376
rect 323 471 374 487
rect 323 437 331 471
rect 365 437 374 471
rect 323 383 374 437
rect 131 326 182 349
rect 323 349 331 383
rect 365 349 374 383
rect 418 478 470 527
rect 418 444 427 478
rect 461 444 470 478
rect 418 410 470 444
rect 418 376 427 410
rect 461 376 470 410
rect 418 360 470 376
rect 514 471 566 487
rect 514 437 523 471
rect 557 437 566 471
rect 514 383 566 437
rect 323 326 374 349
rect 514 349 523 383
rect 557 349 566 383
rect 610 478 687 527
rect 610 444 619 478
rect 653 444 687 478
rect 610 410 687 444
rect 610 376 619 410
rect 653 376 687 410
rect 610 360 687 376
rect 514 326 566 349
rect 21 292 714 326
rect 21 179 55 292
rect 89 249 582 258
rect 89 215 115 249
rect 149 215 193 249
rect 227 215 271 249
rect 305 215 349 249
rect 383 215 427 249
rect 461 215 495 249
rect 529 215 582 249
rect 89 213 582 215
rect 654 179 714 292
rect 21 145 714 179
rect 113 95 182 111
rect 113 61 139 95
rect 173 61 182 95
rect 113 17 182 61
rect 226 106 278 145
rect 226 72 235 106
rect 269 72 278 106
rect 226 56 278 72
rect 322 95 374 111
rect 322 61 331 95
rect 365 61 374 95
rect 322 17 374 61
rect 418 106 469 145
rect 418 72 427 106
rect 461 72 469 106
rect 418 56 469 72
rect 513 95 573 111
rect 513 61 523 95
rect 557 61 573 95
rect 513 17 573 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel corelocali s 230 238 230 238 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 322 238 322 238 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 668 153 702 187 0 FreeSans 400 0 0 0 Y
port 6 nsew
flabel corelocali s 131 221 165 255 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 668 289 702 323 0 FreeSans 400 0 0 0 Y
port 6 nsew
flabel corelocali s 506 238 506 238 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 414 238 414 238 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 668 221 702 255 0 FreeSans 400 0 0 0 Y
port 6 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew
rlabel comment s 0 0 0 0 4 clkinv_4
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1808132
string GDS_START 1801974
<< end >>
