magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 2246 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 94 47 124 177
rect 188 47 218 177
rect 282 47 312 177
rect 386 47 416 177
rect 470 47 500 177
rect 564 47 594 177
rect 658 47 688 177
rect 762 47 792 177
rect 950 47 980 177
rect 1044 47 1074 177
rect 1138 47 1168 177
rect 1242 47 1272 177
rect 1326 47 1356 177
rect 1420 47 1450 177
rect 1514 47 1544 177
rect 1618 47 1648 177
rect 1806 47 1836 177
rect 1900 47 1930 177
rect 1994 47 2024 177
rect 2098 47 2128 177
<< pmoshvt >>
rect 96 297 132 497
rect 190 297 226 497
rect 284 297 320 497
rect 378 297 414 497
rect 472 297 508 497
rect 566 297 602 497
rect 660 297 696 497
rect 754 297 790 497
rect 952 297 988 497
rect 1046 297 1082 497
rect 1140 297 1176 497
rect 1234 297 1270 497
rect 1328 297 1364 497
rect 1422 297 1458 497
rect 1516 297 1552 497
rect 1610 297 1646 497
rect 1808 297 1844 497
rect 1902 297 1938 497
rect 1996 297 2032 497
rect 2090 297 2126 497
<< ndiff >>
rect 38 95 94 177
rect 38 61 50 95
rect 84 61 94 95
rect 38 47 94 61
rect 124 163 188 177
rect 124 129 144 163
rect 178 129 188 163
rect 124 47 188 129
rect 218 95 282 177
rect 218 61 238 95
rect 272 61 282 95
rect 218 47 282 61
rect 312 163 386 177
rect 312 129 332 163
rect 366 129 386 163
rect 312 47 386 129
rect 416 163 470 177
rect 416 129 426 163
rect 460 129 470 163
rect 416 95 470 129
rect 416 61 426 95
rect 460 61 470 95
rect 416 47 470 61
rect 500 95 564 177
rect 500 61 520 95
rect 554 61 564 95
rect 500 47 564 61
rect 594 163 658 177
rect 594 129 614 163
rect 648 129 658 163
rect 594 95 658 129
rect 594 61 614 95
rect 648 61 658 95
rect 594 47 658 61
rect 688 95 762 177
rect 688 61 708 95
rect 742 61 762 95
rect 688 47 762 61
rect 792 163 844 177
rect 792 129 802 163
rect 836 129 844 163
rect 792 95 844 129
rect 792 61 802 95
rect 836 61 844 95
rect 792 47 844 61
rect 898 163 950 177
rect 898 129 906 163
rect 940 129 950 163
rect 898 95 950 129
rect 898 61 906 95
rect 940 61 950 95
rect 898 47 950 61
rect 980 163 1044 177
rect 980 129 1000 163
rect 1034 129 1044 163
rect 980 95 1044 129
rect 980 61 1000 95
rect 1034 61 1044 95
rect 980 47 1044 61
rect 1074 95 1138 177
rect 1074 61 1094 95
rect 1128 61 1138 95
rect 1074 47 1138 61
rect 1168 163 1242 177
rect 1168 129 1188 163
rect 1222 129 1242 163
rect 1168 95 1242 129
rect 1168 61 1188 95
rect 1222 61 1242 95
rect 1168 47 1242 61
rect 1272 95 1326 177
rect 1272 61 1282 95
rect 1316 61 1326 95
rect 1272 47 1326 61
rect 1356 163 1420 177
rect 1356 129 1376 163
rect 1410 129 1420 163
rect 1356 95 1420 129
rect 1356 61 1376 95
rect 1410 61 1420 95
rect 1356 47 1420 61
rect 1450 95 1514 177
rect 1450 61 1470 95
rect 1504 61 1514 95
rect 1450 47 1514 61
rect 1544 163 1618 177
rect 1544 129 1564 163
rect 1598 129 1618 163
rect 1544 95 1618 129
rect 1544 61 1564 95
rect 1598 61 1618 95
rect 1544 47 1618 61
rect 1648 95 1700 177
rect 1648 61 1658 95
rect 1692 61 1700 95
rect 1648 47 1700 61
rect 1754 163 1806 177
rect 1754 129 1762 163
rect 1796 129 1806 163
rect 1754 95 1806 129
rect 1754 61 1762 95
rect 1796 61 1806 95
rect 1754 47 1806 61
rect 1836 165 1900 177
rect 1836 131 1856 165
rect 1890 131 1900 165
rect 1836 47 1900 131
rect 1930 95 1994 177
rect 1930 61 1950 95
rect 1984 61 1994 95
rect 1930 47 1994 61
rect 2024 165 2098 177
rect 2024 131 2044 165
rect 2078 131 2098 165
rect 2024 47 2098 131
rect 2128 95 2180 177
rect 2128 61 2138 95
rect 2172 61 2180 95
rect 2128 47 2180 61
<< pdiff >>
rect 38 477 96 497
rect 38 443 50 477
rect 84 443 96 477
rect 38 409 96 443
rect 38 375 50 409
rect 84 375 96 409
rect 38 341 96 375
rect 38 307 50 341
rect 84 307 96 341
rect 38 297 96 307
rect 132 485 190 497
rect 132 451 144 485
rect 178 451 190 485
rect 132 417 190 451
rect 132 383 144 417
rect 178 383 190 417
rect 132 297 190 383
rect 226 477 284 497
rect 226 443 238 477
rect 272 443 284 477
rect 226 409 284 443
rect 226 375 238 409
rect 272 375 284 409
rect 226 341 284 375
rect 226 307 238 341
rect 272 307 284 341
rect 226 297 284 307
rect 320 485 378 497
rect 320 451 332 485
rect 366 451 378 485
rect 320 297 378 451
rect 414 477 472 497
rect 414 443 426 477
rect 460 443 472 477
rect 414 409 472 443
rect 414 375 426 409
rect 460 375 472 409
rect 414 297 472 375
rect 508 485 566 497
rect 508 451 520 485
rect 554 451 566 485
rect 508 297 566 451
rect 602 477 660 497
rect 602 443 614 477
rect 648 443 660 477
rect 602 409 660 443
rect 602 375 614 409
rect 648 375 660 409
rect 602 297 660 375
rect 696 485 754 497
rect 696 451 708 485
rect 742 451 754 485
rect 696 297 754 451
rect 790 477 844 497
rect 790 443 802 477
rect 836 443 844 477
rect 790 409 844 443
rect 790 375 802 409
rect 836 375 844 409
rect 790 297 844 375
rect 898 477 952 497
rect 898 443 906 477
rect 940 443 952 477
rect 898 409 952 443
rect 898 375 906 409
rect 940 375 952 409
rect 898 297 952 375
rect 988 485 1046 497
rect 988 451 1000 485
rect 1034 451 1046 485
rect 988 297 1046 451
rect 1082 477 1140 497
rect 1082 443 1094 477
rect 1128 443 1140 477
rect 1082 409 1140 443
rect 1082 375 1094 409
rect 1128 375 1140 409
rect 1082 297 1140 375
rect 1176 485 1234 497
rect 1176 451 1188 485
rect 1222 451 1234 485
rect 1176 297 1234 451
rect 1270 477 1328 497
rect 1270 443 1282 477
rect 1316 443 1328 477
rect 1270 409 1328 443
rect 1270 375 1282 409
rect 1316 375 1328 409
rect 1270 297 1328 375
rect 1364 409 1422 497
rect 1364 375 1376 409
rect 1410 375 1422 409
rect 1364 297 1422 375
rect 1458 477 1516 497
rect 1458 443 1470 477
rect 1504 443 1516 477
rect 1458 297 1516 443
rect 1552 409 1610 497
rect 1552 375 1564 409
rect 1598 375 1610 409
rect 1552 297 1610 375
rect 1646 477 1700 497
rect 1646 443 1658 477
rect 1692 443 1700 477
rect 1646 297 1700 443
rect 1754 485 1808 497
rect 1754 451 1762 485
rect 1796 451 1808 485
rect 1754 417 1808 451
rect 1754 383 1762 417
rect 1796 383 1808 417
rect 1754 349 1808 383
rect 1754 315 1762 349
rect 1796 315 1808 349
rect 1754 297 1808 315
rect 1844 485 1902 497
rect 1844 451 1856 485
rect 1890 451 1902 485
rect 1844 417 1902 451
rect 1844 383 1856 417
rect 1890 383 1902 417
rect 1844 297 1902 383
rect 1938 477 1996 497
rect 1938 443 1950 477
rect 1984 443 1996 477
rect 1938 409 1996 443
rect 1938 375 1950 409
rect 1984 375 1996 409
rect 1938 341 1996 375
rect 1938 307 1950 341
rect 1984 307 1996 341
rect 1938 297 1996 307
rect 2032 485 2090 497
rect 2032 451 2044 485
rect 2078 451 2090 485
rect 2032 417 2090 451
rect 2032 383 2044 417
rect 2078 383 2090 417
rect 2032 297 2090 383
rect 2126 485 2180 497
rect 2126 451 2138 485
rect 2172 451 2180 485
rect 2126 417 2180 451
rect 2126 383 2138 417
rect 2172 383 2180 417
rect 2126 349 2180 383
rect 2126 315 2138 349
rect 2172 315 2180 349
rect 2126 297 2180 315
<< ndiffc >>
rect 50 61 84 95
rect 144 129 178 163
rect 238 61 272 95
rect 332 129 366 163
rect 426 129 460 163
rect 426 61 460 95
rect 520 61 554 95
rect 614 129 648 163
rect 614 61 648 95
rect 708 61 742 95
rect 802 129 836 163
rect 802 61 836 95
rect 906 129 940 163
rect 906 61 940 95
rect 1000 129 1034 163
rect 1000 61 1034 95
rect 1094 61 1128 95
rect 1188 129 1222 163
rect 1188 61 1222 95
rect 1282 61 1316 95
rect 1376 129 1410 163
rect 1376 61 1410 95
rect 1470 61 1504 95
rect 1564 129 1598 163
rect 1564 61 1598 95
rect 1658 61 1692 95
rect 1762 129 1796 163
rect 1762 61 1796 95
rect 1856 131 1890 165
rect 1950 61 1984 95
rect 2044 131 2078 165
rect 2138 61 2172 95
<< pdiffc >>
rect 50 443 84 477
rect 50 375 84 409
rect 50 307 84 341
rect 144 451 178 485
rect 144 383 178 417
rect 238 443 272 477
rect 238 375 272 409
rect 238 307 272 341
rect 332 451 366 485
rect 426 443 460 477
rect 426 375 460 409
rect 520 451 554 485
rect 614 443 648 477
rect 614 375 648 409
rect 708 451 742 485
rect 802 443 836 477
rect 802 375 836 409
rect 906 443 940 477
rect 906 375 940 409
rect 1000 451 1034 485
rect 1094 443 1128 477
rect 1094 375 1128 409
rect 1188 451 1222 485
rect 1282 443 1316 477
rect 1282 375 1316 409
rect 1376 375 1410 409
rect 1470 443 1504 477
rect 1564 375 1598 409
rect 1658 443 1692 477
rect 1762 451 1796 485
rect 1762 383 1796 417
rect 1762 315 1796 349
rect 1856 451 1890 485
rect 1856 383 1890 417
rect 1950 443 1984 477
rect 1950 375 1984 409
rect 1950 307 1984 341
rect 2044 451 2078 485
rect 2044 383 2078 417
rect 2138 451 2172 485
rect 2138 383 2172 417
rect 2138 315 2172 349
<< poly >>
rect 96 497 132 523
rect 190 497 226 523
rect 284 497 320 523
rect 378 497 414 523
rect 472 497 508 523
rect 566 497 602 523
rect 660 497 696 523
rect 754 497 790 523
rect 952 497 988 523
rect 1046 497 1082 523
rect 1140 497 1176 523
rect 1234 497 1270 523
rect 1328 497 1364 523
rect 1422 497 1458 523
rect 1516 497 1552 523
rect 1610 497 1646 523
rect 1808 497 1844 523
rect 1902 497 1938 523
rect 1996 497 2032 523
rect 2090 497 2126 523
rect 96 282 132 297
rect 190 282 226 297
rect 284 282 320 297
rect 378 282 414 297
rect 472 282 508 297
rect 566 282 602 297
rect 660 282 696 297
rect 754 282 790 297
rect 952 282 988 297
rect 1046 282 1082 297
rect 1140 282 1176 297
rect 1234 282 1270 297
rect 1328 282 1364 297
rect 1422 282 1458 297
rect 1516 282 1552 297
rect 1610 282 1646 297
rect 1808 282 1844 297
rect 1902 282 1938 297
rect 1996 282 2032 297
rect 2090 282 2126 297
rect 94 265 134 282
rect 188 265 228 282
rect 282 265 322 282
rect 376 265 416 282
rect 94 249 416 265
rect 94 215 114 249
rect 148 215 192 249
rect 226 215 270 249
rect 304 215 348 249
rect 382 215 416 249
rect 94 199 416 215
rect 94 177 124 199
rect 188 177 218 199
rect 282 177 312 199
rect 386 177 416 199
rect 470 265 510 282
rect 564 265 604 282
rect 658 265 698 282
rect 752 265 792 282
rect 470 249 792 265
rect 470 215 493 249
rect 527 215 571 249
rect 605 215 649 249
rect 683 215 727 249
rect 761 215 792 249
rect 470 199 792 215
rect 470 177 500 199
rect 564 177 594 199
rect 658 177 688 199
rect 762 177 792 199
rect 950 265 990 282
rect 1044 265 1084 282
rect 1138 265 1178 282
rect 1232 265 1272 282
rect 950 249 1272 265
rect 950 215 970 249
rect 1004 215 1048 249
rect 1082 215 1126 249
rect 1160 215 1272 249
rect 950 199 1272 215
rect 950 177 980 199
rect 1044 177 1074 199
rect 1138 177 1168 199
rect 1242 177 1272 199
rect 1326 265 1366 282
rect 1420 265 1460 282
rect 1514 265 1554 282
rect 1608 265 1648 282
rect 1326 249 1648 265
rect 1326 215 1349 249
rect 1383 215 1427 249
rect 1461 215 1505 249
rect 1539 215 1583 249
rect 1617 215 1648 249
rect 1326 199 1648 215
rect 1326 177 1356 199
rect 1420 177 1450 199
rect 1514 177 1544 199
rect 1618 177 1648 199
rect 1806 265 1846 282
rect 1900 265 1940 282
rect 1994 265 2034 282
rect 2088 265 2128 282
rect 1806 249 2128 265
rect 1806 215 1823 249
rect 1857 215 1901 249
rect 1935 215 1979 249
rect 2013 215 2057 249
rect 2091 215 2128 249
rect 1806 199 2128 215
rect 1806 177 1836 199
rect 1900 177 1930 199
rect 1994 177 2024 199
rect 2098 177 2128 199
rect 94 21 124 47
rect 188 21 218 47
rect 282 21 312 47
rect 386 21 416 47
rect 470 21 500 47
rect 564 21 594 47
rect 658 21 688 47
rect 762 21 792 47
rect 950 21 980 47
rect 1044 21 1074 47
rect 1138 21 1168 47
rect 1242 21 1272 47
rect 1326 21 1356 47
rect 1420 21 1450 47
rect 1514 21 1544 47
rect 1618 21 1648 47
rect 1806 21 1836 47
rect 1900 21 1930 47
rect 1994 21 2024 47
rect 2098 21 2128 47
<< polycont >>
rect 114 215 148 249
rect 192 215 226 249
rect 270 215 304 249
rect 348 215 382 249
rect 493 215 527 249
rect 571 215 605 249
rect 649 215 683 249
rect 727 215 761 249
rect 970 215 1004 249
rect 1048 215 1082 249
rect 1126 215 1160 249
rect 1349 215 1383 249
rect 1427 215 1461 249
rect 1505 215 1539 249
rect 1583 215 1617 249
rect 1823 215 1857 249
rect 1901 215 1935 249
rect 1979 215 2013 249
rect 2057 215 2091 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 17 477 92 493
rect 17 443 50 477
rect 84 443 92 477
rect 17 409 92 443
rect 17 375 50 409
rect 84 375 92 409
rect 17 341 92 375
rect 136 485 186 527
rect 136 451 144 485
rect 178 451 186 485
rect 136 417 186 451
rect 136 383 144 417
rect 178 383 186 417
rect 136 367 186 383
rect 230 477 280 493
rect 230 443 238 477
rect 272 443 280 477
rect 230 409 280 443
rect 324 485 374 527
rect 324 451 332 485
rect 366 451 374 485
rect 324 435 374 451
rect 418 477 468 493
rect 418 443 426 477
rect 460 443 468 477
rect 230 375 238 409
rect 272 401 280 409
rect 418 409 468 443
rect 512 485 562 527
rect 512 451 520 485
rect 554 451 562 485
rect 512 435 562 451
rect 606 477 656 493
rect 606 443 614 477
rect 648 443 656 477
rect 418 401 426 409
rect 272 375 426 401
rect 460 401 468 409
rect 606 409 656 443
rect 700 485 750 527
rect 700 451 708 485
rect 742 451 750 485
rect 700 435 750 451
rect 794 477 844 493
rect 794 443 802 477
rect 836 443 844 477
rect 606 401 614 409
rect 460 375 614 401
rect 648 401 656 409
rect 794 409 844 443
rect 794 401 802 409
rect 648 375 802 401
rect 836 375 844 409
rect 17 307 50 341
rect 84 323 92 341
rect 230 357 844 375
rect 885 477 948 493
rect 885 443 906 477
rect 940 443 948 477
rect 885 409 948 443
rect 992 485 1042 527
rect 992 451 1000 485
rect 1034 451 1042 485
rect 992 435 1042 451
rect 1086 477 1136 493
rect 1086 443 1094 477
rect 1128 443 1136 477
rect 885 375 906 409
rect 940 401 948 409
rect 1086 409 1136 443
rect 1180 485 1230 527
rect 1180 451 1188 485
rect 1222 451 1230 485
rect 1180 435 1230 451
rect 1274 477 1708 493
rect 1274 443 1282 477
rect 1316 443 1470 477
rect 1504 443 1658 477
rect 1692 443 1708 477
rect 1746 485 1812 493
rect 1746 451 1762 485
rect 1796 451 1812 485
rect 1086 401 1094 409
rect 940 375 1094 401
rect 1128 401 1136 409
rect 1274 409 1316 443
rect 1746 417 1812 451
rect 1746 409 1762 417
rect 1274 401 1282 409
rect 1128 375 1282 401
rect 885 357 1316 375
rect 1350 375 1376 409
rect 1410 375 1564 409
rect 1598 383 1762 409
rect 1796 383 1812 417
rect 1598 375 1812 383
rect 1350 357 1812 375
rect 1848 485 1898 527
rect 1848 451 1856 485
rect 1890 451 1898 485
rect 1848 417 1898 451
rect 1848 383 1856 417
rect 1890 383 1898 417
rect 1848 367 1898 383
rect 1942 477 1992 493
rect 1942 443 1950 477
rect 1984 443 1992 477
rect 1942 409 1992 443
rect 1942 375 1950 409
rect 1984 375 1992 409
rect 230 341 280 357
rect 230 323 238 341
rect 84 307 233 323
rect 272 307 280 341
rect 1746 349 1812 357
rect 17 289 233 307
rect 267 289 280 307
rect 367 289 1254 323
rect 1298 289 1345 323
rect 1379 289 1712 323
rect 1746 315 1762 349
rect 1796 333 1812 349
rect 1942 341 1992 375
rect 2036 485 2086 527
rect 2036 451 2044 485
rect 2078 451 2086 485
rect 2036 417 2086 451
rect 2036 383 2044 417
rect 2078 383 2086 417
rect 2036 367 2086 383
rect 2122 485 2188 493
rect 2122 451 2138 485
rect 2172 451 2188 485
rect 2122 417 2188 451
rect 2122 383 2138 417
rect 2172 383 2188 417
rect 1942 333 1950 341
rect 1796 315 1950 333
rect 1746 307 1950 315
rect 1984 333 1992 341
rect 2122 349 2188 383
rect 2122 333 2138 349
rect 1984 315 2138 333
rect 2172 315 2188 349
rect 1984 307 2188 315
rect 1746 289 2188 307
rect 17 181 64 289
rect 367 255 401 289
rect 1220 255 1254 289
rect 1678 255 1712 289
rect 98 249 401 255
rect 98 215 114 249
rect 148 215 192 249
rect 226 215 270 249
rect 304 215 348 249
rect 382 215 401 249
rect 475 249 1186 255
rect 475 215 493 249
rect 527 215 571 249
rect 605 215 649 249
rect 683 215 727 249
rect 761 215 970 249
rect 1004 215 1048 249
rect 1082 215 1126 249
rect 1160 215 1186 249
rect 1220 249 1634 255
rect 1220 215 1349 249
rect 1383 215 1427 249
rect 1461 215 1505 249
rect 1539 215 1583 249
rect 1617 215 1634 249
rect 1678 249 2107 255
rect 1678 215 1823 249
rect 1857 215 1901 249
rect 1935 215 1979 249
rect 2013 215 2057 249
rect 2091 215 2107 249
rect 2141 181 2188 289
rect 17 163 382 181
rect 17 129 144 163
rect 178 129 332 163
rect 366 129 382 163
rect 426 163 852 181
rect 460 145 614 163
rect 460 129 476 145
rect 426 95 476 129
rect 588 129 614 145
rect 648 145 802 163
rect 648 129 664 145
rect 34 61 50 95
rect 84 61 238 95
rect 272 61 426 95
rect 460 61 476 95
rect 34 51 476 61
rect 520 95 554 111
rect 520 17 554 61
rect 588 95 664 129
rect 776 129 802 145
rect 836 129 852 163
rect 588 61 614 95
rect 648 61 664 95
rect 588 51 664 61
rect 708 95 742 111
rect 708 17 742 61
rect 776 95 852 129
rect 776 61 802 95
rect 836 61 852 95
rect 776 51 852 61
rect 886 163 940 181
rect 886 129 906 163
rect 886 95 940 129
rect 886 61 906 95
rect 886 17 940 61
rect 974 163 1796 181
rect 974 129 1000 163
rect 1034 145 1188 163
rect 1034 129 1050 145
rect 974 95 1050 129
rect 1162 129 1188 145
rect 1222 145 1376 163
rect 1222 129 1238 145
rect 974 61 1000 95
rect 1034 61 1050 95
rect 974 51 1050 61
rect 1094 95 1128 111
rect 1094 17 1128 61
rect 1162 95 1238 129
rect 1350 129 1376 145
rect 1410 145 1564 163
rect 1410 129 1426 145
rect 1162 61 1188 95
rect 1222 61 1238 95
rect 1162 51 1238 61
rect 1282 95 1316 111
rect 1282 17 1316 61
rect 1350 95 1426 129
rect 1538 129 1564 145
rect 1598 147 1762 163
rect 1598 145 1634 147
rect 1598 129 1614 145
rect 1350 61 1376 95
rect 1410 61 1426 95
rect 1350 51 1426 61
rect 1470 95 1504 111
rect 1470 17 1504 61
rect 1538 95 1614 129
rect 1746 129 1762 147
rect 1830 165 2188 181
rect 1830 131 1856 165
rect 1890 131 2044 165
rect 2078 131 2188 165
rect 1538 61 1564 95
rect 1598 61 1614 95
rect 1538 51 1614 61
rect 1658 95 1692 111
rect 1746 95 1796 129
rect 1746 61 1762 95
rect 1796 61 1950 95
rect 1984 61 2138 95
rect 2172 61 2188 95
rect 1658 17 1692 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 233 307 238 323
rect 238 307 267 323
rect 233 289 267 307
rect 1345 289 1379 323
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
<< metal1 >>
rect 0 561 2208 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 0 496 2208 527
rect 211 323 279 329
rect 211 289 233 323
rect 267 320 279 323
rect 1331 323 1401 329
rect 1331 320 1345 323
rect 267 292 1345 320
rect 267 289 279 292
rect 211 283 279 289
rect 1331 289 1345 292
rect 1379 289 1401 323
rect 1331 283 1401 289
rect 0 17 2208 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
rect 0 -48 2208 -17
<< labels >>
flabel corelocali s 2145 221 2179 255 0 FreeSans 400 0 0 0 Y
port 7 nsew
flabel corelocali s 214 221 248 255 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel corelocali s 857 221 891 255 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew
rlabel comment s 0 0 0 0 4 xnor2_4
<< properties >>
string FIXED_BBOX 0 0 2208 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 710770
string GDS_START 695802
<< end >>
