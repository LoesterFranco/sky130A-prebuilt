magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 644 561
rect 103 425 175 527
rect 17 199 66 323
rect 291 379 357 527
rect 103 17 175 97
rect 282 17 354 97
rect 470 119 536 425
rect 570 153 627 323
rect 0 -17 644 17
<< obsli1 >>
rect 17 391 69 493
rect 17 357 175 391
rect 100 265 175 357
rect 209 345 257 493
rect 397 459 627 493
rect 397 345 431 459
rect 209 311 431 345
rect 100 199 436 265
rect 100 165 175 199
rect 17 131 175 165
rect 209 131 436 165
rect 17 51 69 131
rect 209 51 248 131
rect 388 85 436 131
rect 570 357 627 459
rect 570 85 627 119
rect 388 51 627 85
<< metal1 >>
rect 0 496 644 592
rect 0 -48 644 48
<< labels >>
rlabel locali s 570 153 627 323 6 A
port 1 nsew signal input
rlabel locali s 17 199 66 323 6 TE
port 2 nsew signal input
rlabel locali s 470 119 536 425 6 Z
port 3 nsew signal output
rlabel locali s 282 17 354 97 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 103 17 175 97 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 644 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 644 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 291 379 357 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 103 425 175 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 644 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 644 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2918784
string GDS_START 2912596
<< end >>
