magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 391 405 764 421
rect 899 405 1696 421
rect 391 371 1696 405
rect 203 303 806 337
rect 203 266 312 303
rect 80 215 312 266
rect 371 215 706 269
rect 740 199 806 303
rect 942 303 1560 337
rect 942 282 1105 303
rect 840 199 1105 282
rect 1194 215 1428 269
rect 1516 199 1560 303
rect 1596 268 1696 371
rect 1596 165 1632 268
rect 1453 131 1632 165
rect 1453 90 1497 131
rect 1166 54 1497 90
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 18 333 77 527
rect 201 455 277 527
rect 321 455 757 493
rect 121 421 165 438
rect 321 421 357 455
rect 803 439 857 527
rect 977 455 1053 527
rect 1166 455 1242 527
rect 1354 455 1431 527
rect 1631 455 1697 527
rect 121 387 357 421
rect 121 372 165 387
rect 31 159 696 181
rect 31 125 847 159
rect 881 127 1374 163
rect 31 107 71 125
rect 105 17 181 89
rect 225 85 268 125
rect 801 91 847 125
rect 307 17 373 91
rect 489 17 565 89
rect 681 17 757 89
rect 801 51 1094 91
rect 1664 96 1698 119
rect 1546 62 1698 96
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
<< metal1 >>
rect 0 561 1748 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 0 496 1748 527
rect 0 17 1748 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
rect 0 -48 1748 -17
<< obsm1 >>
rect 222 116 280 125
rect 1652 116 1710 125
rect 222 88 1710 116
rect 222 79 280 88
rect 1652 79 1710 88
<< labels >>
rlabel locali s 740 199 806 303 6 A1
port 1 nsew signal input
rlabel locali s 203 303 806 337 6 A1
port 1 nsew signal input
rlabel locali s 203 266 312 303 6 A1
port 1 nsew signal input
rlabel locali s 80 215 312 266 6 A1
port 1 nsew signal input
rlabel locali s 371 215 706 269 6 A2
port 2 nsew signal input
rlabel locali s 1516 199 1560 303 6 B1
port 3 nsew signal input
rlabel locali s 942 303 1560 337 6 B1
port 3 nsew signal input
rlabel locali s 942 282 1105 303 6 B1
port 3 nsew signal input
rlabel locali s 840 199 1105 282 6 B1
port 3 nsew signal input
rlabel locali s 1194 215 1428 269 6 C1
port 4 nsew signal input
rlabel locali s 1596 268 1696 371 6 Y
port 5 nsew signal output
rlabel locali s 1596 165 1632 268 6 Y
port 5 nsew signal output
rlabel locali s 1453 131 1632 165 6 Y
port 5 nsew signal output
rlabel locali s 1453 90 1497 131 6 Y
port 5 nsew signal output
rlabel locali s 1166 54 1497 90 6 Y
port 5 nsew signal output
rlabel locali s 899 405 1696 421 6 Y
port 5 nsew signal output
rlabel locali s 391 405 764 421 6 Y
port 5 nsew signal output
rlabel locali s 391 371 1696 405 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -48 1748 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 1748 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1748 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 979962
string GDS_START 969190
<< end >>
