magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1196 561
rect 114 427 164 527
rect 282 427 332 527
rect 562 427 612 527
rect 925 427 975 527
rect 745 393 787 425
rect 1009 393 1059 425
rect 745 359 1059 393
rect 1093 359 1179 527
rect 1009 325 1059 359
rect 158 289 620 323
rect 158 257 192 289
rect 97 215 192 257
rect 586 257 620 289
rect 251 215 541 255
rect 586 215 791 257
rect 1009 283 1179 325
rect 290 17 324 111
rect 486 17 520 181
rect 654 17 688 111
rect 829 17 863 111
rect 1101 95 1179 283
rect 917 61 1179 95
rect 0 -17 1196 17
<< obsli1 >>
rect 17 393 80 493
rect 198 393 248 493
rect 366 393 416 493
rect 478 459 528 493
rect 478 425 493 459
rect 527 425 528 459
rect 646 459 871 493
rect 646 425 677 459
rect 821 427 871 459
rect 17 391 416 393
rect 17 357 696 391
rect 17 179 63 357
rect 662 325 696 357
rect 662 291 961 325
rect 927 249 961 291
rect 927 215 1059 249
rect 17 129 172 179
rect 206 145 424 181
rect 206 95 256 145
rect 21 51 256 95
rect 358 51 424 145
rect 554 145 1067 181
rect 554 51 620 145
rect 722 51 795 145
rect 1001 129 1067 145
<< obsli1c >>
rect 493 425 527 459
rect 677 425 711 459
<< metal1 >>
rect 0 496 1196 592
rect 0 -48 1196 48
<< obsm1 >>
rect 481 459 539 465
rect 481 425 493 459
rect 527 456 539 459
rect 665 459 723 465
rect 665 456 677 459
rect 527 428 677 456
rect 527 425 539 428
rect 481 419 539 425
rect 665 425 677 428
rect 711 425 723 459
rect 665 419 723 425
<< labels >>
rlabel locali s 251 215 541 255 6 A
port 1 nsew signal input
rlabel locali s 586 257 620 289 6 B
port 2 nsew signal input
rlabel locali s 586 215 791 257 6 B
port 2 nsew signal input
rlabel locali s 158 289 620 323 6 B
port 2 nsew signal input
rlabel locali s 158 257 192 289 6 B
port 2 nsew signal input
rlabel locali s 97 215 192 257 6 B
port 2 nsew signal input
rlabel locali s 1101 95 1179 283 6 Y
port 3 nsew signal output
rlabel locali s 1009 393 1059 425 6 Y
port 3 nsew signal output
rlabel locali s 1009 325 1059 359 6 Y
port 3 nsew signal output
rlabel locali s 1009 283 1179 325 6 Y
port 3 nsew signal output
rlabel locali s 917 61 1179 95 6 Y
port 3 nsew signal output
rlabel locali s 745 393 787 425 6 Y
port 3 nsew signal output
rlabel locali s 745 359 1059 393 6 Y
port 3 nsew signal output
rlabel locali s 829 17 863 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 654 17 688 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 486 17 520 181 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 290 17 324 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 1196 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1196 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 1093 359 1179 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 925 427 975 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 562 427 612 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 282 427 332 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 114 427 164 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 1196 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 1196 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 626992
string GDS_START 618312
<< end >>
