magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 1284 339 1318 493
rect 1472 339 1506 493
rect 1660 339 1725 493
rect 835 289 1725 339
rect 18 211 386 285
rect 430 211 801 285
rect 835 211 1318 255
rect 1352 177 1399 289
rect 1433 211 1717 255
rect 1352 129 1616 177
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 18 379 89 493
rect 133 413 167 527
rect 201 379 277 493
rect 321 413 355 527
rect 389 441 857 493
rect 389 379 465 441
rect 18 319 465 379
rect 509 353 543 407
rect 577 387 653 441
rect 906 407 1240 493
rect 697 373 1240 407
rect 697 353 801 373
rect 509 319 801 353
rect 1352 378 1428 527
rect 1540 378 1616 527
rect 18 143 1318 177
rect 18 51 89 143
rect 133 17 167 109
rect 201 51 277 143
rect 321 17 355 109
rect 389 51 465 143
rect 509 17 543 109
rect 577 51 653 143
rect 697 17 731 109
rect 765 51 841 143
rect 889 17 1028 109
rect 1072 79 1106 143
rect 1158 17 1232 109
rect 1284 95 1318 143
rect 1660 95 1717 177
rect 1284 51 1717 95
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
<< metal1 >>
rect 0 561 1748 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 0 496 1748 527
rect 0 17 1748 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
rect 0 -48 1748 -17
<< labels >>
rlabel locali s 18 211 386 285 6 A1
port 1 nsew signal input
rlabel locali s 430 211 801 285 6 A2
port 2 nsew signal input
rlabel locali s 835 211 1318 255 6 A3
port 3 nsew signal input
rlabel locali s 1433 211 1717 255 6 B1
port 4 nsew signal input
rlabel locali s 1660 339 1725 493 6 Y
port 5 nsew signal output
rlabel locali s 1472 339 1506 493 6 Y
port 5 nsew signal output
rlabel locali s 1352 177 1399 289 6 Y
port 5 nsew signal output
rlabel locali s 1352 129 1616 177 6 Y
port 5 nsew signal output
rlabel locali s 1284 339 1318 493 6 Y
port 5 nsew signal output
rlabel locali s 835 289 1725 339 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -48 1748 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 1748 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1748 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 574094
string GDS_START 559094
<< end >>
