magic
tech sky130A
magscale 1 2
timestamp 1604502705
<< nwell >>
rect -38 332 1478 704
<< pwell >>
rect 0 0 1440 49
<< scnmos >>
rect 89 112 119 222
rect 205 74 235 222
rect 420 98 450 246
rect 538 74 568 202
rect 616 74 646 202
rect 754 81 784 165
rect 832 81 862 165
rect 1030 74 1060 222
rect 1108 74 1138 222
rect 1226 74 1256 222
rect 1314 74 1344 222
<< pmoshvt >>
rect 86 392 116 560
rect 210 392 240 560
rect 412 392 442 560
rect 535 392 565 592
rect 619 392 649 592
rect 726 508 756 592
rect 863 508 893 592
rect 1024 368 1054 592
rect 1114 368 1144 592
rect 1224 368 1254 592
rect 1317 368 1347 592
<< ndiff >>
rect 347 234 420 246
rect 32 184 89 222
rect 32 150 44 184
rect 78 150 89 184
rect 32 112 89 150
rect 119 188 205 222
rect 119 154 146 188
rect 180 154 205 188
rect 119 120 205 154
rect 119 112 146 120
rect 134 86 146 112
rect 180 86 205 120
rect 134 74 205 86
rect 235 196 292 222
rect 235 162 246 196
rect 280 162 292 196
rect 235 120 292 162
rect 235 86 246 120
rect 280 86 292 120
rect 347 200 359 234
rect 393 200 420 234
rect 347 98 420 200
rect 450 202 500 246
rect 450 98 538 202
rect 235 74 292 86
rect 465 82 538 98
rect 465 48 477 82
rect 511 74 538 82
rect 568 74 616 202
rect 646 165 739 202
rect 973 210 1030 222
rect 973 176 985 210
rect 1019 176 1030 210
rect 646 153 754 165
rect 646 119 675 153
rect 709 119 754 153
rect 646 81 754 119
rect 784 81 832 165
rect 862 140 919 165
rect 862 106 873 140
rect 907 106 919 140
rect 862 81 919 106
rect 973 120 1030 176
rect 973 86 985 120
rect 1019 86 1030 120
rect 646 74 696 81
rect 511 48 523 74
rect 973 74 1030 86
rect 1060 74 1108 222
rect 1138 198 1226 222
rect 1138 164 1167 198
rect 1201 164 1226 198
rect 1138 120 1226 164
rect 1138 86 1167 120
rect 1201 86 1226 120
rect 1138 74 1226 86
rect 1256 210 1314 222
rect 1256 176 1267 210
rect 1301 176 1314 210
rect 1256 120 1314 176
rect 1256 86 1267 120
rect 1301 86 1314 120
rect 1256 74 1314 86
rect 1344 142 1413 222
rect 1344 108 1367 142
rect 1401 108 1413 142
rect 1344 74 1413 108
rect 465 36 523 48
<< pdiff >>
rect 134 606 192 618
rect 134 572 146 606
rect 180 572 192 606
rect 460 606 517 618
rect 134 560 192 572
rect 460 572 472 606
rect 506 592 517 606
rect 506 572 535 592
rect 460 560 535 572
rect 27 548 86 560
rect 27 514 39 548
rect 73 514 86 548
rect 27 440 86 514
rect 27 406 39 440
rect 73 406 86 440
rect 27 392 86 406
rect 116 392 210 560
rect 240 438 299 560
rect 240 404 253 438
rect 287 404 299 438
rect 240 392 299 404
rect 353 438 412 560
rect 353 404 365 438
rect 399 404 412 438
rect 353 392 412 404
rect 442 392 535 560
rect 565 392 619 592
rect 649 531 726 592
rect 649 497 662 531
rect 696 508 726 531
rect 756 508 863 592
rect 893 580 1024 592
rect 893 546 936 580
rect 970 546 1024 580
rect 893 508 1024 546
rect 696 497 708 508
rect 649 392 708 497
rect 971 368 1024 508
rect 1054 580 1114 592
rect 1054 546 1067 580
rect 1101 546 1114 580
rect 1054 497 1114 546
rect 1054 463 1067 497
rect 1101 463 1114 497
rect 1054 414 1114 463
rect 1054 380 1067 414
rect 1101 380 1114 414
rect 1054 368 1114 380
rect 1144 582 1224 592
rect 1144 548 1167 582
rect 1201 548 1224 582
rect 1144 514 1224 548
rect 1144 480 1167 514
rect 1201 480 1224 514
rect 1144 446 1224 480
rect 1144 412 1167 446
rect 1201 412 1224 446
rect 1144 368 1224 412
rect 1254 582 1317 592
rect 1254 548 1267 582
rect 1301 548 1317 582
rect 1254 514 1317 548
rect 1254 480 1267 514
rect 1301 480 1317 514
rect 1254 446 1317 480
rect 1254 412 1267 446
rect 1301 412 1317 446
rect 1254 368 1317 412
rect 1347 580 1413 592
rect 1347 546 1367 580
rect 1401 546 1413 580
rect 1347 478 1413 546
rect 1347 444 1367 478
rect 1401 444 1413 478
rect 1347 368 1413 444
<< ndiffc >>
rect 44 150 78 184
rect 146 154 180 188
rect 146 86 180 120
rect 246 162 280 196
rect 246 86 280 120
rect 359 200 393 234
rect 477 48 511 82
rect 985 176 1019 210
rect 675 119 709 153
rect 873 106 907 140
rect 985 86 1019 120
rect 1167 164 1201 198
rect 1167 86 1201 120
rect 1267 176 1301 210
rect 1267 86 1301 120
rect 1367 108 1401 142
<< pdiffc >>
rect 146 572 180 606
rect 472 572 506 606
rect 39 514 73 548
rect 39 406 73 440
rect 253 404 287 438
rect 365 404 399 438
rect 662 497 696 531
rect 936 546 970 580
rect 1067 546 1101 580
rect 1067 463 1101 497
rect 1067 380 1101 414
rect 1167 548 1201 582
rect 1167 480 1201 514
rect 1167 412 1201 446
rect 1267 548 1301 582
rect 1267 480 1301 514
rect 1267 412 1301 446
rect 1367 546 1401 580
rect 1367 444 1401 478
<< poly >>
rect 86 560 116 586
rect 210 560 240 586
rect 412 560 442 586
rect 535 592 565 618
rect 619 592 649 618
rect 726 592 756 618
rect 863 592 893 618
rect 1024 592 1054 618
rect 1114 592 1144 618
rect 1224 592 1254 618
rect 1317 592 1347 618
rect 726 493 756 508
rect 863 493 893 508
rect 723 476 759 493
rect 860 476 896 493
rect 723 460 812 476
rect 723 426 762 460
rect 796 426 812 460
rect 723 410 812 426
rect 860 460 926 476
rect 860 426 876 460
rect 910 426 926 460
rect 860 410 926 426
rect 86 377 116 392
rect 210 377 240 392
rect 412 377 442 392
rect 535 377 565 392
rect 619 377 649 392
rect 83 356 119 377
rect 44 340 119 356
rect 44 306 60 340
rect 94 306 119 340
rect 207 310 243 377
rect 409 350 445 377
rect 532 354 568 377
rect 312 334 445 350
rect 44 290 119 306
rect 89 222 119 290
rect 198 294 264 310
rect 198 260 214 294
rect 248 260 264 294
rect 312 300 328 334
rect 362 314 445 334
rect 502 338 568 354
rect 362 300 450 314
rect 312 284 450 300
rect 502 304 518 338
rect 552 304 568 338
rect 616 362 652 377
rect 616 332 782 362
rect 502 288 568 304
rect 752 318 782 332
rect 752 302 818 318
rect 198 244 264 260
rect 420 246 450 284
rect 205 222 235 244
rect 89 86 119 112
rect 538 202 568 288
rect 610 274 676 290
rect 610 240 626 274
rect 660 240 676 274
rect 752 268 768 302
rect 802 268 818 302
rect 752 252 818 268
rect 610 224 676 240
rect 616 202 646 224
rect 205 48 235 74
rect 420 72 450 98
rect 754 165 784 252
rect 860 210 890 410
rect 1024 353 1054 368
rect 1114 353 1144 368
rect 1224 353 1254 368
rect 1317 353 1347 368
rect 1021 336 1057 353
rect 932 320 1057 336
rect 932 286 948 320
rect 982 300 1057 320
rect 1111 310 1147 353
rect 1221 326 1257 353
rect 1314 326 1350 353
rect 1210 310 1350 326
rect 982 286 1060 300
rect 932 270 1060 286
rect 1030 222 1060 270
rect 1102 294 1168 310
rect 1102 260 1118 294
rect 1152 260 1168 294
rect 1210 276 1226 310
rect 1260 276 1294 310
rect 1328 296 1350 310
rect 1328 276 1344 296
rect 1210 260 1344 276
rect 1102 244 1168 260
rect 1108 222 1138 244
rect 1226 222 1256 260
rect 1314 222 1344 260
rect 832 180 890 210
rect 832 165 862 180
rect 538 48 568 74
rect 616 48 646 74
rect 754 55 784 81
rect 832 55 862 81
rect 1030 48 1060 74
rect 1108 48 1138 74
rect 1226 48 1256 74
rect 1314 48 1344 74
<< polycont >>
rect 762 426 796 460
rect 876 426 910 460
rect 60 306 94 340
rect 214 260 248 294
rect 328 300 362 334
rect 518 304 552 338
rect 626 240 660 274
rect 768 268 802 302
rect 948 286 982 320
rect 1118 260 1152 294
rect 1226 276 1260 310
rect 1294 276 1328 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 130 606 196 649
rect 130 572 146 606
rect 180 572 196 606
rect 23 548 89 564
rect 130 556 196 572
rect 456 606 522 649
rect 456 572 472 606
rect 506 572 522 606
rect 456 556 522 572
rect 578 581 812 615
rect 23 514 39 548
rect 73 522 89 548
rect 73 514 536 522
rect 23 488 536 514
rect 23 440 171 488
rect 23 406 39 440
rect 73 406 171 440
rect 23 390 171 406
rect 25 340 103 356
rect 25 306 60 340
rect 94 306 103 340
rect 25 290 103 306
rect 137 256 171 390
rect 237 438 325 454
rect 237 404 253 438
rect 287 404 325 438
rect 237 388 325 404
rect 365 438 446 454
rect 399 404 446 438
rect 365 388 446 404
rect 291 350 325 388
rect 291 334 378 350
rect 28 222 171 256
rect 205 294 257 310
rect 205 260 214 294
rect 248 260 257 294
rect 205 236 257 260
rect 291 300 328 334
rect 362 300 378 334
rect 291 284 378 300
rect 28 184 94 222
rect 291 202 325 284
rect 412 250 446 388
rect 502 354 536 488
rect 578 422 612 581
rect 646 531 712 547
rect 646 497 662 531
rect 696 497 712 531
rect 646 481 712 497
rect 578 388 644 422
rect 502 338 568 354
rect 502 304 518 338
rect 552 304 568 338
rect 502 288 568 304
rect 610 290 644 388
rect 678 386 712 481
rect 746 460 812 581
rect 890 580 1017 649
rect 890 546 936 580
rect 970 546 1017 580
rect 890 530 1017 546
rect 1051 580 1117 596
rect 1051 546 1067 580
rect 1101 546 1117 580
rect 1051 497 1117 546
rect 1051 476 1067 497
rect 746 426 762 460
rect 796 426 812 460
rect 746 420 812 426
rect 860 463 1067 476
rect 1101 463 1117 497
rect 860 460 1117 463
rect 860 426 876 460
rect 910 426 1117 460
rect 860 420 1117 426
rect 1019 414 1117 420
rect 678 352 985 386
rect 610 274 663 290
rect 610 250 626 274
rect 230 196 325 202
rect 28 150 44 184
rect 78 150 94 184
rect 28 108 94 150
rect 130 154 146 188
rect 180 154 196 188
rect 130 120 196 154
rect 130 86 146 120
rect 180 86 196 120
rect 130 17 196 86
rect 230 162 246 196
rect 280 162 325 196
rect 359 240 626 250
rect 660 240 663 274
rect 359 234 663 240
rect 393 216 663 234
rect 393 200 446 216
rect 359 184 446 200
rect 697 169 731 352
rect 932 320 985 352
rect 765 302 818 318
rect 765 268 768 302
rect 802 268 818 302
rect 932 286 948 320
rect 982 286 985 320
rect 932 270 985 286
rect 1019 380 1067 414
rect 1101 380 1117 414
rect 1151 582 1217 649
rect 1151 548 1167 582
rect 1201 548 1217 582
rect 1151 514 1217 548
rect 1151 480 1167 514
rect 1201 480 1217 514
rect 1151 446 1217 480
rect 1151 412 1167 446
rect 1201 412 1217 446
rect 1251 582 1317 596
rect 1251 548 1267 582
rect 1301 548 1317 582
rect 1251 514 1317 548
rect 1251 480 1267 514
rect 1301 480 1317 514
rect 1251 446 1317 480
rect 1251 412 1267 446
rect 1301 412 1317 446
rect 1351 580 1417 649
rect 1351 546 1367 580
rect 1401 546 1417 580
rect 1351 478 1417 546
rect 1351 444 1367 478
rect 1401 444 1417 478
rect 1351 428 1417 444
rect 1019 378 1117 380
rect 1283 394 1317 412
rect 1019 344 1244 378
rect 1283 360 1415 394
rect 765 252 818 268
rect 230 150 325 162
rect 641 153 743 169
rect 230 120 595 150
rect 230 86 246 120
rect 280 116 595 120
rect 641 119 675 153
rect 709 119 743 153
rect 280 86 325 116
rect 230 70 325 86
rect 561 85 595 116
rect 784 85 818 252
rect 1019 226 1053 344
rect 1210 326 1244 344
rect 1210 310 1335 326
rect 1087 294 1168 310
rect 1087 260 1118 294
rect 1152 260 1168 294
rect 1210 276 1226 310
rect 1260 276 1294 310
rect 1328 276 1335 310
rect 1210 260 1335 276
rect 1087 236 1168 260
rect 1369 226 1415 360
rect 969 210 1053 226
rect 969 176 985 210
rect 1019 176 1053 210
rect 1251 210 1415 226
rect 461 48 477 82
rect 511 48 527 82
rect 561 51 818 85
rect 857 140 923 169
rect 857 106 873 140
rect 907 106 923 140
rect 461 17 527 48
rect 857 17 923 106
rect 969 120 1053 176
rect 969 86 985 120
rect 1019 86 1053 120
rect 969 70 1053 86
rect 1151 198 1217 202
rect 1151 164 1167 198
rect 1201 164 1217 198
rect 1151 120 1217 164
rect 1151 86 1167 120
rect 1201 86 1217 120
rect 1151 17 1217 86
rect 1251 176 1267 210
rect 1301 192 1415 210
rect 1301 176 1317 192
rect 1251 120 1317 176
rect 1251 86 1267 120
rect 1301 86 1317 120
rect 1251 70 1317 86
rect 1351 142 1417 158
rect 1351 108 1367 142
rect 1401 108 1417 142
rect 1351 17 1417 108
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 683 1440 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 0 617 1440 649
rect 0 17 1440 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -49 1440 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dlrtp_2
flabel pwell s 0 0 1440 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 1440 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 1440 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 1440 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 D
port 1 nsew
flabel corelocali s 223 242 257 276 0 FreeSans 340 0 0 0 GATE
port 2 nsew
flabel corelocali s 1087 242 1121 276 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew
flabel corelocali s 1375 242 1409 276 0 FreeSans 340 0 0 0 Q
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 1440 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2945362
string GDS_START 2934372
<< end >>
