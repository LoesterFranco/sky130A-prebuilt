magic
tech sky130A
magscale 1 2
timestamp 1599588238
<< locali >>
rect 25 290 110 356
rect 415 368 661 424
rect 511 234 661 368
rect 697 290 839 356
rect 980 290 1127 356
rect 1177 290 1415 356
rect 1465 290 1607 356
rect 310 200 661 234
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 23 581 279 615
rect 23 390 89 581
rect 123 390 178 547
rect 144 334 178 390
rect 213 492 279 581
rect 325 526 391 649
rect 505 526 571 649
rect 685 530 755 649
rect 809 492 875 596
rect 213 458 875 492
rect 927 458 1019 649
rect 213 388 279 458
rect 809 424 875 458
rect 1053 424 1119 596
rect 1153 458 1219 649
rect 1253 424 1319 596
rect 1353 458 1419 649
rect 1453 424 1519 596
rect 809 390 1519 424
rect 1559 390 1609 649
rect 144 268 477 334
rect 144 250 245 268
rect 22 17 72 250
rect 108 166 245 250
rect 108 132 729 166
rect 763 154 969 230
rect 1005 222 1336 256
rect 1005 154 1057 222
rect 763 140 797 154
rect 108 94 174 132
rect 209 17 275 98
rect 411 17 477 98
rect 611 17 661 98
rect 695 85 729 132
rect 935 120 969 154
rect 1091 120 1157 188
rect 833 85 899 120
rect 695 51 899 85
rect 935 66 1157 120
rect 1200 85 1266 188
rect 1302 119 1336 222
rect 1372 222 1610 256
rect 1372 85 1422 222
rect 1200 51 1422 85
rect 1458 17 1524 188
rect 1558 70 1610 222
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
rlabel locali s 697 290 839 356 6 A1
port 1 nsew signal input
rlabel locali s 980 290 1127 356 6 A2
port 2 nsew signal input
rlabel locali s 1177 290 1415 356 6 A3
port 3 nsew signal input
rlabel locali s 1465 290 1607 356 6 A4
port 4 nsew signal input
rlabel locali s 25 290 110 356 6 B1
port 5 nsew signal input
rlabel locali s 511 234 661 368 6 X
port 6 nsew signal output
rlabel locali s 415 368 661 424 6 X
port 6 nsew signal output
rlabel locali s 310 200 661 234 6 X
port 6 nsew signal output
rlabel metal1 s 0 -49 1632 49 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1632 715 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3781754
string GDS_START 3768376
<< end >>
