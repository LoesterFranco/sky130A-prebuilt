magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 710 704
<< pwell >>
rect 0 0 672 49
<< scnmos >>
rect 84 74 114 222
rect 184 74 214 222
rect 273 74 303 222
rect 370 74 400 222
rect 465 74 495 222
rect 558 74 588 222
<< pmoshvt >>
rect 86 368 116 592
rect 176 368 206 592
rect 276 368 306 592
rect 376 368 406 592
rect 466 368 496 592
rect 556 368 586 592
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 150 184 222
rect 114 116 139 150
rect 173 116 184 150
rect 114 74 184 116
rect 214 210 273 222
rect 214 176 225 210
rect 259 176 273 210
rect 214 120 273 176
rect 214 86 225 120
rect 259 86 273 120
rect 214 74 273 86
rect 303 150 370 222
rect 303 116 325 150
rect 359 116 370 150
rect 303 74 370 116
rect 400 210 465 222
rect 400 176 411 210
rect 445 176 465 210
rect 400 120 465 176
rect 400 86 411 120
rect 445 86 465 120
rect 400 74 465 86
rect 495 193 558 222
rect 495 159 512 193
rect 546 159 558 193
rect 495 74 558 159
rect 588 202 645 222
rect 588 168 599 202
rect 633 168 645 202
rect 588 120 645 168
rect 588 86 599 120
rect 633 86 645 120
rect 588 74 645 86
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 508 86 546
rect 27 474 39 508
rect 73 474 86 508
rect 27 368 86 474
rect 116 580 176 592
rect 116 546 129 580
rect 163 546 176 580
rect 116 508 176 546
rect 116 474 129 508
rect 163 474 176 508
rect 116 368 176 474
rect 206 519 276 592
rect 206 485 229 519
rect 263 485 276 519
rect 206 368 276 485
rect 306 578 376 592
rect 306 544 329 578
rect 363 544 376 578
rect 306 368 376 544
rect 406 578 466 592
rect 406 544 419 578
rect 453 544 466 578
rect 406 368 466 544
rect 496 580 556 592
rect 496 546 509 580
rect 543 546 556 580
rect 496 497 556 546
rect 496 463 509 497
rect 543 463 556 497
rect 496 414 556 463
rect 496 380 509 414
rect 543 380 556 414
rect 496 368 556 380
rect 586 580 645 592
rect 586 546 599 580
rect 633 546 645 580
rect 586 497 645 546
rect 586 463 599 497
rect 633 463 645 497
rect 586 414 645 463
rect 586 380 599 414
rect 633 380 645 414
rect 586 368 645 380
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 139 116 173 150
rect 225 176 259 210
rect 225 86 259 120
rect 325 116 359 150
rect 411 176 445 210
rect 411 86 445 120
rect 512 159 546 193
rect 599 168 633 202
rect 599 86 633 120
<< pdiffc >>
rect 39 546 73 580
rect 39 474 73 508
rect 129 546 163 580
rect 129 474 163 508
rect 229 485 263 519
rect 329 544 363 578
rect 419 544 453 578
rect 509 546 543 580
rect 509 463 543 497
rect 509 380 543 414
rect 599 546 633 580
rect 599 463 633 497
rect 599 380 633 414
<< poly >>
rect 86 592 116 618
rect 176 592 206 618
rect 276 592 306 618
rect 376 592 406 618
rect 466 592 496 618
rect 556 592 586 618
rect 86 353 116 368
rect 176 353 206 368
rect 276 353 306 368
rect 376 353 406 368
rect 466 353 496 368
rect 556 353 586 368
rect 83 336 119 353
rect 173 336 209 353
rect 273 336 309 353
rect 373 336 409 353
rect 53 320 119 336
rect 53 286 69 320
rect 103 286 119 320
rect 53 270 119 286
rect 169 320 309 336
rect 169 286 185 320
rect 219 286 253 320
rect 287 300 309 320
rect 351 320 417 336
rect 287 286 303 300
rect 169 270 303 286
rect 351 286 367 320
rect 401 286 417 320
rect 463 323 499 353
rect 553 323 589 353
rect 463 310 589 323
rect 463 304 647 310
rect 351 270 417 286
rect 465 294 647 304
rect 465 274 597 294
rect 84 222 114 270
rect 184 222 214 270
rect 273 222 303 270
rect 370 222 400 270
rect 465 222 495 274
rect 558 260 597 274
rect 631 260 647 294
rect 558 244 647 260
rect 558 222 588 244
rect 84 48 114 74
rect 184 48 214 74
rect 273 48 303 74
rect 370 48 400 74
rect 465 48 495 74
rect 558 48 588 74
<< polycont >>
rect 69 286 103 320
rect 185 286 219 320
rect 253 286 287 320
rect 367 286 401 320
rect 597 260 631 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 23 580 73 649
rect 23 546 39 580
rect 23 508 73 546
rect 23 474 39 508
rect 23 458 73 474
rect 113 581 379 615
rect 113 580 179 581
rect 113 546 129 580
rect 163 546 179 580
rect 313 578 379 581
rect 113 508 179 546
rect 113 474 129 508
rect 163 474 179 508
rect 113 458 179 474
rect 213 519 279 547
rect 313 544 329 578
rect 363 544 379 578
rect 313 526 379 544
rect 419 578 469 649
rect 453 544 469 578
rect 419 526 469 544
rect 505 580 559 596
rect 505 546 509 580
rect 543 546 559 580
rect 213 485 229 519
rect 263 492 279 519
rect 505 497 559 546
rect 505 492 509 497
rect 263 485 509 492
rect 213 463 509 485
rect 543 463 559 497
rect 213 458 559 463
rect 53 390 455 424
rect 53 320 119 390
rect 53 286 69 320
rect 103 286 119 320
rect 53 270 119 286
rect 169 320 303 356
rect 169 286 185 320
rect 219 286 253 320
rect 287 286 303 320
rect 169 270 303 286
rect 351 320 455 390
rect 351 286 367 320
rect 401 286 455 320
rect 351 270 455 286
rect 505 414 559 458
rect 505 380 509 414
rect 543 380 559 414
rect 505 364 559 380
rect 599 580 649 649
rect 633 546 649 580
rect 599 497 649 546
rect 633 463 649 497
rect 599 414 649 463
rect 633 380 649 414
rect 599 364 649 380
rect 23 210 461 236
rect 505 226 547 364
rect 581 294 647 310
rect 581 260 597 294
rect 631 260 647 294
rect 581 236 647 260
rect 23 176 39 210
rect 73 202 225 210
rect 73 176 89 202
rect 23 120 89 176
rect 259 202 411 210
rect 259 176 275 202
rect 23 86 39 120
rect 73 86 89 120
rect 23 70 89 86
rect 123 150 189 166
rect 123 116 139 150
rect 173 116 189 150
rect 123 17 189 116
rect 225 120 275 176
rect 445 176 461 210
rect 259 86 275 120
rect 225 70 275 86
rect 309 150 375 166
rect 309 116 325 150
rect 359 116 375 150
rect 309 17 375 116
rect 411 120 461 176
rect 495 193 547 226
rect 495 159 512 193
rect 546 159 547 193
rect 495 143 547 159
rect 583 168 599 202
rect 633 168 649 202
rect 445 104 461 120
rect 583 120 649 168
rect 583 104 599 120
rect 445 86 599 104
rect 633 86 649 120
rect 411 70 649 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o21ai_2
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 607 242 641 276 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 511 390 545 424 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 511 464 545 498 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 511 538 545 572 0 FreeSans 340 0 0 0 Y
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 672 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1353620
string GDS_START 1347090
<< end >>
