magic
tech sky130A
magscale 1 2
timestamp 1604502741
<< locali >>
rect 25 291 110 357
rect 167 291 263 357
rect 1541 394 1607 596
rect 1731 394 1797 596
rect 1541 360 1797 394
rect 1157 236 1223 310
rect 1745 282 1797 360
rect 1745 226 1811 282
rect 1573 192 1811 226
rect 1573 70 1623 192
rect 1745 70 1811 192
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 23 391 89 649
rect 197 496 263 567
rect 309 530 432 649
rect 585 496 651 551
rect 197 462 651 496
rect 197 391 331 462
rect 23 17 89 257
rect 123 157 189 257
rect 297 157 331 391
rect 473 347 539 428
rect 585 381 651 462
rect 365 313 651 347
rect 365 191 415 313
rect 585 281 651 313
rect 685 281 741 551
rect 886 415 936 649
rect 976 482 1054 579
rect 1196 516 1262 649
rect 976 448 1291 482
rect 976 381 1054 448
rect 792 347 1054 381
rect 1088 364 1155 414
rect 792 315 858 347
rect 920 281 986 313
rect 449 247 515 279
rect 685 247 986 281
rect 449 213 595 247
rect 461 157 527 179
rect 123 123 527 157
rect 225 17 313 89
rect 461 70 527 123
rect 561 88 595 213
rect 685 188 719 247
rect 1020 213 1054 347
rect 629 122 719 188
rect 753 179 955 213
rect 753 88 787 179
rect 561 54 787 88
rect 821 17 887 145
rect 921 85 955 179
rect 989 119 1055 213
rect 1089 202 1123 364
rect 1257 326 1291 448
rect 1325 394 1391 596
rect 1425 428 1491 649
rect 1647 428 1697 649
rect 1325 360 1507 394
rect 1831 364 1897 649
rect 1473 326 1507 360
rect 1257 260 1406 326
rect 1473 260 1687 326
rect 1473 226 1507 260
rect 1089 85 1167 202
rect 921 51 1167 85
rect 1201 17 1267 202
rect 1365 192 1507 226
rect 1365 70 1431 192
rect 1477 17 1527 158
rect 1659 17 1709 158
rect 1847 17 1897 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
<< metal1 >>
rect 0 683 1920 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 0 617 1920 649
rect 0 17 1920 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
rect 0 -49 1920 -17
<< labels >>
rlabel locali s 167 291 263 357 6 GATE
port 1 nsew signal input
rlabel locali s 1745 282 1797 360 6 GCLK
port 2 nsew signal output
rlabel locali s 1745 226 1811 282 6 GCLK
port 2 nsew signal output
rlabel locali s 1745 70 1811 192 6 GCLK
port 2 nsew signal output
rlabel locali s 1731 394 1797 596 6 GCLK
port 2 nsew signal output
rlabel locali s 1573 192 1811 226 6 GCLK
port 2 nsew signal output
rlabel locali s 1573 70 1623 192 6 GCLK
port 2 nsew signal output
rlabel locali s 1541 394 1607 596 6 GCLK
port 2 nsew signal output
rlabel locali s 1541 360 1797 394 6 GCLK
port 2 nsew signal output
rlabel locali s 25 291 110 357 6 SCE
port 3 nsew signal input
rlabel locali s 1157 236 1223 310 6 CLK
port 4 nsew clock input
rlabel metal1 s 0 -49 1920 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 617 1920 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1920 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 338952
string GDS_START 326072
<< end >>
