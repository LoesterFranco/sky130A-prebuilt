magic
tech sky130A
magscale 1 2
timestamp 1604502729
<< locali >>
rect 486 424 552 547
rect 676 424 742 547
rect 988 424 1054 596
rect 1188 424 1254 596
rect 1509 424 1607 578
rect 486 390 1607 424
rect 25 270 359 356
rect 409 270 839 356
rect 889 270 1127 356
rect 1174 270 1415 356
rect 1473 310 1607 390
rect 1473 236 1509 310
rect 1301 202 1509 236
rect 1301 119 1335 202
rect 1473 119 1509 202
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 26 424 92 596
rect 132 458 166 649
rect 206 424 272 596
rect 312 458 346 649
rect 386 581 842 615
rect 386 424 452 581
rect 26 390 452 424
rect 592 458 642 581
rect 776 458 842 581
rect 888 458 954 649
rect 1088 458 1154 649
rect 1288 458 1458 649
rect 23 202 1153 236
rect 23 70 89 202
rect 123 17 189 168
rect 225 70 275 202
rect 309 17 375 168
rect 411 70 445 202
rect 481 17 547 168
rect 583 70 617 202
rect 653 17 719 168
rect 759 164 981 202
rect 759 70 793 164
rect 1017 130 1051 168
rect 829 85 1051 130
rect 1087 119 1153 202
rect 1199 85 1265 236
rect 1371 85 1437 168
rect 1543 85 1609 236
rect 829 51 1609 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
rlabel locali s 25 270 359 356 6 A1
port 1 nsew signal input
rlabel locali s 409 270 839 356 6 A2
port 2 nsew signal input
rlabel locali s 889 270 1127 356 6 B1
port 3 nsew signal input
rlabel locali s 1174 270 1415 356 6 C1
port 4 nsew signal input
rlabel locali s 1509 424 1607 578 6 Y
port 5 nsew signal output
rlabel locali s 1473 310 1607 390 6 Y
port 5 nsew signal output
rlabel locali s 1473 236 1509 310 6 Y
port 5 nsew signal output
rlabel locali s 1473 119 1509 202 6 Y
port 5 nsew signal output
rlabel locali s 1301 202 1509 236 6 Y
port 5 nsew signal output
rlabel locali s 1301 119 1335 202 6 Y
port 5 nsew signal output
rlabel locali s 1188 424 1254 596 6 Y
port 5 nsew signal output
rlabel locali s 988 424 1054 596 6 Y
port 5 nsew signal output
rlabel locali s 676 424 742 547 6 Y
port 5 nsew signal output
rlabel locali s 486 424 552 547 6 Y
port 5 nsew signal output
rlabel locali s 486 390 1607 424 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -49 1632 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 1632 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1080700
string GDS_START 1066836
<< end >>
