magic
tech sky130A
magscale 1 2
timestamp 1601050082
<< locali >>
rect 327 464 569 498
rect 21 228 82 294
rect 327 294 361 464
rect 184 228 257 294
rect 291 228 361 294
rect 395 224 461 430
rect 503 289 569 464
rect 771 392 847 596
rect 603 224 677 290
rect 813 226 847 392
rect 774 70 847 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 27 362 93 591
rect 127 396 193 649
rect 227 557 637 591
rect 227 362 293 557
rect 27 328 293 362
rect 116 194 150 328
rect 603 358 637 557
rect 671 392 737 649
rect 603 324 779 358
rect 719 270 779 324
rect 40 160 150 194
rect 40 70 106 160
rect 212 122 278 194
rect 312 156 738 190
rect 212 56 636 122
rect 672 17 738 156
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel locali s 603 224 677 290 6 A1
port 1 nsew signal input
rlabel locali s 503 289 569 464 6 A2
port 2 nsew signal input
rlabel locali s 327 464 569 498 6 A2
port 2 nsew signal input
rlabel locali s 327 294 361 464 6 A2
port 2 nsew signal input
rlabel locali s 291 228 361 294 6 A2
port 2 nsew signal input
rlabel locali s 395 224 461 430 6 A3
port 3 nsew signal input
rlabel locali s 184 228 257 294 6 B1
port 4 nsew signal input
rlabel locali s 21 228 82 294 6 C1
port 5 nsew signal input
rlabel locali s 813 226 847 392 6 X
port 6 nsew signal output
rlabel locali s 774 70 847 226 6 X
port 6 nsew signal output
rlabel locali s 771 392 847 596 6 X
port 6 nsew signal output
rlabel metal1 s 0 -49 864 49 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 617 864 715 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 743424
string GDS_START 735572
<< end >>
