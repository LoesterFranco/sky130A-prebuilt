magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 736 561
rect 23 289 73 527
rect 37 17 71 177
rect 118 73 161 493
rect 199 375 359 527
rect 580 323 620 481
rect 654 359 718 527
rect 549 289 620 323
rect 549 265 585 289
rect 287 215 358 265
rect 392 215 485 265
rect 519 215 585 265
rect 654 255 718 323
rect 619 215 718 255
rect 205 17 241 109
rect 583 17 617 105
rect 0 -17 736 17
<< obsli1 >>
rect 438 341 515 493
rect 195 299 515 341
rect 195 179 251 299
rect 195 143 443 179
rect 512 165 718 173
rect 370 129 443 143
rect 478 139 718 165
rect 478 95 546 139
rect 293 59 546 95
rect 651 56 718 139
<< metal1 >>
rect 0 496 736 592
rect 0 -48 736 48
<< labels >>
rlabel locali s 654 255 718 323 6 A1
port 1 nsew signal input
rlabel locali s 619 215 718 255 6 A1
port 1 nsew signal input
rlabel locali s 580 323 620 481 6 A2
port 2 nsew signal input
rlabel locali s 549 289 620 323 6 A2
port 2 nsew signal input
rlabel locali s 549 265 585 289 6 A2
port 2 nsew signal input
rlabel locali s 519 215 585 265 6 A2
port 2 nsew signal input
rlabel locali s 287 215 358 265 6 B1
port 3 nsew signal input
rlabel locali s 392 215 485 265 6 B2
port 4 nsew signal input
rlabel locali s 118 73 161 493 6 X
port 5 nsew signal output
rlabel locali s 583 17 617 105 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 205 17 241 109 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 37 17 71 177 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 736 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 736 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 654 359 718 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 199 375 359 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 23 289 73 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 736 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 736 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1479446
string GDS_START 1472852
<< end >>
