magic
tech sky130A
magscale 1 2
timestamp 1601050039
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 527 47 557 177
rect 611 47 641 177
rect 695 47 725 177
rect 779 47 809 177
<< pmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 447 297 477 497
rect 531 297 561 497
rect 695 297 725 497
rect 779 297 809 497
<< ndiff >>
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 93 163 177
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 161 247 177
rect 193 127 203 161
rect 237 127 247 161
rect 193 93 247 127
rect 193 59 203 93
rect 237 59 247 93
rect 193 47 247 59
rect 277 161 331 177
rect 277 127 287 161
rect 321 127 331 161
rect 277 47 331 127
rect 361 93 417 177
rect 361 59 375 93
rect 409 59 417 93
rect 361 47 417 59
rect 471 93 527 177
rect 471 59 479 93
rect 513 59 527 93
rect 471 47 527 59
rect 557 161 611 177
rect 557 127 567 161
rect 601 127 611 161
rect 557 47 611 127
rect 641 161 695 177
rect 641 127 651 161
rect 685 127 695 161
rect 641 93 695 127
rect 641 59 651 93
rect 685 59 695 93
rect 641 47 695 59
rect 725 161 779 177
rect 725 127 735 161
rect 769 127 779 161
rect 725 47 779 127
rect 809 161 881 177
rect 809 127 835 161
rect 869 127 881 161
rect 809 93 881 127
rect 809 59 835 93
rect 869 59 881 93
rect 809 47 881 59
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 485 163 497
rect 109 451 119 485
rect 153 451 163 485
rect 109 417 163 451
rect 109 383 119 417
rect 153 383 163 417
rect 109 349 163 383
rect 109 315 119 349
rect 153 315 163 349
rect 109 297 163 315
rect 193 485 247 497
rect 193 451 203 485
rect 237 451 247 485
rect 193 417 247 451
rect 193 383 203 417
rect 237 383 247 417
rect 193 297 247 383
rect 277 485 331 497
rect 277 451 287 485
rect 321 451 331 485
rect 277 417 331 451
rect 277 383 287 417
rect 321 383 331 417
rect 277 349 331 383
rect 277 315 287 349
rect 321 315 331 349
rect 277 297 331 315
rect 361 485 447 497
rect 361 451 387 485
rect 421 451 447 485
rect 361 417 447 451
rect 361 383 387 417
rect 421 383 447 417
rect 361 297 447 383
rect 477 485 531 497
rect 477 451 487 485
rect 521 451 531 485
rect 477 417 531 451
rect 477 383 487 417
rect 521 383 531 417
rect 477 349 531 383
rect 477 315 487 349
rect 521 315 531 349
rect 477 297 531 315
rect 561 485 695 497
rect 561 451 615 485
rect 649 451 695 485
rect 561 417 695 451
rect 561 383 615 417
rect 649 383 695 417
rect 561 297 695 383
rect 725 485 779 497
rect 725 451 735 485
rect 769 451 779 485
rect 725 417 779 451
rect 725 383 735 417
rect 769 383 779 417
rect 725 349 779 383
rect 725 315 735 349
rect 769 315 779 349
rect 725 297 779 315
rect 809 485 893 497
rect 809 451 835 485
rect 869 451 893 485
rect 809 417 893 451
rect 809 383 835 417
rect 869 383 893 417
rect 809 349 893 383
rect 809 315 835 349
rect 869 315 893 349
rect 809 297 893 315
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 119 59 153 93
rect 203 127 237 161
rect 203 59 237 93
rect 287 127 321 161
rect 375 59 409 93
rect 479 59 513 93
rect 567 127 601 161
rect 651 127 685 161
rect 651 59 685 93
rect 735 127 769 161
rect 835 127 869 161
rect 835 59 869 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 119 451 153 485
rect 119 383 153 417
rect 119 315 153 349
rect 203 451 237 485
rect 203 383 237 417
rect 287 451 321 485
rect 287 383 321 417
rect 287 315 321 349
rect 387 451 421 485
rect 387 383 421 417
rect 487 451 521 485
rect 487 383 521 417
rect 487 315 521 349
rect 615 451 649 485
rect 615 383 649 417
rect 735 451 769 485
rect 735 383 769 417
rect 735 315 769 349
rect 835 451 869 485
rect 835 383 869 417
rect 835 315 869 349
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 447 497 477 523
rect 531 497 561 523
rect 695 497 725 523
rect 779 497 809 523
rect 79 261 109 297
rect 22 259 109 261
rect 163 259 193 297
rect 22 249 193 259
rect 22 215 38 249
rect 72 215 119 249
rect 153 215 193 249
rect 22 205 193 215
rect 22 203 109 205
rect 79 177 109 203
rect 163 177 193 205
rect 247 259 277 297
rect 331 259 361 297
rect 247 249 361 259
rect 247 215 287 249
rect 321 215 361 249
rect 247 205 361 215
rect 447 259 477 297
rect 531 259 561 297
rect 695 259 725 297
rect 779 261 809 297
rect 779 259 899 261
rect 447 249 641 259
rect 447 215 463 249
rect 497 215 561 249
rect 595 215 641 249
rect 447 205 641 215
rect 247 177 277 205
rect 331 177 361 205
rect 527 177 557 205
rect 611 177 641 205
rect 695 249 899 259
rect 695 215 849 249
rect 883 215 899 249
rect 695 205 899 215
rect 695 177 725 205
rect 779 203 899 205
rect 779 177 809 203
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 527 21 557 47
rect 611 21 641 47
rect 695 21 725 47
rect 779 21 809 47
<< polycont >>
rect 38 215 72 249
rect 119 215 153 249
rect 287 215 321 249
rect 463 215 497 249
rect 561 215 595 249
rect 849 215 883 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 18 485 69 527
rect 18 451 35 485
rect 18 417 69 451
rect 18 383 35 417
rect 18 349 69 383
rect 18 315 35 349
rect 18 299 69 315
rect 103 485 169 493
rect 103 451 119 485
rect 153 451 169 485
rect 103 417 169 451
rect 103 383 119 417
rect 153 383 169 417
rect 103 349 169 383
rect 203 485 237 527
rect 203 417 237 451
rect 203 367 237 383
rect 271 485 337 493
rect 271 451 287 485
rect 321 451 337 485
rect 271 417 337 451
rect 271 383 287 417
rect 321 383 337 417
rect 103 315 119 349
rect 153 333 169 349
rect 271 349 337 383
rect 371 485 437 527
rect 371 451 387 485
rect 421 451 437 485
rect 371 417 437 451
rect 371 383 387 417
rect 421 383 437 417
rect 371 367 437 383
rect 471 485 537 493
rect 471 451 487 485
rect 521 451 537 485
rect 471 417 537 451
rect 471 383 487 417
rect 521 383 537 417
rect 271 333 287 349
rect 153 315 287 333
rect 321 333 337 349
rect 471 349 537 383
rect 599 485 665 527
rect 599 451 615 485
rect 649 451 665 485
rect 599 417 665 451
rect 599 383 615 417
rect 649 383 665 417
rect 599 367 665 383
rect 719 485 785 493
rect 719 451 735 485
rect 769 451 785 485
rect 719 417 785 451
rect 719 383 735 417
rect 769 383 785 417
rect 471 333 487 349
rect 321 315 487 333
rect 521 333 537 349
rect 719 349 785 383
rect 719 333 735 349
rect 521 315 735 333
rect 769 315 785 349
rect 103 289 785 315
rect 819 485 885 527
rect 819 451 835 485
rect 869 451 885 485
rect 819 417 885 451
rect 819 383 835 417
rect 869 383 885 417
rect 819 349 885 383
rect 819 315 835 349
rect 869 315 885 349
rect 819 289 885 315
rect 22 249 169 255
rect 22 215 38 249
rect 72 215 119 249
rect 153 215 169 249
rect 214 249 340 255
rect 214 215 287 249
rect 321 215 340 249
rect 447 249 616 255
rect 447 215 463 249
rect 497 215 561 249
rect 595 215 616 249
rect 674 211 785 289
rect 833 249 899 255
rect 833 215 849 249
rect 883 215 899 249
rect 18 161 237 181
rect 18 127 35 161
rect 69 147 203 161
rect 69 127 85 147
rect 18 93 85 127
rect 187 127 203 147
rect 271 161 617 181
rect 271 127 287 161
rect 321 127 567 161
rect 601 127 617 161
rect 651 161 685 177
rect 719 161 785 211
rect 719 127 735 161
rect 769 127 785 161
rect 819 161 885 181
rect 819 127 835 161
rect 869 127 885 161
rect 18 59 35 93
rect 69 59 85 93
rect 18 51 85 59
rect 119 93 153 109
rect 119 17 153 59
rect 187 93 237 127
rect 651 93 685 127
rect 819 93 885 127
rect 187 59 203 93
rect 237 59 375 93
rect 409 59 425 93
rect 187 51 425 59
rect 463 59 479 93
rect 513 59 651 93
rect 685 59 835 93
rect 869 59 885 93
rect 463 51 885 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel corelocali s 582 221 616 255 0 FreeSans 250 0 0 0 B
port 2 nsew
flabel corelocali s 490 221 524 255 0 FreeSans 250 0 0 0 B
port 2 nsew
flabel corelocali s 857 221 891 255 0 FreeSans 250 0 0 0 A
port 1 nsew
flabel corelocali s 490 289 524 323 0 FreeSans 250 0 0 0 Y
port 9 nsew
flabel corelocali s 582 289 616 323 0 FreeSans 250 0 0 0 Y
port 9 nsew
flabel corelocali s 674 221 708 255 0 FreeSans 250 0 0 0 Y
port 9 nsew
flabel corelocali s 674 289 708 323 0 FreeSans 250 0 0 0 Y
port 9 nsew
flabel corelocali s 122 221 156 255 0 FreeSans 250 0 0 0 D
port 4 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 250 0 0 0 D
port 4 nsew
flabel corelocali s 306 221 340 255 0 FreeSans 250 0 0 0 C
port 3 nsew
flabel corelocali s 214 221 248 255 0 FreeSans 250 0 0 0 C
port 3 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
rlabel comment s 0 0 0 0 4 nand4_2
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1850160
string GDS_START 1841432
string path 0.000 0.000 23.000 0.000 
<< end >>
