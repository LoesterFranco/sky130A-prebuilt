magic
tech sky130A
magscale 1 2
timestamp 1604502693
<< nwell >>
rect -38 261 1970 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 351 47 381 175
rect 446 47 476 119
rect 556 47 586 119
rect 652 47 682 131
rect 766 47 796 131
rect 838 47 868 131
rect 1026 47 1056 131
rect 1098 47 1128 131
rect 1198 47 1228 131
rect 1270 47 1300 131
rect 1342 47 1372 131
rect 1466 47 1496 155
rect 1654 47 1684 177
rect 1738 47 1768 177
rect 1822 47 1852 177
<< pmoshvt >>
rect 79 363 109 491
rect 163 363 193 491
rect 351 329 381 497
rect 448 413 478 497
rect 532 413 562 497
rect 652 413 682 497
rect 758 413 788 497
rect 842 413 872 497
rect 926 413 956 497
rect 998 413 1028 497
rect 1106 413 1136 497
rect 1178 413 1208 497
rect 1366 413 1396 497
rect 1461 329 1491 497
rect 1654 297 1684 497
rect 1738 297 1768 497
rect 1822 297 1852 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 299 93 351 175
rect 299 59 307 93
rect 341 59 351 93
rect 299 47 351 59
rect 381 119 431 175
rect 1416 131 1466 155
rect 601 119 652 131
rect 381 111 446 119
rect 381 77 391 111
rect 425 77 446 111
rect 381 47 446 77
rect 476 93 556 119
rect 476 59 501 93
rect 535 59 556 93
rect 476 47 556 59
rect 586 47 652 119
rect 682 89 766 131
rect 682 55 722 89
rect 756 55 766 89
rect 682 47 766 55
rect 796 47 838 131
rect 868 109 920 131
rect 868 75 878 109
rect 912 75 920 109
rect 868 47 920 75
rect 974 93 1026 131
rect 974 59 982 93
rect 1016 59 1026 93
rect 974 47 1026 59
rect 1056 47 1098 131
rect 1128 95 1198 131
rect 1128 61 1144 95
rect 1178 61 1198 95
rect 1128 47 1198 61
rect 1228 47 1270 131
rect 1300 47 1342 131
rect 1372 113 1466 131
rect 1372 79 1402 113
rect 1436 79 1466 113
rect 1372 47 1466 79
rect 1496 120 1548 155
rect 1496 86 1506 120
rect 1540 86 1548 120
rect 1496 47 1548 86
rect 1602 119 1654 177
rect 1602 85 1610 119
rect 1644 85 1654 119
rect 1602 47 1654 85
rect 1684 161 1738 177
rect 1684 127 1694 161
rect 1728 127 1738 161
rect 1684 93 1738 127
rect 1684 59 1694 93
rect 1728 59 1738 93
rect 1684 47 1738 59
rect 1768 143 1822 177
rect 1768 109 1778 143
rect 1812 109 1822 143
rect 1768 47 1822 109
rect 1852 93 1904 177
rect 1852 59 1862 93
rect 1896 59 1904 93
rect 1852 47 1904 59
<< pdiff >>
rect 27 477 79 491
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 363 79 375
rect 109 461 163 491
rect 109 427 119 461
rect 153 427 163 461
rect 109 363 163 427
rect 193 477 245 491
rect 193 443 203 477
rect 237 443 245 477
rect 193 409 245 443
rect 193 375 203 409
rect 237 375 245 409
rect 193 363 245 375
rect 299 461 351 497
rect 299 427 307 461
rect 341 427 351 461
rect 299 329 351 427
rect 381 477 448 497
rect 381 443 391 477
rect 425 443 448 477
rect 381 413 448 443
rect 478 484 532 497
rect 478 450 488 484
rect 522 450 532 484
rect 478 413 532 450
rect 562 413 652 497
rect 682 485 758 497
rect 682 451 702 485
rect 736 451 758 485
rect 682 413 758 451
rect 788 459 842 497
rect 788 425 798 459
rect 832 425 842 459
rect 788 413 842 425
rect 872 485 926 497
rect 872 451 882 485
rect 916 451 926 485
rect 872 413 926 451
rect 956 413 998 497
rect 1028 483 1106 497
rect 1028 449 1038 483
rect 1072 449 1106 483
rect 1028 413 1106 449
rect 1136 413 1178 497
rect 1208 485 1260 497
rect 1208 451 1218 485
rect 1252 451 1260 485
rect 1208 413 1260 451
rect 1314 459 1366 497
rect 1314 425 1322 459
rect 1356 425 1366 459
rect 1314 413 1366 425
rect 1396 459 1461 497
rect 1396 425 1417 459
rect 1451 425 1461 459
rect 1396 413 1461 425
rect 381 409 433 413
rect 381 375 391 409
rect 425 375 433 409
rect 381 329 433 375
rect 1411 329 1461 413
rect 1491 459 1544 497
rect 1491 425 1502 459
rect 1536 425 1544 459
rect 1491 391 1544 425
rect 1491 357 1502 391
rect 1536 357 1544 391
rect 1491 329 1544 357
rect 1602 485 1654 497
rect 1602 451 1610 485
rect 1644 451 1654 485
rect 1602 417 1654 451
rect 1602 383 1610 417
rect 1644 383 1654 417
rect 1602 349 1654 383
rect 1602 315 1610 349
rect 1644 315 1654 349
rect 1602 297 1654 315
rect 1684 485 1738 497
rect 1684 451 1694 485
rect 1728 451 1738 485
rect 1684 417 1738 451
rect 1684 383 1694 417
rect 1728 383 1738 417
rect 1684 349 1738 383
rect 1684 315 1694 349
rect 1728 315 1738 349
rect 1684 297 1738 315
rect 1768 485 1822 497
rect 1768 451 1778 485
rect 1812 451 1822 485
rect 1768 417 1822 451
rect 1768 383 1778 417
rect 1812 383 1822 417
rect 1768 349 1822 383
rect 1768 315 1778 349
rect 1812 315 1822 349
rect 1768 297 1822 315
rect 1852 485 1904 497
rect 1852 451 1862 485
rect 1896 451 1904 485
rect 1852 408 1904 451
rect 1852 374 1862 408
rect 1896 374 1904 408
rect 1852 297 1904 374
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 307 59 341 93
rect 391 77 425 111
rect 501 59 535 93
rect 722 55 756 89
rect 878 75 912 109
rect 982 59 1016 93
rect 1144 61 1178 95
rect 1402 79 1436 113
rect 1506 86 1540 120
rect 1610 85 1644 119
rect 1694 127 1728 161
rect 1694 59 1728 93
rect 1778 109 1812 143
rect 1862 59 1896 93
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 427 153 461
rect 203 443 237 477
rect 203 375 237 409
rect 307 427 341 461
rect 391 443 425 477
rect 488 450 522 484
rect 702 451 736 485
rect 798 425 832 459
rect 882 451 916 485
rect 1038 449 1072 483
rect 1218 451 1252 485
rect 1322 425 1356 459
rect 1417 425 1451 459
rect 391 375 425 409
rect 1502 425 1536 459
rect 1502 357 1536 391
rect 1610 451 1644 485
rect 1610 383 1644 417
rect 1610 315 1644 349
rect 1694 451 1728 485
rect 1694 383 1728 417
rect 1694 315 1728 349
rect 1778 451 1812 485
rect 1778 383 1812 417
rect 1778 315 1812 349
rect 1862 451 1896 485
rect 1862 374 1896 408
<< poly >>
rect 79 491 109 517
rect 163 491 193 517
rect 351 497 381 523
rect 448 497 478 523
rect 532 497 562 523
rect 652 497 682 523
rect 758 497 788 523
rect 842 497 872 523
rect 926 497 956 523
rect 998 497 1028 523
rect 1106 497 1136 523
rect 1178 497 1208 523
rect 1366 497 1396 523
rect 1461 497 1491 523
rect 1654 497 1684 523
rect 1738 497 1768 523
rect 1822 497 1852 523
rect 79 348 109 363
rect 45 318 109 348
rect 45 280 75 318
rect 21 264 75 280
rect 163 274 193 363
rect 21 230 31 264
rect 65 230 75 264
rect 21 214 75 230
rect 117 264 193 274
rect 351 267 381 329
rect 448 279 478 413
rect 532 375 562 413
rect 652 381 682 413
rect 520 365 586 375
rect 520 331 536 365
rect 570 331 586 365
rect 520 321 586 331
rect 652 365 716 381
rect 652 331 672 365
rect 706 331 716 365
rect 652 315 716 331
rect 117 230 133 264
rect 167 230 193 264
rect 117 220 193 230
rect 45 176 75 214
rect 45 146 109 176
rect 79 131 109 146
rect 163 131 193 220
rect 344 251 398 267
rect 344 217 354 251
rect 388 217 398 251
rect 448 249 586 279
rect 344 201 398 217
rect 556 219 586 249
rect 351 175 381 201
rect 446 191 514 207
rect 446 157 470 191
rect 504 157 514 191
rect 446 141 514 157
rect 556 203 610 219
rect 556 169 566 203
rect 600 169 610 203
rect 556 153 610 169
rect 446 119 476 141
rect 556 119 586 153
rect 652 131 682 315
rect 758 229 788 413
rect 842 313 872 413
rect 926 313 956 413
rect 998 375 1028 413
rect 998 365 1064 375
rect 998 331 1014 365
rect 1048 331 1064 365
rect 998 321 1064 331
rect 830 297 956 313
rect 830 263 840 297
rect 874 263 956 297
rect 1106 291 1136 413
rect 1094 279 1136 291
rect 830 247 956 263
rect 1030 269 1136 279
rect 728 213 788 229
rect 728 179 738 213
rect 772 193 788 213
rect 772 179 796 193
rect 728 163 796 179
rect 766 131 796 163
rect 838 183 868 247
rect 1030 235 1046 269
rect 1080 261 1136 269
rect 1178 365 1208 413
rect 1178 349 1242 365
rect 1178 315 1198 349
rect 1232 315 1242 349
rect 1366 337 1396 413
rect 1178 291 1242 315
rect 1178 261 1300 291
rect 1080 235 1128 261
rect 1030 225 1128 235
rect 838 147 1056 183
rect 838 131 868 147
rect 1026 131 1056 147
rect 1098 131 1128 225
rect 1170 203 1228 219
rect 1170 169 1180 203
rect 1214 169 1228 203
rect 1170 153 1228 169
rect 1198 131 1228 153
rect 1270 131 1300 261
rect 1362 229 1396 337
rect 1461 285 1491 329
rect 1342 213 1396 229
rect 1438 282 1491 285
rect 1654 282 1684 297
rect 1438 269 1684 282
rect 1438 235 1448 269
rect 1482 235 1684 269
rect 1738 265 1768 297
rect 1822 265 1852 297
rect 1438 219 1684 235
rect 1342 179 1352 213
rect 1386 179 1396 213
rect 1342 163 1396 179
rect 1342 131 1372 163
rect 1466 155 1496 219
rect 1654 177 1684 219
rect 1726 249 1852 265
rect 1726 215 1736 249
rect 1770 215 1852 249
rect 1726 199 1852 215
rect 1738 177 1768 199
rect 1822 177 1852 199
rect 79 21 109 47
rect 163 21 193 47
rect 351 21 381 47
rect 446 21 476 47
rect 556 21 586 47
rect 652 21 682 47
rect 766 21 796 47
rect 838 21 868 47
rect 1026 21 1056 47
rect 1098 21 1128 47
rect 1198 21 1228 47
rect 1270 21 1300 47
rect 1342 21 1372 47
rect 1466 21 1496 47
rect 1654 21 1684 47
rect 1738 21 1768 47
rect 1822 21 1852 47
<< polycont >>
rect 31 230 65 264
rect 536 331 570 365
rect 672 331 706 365
rect 133 230 167 264
rect 354 217 388 251
rect 470 157 504 191
rect 566 169 600 203
rect 1014 331 1048 365
rect 840 263 874 297
rect 738 179 772 213
rect 1046 235 1080 269
rect 1198 315 1232 349
rect 1180 169 1214 203
rect 1448 235 1482 269
rect 1352 179 1386 213
rect 1736 215 1770 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 17 477 69 493
rect 17 443 35 477
rect 17 409 69 443
rect 103 461 169 527
rect 103 427 119 461
rect 153 427 169 461
rect 203 477 247 493
rect 237 443 247 477
rect 203 409 247 443
rect 291 461 357 527
rect 291 427 307 461
rect 341 427 357 461
rect 391 477 425 493
rect 686 485 762 527
rect 472 450 488 484
rect 522 450 638 484
rect 686 451 702 485
rect 736 451 762 485
rect 866 485 932 527
rect 798 459 832 475
rect 17 375 35 409
rect 69 391 167 393
rect 69 375 121 391
rect 17 359 121 375
rect 155 357 167 391
rect 17 264 87 325
rect 17 230 31 264
rect 65 230 87 264
rect 17 195 87 230
rect 121 264 167 357
rect 121 230 133 264
rect 121 161 167 230
rect 17 127 167 161
rect 201 375 203 409
rect 237 375 247 409
rect 391 409 425 443
rect 201 187 247 375
rect 201 153 213 187
rect 17 119 69 127
rect 17 85 35 119
rect 201 119 247 153
rect 286 375 391 393
rect 286 359 425 375
rect 286 165 320 359
rect 470 357 489 391
rect 523 365 570 391
rect 523 357 536 365
rect 470 331 536 357
rect 354 251 436 325
rect 388 217 436 251
rect 354 201 436 217
rect 470 315 570 331
rect 470 191 514 315
rect 604 281 638 450
rect 866 451 882 485
rect 916 451 932 485
rect 1184 485 1268 527
rect 1022 449 1038 483
rect 1072 449 1148 483
rect 1184 451 1218 485
rect 1252 451 1268 485
rect 1308 459 1356 475
rect 1022 433 1148 449
rect 798 417 832 425
rect 1114 417 1148 433
rect 1308 425 1322 459
rect 1308 417 1356 425
rect 672 367 942 417
rect 672 365 722 367
rect 706 331 722 365
rect 672 315 722 331
rect 824 297 874 313
rect 824 281 840 297
rect 604 263 840 281
rect 604 247 874 263
rect 604 239 688 247
rect 286 127 425 165
rect 504 157 514 191
rect 470 141 514 157
rect 550 169 566 203
rect 600 187 620 203
rect 550 153 581 169
rect 615 153 620 187
rect 550 129 620 153
rect 201 113 203 119
rect 17 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 237 85 247 119
rect 391 111 425 127
rect 203 69 247 85
rect 103 17 169 59
rect 291 59 307 93
rect 341 59 357 93
rect 654 93 688 239
rect 908 213 942 367
rect 722 179 738 213
rect 772 187 804 213
rect 722 153 765 179
rect 799 153 804 187
rect 722 147 804 153
rect 862 145 942 213
rect 976 391 1080 393
rect 976 365 1041 391
rect 976 331 1014 365
rect 1075 357 1080 391
rect 1048 331 1080 357
rect 1114 383 1356 417
rect 1402 459 1468 527
rect 1694 485 1728 527
rect 1402 425 1417 459
rect 1451 425 1468 459
rect 1402 389 1468 425
rect 1502 459 1536 475
rect 1502 391 1536 425
rect 976 179 1010 331
rect 1044 269 1080 295
rect 1044 255 1046 269
rect 1044 221 1045 255
rect 1114 281 1148 383
rect 1594 451 1610 485
rect 1644 451 1660 485
rect 1594 417 1660 451
rect 1594 383 1610 417
rect 1644 383 1660 417
rect 1502 353 1536 357
rect 1502 349 1576 353
rect 1182 315 1198 349
rect 1232 315 1576 349
rect 1114 269 1498 281
rect 1114 247 1448 269
rect 1079 221 1080 235
rect 1044 213 1080 221
rect 1160 179 1180 203
rect 976 169 1180 179
rect 1214 169 1230 203
rect 976 145 1230 169
rect 862 109 912 145
rect 391 61 425 77
rect 291 17 357 59
rect 485 59 501 93
rect 535 59 688 93
rect 485 53 688 59
rect 722 89 804 105
rect 756 55 804 89
rect 862 75 878 109
rect 862 59 912 75
rect 952 93 1016 109
rect 1264 95 1298 247
rect 1428 235 1448 247
rect 1482 235 1498 269
rect 1332 179 1352 213
rect 1386 201 1402 213
rect 1386 187 1468 201
rect 1386 179 1409 187
rect 1332 153 1409 179
rect 1443 153 1468 187
rect 1332 147 1468 153
rect 1538 136 1576 315
rect 1506 120 1576 136
rect 952 59 982 93
rect 1128 61 1144 95
rect 1178 61 1298 95
rect 1338 79 1402 113
rect 1436 79 1466 113
rect 722 17 804 55
rect 952 17 1016 59
rect 1338 17 1466 79
rect 1540 86 1576 120
rect 1506 70 1576 86
rect 1610 349 1660 383
rect 1644 315 1660 349
rect 1610 265 1660 315
rect 1694 417 1728 451
rect 1694 349 1728 383
rect 1694 299 1728 315
rect 1762 485 1828 492
rect 1762 451 1778 485
rect 1812 451 1828 485
rect 1762 417 1828 451
rect 1762 383 1778 417
rect 1812 383 1828 417
rect 1762 349 1828 383
rect 1862 485 1915 527
rect 1896 451 1915 485
rect 1862 408 1915 451
rect 1896 374 1915 408
rect 1862 357 1915 374
rect 1762 315 1778 349
rect 1812 323 1828 349
rect 1812 315 1915 323
rect 1762 299 1915 315
rect 1795 289 1915 299
rect 1610 249 1770 265
rect 1610 215 1736 249
rect 1610 199 1770 215
rect 1610 119 1644 199
rect 1804 179 1915 289
rect 1798 171 1915 179
rect 1795 165 1915 171
rect 1610 69 1644 85
rect 1678 161 1744 165
rect 1678 127 1694 161
rect 1728 127 1744 161
rect 1678 93 1744 127
rect 1678 59 1694 93
rect 1728 59 1744 93
rect 1678 17 1744 59
rect 1778 153 1915 165
rect 1778 143 1827 153
rect 1812 109 1827 143
rect 1778 53 1827 109
rect 1861 93 1915 119
rect 1861 59 1862 93
rect 1896 59 1915 93
rect 1861 17 1915 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 121 357 155 391
rect 213 153 247 187
rect 489 357 523 391
rect 581 169 600 187
rect 600 169 615 187
rect 581 153 615 169
rect 765 179 772 187
rect 772 179 799 187
rect 765 153 799 179
rect 1041 365 1075 391
rect 1041 357 1048 365
rect 1048 357 1075 365
rect 1045 235 1046 255
rect 1046 235 1079 255
rect 1045 221 1079 235
rect 1409 153 1443 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
rect 109 391 167 397
rect 109 357 121 391
rect 155 388 167 391
rect 477 391 535 397
rect 477 388 489 391
rect 155 360 489 388
rect 155 357 167 360
rect 109 351 167 357
rect 477 357 489 360
rect 523 388 535 391
rect 1029 391 1087 397
rect 1029 388 1041 391
rect 523 360 1041 388
rect 523 357 535 360
rect 477 351 535 357
rect 1029 357 1041 360
rect 1075 357 1087 391
rect 1029 351 1087 357
rect 1033 255 1091 261
rect 1033 252 1045 255
rect 584 224 1045 252
rect 584 193 627 224
rect 1033 221 1045 224
rect 1079 221 1091 255
rect 1033 215 1091 221
rect 201 187 259 193
rect 201 153 213 187
rect 247 184 259 187
rect 569 187 627 193
rect 569 184 581 187
rect 247 156 581 184
rect 247 153 259 156
rect 201 147 259 153
rect 569 153 581 156
rect 615 153 627 187
rect 569 147 627 153
rect 753 187 811 193
rect 753 153 765 187
rect 799 184 811 187
rect 1397 187 1455 193
rect 1397 184 1409 187
rect 799 156 1409 184
rect 799 153 811 156
rect 753 147 811 153
rect 1397 153 1409 156
rect 1443 153 1455 187
rect 1397 147 1455 153
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< labels >>
flabel corelocali s 1869 153 1903 187 0 FreeSans 400 0 0 0 Q
port 8 nsew
flabel corelocali s 1869 289 1903 323 0 FreeSans 400 0 0 0 Q
port 8 nsew
flabel corelocali s 1869 221 1903 255 0 FreeSans 400 0 0 0 Q
port 8 nsew
flabel corelocali s 397 289 431 323 0 FreeSans 200 0 0 0 D
port 2 nsew
flabel corelocali s 397 221 431 255 0 FreeSans 200 0 0 0 D
port 2 nsew
flabel corelocali s 29 527 63 561 3 FreeSans 400 0 0 0 VPWR
port 7 nsew
flabel corelocali s 1779 425 1813 459 0 FreeSans 400 0 0 0 Q
port 8 nsew
flabel corelocali s 1779 357 1813 391 0 FreeSans 400 0 0 0 Q
port 8 nsew
flabel corelocali s 1779 85 1813 119 0 FreeSans 400 0 0 0 Q
port 8 nsew
flabel corelocali s 765 153 799 187 0 FreeSans 400 0 0 0 SET_B
port 3 nsew
flabel corelocali s 29 289 63 323 0 FreeSans 400 0 0 0 CLK
port 1 nsew
flabel corelocali s 29 221 63 255 0 FreeSans 400 0 0 0 CLK
port 1 nsew
flabel corelocali s 29 -17 63 17 3 FreeSans 400 0 0 0 VGND
port 4 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel nbase s 46 544 46 544 3 FreeSans 400 0 0 0 VPB
port 6 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel pwell s 46 0 46 0 3 FreeSans 400 0 0 0 VNB
port 5 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
rlabel comment s 0 0 0 0 4 dfstp_2
<< properties >>
string FIXED_BBOX 0 0 1932 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2476390
string GDS_START 2460278
<< end >>
