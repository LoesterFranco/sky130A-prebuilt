magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1288 561
rect 18 375 85 527
rect 119 341 156 493
rect 190 375 256 527
rect 290 341 328 493
rect 362 367 412 527
rect 924 455 990 527
rect 1118 455 1184 527
rect 17 299 328 341
rect 17 175 68 299
rect 525 289 835 340
rect 525 265 561 289
rect 17 127 405 175
rect 197 123 405 127
rect 508 197 561 265
rect 595 197 729 255
rect 769 197 835 289
rect 899 302 1169 340
rect 899 204 965 302
rect 1007 204 1076 266
rect 1127 264 1169 302
rect 1127 204 1245 264
rect 97 17 163 93
rect 197 51 235 123
rect 269 17 335 89
rect 369 51 405 123
rect 444 17 511 89
rect 628 17 694 89
rect 838 17 912 89
rect 1203 17 1269 161
rect 0 -17 1288 17
<< obsli1 >>
rect 464 442 890 493
rect 824 421 890 442
rect 1032 421 1084 493
rect 1218 421 1269 493
rect 456 374 702 408
rect 824 376 1269 421
rect 456 335 491 374
rect 437 301 491 335
rect 437 265 474 301
rect 105 209 474 265
rect 439 161 474 209
rect 1203 307 1269 376
rect 439 123 1098 161
rect 545 51 594 123
rect 728 51 804 123
rect 1032 55 1098 123
<< metal1 >>
rect 0 496 1288 592
rect 0 -48 1288 48
<< labels >>
rlabel locali s 1007 204 1076 266 6 A1
port 1 nsew signal input
rlabel locali s 1127 264 1169 302 6 A2
port 2 nsew signal input
rlabel locali s 1127 204 1245 264 6 A2
port 2 nsew signal input
rlabel locali s 899 302 1169 340 6 A2
port 2 nsew signal input
rlabel locali s 899 204 965 302 6 A2
port 2 nsew signal input
rlabel locali s 769 197 835 289 6 B1
port 3 nsew signal input
rlabel locali s 525 289 835 340 6 B1
port 3 nsew signal input
rlabel locali s 525 265 561 289 6 B1
port 3 nsew signal input
rlabel locali s 508 197 561 265 6 B1
port 3 nsew signal input
rlabel locali s 595 197 729 255 6 C1
port 4 nsew signal input
rlabel locali s 369 51 405 123 6 X
port 5 nsew signal output
rlabel locali s 290 341 328 493 6 X
port 5 nsew signal output
rlabel locali s 197 123 405 127 6 X
port 5 nsew signal output
rlabel locali s 197 51 235 123 6 X
port 5 nsew signal output
rlabel locali s 119 341 156 493 6 X
port 5 nsew signal output
rlabel locali s 17 299 328 341 6 X
port 5 nsew signal output
rlabel locali s 17 175 68 299 6 X
port 5 nsew signal output
rlabel locali s 17 127 405 175 6 X
port 5 nsew signal output
rlabel locali s 1203 17 1269 161 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 838 17 912 89 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 628 17 694 89 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 444 17 511 89 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 269 17 335 89 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 97 17 163 93 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 1288 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1288 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1118 455 1184 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 924 455 990 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 362 367 412 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 190 375 256 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 18 375 85 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 1288 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 1288 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1288 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3934994
string GDS_START 3925934
<< end >>
