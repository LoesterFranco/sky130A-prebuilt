magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 17 199 66 323
rect 1074 323 1150 425
rect 1262 323 1338 425
rect 1450 323 1526 425
rect 1638 323 1714 425
rect 1074 289 1714 323
rect 1074 170 1160 289
rect 1204 204 1810 255
rect 1074 127 1819 170
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 17 391 69 493
rect 103 425 185 527
rect 17 357 185 391
rect 100 265 185 357
rect 235 345 277 493
rect 321 379 387 527
rect 431 345 465 493
rect 509 379 575 527
rect 619 345 653 493
rect 697 379 763 527
rect 807 345 841 493
rect 885 379 951 527
rect 995 459 1819 493
rect 995 345 1040 459
rect 235 311 1040 345
rect 1194 357 1228 459
rect 1382 357 1416 459
rect 1570 357 1604 459
rect 1758 289 1819 459
rect 100 199 1040 265
rect 100 165 149 199
rect 17 131 149 165
rect 227 131 1040 165
rect 17 51 69 131
rect 103 17 179 97
rect 227 51 261 131
rect 295 17 371 97
rect 415 51 449 131
rect 483 17 559 97
rect 603 51 637 131
rect 671 17 747 97
rect 791 51 825 131
rect 859 17 937 97
rect 971 93 1040 131
rect 971 51 1819 93
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
<< metal1 >>
rect 0 561 1840 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 0 496 1840 527
rect 0 17 1840 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
rect 0 -48 1840 -17
<< labels >>
rlabel locali s 1204 204 1810 255 6 A
port 1 nsew signal input
rlabel locali s 17 199 66 323 6 TE
port 2 nsew signal input
rlabel locali s 1638 323 1714 425 6 Z
port 3 nsew signal output
rlabel locali s 1450 323 1526 425 6 Z
port 3 nsew signal output
rlabel locali s 1262 323 1338 425 6 Z
port 3 nsew signal output
rlabel locali s 1074 323 1150 425 6 Z
port 3 nsew signal output
rlabel locali s 1074 289 1714 323 6 Z
port 3 nsew signal output
rlabel locali s 1074 170 1160 289 6 Z
port 3 nsew signal output
rlabel locali s 1074 127 1819 170 6 Z
port 3 nsew signal output
rlabel metal1 s 0 -48 1840 48 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 496 1840 592 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1840 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2071196
string GDS_START 2057916
<< end >>
