magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 167 289 301 356
rect 359 289 455 356
rect 489 303 647 356
rect 763 378 829 596
rect 963 378 1029 596
rect 763 356 1029 378
rect 763 344 1127 356
rect 993 310 1127 344
rect 993 201 1027 310
rect 798 167 1027 201
rect 798 66 848 167
rect 993 70 1027 167
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 23 383 89 649
rect 123 581 379 615
rect 123 390 173 581
rect 213 424 279 547
rect 313 458 379 581
rect 413 458 479 649
rect 513 424 579 559
rect 627 460 723 649
rect 213 390 715 424
rect 681 310 715 390
rect 863 412 929 649
rect 1063 390 1129 649
rect 681 269 959 310
rect 23 255 89 257
rect 23 221 478 255
rect 23 121 89 221
rect 123 17 190 187
rect 226 121 276 221
rect 312 17 378 187
rect 412 87 478 221
rect 514 235 959 269
rect 514 121 564 235
rect 600 87 666 201
rect 412 53 666 87
rect 712 17 762 201
rect 884 17 957 133
rect 1063 17 1129 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
rlabel locali s 359 289 455 356 6 A1
port 1 nsew signal input
rlabel locali s 167 289 301 356 6 A2
port 2 nsew signal input
rlabel locali s 489 303 647 356 6 B1
port 3 nsew signal input
rlabel locali s 993 310 1127 344 6 X
port 4 nsew signal output
rlabel locali s 993 201 1027 310 6 X
port 4 nsew signal output
rlabel locali s 993 70 1027 167 6 X
port 4 nsew signal output
rlabel locali s 963 378 1029 596 6 X
port 4 nsew signal output
rlabel locali s 798 167 1027 201 6 X
port 4 nsew signal output
rlabel locali s 798 66 848 167 6 X
port 4 nsew signal output
rlabel locali s 763 378 829 596 6 X
port 4 nsew signal output
rlabel locali s 763 356 1029 378 6 X
port 4 nsew signal output
rlabel locali s 763 344 1127 356 6 X
port 4 nsew signal output
rlabel metal1 s 0 -49 1152 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 617 1152 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1053078
string GDS_START 1043364
<< end >>
