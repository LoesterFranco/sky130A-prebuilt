magic
tech sky130A
magscale 1 2
timestamp 1601050047
<< nwell >>
rect -38 332 806 704
<< pwell >>
rect 0 0 768 49
<< scpmos >>
rect 86 404 116 572
rect 210 404 240 572
rect 536 368 566 592
rect 620 368 650 592
<< nmoslvt >>
rect 109 74 139 184
rect 199 74 229 184
rect 539 74 569 222
rect 617 74 647 222
<< ndiff >>
rect 52 146 109 184
rect 52 112 64 146
rect 98 112 109 146
rect 52 74 109 112
rect 139 146 199 184
rect 139 112 152 146
rect 186 112 199 146
rect 139 74 199 112
rect 229 146 282 184
rect 229 112 240 146
rect 274 112 282 146
rect 229 74 282 112
rect 482 124 539 222
rect 482 90 494 124
rect 528 90 539 124
rect 482 74 539 90
rect 569 74 617 222
rect 647 210 704 222
rect 647 176 658 210
rect 692 176 704 210
rect 647 120 704 176
rect 647 86 658 120
rect 692 86 704 120
rect 647 74 704 86
<< pdiff >>
rect 134 602 192 614
rect 134 572 146 602
rect 27 560 86 572
rect 27 526 39 560
rect 73 526 86 560
rect 27 450 86 526
rect 27 416 39 450
rect 73 416 86 450
rect 27 404 86 416
rect 116 568 146 572
rect 180 572 192 602
rect 180 568 210 572
rect 116 404 210 568
rect 240 450 301 572
rect 240 416 254 450
rect 288 416 301 450
rect 240 404 301 416
rect 477 580 536 592
rect 477 546 489 580
rect 523 546 536 580
rect 477 512 536 546
rect 477 478 489 512
rect 523 478 536 512
rect 477 444 536 478
rect 477 410 489 444
rect 523 410 536 444
rect 477 368 536 410
rect 566 368 620 592
rect 650 580 709 592
rect 650 546 663 580
rect 697 546 709 580
rect 650 497 709 546
rect 650 463 663 497
rect 697 463 709 497
rect 650 414 709 463
rect 650 380 663 414
rect 697 380 709 414
rect 650 368 709 380
<< ndiffc >>
rect 64 112 98 146
rect 152 112 186 146
rect 240 112 274 146
rect 494 90 528 124
rect 658 176 692 210
rect 658 86 692 120
<< pdiffc >>
rect 39 526 73 560
rect 39 416 73 450
rect 146 568 180 602
rect 254 416 288 450
rect 489 546 523 580
rect 489 478 523 512
rect 489 410 523 444
rect 663 546 697 580
rect 663 463 697 497
rect 663 380 697 414
<< poly >>
rect 86 572 116 598
rect 210 572 240 598
rect 373 586 439 602
rect 536 592 566 618
rect 620 592 650 618
rect 373 552 389 586
rect 423 552 439 586
rect 373 518 439 552
rect 373 484 389 518
rect 423 484 439 518
rect 373 468 439 484
rect 86 389 116 404
rect 210 389 240 404
rect 83 366 119 389
rect 207 366 243 389
rect 83 350 151 366
rect 83 316 101 350
rect 135 316 151 350
rect 83 300 151 316
rect 199 350 335 366
rect 199 316 217 350
rect 251 316 285 350
rect 319 316 335 350
rect 409 353 439 468
rect 536 353 566 368
rect 620 353 650 368
rect 409 323 569 353
rect 617 330 653 353
rect 199 300 335 316
rect 617 314 683 330
rect 109 184 139 300
rect 199 184 229 300
rect 374 265 569 281
rect 374 231 390 265
rect 424 237 569 265
rect 424 231 440 237
rect 374 215 440 231
rect 539 222 569 237
rect 617 280 633 314
rect 667 280 683 314
rect 617 264 683 280
rect 617 222 647 264
rect 109 48 139 74
rect 199 48 229 74
rect 539 48 569 74
rect 617 48 647 74
<< polycont >>
rect 389 552 423 586
rect 389 484 423 518
rect 101 316 135 350
rect 217 316 251 350
rect 285 316 319 350
rect 390 231 424 265
rect 633 280 667 314
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 130 602 196 649
rect 17 560 89 576
rect 17 526 39 560
rect 73 526 89 560
rect 130 568 146 602
rect 180 568 196 602
rect 130 552 196 568
rect 373 586 439 602
rect 373 552 389 586
rect 423 552 439 586
rect 17 450 89 526
rect 373 518 439 552
rect 17 416 39 450
rect 73 416 89 450
rect 17 400 89 416
rect 133 484 389 518
rect 423 484 439 518
rect 17 264 51 400
rect 133 366 167 484
rect 373 468 439 484
rect 473 580 539 649
rect 473 546 489 580
rect 523 546 539 580
rect 473 512 539 546
rect 473 478 489 512
rect 523 478 539 512
rect 237 416 254 450
rect 288 434 339 450
rect 473 444 539 478
rect 288 416 427 434
rect 237 400 427 416
rect 473 410 489 444
rect 523 410 539 444
rect 647 580 751 596
rect 647 546 663 580
rect 697 546 751 580
rect 647 497 751 546
rect 647 463 663 497
rect 697 463 751 497
rect 647 414 751 463
rect 393 376 427 400
rect 647 380 663 414
rect 697 380 751 414
rect 85 350 167 366
rect 85 316 101 350
rect 135 316 167 350
rect 85 300 167 316
rect 201 350 359 366
rect 201 316 217 350
rect 251 316 285 350
rect 319 316 359 350
rect 393 342 613 376
rect 647 364 751 380
rect 201 300 359 316
rect 492 330 613 342
rect 492 314 683 330
rect 492 280 633 314
rect 667 280 683 314
rect 374 265 440 268
rect 374 264 390 265
rect 17 231 390 264
rect 424 231 440 265
rect 17 230 440 231
rect 492 264 683 280
rect 17 146 106 230
rect 492 196 532 264
rect 717 226 751 364
rect 17 112 64 146
rect 98 112 106 146
rect 17 91 106 112
rect 140 146 197 170
rect 140 112 152 146
rect 186 112 197 146
rect 140 17 197 112
rect 231 162 532 196
rect 642 210 751 226
rect 642 176 658 210
rect 692 176 751 210
rect 231 146 290 162
rect 231 112 240 146
rect 274 112 290 146
rect 231 91 290 112
rect 478 124 544 128
rect 478 90 494 124
rect 528 90 544 124
rect 478 17 544 90
rect 642 120 751 176
rect 642 86 658 120
rect 692 86 751 120
rect 642 70 751 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel comment s 0 0 0 0 4 ebufn_1
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 703 94 737 128 0 FreeSans 340 0 0 0 Z
port 7 nsew
flabel corelocali s 703 168 737 202 0 FreeSans 340 0 0 0 Z
port 7 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 TE_B
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 768 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 2431750
string GDS_START 2425360
<< end >>
