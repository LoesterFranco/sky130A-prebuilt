magic
tech sky130A
magscale 1 2
timestamp 1604502705
<< nwell >>
rect -38 332 1094 704
<< pwell >>
rect 0 0 1056 49
<< scnmos >>
rect 121 74 151 222
rect 199 74 229 222
rect 397 74 427 222
rect 526 74 556 222
rect 612 74 642 222
rect 731 74 761 222
rect 821 74 851 222
rect 942 74 972 222
<< pmoshvt >>
rect 103 368 133 568
rect 202 368 232 568
rect 394 368 424 592
rect 484 368 514 592
rect 608 368 638 592
rect 734 368 764 592
rect 824 368 854 592
rect 924 368 954 592
<< ndiff >>
rect 71 130 121 222
rect 27 118 121 130
rect 27 84 49 118
rect 83 84 121 118
rect 27 74 121 84
rect 151 74 199 222
rect 229 177 286 222
rect 347 180 397 222
rect 229 143 240 177
rect 274 143 286 177
rect 229 97 286 143
rect 340 160 397 180
rect 340 126 352 160
rect 386 126 397 160
rect 340 107 397 126
rect 229 74 279 97
rect 347 74 397 107
rect 427 100 526 222
rect 427 74 459 100
rect 27 72 95 74
rect 442 66 459 74
rect 493 74 526 100
rect 556 188 612 222
rect 556 154 567 188
rect 601 154 612 188
rect 556 120 612 154
rect 556 86 567 120
rect 601 86 612 120
rect 556 74 612 86
rect 642 84 731 222
rect 642 74 669 84
rect 493 66 511 74
rect 442 54 511 66
rect 657 50 669 74
rect 703 74 731 84
rect 761 152 821 222
rect 761 118 772 152
rect 806 118 821 152
rect 761 74 821 118
rect 851 84 942 222
rect 851 74 879 84
rect 703 50 716 74
rect 657 38 716 50
rect 866 50 879 74
rect 913 74 942 84
rect 972 180 1022 222
rect 972 152 1029 180
rect 972 118 983 152
rect 1017 118 1029 152
rect 972 74 1029 118
rect 913 50 927 74
rect 866 38 927 50
<< pdiff >>
rect 27 582 85 594
rect 27 548 39 582
rect 73 568 85 582
rect 250 592 371 594
rect 532 598 590 610
rect 532 592 544 598
rect 250 582 394 592
rect 250 568 258 582
rect 73 548 103 568
rect 27 368 103 548
rect 133 414 202 568
rect 133 380 150 414
rect 184 380 202 414
rect 133 368 202 380
rect 232 548 258 568
rect 292 548 341 582
rect 375 548 394 582
rect 232 368 394 548
rect 424 582 484 592
rect 424 548 437 582
rect 471 548 484 582
rect 424 514 484 548
rect 424 480 437 514
rect 471 480 484 514
rect 424 446 484 480
rect 424 412 437 446
rect 471 412 484 446
rect 424 368 484 412
rect 514 564 544 592
rect 578 592 590 598
rect 656 598 716 610
rect 656 592 669 598
rect 578 564 608 592
rect 514 368 608 564
rect 638 564 669 592
rect 703 592 716 598
rect 703 564 734 592
rect 638 368 734 564
rect 764 530 824 592
rect 764 496 777 530
rect 811 496 824 530
rect 764 368 824 496
rect 854 582 924 592
rect 854 548 877 582
rect 911 548 924 582
rect 854 514 924 548
rect 854 480 877 514
rect 911 480 924 514
rect 854 368 924 480
rect 954 582 1023 592
rect 954 548 977 582
rect 1011 548 1023 582
rect 954 514 1023 548
rect 954 480 977 514
rect 1011 480 1023 514
rect 954 368 1023 480
<< ndiffc >>
rect 49 84 83 118
rect 240 143 274 177
rect 352 126 386 160
rect 459 66 493 100
rect 567 154 601 188
rect 567 86 601 120
rect 669 50 703 84
rect 772 118 806 152
rect 879 50 913 84
rect 983 118 1017 152
<< pdiffc >>
rect 39 548 73 582
rect 150 380 184 414
rect 258 548 292 582
rect 341 548 375 582
rect 437 548 471 582
rect 437 480 471 514
rect 437 412 471 446
rect 544 564 578 598
rect 669 564 703 598
rect 777 496 811 530
rect 877 548 911 582
rect 877 480 911 514
rect 977 548 1011 582
rect 977 480 1011 514
<< poly >>
rect 103 568 133 594
rect 202 568 232 594
rect 394 592 424 618
rect 484 592 514 618
rect 608 592 638 618
rect 734 592 764 618
rect 824 592 854 618
rect 924 592 954 618
rect 103 353 133 368
rect 202 353 232 368
rect 394 353 424 368
rect 484 353 514 368
rect 608 353 638 368
rect 734 353 764 368
rect 824 353 854 368
rect 924 353 954 368
rect 100 310 136 353
rect 199 336 235 353
rect 199 320 335 336
rect 85 294 151 310
rect 85 260 101 294
rect 135 260 151 294
rect 85 244 151 260
rect 121 222 151 244
rect 199 286 285 320
rect 319 286 335 320
rect 391 310 427 353
rect 481 310 517 353
rect 199 270 335 286
rect 383 294 517 310
rect 199 222 229 270
rect 383 260 399 294
rect 433 260 467 294
rect 501 274 517 294
rect 605 310 641 353
rect 731 310 767 353
rect 821 310 857 353
rect 921 336 957 353
rect 905 320 972 336
rect 605 294 671 310
rect 501 260 556 274
rect 383 244 556 260
rect 605 260 621 294
rect 655 260 671 294
rect 605 244 671 260
rect 731 294 851 310
rect 731 260 801 294
rect 835 260 851 294
rect 905 286 921 320
rect 955 286 972 320
rect 905 270 972 286
rect 731 244 851 260
rect 397 222 427 244
rect 526 222 556 244
rect 612 222 642 244
rect 731 222 761 244
rect 821 222 851 244
rect 942 222 972 270
rect 121 48 151 74
rect 199 48 229 74
rect 397 48 427 74
rect 526 48 556 74
rect 612 48 642 74
rect 731 48 761 74
rect 821 48 851 74
rect 942 48 972 74
<< polycont >>
rect 101 260 135 294
rect 285 286 319 320
rect 399 260 433 294
rect 467 260 501 294
rect 621 260 655 294
rect 801 260 835 294
rect 921 286 955 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 23 582 89 649
rect 23 548 39 582
rect 73 548 89 582
rect 23 532 89 548
rect 246 582 375 649
rect 528 598 594 649
rect 246 548 258 582
rect 292 548 341 582
rect 246 532 375 548
rect 409 582 487 596
rect 409 548 437 582
rect 471 548 487 582
rect 528 564 544 598
rect 578 564 594 598
rect 528 548 594 564
rect 652 598 927 615
rect 652 564 669 598
rect 703 582 927 598
rect 703 581 877 582
rect 703 564 720 581
rect 652 548 720 564
rect 861 548 877 581
rect 911 548 927 582
rect 409 514 487 548
rect 761 530 827 547
rect 761 514 777 530
rect 409 498 437 514
rect 17 480 437 498
rect 471 496 777 514
rect 811 496 827 530
rect 471 480 827 496
rect 861 514 927 548
rect 861 480 877 514
rect 911 480 927 514
rect 961 582 1027 649
rect 961 548 977 582
rect 1011 548 1027 582
rect 961 514 1027 548
rect 961 480 977 514
rect 1011 480 1027 514
rect 17 464 487 480
rect 17 202 51 464
rect 409 446 487 464
rect 130 414 235 430
rect 130 380 150 414
rect 184 380 235 414
rect 409 412 437 446
rect 471 412 487 446
rect 521 412 1039 446
rect 130 364 235 380
rect 521 378 555 412
rect 85 294 167 310
rect 85 260 101 294
rect 135 276 167 294
rect 85 242 127 260
rect 161 242 167 276
rect 85 236 167 242
rect 201 236 235 364
rect 269 344 555 378
rect 605 344 935 378
rect 269 320 335 344
rect 269 286 285 320
rect 319 286 335 320
rect 605 310 671 344
rect 889 336 935 344
rect 889 320 971 336
rect 269 270 335 286
rect 383 294 517 310
rect 383 260 399 294
rect 433 260 467 294
rect 501 260 517 294
rect 383 236 517 260
rect 601 294 671 310
rect 601 276 621 294
rect 601 242 607 276
rect 655 260 671 294
rect 641 242 671 260
rect 601 236 671 242
rect 785 294 851 310
rect 785 260 801 294
rect 835 260 851 294
rect 889 286 921 320
rect 955 286 971 320
rect 889 270 971 286
rect 785 236 851 260
rect 1005 236 1039 412
rect 201 202 517 236
rect 785 202 1039 236
rect 17 168 167 202
rect 23 118 99 134
rect 23 84 49 118
rect 83 84 99 118
rect 23 17 99 84
rect 133 85 167 168
rect 201 177 290 202
rect 201 143 240 177
rect 274 143 290 177
rect 551 188 617 202
rect 551 168 567 188
rect 201 127 290 143
rect 336 160 567 168
rect 336 126 352 160
rect 386 154 567 160
rect 601 168 617 188
rect 601 154 1033 168
rect 386 152 1033 154
rect 386 134 772 152
rect 386 126 402 134
rect 336 119 402 126
rect 551 120 617 134
rect 438 85 459 100
rect 133 66 459 85
rect 493 66 515 100
rect 551 86 567 120
rect 601 86 617 120
rect 756 118 772 134
rect 806 134 983 152
rect 806 118 822 134
rect 551 70 617 86
rect 653 84 720 100
rect 756 98 822 118
rect 967 118 983 134
rect 1017 118 1033 152
rect 133 51 515 66
rect 653 50 669 84
rect 703 50 720 84
rect 653 17 720 50
rect 862 84 931 100
rect 967 98 1033 118
rect 862 50 879 84
rect 913 50 931 84
rect 862 17 931 50
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 127 260 135 276
rect 135 260 161 276
rect 127 242 161 260
rect 607 260 621 276
rect 621 260 641 276
rect 607 242 641 260
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 683 1056 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 0 617 1056 649
rect 115 276 173 282
rect 115 242 127 276
rect 161 273 173 276
rect 595 276 653 282
rect 595 273 607 276
rect 161 245 607 273
rect 161 242 173 245
rect 115 236 173 242
rect 595 242 607 245
rect 641 242 653 276
rect 595 236 653 242
rect 0 17 1056 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -49 1056 -17
<< labels >>
rlabel comment s 0 0 0 0 4 xnor2_2
flabel pwell s 0 0 1056 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 0 617 1056 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 0 617 1056 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 1056 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 415 464 449 498 0 FreeSans 340 0 0 0 Y
port 7 nsew
flabel corelocali s 415 538 449 572 0 FreeSans 340 0 0 0 Y
port 7 nsew
flabel corelocali s 799 242 833 276 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 A
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 1056 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 589988
string GDS_START 581694
<< end >>
