magic
tech sky130A
magscale 1 2
timestamp 1599588232
<< locali >>
rect 120 394 186 596
rect 20 360 186 394
rect 20 226 67 360
rect 20 192 171 226
rect 121 70 171 192
rect 273 252 353 356
rect 387 290 455 356
rect 491 290 552 356
rect 654 236 739 310
rect 773 236 839 310
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 30 428 80 649
rect 226 390 276 649
rect 313 424 363 596
rect 403 458 469 649
rect 507 581 737 615
rect 507 480 557 581
rect 597 446 663 547
rect 508 424 663 446
rect 313 412 663 424
rect 703 412 737 581
rect 313 390 546 412
rect 777 378 843 596
rect 105 260 239 326
rect 35 17 85 158
rect 205 218 239 260
rect 586 344 843 378
rect 586 226 620 344
rect 404 218 620 226
rect 205 202 620 218
rect 205 184 844 202
rect 404 168 844 184
rect 207 17 312 150
rect 404 70 578 168
rect 670 17 744 134
rect 778 70 844 168
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel locali s 387 290 455 356 6 A1
port 1 nsew signal input
rlabel locali s 273 252 353 356 6 A2
port 2 nsew signal input
rlabel locali s 491 290 552 356 6 B1
port 3 nsew signal input
rlabel locali s 654 236 739 310 6 B2
port 4 nsew signal input
rlabel locali s 773 236 839 310 6 C1
port 5 nsew signal input
rlabel locali s 121 70 171 192 6 X
port 6 nsew signal output
rlabel locali s 120 394 186 596 6 X
port 6 nsew signal output
rlabel locali s 20 360 186 394 6 X
port 6 nsew signal output
rlabel locali s 20 226 67 360 6 X
port 6 nsew signal output
rlabel locali s 20 192 171 226 6 X
port 6 nsew signal output
rlabel metal1 s 0 -49 864 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 8 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 9 nsew power bidirectional
rlabel metal1 s 0 617 864 715 6 VPWR
port 10 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3514488
string GDS_START 3506170
<< end >>
