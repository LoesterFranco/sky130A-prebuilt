magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 1510 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 99 47 129 177
rect 307 47 337 177
rect 401 47 431 177
rect 495 47 525 177
rect 589 47 619 177
rect 673 47 703 177
rect 767 47 797 177
rect 861 47 891 177
rect 965 47 995 177
rect 1049 47 1079 177
rect 1143 47 1173 177
rect 1237 47 1267 177
rect 1341 47 1371 177
<< pmoshvt >>
rect 91 297 127 497
rect 185 297 221 497
rect 279 297 315 497
rect 373 297 409 497
rect 467 297 503 497
rect 675 297 711 497
rect 769 297 805 497
rect 863 297 899 497
rect 957 297 993 497
rect 1051 297 1087 497
rect 1145 297 1181 497
rect 1239 297 1275 497
rect 1333 297 1369 497
<< ndiff >>
rect 33 163 99 177
rect 33 129 45 163
rect 79 129 99 163
rect 33 95 99 129
rect 33 61 45 95
rect 79 61 99 95
rect 33 47 99 61
rect 129 163 181 177
rect 129 129 139 163
rect 173 129 181 163
rect 129 95 181 129
rect 129 61 139 95
rect 173 61 181 95
rect 129 47 181 61
rect 245 95 307 177
rect 245 61 253 95
rect 287 61 307 95
rect 245 47 307 61
rect 337 163 401 177
rect 337 129 347 163
rect 381 129 401 163
rect 337 47 401 129
rect 431 95 495 177
rect 431 61 441 95
rect 475 61 495 95
rect 431 47 495 61
rect 525 163 589 177
rect 525 129 535 163
rect 569 129 589 163
rect 525 47 589 129
rect 619 163 673 177
rect 619 129 629 163
rect 663 129 673 163
rect 619 95 673 129
rect 619 61 629 95
rect 663 61 673 95
rect 619 47 673 61
rect 703 95 767 177
rect 703 61 723 95
rect 757 61 767 95
rect 703 47 767 61
rect 797 163 861 177
rect 797 129 817 163
rect 851 129 861 163
rect 797 95 861 129
rect 797 61 817 95
rect 851 61 861 95
rect 797 47 861 61
rect 891 95 965 177
rect 891 61 911 95
rect 945 61 965 95
rect 891 47 965 61
rect 995 163 1049 177
rect 995 129 1005 163
rect 1039 129 1049 163
rect 995 95 1049 129
rect 995 61 1005 95
rect 1039 61 1049 95
rect 995 47 1049 61
rect 1079 95 1143 177
rect 1079 61 1099 95
rect 1133 61 1143 95
rect 1079 47 1143 61
rect 1173 163 1237 177
rect 1173 129 1193 163
rect 1227 129 1237 163
rect 1173 95 1237 129
rect 1173 61 1193 95
rect 1227 61 1237 95
rect 1173 47 1237 61
rect 1267 95 1341 177
rect 1267 61 1287 95
rect 1321 61 1341 95
rect 1267 47 1341 61
rect 1371 163 1423 177
rect 1371 129 1381 163
rect 1415 129 1423 163
rect 1371 95 1423 129
rect 1371 61 1381 95
rect 1415 61 1423 95
rect 1371 47 1423 61
<< pdiff >>
rect 33 477 91 497
rect 33 443 45 477
rect 79 443 91 477
rect 33 409 91 443
rect 33 375 45 409
rect 79 375 91 409
rect 33 341 91 375
rect 33 307 45 341
rect 79 307 91 341
rect 33 297 91 307
rect 127 477 185 497
rect 127 443 139 477
rect 173 443 185 477
rect 127 409 185 443
rect 127 375 139 409
rect 173 375 185 409
rect 127 297 185 375
rect 221 477 279 497
rect 221 443 233 477
rect 267 443 279 477
rect 221 409 279 443
rect 221 375 233 409
rect 267 375 279 409
rect 221 341 279 375
rect 221 307 233 341
rect 267 307 279 341
rect 221 297 279 307
rect 315 477 373 497
rect 315 443 327 477
rect 361 443 373 477
rect 315 409 373 443
rect 315 375 327 409
rect 361 375 373 409
rect 315 297 373 375
rect 409 477 467 497
rect 409 443 421 477
rect 455 443 467 477
rect 409 409 467 443
rect 409 375 421 409
rect 455 375 467 409
rect 409 341 467 375
rect 409 307 421 341
rect 455 307 467 341
rect 409 297 467 307
rect 503 477 557 497
rect 503 443 515 477
rect 549 443 557 477
rect 503 409 557 443
rect 503 375 515 409
rect 549 375 557 409
rect 503 297 557 375
rect 621 477 675 497
rect 621 443 629 477
rect 663 443 675 477
rect 621 409 675 443
rect 621 375 629 409
rect 663 375 675 409
rect 621 297 675 375
rect 711 409 769 497
rect 711 375 723 409
rect 757 375 769 409
rect 711 341 769 375
rect 711 307 723 341
rect 757 307 769 341
rect 711 297 769 307
rect 805 477 863 497
rect 805 443 817 477
rect 851 443 863 477
rect 805 409 863 443
rect 805 375 817 409
rect 851 375 863 409
rect 805 297 863 375
rect 899 409 957 497
rect 899 375 911 409
rect 945 375 957 409
rect 899 341 957 375
rect 899 307 911 341
rect 945 307 957 341
rect 899 297 957 307
rect 993 477 1051 497
rect 993 443 1005 477
rect 1039 443 1051 477
rect 993 409 1051 443
rect 993 375 1005 409
rect 1039 375 1051 409
rect 993 341 1051 375
rect 993 307 1005 341
rect 1039 307 1051 341
rect 993 297 1051 307
rect 1087 477 1145 497
rect 1087 443 1099 477
rect 1133 443 1145 477
rect 1087 409 1145 443
rect 1087 375 1099 409
rect 1133 375 1145 409
rect 1087 297 1145 375
rect 1181 477 1239 497
rect 1181 443 1193 477
rect 1227 443 1239 477
rect 1181 409 1239 443
rect 1181 375 1193 409
rect 1227 375 1239 409
rect 1181 341 1239 375
rect 1181 307 1193 341
rect 1227 307 1239 341
rect 1181 297 1239 307
rect 1275 477 1333 497
rect 1275 443 1287 477
rect 1321 443 1333 477
rect 1275 409 1333 443
rect 1275 375 1287 409
rect 1321 375 1333 409
rect 1275 297 1333 375
rect 1369 477 1427 497
rect 1369 443 1381 477
rect 1415 443 1427 477
rect 1369 409 1427 443
rect 1369 375 1381 409
rect 1415 375 1427 409
rect 1369 341 1427 375
rect 1369 307 1381 341
rect 1415 307 1427 341
rect 1369 297 1427 307
<< ndiffc >>
rect 45 129 79 163
rect 45 61 79 95
rect 139 129 173 163
rect 139 61 173 95
rect 253 61 287 95
rect 347 129 381 163
rect 441 61 475 95
rect 535 129 569 163
rect 629 129 663 163
rect 629 61 663 95
rect 723 61 757 95
rect 817 129 851 163
rect 817 61 851 95
rect 911 61 945 95
rect 1005 129 1039 163
rect 1005 61 1039 95
rect 1099 61 1133 95
rect 1193 129 1227 163
rect 1193 61 1227 95
rect 1287 61 1321 95
rect 1381 129 1415 163
rect 1381 61 1415 95
<< pdiffc >>
rect 45 443 79 477
rect 45 375 79 409
rect 45 307 79 341
rect 139 443 173 477
rect 139 375 173 409
rect 233 443 267 477
rect 233 375 267 409
rect 233 307 267 341
rect 327 443 361 477
rect 327 375 361 409
rect 421 443 455 477
rect 421 375 455 409
rect 421 307 455 341
rect 515 443 549 477
rect 515 375 549 409
rect 629 443 663 477
rect 629 375 663 409
rect 723 375 757 409
rect 723 307 757 341
rect 817 443 851 477
rect 817 375 851 409
rect 911 375 945 409
rect 911 307 945 341
rect 1005 443 1039 477
rect 1005 375 1039 409
rect 1005 307 1039 341
rect 1099 443 1133 477
rect 1099 375 1133 409
rect 1193 443 1227 477
rect 1193 375 1227 409
rect 1193 307 1227 341
rect 1287 443 1321 477
rect 1287 375 1321 409
rect 1381 443 1415 477
rect 1381 375 1415 409
rect 1381 307 1415 341
<< poly >>
rect 91 497 127 523
rect 185 497 221 523
rect 279 497 315 523
rect 373 497 409 523
rect 467 497 503 523
rect 675 497 711 523
rect 769 497 805 523
rect 863 497 899 523
rect 957 497 993 523
rect 1051 497 1087 523
rect 1145 497 1181 523
rect 1239 497 1275 523
rect 1333 497 1369 523
rect 91 282 127 297
rect 185 282 221 297
rect 279 282 315 297
rect 373 282 409 297
rect 467 282 503 297
rect 675 282 711 297
rect 769 282 805 297
rect 863 282 899 297
rect 957 282 993 297
rect 1051 282 1087 297
rect 1145 282 1181 297
rect 1239 282 1275 297
rect 1333 282 1369 297
rect 89 265 129 282
rect 42 249 129 265
rect 42 215 52 249
rect 86 215 129 249
rect 42 199 129 215
rect 183 265 223 282
rect 277 265 317 282
rect 371 265 411 282
rect 465 265 505 282
rect 673 265 713 282
rect 767 265 807 282
rect 861 265 901 282
rect 955 265 995 282
rect 183 249 619 265
rect 183 215 199 249
rect 233 215 277 249
rect 311 215 355 249
rect 389 215 433 249
rect 467 215 619 249
rect 183 199 619 215
rect 99 177 129 199
rect 307 177 337 199
rect 401 177 431 199
rect 495 177 525 199
rect 589 177 619 199
rect 673 249 995 265
rect 673 215 689 249
rect 723 215 767 249
rect 801 215 845 249
rect 879 215 923 249
rect 957 215 995 249
rect 673 199 995 215
rect 673 177 703 199
rect 767 177 797 199
rect 861 177 891 199
rect 965 177 995 199
rect 1049 265 1089 282
rect 1143 265 1183 282
rect 1237 265 1277 282
rect 1331 265 1371 282
rect 1049 249 1371 265
rect 1049 215 1059 249
rect 1093 215 1137 249
rect 1171 215 1215 249
rect 1249 215 1293 249
rect 1327 215 1371 249
rect 1049 199 1371 215
rect 1049 177 1079 199
rect 1143 177 1173 199
rect 1237 177 1267 199
rect 1341 177 1371 199
rect 99 21 129 47
rect 307 21 337 47
rect 401 21 431 47
rect 495 21 525 47
rect 589 21 619 47
rect 673 21 703 47
rect 767 21 797 47
rect 861 21 891 47
rect 965 21 995 47
rect 1049 21 1079 47
rect 1143 21 1173 47
rect 1237 21 1267 47
rect 1341 21 1371 47
<< polycont >>
rect 52 215 86 249
rect 199 215 233 249
rect 277 215 311 249
rect 355 215 389 249
rect 433 215 467 249
rect 689 215 723 249
rect 767 215 801 249
rect 845 215 879 249
rect 923 215 957 249
rect 1059 215 1093 249
rect 1137 215 1171 249
rect 1215 215 1249 249
rect 1293 215 1327 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 29 477 95 487
rect 29 443 45 477
rect 79 443 95 477
rect 29 409 95 443
rect 29 375 45 409
rect 79 375 95 409
rect 29 341 95 375
rect 139 477 173 527
rect 139 409 173 443
rect 139 359 173 375
rect 207 477 275 493
rect 207 443 233 477
rect 267 443 275 477
rect 207 409 275 443
rect 207 375 233 409
rect 267 375 275 409
rect 29 307 45 341
rect 79 325 95 341
rect 207 341 275 375
rect 319 477 369 527
rect 319 443 327 477
rect 361 443 369 477
rect 319 409 369 443
rect 319 375 327 409
rect 361 375 369 409
rect 319 359 369 375
rect 413 477 463 493
rect 413 443 421 477
rect 455 443 463 477
rect 413 409 463 443
rect 413 375 421 409
rect 455 375 463 409
rect 79 307 170 325
rect 29 291 170 307
rect 207 307 233 341
rect 267 325 275 341
rect 413 341 463 375
rect 507 477 557 527
rect 507 443 515 477
rect 549 443 557 477
rect 507 409 557 443
rect 507 375 515 409
rect 549 375 557 409
rect 507 359 557 375
rect 605 477 1047 493
rect 605 443 629 477
rect 663 459 817 477
rect 663 443 671 459
rect 605 409 671 443
rect 809 443 817 459
rect 851 459 1005 477
rect 851 443 859 459
rect 605 375 629 409
rect 663 375 671 409
rect 605 359 671 375
rect 715 409 765 425
rect 715 375 723 409
rect 757 375 765 409
rect 413 325 421 341
rect 267 307 421 325
rect 455 325 463 341
rect 715 341 765 375
rect 809 409 859 443
rect 997 443 1005 459
rect 1039 443 1047 477
rect 809 375 817 409
rect 851 375 859 409
rect 809 359 859 375
rect 903 409 953 425
rect 903 375 911 409
rect 945 375 953 409
rect 715 325 723 341
rect 455 307 723 325
rect 757 325 765 341
rect 903 341 953 375
rect 903 325 911 341
rect 757 307 911 325
rect 945 307 953 341
rect 207 291 953 307
rect 997 409 1047 443
rect 997 375 1005 409
rect 1039 375 1047 409
rect 997 341 1047 375
rect 1091 477 1141 527
rect 1091 443 1099 477
rect 1133 443 1141 477
rect 1091 409 1141 443
rect 1091 375 1099 409
rect 1133 375 1141 409
rect 1091 359 1141 375
rect 1185 477 1235 493
rect 1185 443 1193 477
rect 1227 443 1235 477
rect 1185 409 1235 443
rect 1185 375 1193 409
rect 1227 375 1235 409
rect 997 307 1005 341
rect 1039 325 1047 341
rect 1185 341 1235 375
rect 1279 477 1329 527
rect 1279 443 1287 477
rect 1321 443 1329 477
rect 1279 409 1329 443
rect 1279 375 1287 409
rect 1321 375 1329 409
rect 1279 359 1329 375
rect 1373 477 1423 493
rect 1373 443 1381 477
rect 1415 443 1423 477
rect 1373 409 1423 443
rect 1373 375 1381 409
rect 1415 375 1423 409
rect 1185 325 1193 341
rect 1039 307 1193 325
rect 1227 325 1235 341
rect 1373 341 1423 375
rect 1373 325 1381 341
rect 1227 307 1381 325
rect 1415 307 1423 341
rect 997 291 1423 307
rect 136 257 170 291
rect 539 289 953 291
rect 17 249 102 257
rect 17 215 52 249
rect 86 215 102 249
rect 136 249 505 257
rect 136 215 199 249
rect 233 215 277 249
rect 311 215 355 249
rect 389 215 433 249
rect 467 215 505 249
rect 539 215 639 289
rect 673 249 995 255
rect 673 215 689 249
rect 723 215 767 249
rect 801 215 845 249
rect 879 215 923 249
rect 957 215 995 249
rect 1029 249 1450 257
rect 1029 215 1059 249
rect 1093 215 1137 249
rect 1171 215 1215 249
rect 1249 215 1293 249
rect 1327 215 1450 249
rect 136 179 189 215
rect 45 163 79 179
rect 45 95 79 129
rect 45 17 79 61
rect 113 163 189 179
rect 539 163 585 215
rect 113 129 139 163
rect 173 129 189 163
rect 304 129 347 163
rect 381 129 535 163
rect 569 129 585 163
rect 629 163 1431 181
rect 663 145 817 163
rect 663 129 679 145
rect 113 95 189 129
rect 629 95 679 129
rect 791 129 817 145
rect 851 145 1005 163
rect 851 129 867 145
rect 113 61 139 95
rect 173 61 189 95
rect 236 61 253 95
rect 287 61 441 95
rect 475 61 629 95
rect 663 61 679 95
rect 723 95 757 111
rect 113 58 189 61
rect 723 17 757 61
rect 791 95 867 129
rect 979 129 1005 145
rect 1039 145 1193 163
rect 1039 129 1055 145
rect 791 61 817 95
rect 851 61 867 95
rect 791 51 867 61
rect 911 95 945 111
rect 911 17 945 61
rect 979 95 1055 129
rect 1167 129 1193 145
rect 1227 145 1381 163
rect 1227 129 1243 145
rect 979 61 1005 95
rect 1039 61 1055 95
rect 979 51 1055 61
rect 1099 95 1133 111
rect 1099 17 1133 61
rect 1167 95 1243 129
rect 1355 129 1381 145
rect 1415 129 1431 163
rect 1167 61 1193 95
rect 1227 61 1243 95
rect 1167 51 1243 61
rect 1287 95 1321 111
rect 1287 17 1321 61
rect 1355 95 1431 129
rect 1355 61 1381 95
rect 1415 61 1431 95
rect 1355 51 1431 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< labels >>
flabel corelocali s 539 289 573 323 0 FreeSans 400 0 0 0 Y
port 8 nsew
flabel corelocali s 75 238 75 238 0 FreeSans 400 0 0 0 B1_N
port 3 nsew
flabel corelocali s 1058 238 1058 238 0 FreeSans 400 0 0 0 A1
port 1 nsew
flabel corelocali s 782 238 782 238 0 FreeSans 400 0 0 0 A2
port 2 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
rlabel comment s 0 0 0 0 4 o21bai_4
<< properties >>
string FIXED_BBOX 0 0 1472 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1047426
string GDS_START 1036122
<< end >>
