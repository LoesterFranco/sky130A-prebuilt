magic
tech sky130A
magscale 1 2
timestamp 1604502729
<< locali >>
rect 25 200 103 434
rect 409 328 455 356
rect 359 262 455 328
rect 1945 377 2085 596
rect 2033 226 2085 377
rect 2033 70 2099 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 21 504 71 649
rect 111 504 177 596
rect 217 530 267 649
rect 397 536 463 649
rect 877 548 943 649
rect 137 496 177 504
rect 602 502 652 545
rect 301 496 652 502
rect 137 468 652 496
rect 692 514 758 545
rect 692 480 1050 514
rect 137 462 335 468
rect 137 166 171 462
rect 602 446 652 468
rect 205 424 257 428
rect 205 390 223 424
rect 205 226 257 390
rect 291 362 373 428
rect 503 378 553 434
rect 602 412 751 446
rect 291 228 325 362
rect 503 344 683 378
rect 573 312 683 344
rect 489 228 539 310
rect 291 194 539 228
rect 26 132 171 166
rect 26 74 92 132
rect 206 17 256 166
rect 291 70 368 194
rect 573 160 607 312
rect 717 278 751 412
rect 402 17 468 160
rect 502 100 607 160
rect 641 244 751 278
rect 641 134 691 244
rect 785 210 819 480
rect 923 464 1050 480
rect 725 134 819 210
rect 853 215 889 425
rect 923 315 957 464
rect 991 424 1057 430
rect 1025 390 1057 424
rect 991 359 1057 390
rect 1096 349 1162 649
rect 1196 373 1262 551
rect 1296 495 1527 561
rect 923 249 1130 315
rect 1196 226 1230 373
rect 1296 337 1330 495
rect 1164 215 1230 226
rect 853 181 1230 215
rect 853 113 1130 147
rect 1164 133 1230 181
rect 1264 303 1330 337
rect 1264 169 1298 303
rect 1393 269 1459 461
rect 1493 337 1527 495
rect 1561 489 1627 649
rect 1664 489 1737 581
rect 1561 424 1669 451
rect 1561 390 1567 424
rect 1601 390 1669 424
rect 1561 384 1669 390
rect 1703 405 1737 489
rect 1771 439 1837 649
rect 1703 371 1838 405
rect 1493 303 1770 337
rect 1704 271 1770 303
rect 1338 203 1484 269
rect 1518 237 1584 269
rect 1804 237 1838 371
rect 1877 343 1911 581
rect 1877 277 1987 343
rect 1518 203 1838 237
rect 1264 119 1416 169
rect 853 100 887 113
rect 502 66 887 100
rect 1096 85 1130 113
rect 1450 85 1484 203
rect 983 17 1062 79
rect 1096 51 1484 85
rect 1549 17 1615 169
rect 1723 77 1789 203
rect 1835 17 1885 169
rect 1921 70 1987 277
rect 2119 364 2185 649
rect 2135 17 2185 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 223 390 257 424
rect 991 390 1025 424
rect 1567 390 1601 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
<< metal1 >>
rect 0 683 2208 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 0 617 2208 649
rect 211 424 269 430
rect 211 390 223 424
rect 257 421 269 424
rect 979 424 1037 430
rect 979 421 991 424
rect 257 393 991 421
rect 257 390 269 393
rect 211 384 269 390
rect 979 390 991 393
rect 1025 421 1037 424
rect 1555 424 1613 430
rect 1555 421 1567 424
rect 1025 393 1567 421
rect 1025 390 1037 393
rect 979 384 1037 390
rect 1555 390 1567 393
rect 1601 390 1613 424
rect 1555 384 1613 390
rect 0 17 2208 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
rect 0 -49 2208 -17
<< labels >>
rlabel locali s 25 200 103 434 6 D
port 1 nsew signal input
rlabel locali s 2033 226 2085 377 6 Q
port 2 nsew signal output
rlabel locali s 2033 70 2099 226 6 Q
port 2 nsew signal output
rlabel locali s 1945 377 2085 596 6 Q
port 2 nsew signal output
rlabel metal1 s 1555 421 1613 430 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 1555 384 1613 393 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 979 421 1037 430 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 979 384 1037 393 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 211 421 269 430 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 211 393 1613 421 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 211 384 269 393 6 RESET_B
port 3 nsew signal input
rlabel locali s 409 328 455 356 6 CLK
port 4 nsew clock input
rlabel locali s 359 262 455 328 6 CLK
port 4 nsew clock input
rlabel metal1 s 0 -49 2208 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 617 2208 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2208 666
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 2960208
string GDS_START 2943866
<< end >>
