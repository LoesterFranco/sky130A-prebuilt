magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 90 93 120 177
rect 311 47 341 177
rect 405 47 435 177
rect 489 47 519 177
rect 593 47 623 177
rect 677 47 707 177
rect 781 47 811 177
<< pmoshvt >>
rect 82 297 118 381
rect 189 297 225 497
rect 283 297 319 497
rect 491 297 527 497
rect 585 297 621 497
rect 679 297 715 497
rect 773 297 809 497
<< ndiff >>
rect 28 149 90 177
rect 28 115 36 149
rect 70 115 90 149
rect 28 93 90 115
rect 120 149 172 177
rect 120 115 130 149
rect 164 115 172 149
rect 120 93 172 115
rect 226 163 311 177
rect 226 129 234 163
rect 268 129 311 163
rect 226 95 311 129
rect 226 61 234 95
rect 268 61 311 95
rect 226 47 311 61
rect 341 163 405 177
rect 341 129 351 163
rect 385 129 405 163
rect 341 47 405 129
rect 435 163 489 177
rect 435 129 445 163
rect 479 129 489 163
rect 435 95 489 129
rect 435 61 445 95
rect 479 61 489 95
rect 435 47 489 61
rect 519 95 593 177
rect 519 61 539 95
rect 573 61 593 95
rect 519 47 593 61
rect 623 163 677 177
rect 623 129 633 163
rect 667 129 677 163
rect 623 95 677 129
rect 623 61 633 95
rect 667 61 677 95
rect 623 47 677 61
rect 707 95 781 177
rect 707 61 727 95
rect 761 61 781 95
rect 707 47 781 61
rect 811 163 867 177
rect 811 129 821 163
rect 855 129 867 163
rect 811 95 867 129
rect 811 61 821 95
rect 855 61 867 95
rect 811 47 867 61
<< pdiff >>
rect 135 477 189 497
rect 135 443 143 477
rect 177 443 189 477
rect 135 409 189 443
rect 135 381 143 409
rect 28 362 82 381
rect 28 328 36 362
rect 70 328 82 362
rect 28 297 82 328
rect 118 375 143 381
rect 177 375 189 409
rect 118 297 189 375
rect 225 477 283 497
rect 225 443 237 477
rect 271 443 283 477
rect 225 409 283 443
rect 225 375 237 409
rect 271 375 283 409
rect 225 341 283 375
rect 225 307 237 341
rect 271 307 283 341
rect 225 297 283 307
rect 319 477 373 497
rect 319 443 331 477
rect 365 443 373 477
rect 319 409 373 443
rect 319 375 331 409
rect 365 375 373 409
rect 319 297 373 375
rect 437 477 491 497
rect 437 443 445 477
rect 479 443 491 477
rect 437 409 491 443
rect 437 375 445 409
rect 479 375 491 409
rect 437 297 491 375
rect 527 409 585 497
rect 527 375 539 409
rect 573 375 585 409
rect 527 341 585 375
rect 527 307 539 341
rect 573 307 585 341
rect 527 297 585 307
rect 621 477 679 497
rect 621 443 633 477
rect 667 443 679 477
rect 621 409 679 443
rect 621 375 633 409
rect 667 375 679 409
rect 621 341 679 375
rect 621 307 633 341
rect 667 307 679 341
rect 621 297 679 307
rect 715 485 773 497
rect 715 451 727 485
rect 761 451 773 485
rect 715 417 773 451
rect 715 383 727 417
rect 761 383 773 417
rect 715 297 773 383
rect 809 477 867 497
rect 809 443 821 477
rect 855 443 867 477
rect 809 409 867 443
rect 809 375 821 409
rect 855 375 867 409
rect 809 341 867 375
rect 809 307 821 341
rect 855 307 867 341
rect 809 297 867 307
<< ndiffc >>
rect 36 115 70 149
rect 130 115 164 149
rect 234 129 268 163
rect 234 61 268 95
rect 351 129 385 163
rect 445 129 479 163
rect 445 61 479 95
rect 539 61 573 95
rect 633 129 667 163
rect 633 61 667 95
rect 727 61 761 95
rect 821 129 855 163
rect 821 61 855 95
<< pdiffc >>
rect 143 443 177 477
rect 36 328 70 362
rect 143 375 177 409
rect 237 443 271 477
rect 237 375 271 409
rect 237 307 271 341
rect 331 443 365 477
rect 331 375 365 409
rect 445 443 479 477
rect 445 375 479 409
rect 539 375 573 409
rect 539 307 573 341
rect 633 443 667 477
rect 633 375 667 409
rect 633 307 667 341
rect 727 451 761 485
rect 727 383 761 417
rect 821 443 855 477
rect 821 375 855 409
rect 821 307 855 341
<< poly >>
rect 189 497 225 523
rect 283 497 319 523
rect 491 497 527 523
rect 585 497 621 523
rect 679 497 715 523
rect 773 497 809 523
rect 82 381 118 407
rect 82 282 118 297
rect 189 282 225 297
rect 283 282 319 297
rect 491 282 527 297
rect 585 282 621 297
rect 679 282 715 297
rect 773 282 809 297
rect 80 265 120 282
rect 35 249 120 265
rect 35 215 54 249
rect 88 215 120 249
rect 35 199 120 215
rect 187 265 227 282
rect 281 265 321 282
rect 489 265 529 282
rect 583 265 623 282
rect 187 249 435 265
rect 187 215 218 249
rect 252 215 435 249
rect 187 199 435 215
rect 90 177 120 199
rect 311 177 341 199
rect 405 177 435 199
rect 489 249 623 265
rect 489 215 539 249
rect 573 215 623 249
rect 489 199 623 215
rect 489 177 519 199
rect 593 177 623 199
rect 677 265 717 282
rect 771 265 811 282
rect 677 249 811 265
rect 677 215 738 249
rect 772 215 811 249
rect 677 199 811 215
rect 677 177 707 199
rect 781 177 811 199
rect 90 67 120 93
rect 311 21 341 47
rect 405 21 435 47
rect 489 21 519 47
rect 593 21 623 47
rect 677 21 707 47
rect 781 21 811 47
<< polycont >>
rect 54 215 88 249
rect 218 215 252 249
rect 539 215 573 249
rect 738 215 772 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 127 477 193 527
rect 127 443 143 477
rect 177 443 193 477
rect 127 409 193 443
rect 36 362 70 383
rect 127 375 143 409
rect 177 375 193 409
rect 237 477 271 493
rect 237 409 271 443
rect 237 341 271 375
rect 324 477 374 527
rect 324 443 331 477
rect 365 443 374 477
rect 324 409 374 443
rect 324 375 331 409
rect 365 375 374 409
rect 324 359 374 375
rect 421 477 667 493
rect 421 443 445 477
rect 479 459 633 477
rect 479 443 487 459
rect 421 409 487 443
rect 421 375 445 409
rect 479 375 487 409
rect 421 359 487 375
rect 531 409 580 425
rect 531 375 539 409
rect 573 375 580 409
rect 70 328 183 333
rect 36 299 183 328
rect 17 249 96 265
rect 17 215 54 249
rect 88 215 96 249
rect 17 199 96 215
rect 130 249 183 299
rect 531 341 580 375
rect 531 323 539 341
rect 271 307 539 323
rect 573 307 580 341
rect 237 289 580 307
rect 633 409 667 443
rect 633 341 667 375
rect 701 485 777 527
rect 701 451 727 485
rect 761 451 777 485
rect 701 417 777 451
rect 701 383 727 417
rect 761 383 777 417
rect 701 367 777 383
rect 821 477 876 493
rect 855 443 876 477
rect 821 409 876 443
rect 855 375 876 409
rect 821 341 876 375
rect 667 307 821 333
rect 855 307 876 341
rect 633 291 876 307
rect 130 215 218 249
rect 252 215 268 249
rect 36 149 70 165
rect 36 17 70 115
rect 130 149 164 215
rect 130 89 164 115
rect 212 163 268 181
rect 212 129 234 163
rect 302 163 401 289
rect 435 249 678 255
rect 435 215 539 249
rect 573 215 678 249
rect 722 249 891 255
rect 722 215 738 249
rect 772 215 891 249
rect 302 129 351 163
rect 385 129 401 163
rect 445 163 876 181
rect 479 145 633 163
rect 479 129 495 145
rect 212 95 268 129
rect 445 95 495 129
rect 607 129 633 145
rect 667 145 821 163
rect 667 129 683 145
rect 212 61 234 95
rect 268 61 445 95
rect 479 61 495 95
rect 212 51 495 61
rect 539 95 573 111
rect 539 17 573 61
rect 607 95 683 129
rect 795 129 821 145
rect 855 129 876 163
rect 607 61 633 95
rect 667 61 683 95
rect 607 51 683 61
rect 727 95 761 111
rect 727 17 761 61
rect 795 95 876 129
rect 795 61 821 95
rect 855 61 876 95
rect 795 53 876 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel corelocali s 72 238 72 238 0 FreeSans 200 0 0 0 B1_N
port 3 nsew
flabel corelocali s 355 277 355 277 0 FreeSans 400 0 0 0 Y
port 8 nsew
flabel corelocali s 539 221 573 255 0 FreeSans 400 180 0 0 A2
port 2 nsew
flabel corelocali s 743 221 777 255 0 FreeSans 400 180 0 0 A1
port 1 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
rlabel comment s 0 0 0 0 4 o21bai_2
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1054894
string GDS_START 1047486
<< end >>
