magic
tech sky130A
magscale 1 2
timestamp 1601050088
<< locali >>
rect 85 196 165 398
rect 307 264 373 356
rect 889 236 957 302
rect 991 236 1074 349
rect 1291 236 1415 310
rect 3013 430 3057 596
rect 3194 430 3237 596
rect 3013 364 3335 430
rect 3033 268 3335 364
rect 3015 218 3335 268
rect 3015 112 3065 218
rect 3199 115 3240 218
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3360 683
rect 17 492 99 596
rect 207 526 257 649
rect 291 581 461 615
rect 291 492 325 581
rect 17 458 325 492
rect 17 162 51 458
rect 359 424 393 547
rect 427 492 461 581
rect 495 526 545 649
rect 647 492 697 595
rect 427 458 697 492
rect 199 390 473 424
rect 199 230 265 390
rect 423 304 473 390
rect 507 304 611 370
rect 663 269 697 458
rect 570 235 697 269
rect 731 581 960 615
rect 731 459 787 581
rect 199 196 370 230
rect 17 68 110 162
rect 208 17 274 162
rect 320 109 370 196
rect 406 17 472 201
rect 570 109 636 235
rect 731 201 765 459
rect 821 451 892 547
rect 926 485 960 581
rect 994 519 1044 649
rect 1146 501 1212 587
rect 1252 535 1318 649
rect 1522 535 1588 649
rect 1631 501 1766 596
rect 1800 504 1872 596
rect 1992 546 2058 649
rect 2199 546 2265 649
rect 1146 485 1665 501
rect 926 467 1665 485
rect 926 451 1240 467
rect 821 417 855 451
rect 670 135 765 201
rect 799 383 1172 417
rect 799 202 855 383
rect 1116 283 1172 383
rect 1206 249 1240 451
rect 1342 357 1498 433
rect 1111 215 1240 249
rect 799 121 917 202
rect 799 51 855 121
rect 953 17 1019 202
rect 1111 121 1177 215
rect 1449 202 1483 357
rect 1544 330 1578 467
rect 1699 433 1766 467
rect 1612 399 1766 433
rect 1612 364 1733 399
rect 1544 296 1665 330
rect 1222 17 1272 181
rect 1308 168 1483 202
rect 1308 70 1374 168
rect 1419 17 1485 134
rect 1521 85 1571 226
rect 1615 119 1665 296
rect 1699 85 1733 364
rect 1800 360 1834 504
rect 1906 478 2459 512
rect 1906 466 1940 478
rect 1868 400 1940 466
rect 2095 394 2185 444
rect 1767 326 2117 360
rect 1767 119 1801 326
rect 2051 308 2117 326
rect 2151 306 2185 394
rect 1943 274 2009 281
rect 2151 274 2295 306
rect 1835 206 1901 251
rect 1943 240 2295 274
rect 2337 272 2391 360
rect 2425 351 2459 478
rect 2493 385 2579 596
rect 2667 530 2775 649
rect 2809 470 2879 596
rect 2631 436 2879 470
rect 2631 419 2697 436
rect 2745 385 2811 398
rect 2545 351 2811 385
rect 2425 306 2511 351
rect 2553 272 2619 317
rect 1835 172 2086 206
rect 1835 85 1901 172
rect 1521 51 1901 85
rect 1968 17 2018 138
rect 2052 85 2086 172
rect 2120 119 2154 240
rect 2337 238 2619 272
rect 2337 206 2371 238
rect 2188 172 2371 206
rect 2653 204 2811 351
rect 2407 198 2811 204
rect 2188 85 2222 172
rect 2407 170 2687 198
rect 2745 196 2811 198
rect 2845 356 2879 436
rect 2913 390 2979 649
rect 3093 464 3159 649
rect 3273 464 3339 649
rect 2845 310 2951 356
rect 2052 51 2222 85
rect 2256 17 2306 138
rect 2407 70 2473 170
rect 2845 162 2879 310
rect 2571 17 2767 136
rect 2801 70 2879 162
rect 2913 17 2979 268
rect 3099 17 3165 184
rect 3274 17 3340 184
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3360 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 3199 649 3233 683
rect 3295 649 3329 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
<< metal1 >>
rect 0 683 3360 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3360 683
rect 0 617 3360 649
rect 0 17 3360 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3360 17
rect 0 -49 3360 -17
<< obsm1 >>
rect 499 347 557 356
rect 2899 347 2957 356
rect 499 319 2957 347
rect 499 310 557 319
rect 2899 310 2957 319
<< labels >>
rlabel locali s 85 196 165 398 6 D
port 1 nsew signal input
rlabel locali s 307 264 373 356 6 DE
port 2 nsew signal input
rlabel locali s 3199 115 3240 218 6 Q
port 3 nsew signal output
rlabel locali s 3194 430 3237 596 6 Q
port 3 nsew signal output
rlabel locali s 3033 268 3335 364 6 Q
port 3 nsew signal output
rlabel locali s 3015 218 3335 268 6 Q
port 3 nsew signal output
rlabel locali s 3015 112 3065 218 6 Q
port 3 nsew signal output
rlabel locali s 3013 430 3057 596 6 Q
port 3 nsew signal output
rlabel locali s 3013 364 3335 430 6 Q
port 3 nsew signal output
rlabel locali s 991 236 1074 349 6 SCD
port 4 nsew signal input
rlabel locali s 889 236 957 302 6 SCE
port 5 nsew signal input
rlabel locali s 1291 236 1415 310 6 CLK
port 6 nsew clock input
rlabel metal1 s 0 -49 3360 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 617 3360 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 3360 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 492310
string GDS_START 469782
<< end >>
