magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 736 561
rect 17 293 76 527
rect 110 367 198 493
rect 110 259 172 367
rect 233 357 296 527
rect 17 215 172 259
rect 17 17 76 181
rect 110 165 172 215
rect 398 265 438 425
rect 274 199 352 255
rect 389 199 438 265
rect 478 199 528 425
rect 651 367 718 527
rect 571 199 651 265
rect 110 53 198 165
rect 232 17 322 165
rect 424 17 508 97
rect 0 -17 736 17
<< obsli1 >>
rect 330 459 616 493
rect 330 323 364 459
rect 206 289 364 323
rect 206 199 240 289
rect 566 333 616 459
rect 566 299 719 333
rect 685 165 719 299
rect 356 131 588 165
rect 356 51 390 131
rect 542 51 588 131
rect 622 51 719 165
<< metal1 >>
rect 0 496 736 592
rect 0 -48 736 48
<< labels >>
rlabel locali s 274 199 352 255 6 A1
port 1 nsew signal input
rlabel locali s 398 265 438 425 6 A2
port 2 nsew signal input
rlabel locali s 389 199 438 265 6 A2
port 2 nsew signal input
rlabel locali s 478 199 528 425 6 A3
port 3 nsew signal input
rlabel locali s 571 199 651 265 6 B1
port 4 nsew signal input
rlabel locali s 110 367 198 493 6 X
port 5 nsew signal output
rlabel locali s 110 259 172 367 6 X
port 5 nsew signal output
rlabel locali s 110 165 172 215 6 X
port 5 nsew signal output
rlabel locali s 110 53 198 165 6 X
port 5 nsew signal output
rlabel locali s 17 215 172 259 6 X
port 5 nsew signal output
rlabel locali s 424 17 508 97 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 232 17 322 165 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 17 17 76 181 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 736 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 736 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 651 367 718 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 233 357 296 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 17 293 76 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 736 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 736 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 822864
string GDS_START 815598
<< end >>
