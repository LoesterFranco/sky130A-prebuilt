magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 506 347 558 492
rect 698 347 750 492
rect 890 347 942 492
rect 1082 347 1134 492
rect 1271 347 1323 492
rect 1463 347 1515 492
rect 1655 347 1707 492
rect 506 344 1707 347
rect 1849 344 1907 492
rect 506 299 2005 344
rect 17 153 80 265
rect 1752 181 2005 299
rect 506 147 2005 181
rect 506 56 558 147
rect 698 56 750 147
rect 890 56 942 147
rect 1069 56 1134 147
rect 1271 56 1323 147
rect 1463 56 1515 147
rect 1655 56 1707 147
rect 1849 56 1901 147
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 19 365 78 527
rect 124 265 173 493
rect 218 365 270 527
rect 410 526 1805 527
rect 316 265 366 492
rect 410 367 462 526
rect 602 381 654 526
rect 794 381 846 526
rect 986 381 1038 526
rect 1178 381 1227 526
rect 1370 381 1419 526
rect 1562 381 1611 526
rect 1754 381 1805 526
rect 1951 378 2005 527
rect 124 215 1708 265
rect 17 17 78 119
rect 124 53 174 215
rect 218 17 270 122
rect 316 53 366 215
rect 410 17 462 129
rect 602 17 654 113
rect 794 17 846 113
rect 986 17 1035 113
rect 1178 17 1227 113
rect 1369 17 1419 113
rect 1561 17 1611 113
rect 1753 17 1805 113
rect 1945 17 2005 113
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
<< metal1 >>
rect 0 561 2024 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 0 496 2024 527
rect 0 17 2024 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
rect 0 -48 2024 -17
<< labels >>
rlabel locali s 17 153 80 265 6 A
port 1 nsew signal input
rlabel locali s 1849 344 1907 492 6 X
port 2 nsew signal output
rlabel locali s 1849 56 1901 147 6 X
port 2 nsew signal output
rlabel locali s 1752 181 2005 299 6 X
port 2 nsew signal output
rlabel locali s 1655 347 1707 492 6 X
port 2 nsew signal output
rlabel locali s 1655 56 1707 147 6 X
port 2 nsew signal output
rlabel locali s 1463 347 1515 492 6 X
port 2 nsew signal output
rlabel locali s 1463 56 1515 147 6 X
port 2 nsew signal output
rlabel locali s 1271 347 1323 492 6 X
port 2 nsew signal output
rlabel locali s 1271 56 1323 147 6 X
port 2 nsew signal output
rlabel locali s 1082 347 1134 492 6 X
port 2 nsew signal output
rlabel locali s 1069 56 1134 147 6 X
port 2 nsew signal output
rlabel locali s 890 347 942 492 6 X
port 2 nsew signal output
rlabel locali s 890 56 942 147 6 X
port 2 nsew signal output
rlabel locali s 698 347 750 492 6 X
port 2 nsew signal output
rlabel locali s 698 56 750 147 6 X
port 2 nsew signal output
rlabel locali s 506 347 558 492 6 X
port 2 nsew signal output
rlabel locali s 506 344 1707 347 6 X
port 2 nsew signal output
rlabel locali s 506 299 2005 344 6 X
port 2 nsew signal output
rlabel locali s 506 147 2005 181 6 X
port 2 nsew signal output
rlabel locali s 506 56 558 147 6 X
port 2 nsew signal output
rlabel metal1 s 0 -48 2024 48 8 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 496 2024 592 6 VPWR
port 4 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2024 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1760850
string GDS_START 1747394
<< end >>
