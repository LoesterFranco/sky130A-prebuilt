magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 552 561
rect 119 367 167 527
rect 18 215 94 263
rect 203 323 237 493
rect 271 367 337 527
rect 371 323 405 493
rect 203 289 405 323
rect 439 297 505 527
rect 306 181 405 289
rect 203 147 405 181
rect 105 17 153 113
rect 203 51 237 147
rect 271 17 337 113
rect 371 51 405 147
rect 439 17 505 177
rect 0 -17 552 17
<< obsli1 >>
rect 19 331 85 493
rect 19 297 162 331
rect 128 249 162 297
rect 128 215 228 249
rect 128 181 162 215
rect 35 147 162 181
rect 35 51 69 147
<< metal1 >>
rect 0 496 552 592
rect 0 -48 552 48
<< labels >>
rlabel locali s 18 215 94 263 6 A
port 1 nsew signal input
rlabel locali s 371 323 405 493 6 X
port 2 nsew signal output
rlabel locali s 371 51 405 147 6 X
port 2 nsew signal output
rlabel locali s 306 181 405 289 6 X
port 2 nsew signal output
rlabel locali s 203 323 237 493 6 X
port 2 nsew signal output
rlabel locali s 203 289 405 323 6 X
port 2 nsew signal output
rlabel locali s 203 147 405 181 6 X
port 2 nsew signal output
rlabel locali s 203 51 237 147 6 X
port 2 nsew signal output
rlabel locali s 439 17 505 177 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 271 17 337 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 105 17 153 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 0 -17 552 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 552 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 439 297 505 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 271 367 337 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 119 367 167 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 0 527 552 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 496 552 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 552 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3041342
string GDS_START 3035994
<< end >>
