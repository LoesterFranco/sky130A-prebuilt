magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 25 291 263 357
rect 313 291 455 357
rect 1244 364 1511 430
rect 1442 226 1511 364
rect 1270 176 1511 226
rect 1270 70 1320 176
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 21 425 77 593
rect 111 459 161 649
rect 201 581 447 615
rect 201 425 251 581
rect 21 391 251 425
rect 291 425 347 547
rect 381 459 447 581
rect 495 481 561 649
rect 675 501 741 649
rect 886 532 952 649
rect 1098 532 1189 649
rect 1335 532 1401 649
rect 1515 532 1581 649
rect 780 467 1579 498
rect 617 464 1579 467
rect 617 447 814 464
rect 585 433 814 447
rect 585 425 651 433
rect 291 391 651 425
rect 991 399 1210 430
rect 500 381 651 391
rect 500 257 534 381
rect 780 364 1210 399
rect 780 349 846 364
rect 780 347 814 349
rect 615 315 814 347
rect 1176 330 1210 364
rect 615 281 856 315
rect 23 223 434 257
rect 23 121 73 223
rect 109 17 159 189
rect 196 121 246 223
rect 282 17 332 189
rect 368 87 434 223
rect 468 121 534 257
rect 568 87 634 247
rect 368 53 634 87
rect 704 97 756 247
rect 790 131 856 281
rect 890 285 1142 319
rect 890 97 956 285
rect 704 63 956 97
rect 990 17 1056 251
rect 1092 115 1142 285
rect 1176 264 1391 330
rect 1545 330 1579 464
rect 1615 430 1661 596
rect 1695 464 1761 649
rect 1815 430 1881 596
rect 1927 464 1993 649
rect 1615 424 1999 430
rect 1615 390 1759 424
rect 1793 390 1951 424
rect 1985 390 1999 424
rect 1615 364 1999 390
rect 1545 264 1929 330
rect 1965 230 1999 364
rect 1184 17 1234 226
rect 1630 196 1999 230
rect 1356 17 1422 142
rect 1528 17 1594 142
rect 1630 70 1680 196
rect 1714 17 1780 162
rect 1814 70 1880 196
rect 1916 17 1977 162
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 1759 390 1793 424
rect 1951 390 1985 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 1747 424 1805 430
rect 1747 390 1759 424
rect 1793 421 1805 424
rect 1939 424 1997 430
rect 1939 421 1951 424
rect 1793 393 1951 421
rect 1793 390 1805 393
rect 1747 384 1805 390
rect 1939 390 1951 393
rect 1985 390 1997 424
rect 1939 384 1997 390
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
rlabel locali s 25 291 263 357 6 A
port 1 nsew signal input
rlabel locali s 313 291 455 357 6 B
port 2 nsew signal input
rlabel locali s 1442 226 1511 364 6 COUT
port 3 nsew signal output
rlabel locali s 1270 176 1511 226 6 COUT
port 3 nsew signal output
rlabel locali s 1270 70 1320 176 6 COUT
port 3 nsew signal output
rlabel locali s 1244 364 1511 430 6 COUT
port 3 nsew signal output
rlabel metal1 s 1939 421 1997 430 6 SUM
port 4 nsew signal output
rlabel metal1 s 1939 384 1997 393 6 SUM
port 4 nsew signal output
rlabel metal1 s 1747 421 1805 430 6 SUM
port 4 nsew signal output
rlabel metal1 s 1747 393 1997 421 6 SUM
port 4 nsew signal output
rlabel metal1 s 1747 384 1805 393 6 SUM
port 4 nsew signal output
rlabel metal1 s 0 -49 2016 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 617 2016 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2016 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1918194
string GDS_START 1903074
<< end >>
