magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 285 2614 582
rect -38 261 424 285
rect 891 261 2614 285
<< pwell >>
rect 43 -2 47 3
<< scnmos >>
rect 89 47 119 177
rect 183 47 213 177
rect 393 66 423 150
rect 601 119 631 203
rect 693 119 723 203
rect 799 66 899 150
rect 973 66 1009 150
rect 1182 47 1212 119
rect 1292 47 1322 119
rect 1398 47 1428 131
rect 1480 47 1510 131
rect 1632 47 1662 175
rect 1727 47 1757 119
rect 1836 47 1866 119
rect 1972 47 2002 131
rect 2127 47 2157 131
rect 2223 47 2253 131
rect 2435 47 2465 177
<< pmoshvt >>
rect 81 297 117 497
rect 178 297 214 497
rect 488 389 524 497
rect 582 389 618 497
rect 664 389 700 497
rect 834 389 870 497
rect 943 389 979 497
rect 1166 413 1202 497
rect 1288 413 1324 497
rect 1382 413 1418 497
rect 1506 413 1542 497
rect 1714 329 1750 497
rect 1819 413 1855 497
rect 1915 413 1951 497
rect 2017 413 2053 497
rect 2129 413 2165 497
rect 2229 413 2265 497
rect 2427 297 2463 497
<< ndiff >>
rect 27 119 89 177
rect 27 85 35 119
rect 69 85 89 119
rect 27 47 89 85
rect 119 93 183 177
rect 119 59 129 93
rect 163 59 183 93
rect 119 47 183 59
rect 213 119 265 177
rect 539 165 601 203
rect 213 85 223 119
rect 257 85 265 119
rect 213 47 265 85
rect 331 129 393 150
rect 331 95 339 129
rect 373 95 393 129
rect 331 66 393 95
rect 423 112 475 150
rect 539 131 547 165
rect 581 131 601 165
rect 539 119 601 131
rect 631 119 693 203
rect 723 195 784 203
rect 723 161 733 195
rect 767 161 784 195
rect 723 150 784 161
rect 723 119 799 150
rect 423 78 433 112
rect 467 78 475 112
rect 423 66 475 78
rect 738 66 799 119
rect 899 66 973 150
rect 1009 108 1066 150
rect 1572 131 1632 175
rect 1348 119 1398 131
rect 1009 74 1020 108
rect 1054 74 1066 108
rect 1009 66 1066 74
rect 1120 101 1182 119
rect 1120 67 1128 101
rect 1162 67 1182 101
rect 1120 47 1182 67
rect 1212 95 1292 119
rect 1212 61 1238 95
rect 1272 61 1292 95
rect 1212 47 1292 61
rect 1322 47 1398 119
rect 1428 47 1480 131
rect 1510 93 1632 131
rect 1510 59 1554 93
rect 1588 59 1632 93
rect 1510 47 1632 59
rect 1662 119 1712 175
rect 1901 119 1972 131
rect 1662 89 1727 119
rect 1662 55 1672 89
rect 1706 55 1727 89
rect 1662 47 1727 55
rect 1757 93 1836 119
rect 1757 59 1772 93
rect 1806 59 1836 93
rect 1757 47 1836 59
rect 1866 47 1972 119
rect 2002 89 2127 131
rect 2002 55 2022 89
rect 2056 55 2127 89
rect 2002 47 2127 55
rect 2157 47 2223 131
rect 2253 93 2318 131
rect 2253 59 2272 93
rect 2306 59 2318 93
rect 2253 47 2318 59
rect 2373 93 2435 177
rect 2373 59 2381 93
rect 2415 59 2435 93
rect 2373 47 2435 59
rect 2465 143 2526 177
rect 2465 109 2484 143
rect 2518 109 2526 143
rect 2465 47 2526 109
<< pdiff >>
rect 1435 505 1485 517
rect 1435 497 1443 505
rect 27 477 81 497
rect 27 443 35 477
rect 69 443 81 477
rect 27 409 81 443
rect 27 375 35 409
rect 69 375 81 409
rect 27 297 81 375
rect 117 461 178 497
rect 117 427 132 461
rect 166 427 178 461
rect 117 297 178 427
rect 214 477 269 497
rect 214 443 227 477
rect 261 443 269 477
rect 214 409 269 443
rect 214 375 227 409
rect 261 375 269 409
rect 406 461 488 497
rect 406 427 442 461
rect 476 427 488 461
rect 406 389 488 427
rect 524 485 582 497
rect 524 451 536 485
rect 570 451 582 485
rect 524 389 582 451
rect 618 389 664 497
rect 700 477 834 497
rect 700 443 774 477
rect 808 443 834 477
rect 700 389 834 443
rect 870 389 943 497
rect 979 489 1037 497
rect 979 455 991 489
rect 1025 455 1037 489
rect 979 389 1037 455
rect 1091 471 1166 497
rect 1091 437 1120 471
rect 1154 437 1166 471
rect 1091 413 1166 437
rect 1202 483 1288 497
rect 1202 449 1242 483
rect 1276 449 1288 483
rect 1202 413 1288 449
rect 1324 459 1382 497
rect 1324 425 1336 459
rect 1370 425 1382 459
rect 1324 413 1382 425
rect 1418 471 1443 497
rect 1477 497 1485 505
rect 1477 471 1506 497
rect 1418 413 1506 471
rect 1542 459 1596 497
rect 1542 425 1554 459
rect 1588 425 1596 459
rect 1542 413 1596 425
rect 1650 485 1714 497
rect 1650 451 1668 485
rect 1702 451 1714 485
rect 214 297 269 375
rect 1650 329 1714 451
rect 1750 477 1819 497
rect 1750 443 1763 477
rect 1797 443 1819 477
rect 1750 413 1819 443
rect 1855 484 1915 497
rect 1855 450 1869 484
rect 1903 450 1915 484
rect 1855 413 1915 450
rect 1951 413 2017 497
rect 2053 489 2129 497
rect 2053 455 2083 489
rect 2117 455 2129 489
rect 2053 413 2129 455
rect 2165 459 2229 497
rect 2165 425 2182 459
rect 2216 425 2229 459
rect 2165 413 2229 425
rect 2265 485 2319 497
rect 2265 451 2277 485
rect 2311 451 2319 485
rect 2265 413 2319 451
rect 2373 485 2427 497
rect 2373 451 2381 485
rect 2415 451 2427 485
rect 2373 417 2427 451
rect 1750 329 1802 413
rect 2373 383 2381 417
rect 2415 383 2427 417
rect 2373 349 2427 383
rect 2373 315 2381 349
rect 2415 315 2427 349
rect 2373 297 2427 315
rect 2463 449 2526 497
rect 2463 415 2484 449
rect 2518 415 2526 449
rect 2463 381 2526 415
rect 2463 347 2484 381
rect 2518 347 2526 381
rect 2463 297 2526 347
<< ndiffc >>
rect 35 85 69 119
rect 129 59 163 93
rect 223 85 257 119
rect 339 95 373 129
rect 547 131 581 165
rect 733 161 767 195
rect 433 78 467 112
rect 1020 74 1054 108
rect 1128 67 1162 101
rect 1238 61 1272 95
rect 1554 59 1588 93
rect 1672 55 1706 89
rect 1772 59 1806 93
rect 2022 55 2056 89
rect 2272 59 2306 93
rect 2381 59 2415 93
rect 2484 109 2518 143
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 132 427 166 461
rect 227 443 261 477
rect 227 375 261 409
rect 442 427 476 461
rect 536 451 570 485
rect 774 443 808 477
rect 991 455 1025 489
rect 1120 437 1154 471
rect 1242 449 1276 483
rect 1336 425 1370 459
rect 1443 471 1477 505
rect 1554 425 1588 459
rect 1668 451 1702 485
rect 1763 443 1797 477
rect 1869 450 1903 484
rect 2083 455 2117 489
rect 2182 425 2216 459
rect 2277 451 2311 485
rect 2381 451 2415 485
rect 2381 383 2415 417
rect 2381 315 2415 349
rect 2484 415 2518 449
rect 2484 347 2518 381
<< poly >>
rect 81 497 117 523
rect 178 497 214 523
rect 488 497 524 523
rect 582 497 618 523
rect 664 497 700 523
rect 834 497 870 523
rect 943 497 979 523
rect 1166 497 1202 523
rect 1288 497 1324 523
rect 1382 497 1418 523
rect 1506 497 1542 523
rect 1714 497 1750 523
rect 1819 497 1855 523
rect 1915 497 1951 523
rect 2017 497 2053 523
rect 2129 497 2165 523
rect 2229 497 2265 523
rect 2427 497 2463 523
rect 1166 398 1202 413
rect 1288 398 1324 413
rect 1382 398 1418 413
rect 1506 398 1542 413
rect 488 374 524 389
rect 582 374 618 389
rect 664 374 700 389
rect 834 374 870 389
rect 943 374 979 389
rect 1164 375 1204 398
rect 486 357 526 374
rect 580 357 620 374
rect 393 327 620 357
rect 662 357 702 374
rect 662 341 723 357
rect 81 282 117 297
rect 178 282 214 297
rect 393 295 423 327
rect 79 269 119 282
rect 21 249 119 269
rect 176 265 216 282
rect 312 279 423 295
rect 662 307 672 341
rect 706 307 723 341
rect 662 291 723 307
rect 21 215 31 249
rect 65 215 119 249
rect 21 199 119 215
rect 161 249 225 265
rect 161 215 171 249
rect 205 215 225 249
rect 312 245 344 279
rect 378 245 423 279
rect 312 229 423 245
rect 161 199 225 215
rect 89 177 119 199
rect 183 177 213 199
rect 393 150 423 229
rect 486 275 562 285
rect 486 241 512 275
rect 546 248 562 275
rect 546 241 631 248
rect 486 218 631 241
rect 601 203 631 218
rect 693 203 723 291
rect 832 338 872 374
rect 941 340 981 374
rect 1148 365 1224 375
rect 832 321 899 338
rect 832 287 853 321
rect 887 287 899 321
rect 832 268 899 287
rect 941 324 1009 340
rect 941 290 957 324
rect 991 290 1009 324
rect 1148 331 1164 365
rect 1198 331 1224 365
rect 1148 321 1224 331
rect 941 274 1009 290
rect 1286 279 1326 398
rect 1380 371 1420 398
rect 1380 353 1462 371
rect 1380 319 1408 353
rect 1442 319 1462 353
rect 1380 303 1462 319
rect 799 150 899 176
rect 973 150 1009 274
rect 1081 263 1326 279
rect 1081 229 1096 263
rect 1130 249 1326 263
rect 1130 229 1144 249
rect 1081 213 1144 229
rect 1114 164 1144 213
rect 1258 191 1322 207
rect 601 93 631 119
rect 693 93 723 119
rect 1114 134 1212 164
rect 1258 157 1268 191
rect 1302 157 1322 191
rect 1258 141 1322 157
rect 1182 119 1212 134
rect 1292 119 1322 141
rect 1398 131 1428 303
rect 1504 225 1544 398
rect 1819 398 1855 413
rect 1915 398 1951 413
rect 2017 398 2053 413
rect 2129 398 2165 413
rect 2229 398 2265 413
rect 1714 314 1750 329
rect 1622 284 1752 314
rect 1622 267 1662 284
rect 1480 209 1544 225
rect 1480 175 1490 209
rect 1524 175 1544 209
rect 1586 251 1662 267
rect 1817 274 1857 398
rect 1913 383 1953 398
rect 1913 382 1963 383
rect 1899 366 1963 382
rect 1899 332 1909 366
rect 1943 332 1963 366
rect 1899 316 1963 332
rect 1817 252 1891 274
rect 1586 217 1596 251
rect 1630 217 1662 251
rect 1586 201 1662 217
rect 1836 239 1891 252
rect 1632 175 1662 201
rect 1727 191 1794 207
rect 1480 151 1544 175
rect 1480 131 1510 151
rect 393 51 423 66
rect 799 51 899 66
rect 89 21 119 47
rect 183 21 213 47
rect 393 21 899 51
rect 973 40 1009 66
rect 1727 157 1750 191
rect 1784 157 1794 191
rect 1727 141 1794 157
rect 1836 205 1847 239
rect 1881 205 1891 239
rect 1836 189 1891 205
rect 2015 229 2055 398
rect 2127 263 2167 398
rect 2227 365 2267 398
rect 2209 349 2275 365
rect 2209 315 2219 349
rect 2253 315 2275 349
rect 2209 301 2275 315
rect 2211 300 2275 301
rect 2213 299 2275 300
rect 2127 247 2188 263
rect 2015 213 2084 229
rect 2015 193 2030 213
rect 1727 119 1757 141
rect 1836 119 1866 189
rect 1972 179 2030 193
rect 2064 179 2084 213
rect 1972 163 2084 179
rect 2127 213 2137 247
rect 2171 213 2188 247
rect 2127 197 2188 213
rect 1972 131 2002 163
rect 2127 131 2157 197
rect 2235 170 2275 299
rect 2427 282 2463 297
rect 2425 265 2465 282
rect 2397 249 2465 265
rect 2397 215 2407 249
rect 2441 215 2465 249
rect 2397 199 2465 215
rect 2435 177 2465 199
rect 2223 146 2275 170
rect 2223 131 2253 146
rect 1182 21 1212 47
rect 1292 21 1322 47
rect 1398 21 1428 47
rect 1480 21 1510 47
rect 1632 21 1662 47
rect 1727 21 1757 47
rect 1836 21 1866 47
rect 1972 21 2002 47
rect 2127 21 2157 47
rect 2223 21 2253 47
rect 2435 21 2465 47
<< polycont >>
rect 672 307 706 341
rect 31 215 65 249
rect 171 215 205 249
rect 344 245 378 279
rect 512 241 546 275
rect 853 287 887 321
rect 957 290 991 324
rect 1164 331 1198 365
rect 1408 319 1442 353
rect 1096 229 1130 263
rect 1268 157 1302 191
rect 1490 175 1524 209
rect 1909 332 1943 366
rect 1596 217 1630 251
rect 1750 157 1784 191
rect 1847 205 1881 239
rect 2219 315 2253 349
rect 2030 179 2064 213
rect 2137 213 2171 247
rect 2407 215 2441 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2576 561
rect 18 477 69 493
rect 18 443 35 477
rect 18 409 69 443
rect 106 461 182 527
rect 106 427 132 461
rect 166 427 182 461
rect 227 477 273 493
rect 520 485 586 527
rect 261 443 273 477
rect 18 375 35 409
rect 227 409 273 443
rect 69 375 183 393
rect 18 359 183 375
rect 28 249 98 325
rect 28 215 31 249
rect 65 215 98 249
rect 28 195 98 215
rect 142 265 183 359
rect 261 357 273 409
rect 422 461 476 480
rect 422 427 442 461
rect 520 451 536 485
rect 570 451 586 485
rect 422 417 476 427
rect 422 383 546 417
rect 227 346 273 357
rect 142 255 205 265
rect 142 215 171 255
rect 142 199 205 215
rect 142 161 177 199
rect 19 127 177 161
rect 239 135 273 346
rect 317 279 444 349
rect 317 245 344 279
rect 378 267 444 279
rect 495 275 546 383
rect 378 245 398 267
rect 317 214 398 245
rect 495 241 512 275
rect 624 341 731 493
rect 624 307 672 341
rect 706 307 731 341
rect 624 271 731 307
rect 774 477 808 493
rect 971 489 1041 527
rect 1427 505 1493 527
rect 971 455 991 489
rect 1025 455 1041 489
rect 1096 471 1170 487
rect 774 421 808 443
rect 1096 437 1120 471
rect 1154 437 1170 471
rect 1219 483 1292 493
rect 1219 449 1242 483
rect 1276 449 1292 483
rect 1096 421 1130 437
rect 1219 427 1292 449
rect 774 387 1130 421
rect 495 237 546 241
rect 495 233 689 237
rect 453 199 689 233
rect 774 215 809 387
rect 453 180 487 199
rect 19 119 69 127
rect 19 85 35 119
rect 223 119 273 135
rect 19 69 69 85
rect 103 59 129 93
rect 163 59 179 93
rect 257 85 273 119
rect 223 69 273 85
rect 339 146 487 180
rect 339 129 373 146
rect 531 131 547 165
rect 581 131 607 165
rect 339 79 373 95
rect 407 78 433 112
rect 467 78 483 112
rect 103 17 179 59
rect 407 17 483 78
rect 531 17 607 131
rect 655 85 689 199
rect 733 195 809 215
rect 767 161 809 195
rect 733 135 809 161
rect 853 321 887 337
rect 853 85 887 287
rect 922 324 991 340
rect 922 290 957 324
rect 922 142 991 290
rect 1028 179 1062 387
rect 1164 365 1190 391
rect 1198 331 1224 357
rect 1164 315 1224 331
rect 1096 263 1130 279
rect 1096 213 1130 221
rect 1180 207 1224 315
rect 1258 277 1292 427
rect 1336 459 1370 475
rect 1427 471 1443 505
rect 1477 471 1493 505
rect 1630 485 1714 527
rect 1336 421 1370 425
rect 1554 459 1588 475
rect 1630 451 1668 485
rect 1702 451 1714 485
rect 1630 435 1714 451
rect 1763 477 1797 493
rect 1554 421 1588 425
rect 1336 387 1588 421
rect 1763 401 1797 443
rect 1839 484 2043 493
rect 1839 450 1869 484
rect 1903 450 2043 484
rect 1839 425 2043 450
rect 2083 489 2133 527
rect 2117 455 2133 489
rect 2251 485 2327 527
rect 2083 439 2133 455
rect 2182 459 2216 475
rect 1646 367 1797 401
rect 1646 353 1708 367
rect 1392 319 1408 353
rect 1442 319 1708 353
rect 1837 366 1913 391
rect 1837 333 1909 366
rect 1947 357 1969 391
rect 1258 251 1630 277
rect 1258 243 1596 251
rect 1180 191 1330 207
rect 1028 143 1144 179
rect 655 51 887 85
rect 1001 74 1020 108
rect 1054 74 1070 108
rect 1001 17 1070 74
rect 1110 101 1144 143
rect 1180 157 1268 191
rect 1302 157 1330 191
rect 1180 141 1330 157
rect 1110 67 1128 101
rect 1162 67 1178 101
rect 1368 95 1402 243
rect 1446 187 1490 209
rect 1524 187 1562 209
rect 1596 201 1630 217
rect 1446 153 1451 187
rect 1485 175 1490 187
rect 1485 153 1523 175
rect 1557 153 1562 187
rect 1674 167 1708 319
rect 1222 61 1238 95
rect 1272 61 1402 95
rect 1538 93 1604 109
rect 1538 59 1554 93
rect 1588 59 1604 93
rect 1538 17 1604 59
rect 1646 89 1708 167
rect 1742 332 1909 333
rect 1943 332 1969 357
rect 2008 349 2043 425
rect 2251 451 2277 485
rect 2311 451 2327 485
rect 2381 485 2438 527
rect 2415 451 2438 485
rect 2182 417 2216 425
rect 2381 417 2438 451
rect 2182 383 2346 417
rect 1742 299 1889 332
rect 2008 315 2219 349
rect 2253 315 2274 349
rect 1742 191 1794 299
rect 2008 297 2057 315
rect 1742 157 1750 191
rect 1784 157 1794 191
rect 1847 255 1881 265
rect 1847 184 1881 205
rect 1934 263 2057 297
rect 2312 265 2346 383
rect 2415 383 2438 417
rect 2381 349 2438 383
rect 2415 315 2438 349
rect 2381 299 2438 315
rect 2484 449 2557 465
rect 2518 415 2557 449
rect 2484 381 2557 415
rect 2518 347 2557 381
rect 1742 141 1794 157
rect 1934 107 1978 263
rect 2120 247 2274 255
rect 2030 213 2074 229
rect 2120 213 2137 247
rect 2171 213 2274 247
rect 2064 179 2074 213
rect 2030 173 2074 179
rect 2213 187 2274 213
rect 2030 139 2146 173
rect 1756 93 1978 107
rect 1646 55 1672 89
rect 1706 55 1722 89
rect 1756 59 1772 93
rect 1806 59 1978 93
rect 1756 51 1978 59
rect 2022 89 2066 105
rect 2056 55 2066 89
rect 2112 93 2146 139
rect 2213 153 2235 187
rect 2269 153 2274 187
rect 2213 127 2274 153
rect 2312 249 2441 265
rect 2312 215 2407 249
rect 2312 199 2441 215
rect 2312 93 2347 199
rect 2484 143 2557 347
rect 2112 59 2272 93
rect 2306 59 2347 93
rect 2381 93 2438 142
rect 2415 59 2438 93
rect 2022 17 2066 55
rect 2381 17 2438 59
rect 2518 109 2557 143
rect 2484 53 2557 109
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2576 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 227 375 261 391
rect 227 357 261 375
rect 171 249 205 255
rect 171 221 205 249
rect 1190 365 1224 391
rect 1190 357 1198 365
rect 1198 357 1224 365
rect 1096 229 1130 255
rect 1096 221 1130 229
rect 1913 366 1947 391
rect 1913 357 1943 366
rect 1943 357 1947 366
rect 1451 153 1485 187
rect 1523 175 1524 187
rect 1524 175 1557 187
rect 1523 153 1557 175
rect 1847 239 1881 255
rect 1847 221 1881 239
rect 2235 153 2269 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
<< metal1 >>
rect 0 561 2576 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2576 561
rect 0 496 2576 527
rect 214 391 274 397
rect 214 357 227 391
rect 261 388 274 391
rect 1178 391 1236 397
rect 1178 388 1190 391
rect 261 360 1190 388
rect 261 357 274 360
rect 214 351 274 357
rect 1178 357 1190 360
rect 1224 388 1236 391
rect 1900 391 1959 397
rect 1900 388 1913 391
rect 1224 360 1913 388
rect 1224 357 1236 360
rect 1178 351 1236 357
rect 1900 357 1913 360
rect 1947 357 1959 391
rect 1900 351 1959 357
rect 159 255 217 261
rect 159 221 171 255
rect 205 252 217 255
rect 1084 255 1142 261
rect 1084 252 1096 255
rect 205 224 1096 252
rect 205 221 217 224
rect 159 215 217 221
rect 1084 221 1096 224
rect 1130 252 1142 255
rect 1831 255 1893 261
rect 1831 252 1847 255
rect 1130 224 1847 252
rect 1130 221 1142 224
rect 1084 215 1142 221
rect 1831 221 1847 224
rect 1881 221 1893 255
rect 1831 215 1893 221
rect 1429 187 1580 193
rect 1429 153 1451 187
rect 1485 153 1523 187
rect 1557 184 1580 187
rect 2223 187 2281 193
rect 2223 184 2235 187
rect 1557 156 2235 184
rect 1557 153 1580 156
rect 1429 147 1580 153
rect 2223 153 2235 156
rect 2269 153 2281 187
rect 2223 147 2281 153
rect 0 17 2576 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2576 17
rect 0 -48 2576 -17
<< labels >>
rlabel comment s 0 0 0 0 4 sdfrtp_1
flabel nbase s 34 528 63 556 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel pwell s 43 -2 47 3 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel metal1 s 39 -10 57 7 0 FreeSans 200 0 0 0 VGND
port 6 nsew
flabel metal1 s 31 534 63 554 0 FreeSans 200 0 0 0 VPWR
port 9 nsew
flabel metal1 s 2237 153 2271 187 0 FreeSans 200 0 0 0 RESET_B
port 3 nsew
flabel corelocali s 2513 85 2547 119 0 FreeSans 400 0 0 0 Q
port 10 nsew
flabel corelocali s 2513 289 2547 323 0 FreeSans 400 0 0 0 Q
port 10 nsew
flabel corelocali s 2513 357 2547 391 0 FreeSans 400 0 0 0 Q
port 10 nsew
flabel corelocali s 2513 425 2547 459 0 FreeSans 400 0 0 0 Q
port 10 nsew
flabel corelocali s 30 289 64 323 0 FreeSans 400 0 0 0 CLK
port 1 nsew
flabel corelocali s 31 221 65 255 0 FreeSans 400 0 0 0 CLK
port 1 nsew
flabel corelocali s 671 289 705 323 0 FreeSans 200 0 0 0 D
port 2 nsew
flabel corelocali s 947 289 983 323 0 FreeSans 200 0 0 0 SCD
port 4 nsew
flabel corelocali s 391 289 425 323 0 FreeSans 200 0 0 0 SCE
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 2576 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 64666
string GDS_START 46514
<< end >>
