magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 1190 704
<< pwell >>
rect 0 0 1152 49
<< scnmos >>
rect 91 74 121 222
rect 177 74 207 222
rect 263 74 293 222
rect 349 74 379 222
rect 447 94 477 222
rect 533 94 563 222
rect 753 74 783 202
rect 839 74 869 202
rect 925 74 955 202
rect 1011 74 1041 202
<< pmoshvt >>
rect 94 368 124 592
rect 184 368 214 592
rect 274 368 304 592
rect 364 368 394 592
rect 558 392 588 592
rect 648 392 678 592
rect 738 392 768 592
rect 828 392 858 592
rect 918 392 948 592
rect 1008 392 1038 592
<< ndiff >>
rect 34 142 91 222
rect 34 108 46 142
rect 80 108 91 142
rect 34 74 91 108
rect 121 210 177 222
rect 121 176 132 210
rect 166 176 177 210
rect 121 120 177 176
rect 121 86 132 120
rect 166 86 177 120
rect 121 74 177 86
rect 207 142 263 222
rect 207 108 218 142
rect 252 108 263 142
rect 207 74 263 108
rect 293 210 349 222
rect 293 176 304 210
rect 338 176 349 210
rect 293 120 349 176
rect 293 86 304 120
rect 338 86 349 120
rect 293 74 349 86
rect 379 158 447 222
rect 379 124 390 158
rect 424 124 447 158
rect 379 94 447 124
rect 477 210 533 222
rect 477 176 488 210
rect 522 176 533 210
rect 477 140 533 176
rect 477 106 488 140
rect 522 106 533 140
rect 477 94 533 106
rect 563 169 616 222
rect 563 135 574 169
rect 608 135 616 169
rect 563 94 616 135
rect 700 188 753 202
rect 700 154 708 188
rect 742 154 753 188
rect 700 120 753 154
rect 379 74 432 94
rect 700 86 708 120
rect 742 86 753 120
rect 700 74 753 86
rect 783 169 839 202
rect 783 135 794 169
rect 828 135 839 169
rect 783 74 839 135
rect 869 190 925 202
rect 869 156 880 190
rect 914 156 925 190
rect 869 120 925 156
rect 869 86 880 120
rect 914 86 925 120
rect 869 74 925 86
rect 955 134 1011 202
rect 955 100 966 134
rect 1000 100 1011 134
rect 955 74 1011 100
rect 1041 190 1094 202
rect 1041 156 1052 190
rect 1086 156 1094 190
rect 1041 120 1094 156
rect 1041 86 1052 120
rect 1086 86 1094 120
rect 1041 74 1094 86
<< pdiff >>
rect 39 580 94 592
rect 39 546 47 580
rect 81 546 94 580
rect 39 462 94 546
rect 39 428 47 462
rect 81 428 94 462
rect 39 368 94 428
rect 124 580 184 592
rect 124 546 137 580
rect 171 546 184 580
rect 124 497 184 546
rect 124 463 137 497
rect 171 463 184 497
rect 124 414 184 463
rect 124 380 137 414
rect 171 380 184 414
rect 124 368 184 380
rect 214 580 274 592
rect 214 546 227 580
rect 261 546 274 580
rect 214 478 274 546
rect 214 444 227 478
rect 261 444 274 478
rect 214 368 274 444
rect 304 580 364 592
rect 304 546 317 580
rect 351 546 364 580
rect 304 497 364 546
rect 304 463 317 497
rect 351 463 364 497
rect 304 414 364 463
rect 304 380 317 414
rect 351 380 364 414
rect 304 368 364 380
rect 394 580 449 592
rect 394 546 407 580
rect 441 546 449 580
rect 394 510 449 546
rect 394 476 407 510
rect 441 476 449 510
rect 394 440 449 476
rect 394 406 407 440
rect 441 406 449 440
rect 394 368 449 406
rect 503 580 558 592
rect 503 546 511 580
rect 545 546 558 580
rect 503 510 558 546
rect 503 476 511 510
rect 545 476 558 510
rect 503 440 558 476
rect 503 406 511 440
rect 545 406 558 440
rect 503 392 558 406
rect 588 531 648 592
rect 588 497 601 531
rect 635 497 648 531
rect 588 442 648 497
rect 588 408 601 442
rect 635 408 648 442
rect 588 392 648 408
rect 678 580 738 592
rect 678 546 691 580
rect 725 546 738 580
rect 678 510 738 546
rect 678 476 691 510
rect 725 476 738 510
rect 678 440 738 476
rect 678 406 691 440
rect 725 406 738 440
rect 678 392 738 406
rect 768 580 828 592
rect 768 546 781 580
rect 815 546 828 580
rect 768 508 828 546
rect 768 474 781 508
rect 815 474 828 508
rect 768 392 828 474
rect 858 580 918 592
rect 858 546 871 580
rect 905 546 918 580
rect 858 510 918 546
rect 858 476 871 510
rect 905 476 918 510
rect 858 440 918 476
rect 858 406 871 440
rect 905 406 918 440
rect 858 392 918 406
rect 948 580 1008 592
rect 948 546 961 580
rect 995 546 1008 580
rect 948 508 1008 546
rect 948 474 961 508
rect 995 474 1008 508
rect 948 392 1008 474
rect 1038 580 1093 592
rect 1038 546 1051 580
rect 1085 546 1093 580
rect 1038 509 1093 546
rect 1038 475 1051 509
rect 1085 475 1093 509
rect 1038 438 1093 475
rect 1038 404 1051 438
rect 1085 404 1093 438
rect 1038 392 1093 404
<< ndiffc >>
rect 46 108 80 142
rect 132 176 166 210
rect 132 86 166 120
rect 218 108 252 142
rect 304 176 338 210
rect 304 86 338 120
rect 390 124 424 158
rect 488 176 522 210
rect 488 106 522 140
rect 574 135 608 169
rect 708 154 742 188
rect 708 86 742 120
rect 794 135 828 169
rect 880 156 914 190
rect 880 86 914 120
rect 966 100 1000 134
rect 1052 156 1086 190
rect 1052 86 1086 120
<< pdiffc >>
rect 47 546 81 580
rect 47 428 81 462
rect 137 546 171 580
rect 137 463 171 497
rect 137 380 171 414
rect 227 546 261 580
rect 227 444 261 478
rect 317 546 351 580
rect 317 463 351 497
rect 317 380 351 414
rect 407 546 441 580
rect 407 476 441 510
rect 407 406 441 440
rect 511 546 545 580
rect 511 476 545 510
rect 511 406 545 440
rect 601 497 635 531
rect 601 408 635 442
rect 691 546 725 580
rect 691 476 725 510
rect 691 406 725 440
rect 781 546 815 580
rect 781 474 815 508
rect 871 546 905 580
rect 871 476 905 510
rect 871 406 905 440
rect 961 546 995 580
rect 961 474 995 508
rect 1051 546 1085 580
rect 1051 475 1085 509
rect 1051 404 1085 438
<< poly >>
rect 94 592 124 618
rect 184 592 214 618
rect 274 592 304 618
rect 364 592 394 618
rect 558 592 588 618
rect 648 592 678 618
rect 738 592 768 618
rect 828 592 858 618
rect 918 592 948 618
rect 1008 592 1038 618
rect 558 377 588 392
rect 648 377 678 392
rect 738 377 768 392
rect 828 377 858 392
rect 918 377 948 392
rect 1008 377 1038 392
rect 94 353 124 368
rect 184 353 214 368
rect 274 353 304 368
rect 364 353 394 368
rect 555 353 591 377
rect 645 353 681 377
rect 91 326 127 353
rect 181 326 217 353
rect 271 326 307 353
rect 361 326 397 353
rect 91 310 397 326
rect 91 276 143 310
rect 177 276 211 310
rect 245 276 279 310
rect 313 276 347 310
rect 381 276 397 310
rect 91 260 397 276
rect 447 337 681 353
rect 447 303 501 337
rect 535 303 681 337
rect 447 287 681 303
rect 735 356 771 377
rect 825 356 861 377
rect 735 340 861 356
rect 735 306 751 340
rect 785 320 861 340
rect 785 306 869 320
rect 735 290 869 306
rect 91 222 121 260
rect 177 222 207 260
rect 263 222 293 260
rect 349 222 379 260
rect 447 222 477 287
rect 533 222 563 287
rect 753 202 783 290
rect 839 202 869 290
rect 915 318 951 377
rect 1005 318 1041 377
rect 915 302 1041 318
rect 915 268 931 302
rect 965 268 1041 302
rect 915 252 1041 268
rect 925 202 955 252
rect 1011 202 1041 252
rect 91 48 121 74
rect 177 48 207 74
rect 263 48 293 74
rect 349 48 379 74
rect 447 68 477 94
rect 533 68 563 94
rect 753 48 783 74
rect 839 48 869 74
rect 925 48 955 74
rect 1011 48 1041 74
<< polycont >>
rect 143 276 177 310
rect 211 276 245 310
rect 279 276 313 310
rect 347 276 381 310
rect 501 303 535 337
rect 751 306 785 340
rect 931 268 965 302
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 31 580 97 649
rect 31 546 47 580
rect 81 546 97 580
rect 31 462 97 546
rect 31 428 47 462
rect 81 428 97 462
rect 137 580 171 596
rect 137 497 171 546
rect 137 414 171 463
rect 211 580 261 649
rect 211 546 227 580
rect 211 478 261 546
rect 211 444 227 478
rect 211 428 261 444
rect 301 580 367 596
rect 301 546 317 580
rect 351 546 367 580
rect 301 497 367 546
rect 301 463 317 497
rect 351 463 367 497
rect 25 380 137 394
rect 301 414 367 463
rect 301 394 317 414
rect 171 380 317 394
rect 351 380 367 414
rect 407 580 457 649
rect 441 546 457 580
rect 407 510 457 546
rect 441 476 457 510
rect 407 440 457 476
rect 441 406 457 440
rect 407 390 457 406
rect 495 581 725 615
rect 495 580 545 581
rect 495 546 511 580
rect 691 580 725 581
rect 495 510 545 546
rect 495 476 511 510
rect 495 440 545 476
rect 495 406 511 440
rect 495 390 545 406
rect 585 531 651 547
rect 585 497 601 531
rect 635 497 651 531
rect 585 442 651 497
rect 585 408 601 442
rect 635 408 651 442
rect 25 360 367 380
rect 25 226 71 360
rect 485 337 551 356
rect 127 310 441 326
rect 127 276 143 310
rect 177 276 211 310
rect 245 276 279 310
rect 313 276 347 310
rect 381 276 441 310
rect 485 303 501 337
rect 535 303 551 337
rect 485 287 551 303
rect 127 260 441 276
rect 374 253 441 260
rect 585 256 651 408
rect 691 510 725 546
rect 691 440 725 476
rect 765 580 815 649
rect 765 546 781 580
rect 765 508 815 546
rect 765 474 781 508
rect 765 458 815 474
rect 855 580 905 596
rect 855 546 871 580
rect 855 510 905 546
rect 855 476 871 510
rect 855 440 905 476
rect 945 580 1011 649
rect 945 546 961 580
rect 995 546 1011 580
rect 945 508 1011 546
rect 945 474 961 508
rect 995 474 1011 508
rect 945 458 1011 474
rect 1051 580 1101 596
rect 1085 546 1101 580
rect 1051 509 1101 546
rect 1085 475 1101 509
rect 855 424 871 440
rect 725 406 871 424
rect 1051 438 1101 475
rect 905 406 1051 424
rect 691 404 1051 406
rect 1085 404 1101 438
rect 691 390 1101 404
rect 1051 388 1101 390
rect 697 340 839 356
rect 697 306 751 340
rect 785 306 839 340
rect 697 290 839 306
rect 889 302 981 356
rect 889 268 931 302
rect 965 268 981 302
rect 585 253 844 256
rect 25 210 338 226
rect 374 222 844 253
rect 889 252 981 268
rect 374 219 651 222
rect 25 192 132 210
rect 166 192 304 210
rect 30 142 96 158
rect 30 108 46 142
rect 80 108 96 142
rect 30 17 96 108
rect 132 120 166 176
rect 288 176 304 192
rect 472 210 522 219
rect 132 70 166 86
rect 202 142 252 158
rect 202 108 218 142
rect 202 17 252 108
rect 288 120 338 176
rect 288 86 304 120
rect 288 70 338 86
rect 374 158 424 185
rect 374 124 390 158
rect 374 17 424 124
rect 472 176 488 210
rect 472 140 522 176
rect 472 106 488 140
rect 472 90 522 106
rect 558 169 624 185
rect 558 135 574 169
rect 608 135 624 169
rect 558 17 624 135
rect 692 154 708 188
rect 742 154 758 188
rect 692 120 758 154
rect 692 86 708 120
rect 742 86 758 120
rect 792 169 844 222
rect 792 135 794 169
rect 828 135 844 169
rect 792 119 844 135
rect 880 190 1102 218
rect 914 184 1052 190
rect 880 120 914 156
rect 1086 156 1102 190
rect 692 85 758 86
rect 880 85 914 86
rect 692 51 914 85
rect 950 134 1016 150
rect 950 100 966 134
rect 1000 100 1016 134
rect 950 17 1016 100
rect 1052 120 1102 156
rect 1086 86 1102 120
rect 1052 70 1102 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a21o_4
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 1152 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3998366
string GDS_START 3988526
<< end >>
