magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 409 514 487 596
rect 761 514 827 547
rect 409 498 827 514
rect 17 480 827 498
rect 17 464 487 480
rect 17 202 51 464
rect 409 412 487 464
rect 521 412 1039 446
rect 521 378 555 412
rect 269 344 555 378
rect 269 270 335 344
rect 785 236 851 310
rect 1005 236 1039 412
rect 785 202 1039 236
rect 17 168 167 202
rect 133 85 167 168
rect 438 85 515 100
rect 133 51 515 85
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 23 532 89 649
rect 246 532 375 649
rect 528 548 594 649
rect 652 581 927 615
rect 652 548 720 581
rect 861 480 927 581
rect 961 480 1027 649
rect 130 364 235 430
rect 85 276 167 310
rect 85 242 127 276
rect 161 242 167 276
rect 85 236 167 242
rect 201 236 235 364
rect 605 344 935 378
rect 605 310 671 344
rect 889 336 935 344
rect 383 236 517 310
rect 601 276 671 310
rect 601 242 607 276
rect 641 242 671 276
rect 601 236 671 242
rect 889 270 971 336
rect 201 202 517 236
rect 23 17 99 134
rect 201 127 290 202
rect 551 168 617 202
rect 336 134 1033 168
rect 336 119 402 134
rect 551 70 617 134
rect 653 17 720 100
rect 756 98 822 134
rect 862 17 931 100
rect 967 98 1033 134
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 127 242 161 276
rect 607 242 641 276
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 683 1056 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 0 617 1056 649
rect 115 276 173 282
rect 115 242 127 276
rect 161 273 173 276
rect 595 276 653 282
rect 595 273 607 276
rect 161 245 607 273
rect 161 242 173 245
rect 115 236 173 242
rect 595 242 607 245
rect 641 242 653 276
rect 595 236 653 242
rect 0 17 1056 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -49 1056 -17
<< labels >>
rlabel metal1 s 595 273 653 282 6 A
port 1 nsew signal input
rlabel metal1 s 595 236 653 245 6 A
port 1 nsew signal input
rlabel metal1 s 115 273 173 282 6 A
port 1 nsew signal input
rlabel metal1 s 115 245 653 273 6 A
port 1 nsew signal input
rlabel metal1 s 115 236 173 245 6 A
port 1 nsew signal input
rlabel locali s 1005 236 1039 412 6 B
port 2 nsew signal input
rlabel locali s 785 236 851 310 6 B
port 2 nsew signal input
rlabel locali s 785 202 1039 236 6 B
port 2 nsew signal input
rlabel locali s 521 412 1039 446 6 B
port 2 nsew signal input
rlabel locali s 521 378 555 412 6 B
port 2 nsew signal input
rlabel locali s 269 344 555 378 6 B
port 2 nsew signal input
rlabel locali s 269 270 335 344 6 B
port 2 nsew signal input
rlabel locali s 761 514 827 547 6 Y
port 3 nsew signal output
rlabel locali s 438 85 515 100 6 Y
port 3 nsew signal output
rlabel locali s 409 514 487 596 6 Y
port 3 nsew signal output
rlabel locali s 409 498 827 514 6 Y
port 3 nsew signal output
rlabel locali s 409 412 487 464 6 Y
port 3 nsew signal output
rlabel locali s 133 85 167 168 6 Y
port 3 nsew signal output
rlabel locali s 133 51 515 85 6 Y
port 3 nsew signal output
rlabel locali s 17 480 827 498 6 Y
port 3 nsew signal output
rlabel locali s 17 464 487 480 6 Y
port 3 nsew signal output
rlabel locali s 17 202 51 464 6 Y
port 3 nsew signal output
rlabel locali s 17 168 167 202 6 Y
port 3 nsew signal output
rlabel metal1 s 0 -49 1056 49 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1056 715 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1056 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 589988
string GDS_START 581694
<< end >>
