magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 184 561
rect 17 51 167 493
rect 0 -17 184 17
<< metal1 >>
rect 0 496 184 592
rect 0 -48 184 48
<< labels >>
rlabel locali s 17 51 167 493 6 DIODE
port 1 nsew signal input
rlabel locali s 0 -17 184 17 8 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 184 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel locali s 0 527 184 561 6 VPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 0 496 184 592 6 VPWR
port 3 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 184 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2565610
string GDS_START 2562180
<< end >>
