magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 135 351 169 437
rect 327 351 377 437
rect 29 317 377 351
rect 29 157 136 317
rect 500 199 581 305
rect 789 302 1087 336
rect 789 255 834 302
rect 1027 258 1087 302
rect 745 202 834 255
rect 868 202 993 255
rect 1027 211 1120 258
rect 29 123 377 157
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 23 387 89 527
rect 205 387 281 527
rect 413 303 463 527
rect 531 459 753 493
rect 531 339 565 459
rect 170 199 460 265
rect 426 157 460 199
rect 625 168 659 425
rect 717 404 753 459
rect 787 455 863 527
rect 907 404 941 493
rect 975 455 1051 527
rect 1106 404 1172 479
rect 717 370 1172 404
rect 717 289 753 370
rect 1121 292 1172 370
rect 625 157 953 168
rect 426 134 953 157
rect 426 123 659 134
rect 21 17 89 89
rect 205 17 281 89
rect 422 17 577 89
rect 625 51 659 123
rect 711 17 777 89
rect 897 81 953 134
rect 1089 17 1145 177
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
rlabel locali s 868 202 993 255 6 A1
port 1 nsew signal input
rlabel locali s 1027 258 1087 302 6 A2
port 2 nsew signal input
rlabel locali s 1027 211 1120 258 6 A2
port 2 nsew signal input
rlabel locali s 789 302 1087 336 6 A2
port 2 nsew signal input
rlabel locali s 789 255 834 302 6 A2
port 2 nsew signal input
rlabel locali s 745 202 834 255 6 A2
port 2 nsew signal input
rlabel locali s 500 199 581 305 6 B1
port 3 nsew signal input
rlabel locali s 327 351 377 437 6 X
port 4 nsew signal output
rlabel locali s 135 351 169 437 6 X
port 4 nsew signal output
rlabel locali s 29 317 377 351 6 X
port 4 nsew signal output
rlabel locali s 29 157 136 317 6 X
port 4 nsew signal output
rlabel locali s 29 123 377 157 6 X
port 4 nsew signal output
rlabel metal1 s 0 -48 1196 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 1196 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1194602
string GDS_START 1186030
<< end >>
