magic
tech sky130A
magscale 1 2
timestamp 1601050088
<< locali >>
rect 25 249 167 356
rect 333 390 530 424
rect 333 315 367 390
rect 496 383 530 390
rect 496 378 924 383
rect 496 356 1217 378
rect 269 252 367 315
rect 496 349 1319 356
rect 496 249 562 349
rect 790 252 856 349
rect 890 344 1319 349
rect 1183 310 1319 344
rect 1449 402 1515 596
rect 1639 402 1705 596
rect 1449 368 1705 402
rect 1183 252 1268 310
rect 1657 234 1705 368
rect 1829 398 1895 596
rect 2019 398 2087 596
rect 1829 364 2087 398
rect 2033 310 2087 364
rect 1453 184 1723 234
rect 2033 230 2085 310
rect 1861 196 2085 230
rect 1861 78 1911 196
rect 2033 78 2085 196
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 23 451 89 596
rect 129 485 163 649
rect 197 526 401 592
rect 197 451 231 526
rect 442 492 508 551
rect 23 417 231 451
rect 265 458 508 492
rect 23 390 89 417
rect 265 383 299 458
rect 201 349 299 383
rect 634 417 700 649
rect 734 451 800 551
rect 834 485 914 649
rect 948 451 1014 551
rect 734 417 1014 451
rect 1048 446 1114 551
rect 1359 458 1409 649
rect 1048 424 1285 446
rect 1048 412 1415 424
rect 1251 390 1415 412
rect 201 218 235 349
rect 401 276 455 356
rect 401 242 415 276
rect 449 242 455 276
rect 601 276 748 315
rect 401 236 455 242
rect 601 242 607 276
rect 641 252 748 276
rect 1381 334 1415 390
rect 1555 436 1605 649
rect 641 242 643 252
rect 601 236 643 242
rect 986 244 1052 310
rect 1086 276 1149 310
rect 986 218 1051 244
rect 1086 242 1087 276
rect 1121 242 1149 276
rect 1381 268 1621 334
rect 1086 236 1149 242
rect 1381 218 1415 268
rect 1745 364 1795 649
rect 1935 432 1985 649
rect 2125 364 2175 649
rect 1793 264 1991 330
rect 23 150 89 215
rect 201 202 367 218
rect 677 202 1051 218
rect 1183 202 1415 218
rect 201 184 1051 202
rect 333 168 711 184
rect 23 134 299 150
rect 23 116 393 134
rect 23 70 89 116
rect 125 17 231 82
rect 265 70 393 116
rect 427 70 493 168
rect 635 17 701 134
rect 745 116 983 150
rect 745 70 795 116
rect 831 17 897 82
rect 933 70 983 116
rect 1017 85 1051 184
rect 1085 184 1415 202
rect 1085 168 1217 184
rect 1085 119 1135 168
rect 1793 150 1827 264
rect 1251 116 1827 150
rect 1251 85 1285 116
rect 1017 51 1285 85
rect 1351 17 1417 82
rect 1555 17 1621 82
rect 1759 17 1825 82
rect 1947 17 1997 162
rect 2119 17 2185 234
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 415 242 449 276
rect 607 242 641 276
rect 1087 242 1121 276
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
<< metal1 >>
rect 0 683 2208 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 0 617 2208 649
rect 403 276 461 282
rect 403 242 415 276
rect 449 273 461 276
rect 595 276 653 282
rect 595 273 607 276
rect 449 245 607 273
rect 449 242 461 245
rect 403 236 461 242
rect 595 242 607 245
rect 641 273 653 276
rect 1075 276 1133 282
rect 1075 273 1087 276
rect 641 245 1087 273
rect 641 242 653 245
rect 595 236 653 242
rect 1075 242 1087 245
rect 1121 242 1133 276
rect 1075 236 1133 242
rect 0 17 2208 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
rect 0 -49 2208 -17
<< labels >>
rlabel locali s 25 249 167 356 6 A
port 1 nsew signal input
rlabel locali s 1183 310 1319 344 6 B
port 2 nsew signal input
rlabel locali s 1183 252 1268 310 6 B
port 2 nsew signal input
rlabel locali s 890 344 1319 349 6 B
port 2 nsew signal input
rlabel locali s 790 252 856 349 6 B
port 2 nsew signal input
rlabel locali s 496 383 530 390 6 B
port 2 nsew signal input
rlabel locali s 496 378 924 383 6 B
port 2 nsew signal input
rlabel locali s 496 356 1217 378 6 B
port 2 nsew signal input
rlabel locali s 496 349 1319 356 6 B
port 2 nsew signal input
rlabel locali s 496 249 562 349 6 B
port 2 nsew signal input
rlabel locali s 333 390 530 424 6 B
port 2 nsew signal input
rlabel locali s 333 315 367 390 6 B
port 2 nsew signal input
rlabel locali s 269 252 367 315 6 B
port 2 nsew signal input
rlabel metal1 s 1075 273 1133 282 6 CIN
port 3 nsew signal input
rlabel metal1 s 1075 236 1133 245 6 CIN
port 3 nsew signal input
rlabel metal1 s 595 273 653 282 6 CIN
port 3 nsew signal input
rlabel metal1 s 595 236 653 245 6 CIN
port 3 nsew signal input
rlabel metal1 s 403 273 461 282 6 CIN
port 3 nsew signal input
rlabel metal1 s 403 245 1133 273 6 CIN
port 3 nsew signal input
rlabel metal1 s 403 236 461 245 6 CIN
port 3 nsew signal input
rlabel locali s 2033 310 2087 364 6 COUT
port 4 nsew signal output
rlabel locali s 2033 230 2085 310 6 COUT
port 4 nsew signal output
rlabel locali s 2033 78 2085 196 6 COUT
port 4 nsew signal output
rlabel locali s 2019 398 2087 596 6 COUT
port 4 nsew signal output
rlabel locali s 1861 196 2085 230 6 COUT
port 4 nsew signal output
rlabel locali s 1861 78 1911 196 6 COUT
port 4 nsew signal output
rlabel locali s 1829 398 1895 596 6 COUT
port 4 nsew signal output
rlabel locali s 1829 364 2087 398 6 COUT
port 4 nsew signal output
rlabel locali s 1657 234 1705 368 6 SUM
port 5 nsew signal output
rlabel locali s 1639 402 1705 596 6 SUM
port 5 nsew signal output
rlabel locali s 1453 184 1723 234 6 SUM
port 5 nsew signal output
rlabel locali s 1449 402 1515 596 6 SUM
port 5 nsew signal output
rlabel locali s 1449 368 1705 402 6 SUM
port 5 nsew signal output
rlabel metal1 s 0 -49 2208 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 2208 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2208 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 2445280
string GDS_START 2429006
<< end >>
