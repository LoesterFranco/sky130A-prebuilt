magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 644 561
rect 17 299 69 527
rect 108 417 346 483
rect 382 367 438 527
rect 480 299 526 493
rect 17 215 85 265
rect 492 152 526 299
rect 560 292 611 527
rect 118 17 264 113
rect 366 17 442 97
rect 480 83 526 152
rect 560 17 611 185
rect 0 -17 644 17
<< obsli1 >>
rect 119 265 153 377
rect 197 333 281 383
rect 197 299 446 333
rect 412 265 446 299
rect 119 199 266 265
rect 412 199 458 265
rect 119 181 168 199
rect 21 147 168 181
rect 412 165 446 199
rect 21 53 84 147
rect 298 131 446 165
rect 298 61 332 131
<< metal1 >>
rect 0 496 644 592
rect 0 -48 644 48
<< labels >>
rlabel locali s 108 417 346 483 6 A
port 1 nsew signal input
rlabel locali s 17 215 85 265 6 B_N
port 2 nsew signal input
rlabel locali s 492 152 526 299 6 X
port 3 nsew signal output
rlabel locali s 480 299 526 493 6 X
port 3 nsew signal output
rlabel locali s 480 83 526 152 6 X
port 3 nsew signal output
rlabel locali s 560 17 611 185 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 366 17 442 97 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 118 17 264 113 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 644 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 644 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 560 292 611 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 382 367 438 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 17 299 69 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 644 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 644 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1019650
string GDS_START 1014186
<< end >>
