magic
tech sky130A
magscale 1 2
timestamp 1599588201
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 79 47 109 177
rect 267 47 297 177
rect 351 47 381 177
rect 451 47 481 177
rect 535 47 565 177
<< pmoshvt >>
rect 83 297 113 497
rect 262 297 292 497
rect 339 297 369 497
rect 463 297 493 497
rect 535 297 565 497
<< ndiff >>
rect 27 136 79 177
rect 27 102 35 136
rect 69 102 79 136
rect 27 47 79 102
rect 109 93 161 177
rect 109 59 119 93
rect 153 59 161 93
rect 109 47 161 59
rect 215 95 267 177
rect 215 61 223 95
rect 257 61 267 95
rect 215 47 267 61
rect 297 163 351 177
rect 297 129 307 163
rect 341 129 351 163
rect 297 47 351 129
rect 381 163 451 177
rect 381 129 407 163
rect 441 129 451 163
rect 381 95 451 129
rect 381 61 407 95
rect 441 61 451 95
rect 381 47 451 61
rect 481 89 535 177
rect 481 55 491 89
rect 525 55 535 89
rect 481 47 535 55
rect 565 163 617 177
rect 565 129 575 163
rect 609 129 617 163
rect 565 95 617 129
rect 565 61 575 95
rect 609 61 617 95
rect 565 47 617 61
<< pdiff >>
rect 27 477 83 497
rect 27 443 39 477
rect 73 443 83 477
rect 27 409 83 443
rect 27 375 39 409
rect 73 375 83 409
rect 27 341 83 375
rect 27 307 39 341
rect 73 307 83 341
rect 27 297 83 307
rect 113 477 262 497
rect 113 443 127 477
rect 161 443 218 477
rect 252 443 262 477
rect 113 409 262 443
rect 113 375 127 409
rect 161 375 218 409
rect 252 375 262 409
rect 113 297 262 375
rect 292 297 339 497
rect 369 477 463 497
rect 369 443 379 477
rect 413 443 463 477
rect 369 409 463 443
rect 369 375 379 409
rect 413 375 463 409
rect 369 341 463 375
rect 369 307 379 341
rect 413 307 463 341
rect 369 297 463 307
rect 493 297 535 497
rect 565 485 617 497
rect 565 451 575 485
rect 609 451 617 485
rect 565 417 617 451
rect 565 383 575 417
rect 609 383 617 417
rect 565 349 617 383
rect 565 315 575 349
rect 609 315 617 349
rect 565 297 617 315
<< ndiffc >>
rect 35 102 69 136
rect 119 59 153 93
rect 223 61 257 95
rect 307 129 341 163
rect 407 129 441 163
rect 407 61 441 95
rect 491 55 525 89
rect 575 129 609 163
rect 575 61 609 95
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 127 443 161 477
rect 218 443 252 477
rect 127 375 161 409
rect 218 375 252 409
rect 379 443 413 477
rect 379 375 413 409
rect 379 307 413 341
rect 575 451 609 485
rect 575 383 609 417
rect 575 315 609 349
<< poly >>
rect 83 497 113 523
rect 262 497 292 523
rect 339 497 369 523
rect 463 497 493 523
rect 535 497 565 523
rect 83 265 113 297
rect 262 265 292 297
rect 78 249 165 265
rect 78 215 121 249
rect 155 215 165 249
rect 78 199 165 215
rect 207 264 292 265
rect 339 265 369 297
rect 463 265 493 297
rect 207 249 297 264
rect 207 215 217 249
rect 251 215 297 249
rect 207 199 297 215
rect 339 249 393 265
rect 339 215 349 249
rect 383 215 393 249
rect 339 199 393 215
rect 435 249 493 265
rect 435 215 449 249
rect 483 215 493 249
rect 435 199 493 215
rect 535 265 565 297
rect 535 249 603 265
rect 535 215 550 249
rect 584 215 603 249
rect 535 199 603 215
rect 79 177 109 199
rect 267 177 297 199
rect 351 177 381 199
rect 451 177 481 199
rect 535 177 565 199
rect 79 21 109 47
rect 267 21 297 47
rect 351 21 381 47
rect 451 21 481 47
rect 535 21 565 47
<< polycont >>
rect 121 215 155 249
rect 217 215 251 249
rect 349 215 383 249
rect 449 215 483 249
rect 550 215 584 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 17 477 73 493
rect 17 443 39 477
rect 17 409 73 443
rect 17 375 39 409
rect 111 477 268 527
rect 111 443 127 477
rect 161 443 218 477
rect 252 443 268 477
rect 111 409 268 443
rect 111 375 127 409
rect 161 375 218 409
rect 252 375 268 409
rect 347 477 424 493
rect 563 485 627 527
rect 347 443 379 477
rect 413 443 424 477
rect 347 409 424 443
rect 347 375 379 409
rect 413 375 424 409
rect 17 341 73 375
rect 347 361 424 375
rect 347 341 429 361
rect 17 307 39 341
rect 17 136 73 307
rect 107 307 379 341
rect 413 307 429 341
rect 489 323 529 481
rect 107 299 429 307
rect 107 249 162 299
rect 463 289 529 323
rect 563 451 575 485
rect 609 451 627 485
rect 563 417 627 451
rect 563 383 575 417
rect 609 383 627 417
rect 563 349 627 383
rect 563 315 575 349
rect 609 315 627 349
rect 563 291 627 315
rect 463 265 499 289
rect 107 215 121 249
rect 155 215 162 249
rect 196 249 267 265
rect 196 215 217 249
rect 251 215 267 249
rect 306 249 399 265
rect 306 215 349 249
rect 383 215 399 249
rect 433 249 499 265
rect 433 215 449 249
rect 483 215 499 249
rect 534 249 627 255
rect 534 215 550 249
rect 584 215 627 249
rect 107 179 162 215
rect 107 163 357 179
rect 107 143 307 163
rect 17 102 35 136
rect 69 102 73 136
rect 284 129 307 143
rect 341 129 357 163
rect 391 163 627 173
rect 391 129 407 163
rect 441 139 575 163
rect 441 129 457 139
rect 17 73 73 102
rect 119 93 153 109
rect 391 95 457 129
rect 559 129 575 139
rect 609 129 627 163
rect 207 61 223 95
rect 257 61 407 95
rect 441 61 457 95
rect 207 59 457 61
rect 491 89 525 105
rect 119 17 153 59
rect 559 95 627 129
rect 559 61 575 95
rect 609 61 627 95
rect 559 56 627 61
rect 491 17 525 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel corelocali s 489 357 523 391 0 FreeSans 400 0 0 0 A2
port 2 nsew
flabel corelocali s 29 425 63 459 0 FreeSans 400 0 0 0 X
port 9 nsew
flabel corelocali s 213 221 247 255 0 FreeSans 400 0 0 0 B1
port 3 nsew
flabel corelocali s 581 221 615 255 0 FreeSans 400 0 0 0 A1
port 1 nsew
flabel corelocali s 310 221 344 255 0 FreeSans 400 0 0 0 B2
port 4 nsew
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
rlabel comment s 0 0 0 0 4 o22a_1
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1472796
string GDS_START 1466778
string path 0.000 0.000 3.220 0.000 
<< end >>
