magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 3036 561
rect 103 427 169 527
rect 17 195 87 325
rect 286 377 357 527
rect 659 443 728 527
rect 103 17 169 93
rect 283 205 339 337
rect 387 219 431 339
rect 387 153 467 219
rect 765 265 805 475
rect 286 17 341 127
rect 387 69 429 153
rect 674 17 740 89
rect 1141 441 1217 527
rect 1435 383 1501 527
rect 1924 451 2000 527
rect 1177 193 1243 213
rect 1177 147 1259 193
rect 2188 451 2482 527
rect 1177 17 1211 105
rect 1951 147 2026 213
rect 2516 326 2566 493
rect 2318 219 2414 265
rect 1529 17 1595 93
rect 1912 17 1964 105
rect 2416 17 2482 161
rect 2532 143 2566 326
rect 2600 299 2647 527
rect 2790 353 2849 527
rect 2883 289 2933 493
rect 2967 299 3015 527
rect 2516 51 2566 143
rect 2600 17 2647 177
rect 2892 165 2933 289
rect 2790 17 2849 109
rect 2883 51 2933 165
rect 2967 17 3015 177
rect 0 -17 3036 17
<< obsli1 >>
rect 34 393 69 493
rect 34 359 167 393
rect 121 187 167 359
rect 34 153 121 161
rect 155 153 167 187
rect 34 127 167 153
rect 203 391 247 493
rect 203 357 213 391
rect 443 375 515 477
rect 579 381 613 493
rect 34 69 69 127
rect 203 69 247 357
rect 481 281 515 375
rect 549 349 613 381
rect 549 315 729 349
rect 481 255 615 281
rect 481 250 581 255
rect 487 247 581 250
rect 512 221 581 247
rect 512 215 615 221
rect 695 219 729 315
rect 846 255 891 493
rect 927 450 1093 484
rect 846 221 857 255
rect 512 119 546 215
rect 695 159 754 219
rect 463 53 546 119
rect 591 153 754 159
rect 591 125 729 153
rect 591 61 625 125
rect 846 61 891 221
rect 925 357 949 391
rect 983 357 1025 391
rect 925 315 1025 357
rect 925 141 969 315
rect 1059 281 1093 450
rect 1277 407 1311 475
rect 1127 357 1397 407
rect 1710 450 1876 484
rect 1672 391 1719 397
rect 1127 315 1177 357
rect 1279 281 1329 297
rect 1059 247 1329 281
rect 1059 239 1143 247
rect 1005 187 1075 203
rect 1005 153 1041 187
rect 1005 129 1075 153
rect 1109 93 1143 239
rect 1285 231 1329 247
rect 1363 213 1397 357
rect 1672 357 1685 391
rect 1431 323 1632 331
rect 1431 289 1593 323
rect 1627 289 1632 323
rect 1672 315 1719 357
rect 1431 283 1632 289
rect 1431 247 1497 283
rect 1767 261 1808 381
rect 1684 255 1808 261
rect 1559 213 1625 247
rect 1363 179 1625 213
rect 1684 221 1685 255
rect 1719 225 1808 255
rect 1842 281 1876 450
rect 2048 417 2082 475
rect 1910 383 2482 417
rect 1910 315 1960 383
rect 1842 247 2112 281
rect 1719 221 1741 225
rect 1363 153 1407 179
rect 1341 119 1407 153
rect 940 53 1143 93
rect 1245 85 1311 101
rect 1441 85 1475 143
rect 1684 141 1741 221
rect 1842 93 1876 247
rect 2068 215 2112 247
rect 2146 156 2182 383
rect 2116 119 2182 156
rect 2216 323 2385 349
rect 2216 289 2237 323
rect 2271 315 2385 323
rect 2216 185 2271 289
rect 2448 265 2482 383
rect 2448 199 2496 265
rect 2216 151 2369 185
rect 1245 51 1475 85
rect 1723 53 1876 93
rect 2016 85 2082 109
rect 2216 85 2250 117
rect 2016 51 2250 85
rect 2324 53 2369 151
rect 2691 265 2754 483
rect 2691 199 2858 265
rect 2691 51 2754 199
<< obsli1c >>
rect 121 153 155 187
rect 213 357 247 391
rect 581 221 615 255
rect 857 221 891 255
rect 949 357 983 391
rect 1041 153 1075 187
rect 1685 357 1719 391
rect 1593 289 1627 323
rect 1685 221 1719 255
rect 2237 289 2271 323
<< metal1 >>
rect 0 496 3036 592
rect 1213 184 1271 193
rect 1949 184 2007 193
rect 1213 156 2007 184
rect 1213 147 1271 156
rect 1949 147 2007 156
rect 0 -48 3036 48
<< obsm1 >>
rect 201 391 259 397
rect 201 357 213 391
rect 247 388 259 391
rect 937 391 995 397
rect 937 388 949 391
rect 247 360 949 388
rect 247 357 259 360
rect 201 351 259 357
rect 937 357 949 360
rect 983 388 995 391
rect 1673 391 1731 397
rect 1673 388 1685 391
rect 983 360 1685 388
rect 983 357 995 360
rect 937 351 995 357
rect 1673 357 1685 360
rect 1719 357 1731 391
rect 1673 351 1731 357
rect 1581 323 1639 329
rect 1581 289 1593 323
rect 1627 320 1639 323
rect 2225 323 2283 329
rect 2225 320 2237 323
rect 1627 292 2237 320
rect 1627 289 1639 292
rect 1581 283 1639 289
rect 2225 289 2237 292
rect 2271 289 2283 323
rect 2225 283 2283 289
rect 569 255 627 261
rect 569 221 581 255
rect 615 252 627 255
rect 845 255 903 261
rect 845 252 857 255
rect 615 224 857 252
rect 615 221 627 224
rect 569 215 627 221
rect 845 221 857 224
rect 891 221 903 255
rect 1673 255 1731 261
rect 1673 252 1685 255
rect 845 215 903 221
rect 1044 224 1685 252
rect 1044 193 1087 224
rect 1673 221 1685 224
rect 1719 221 1731 255
rect 1673 215 1731 221
rect 109 187 167 193
rect 109 153 121 187
rect 155 184 167 187
rect 1029 187 1087 193
rect 1029 184 1041 187
rect 155 156 1041 184
rect 155 153 167 156
rect 109 147 167 153
rect 1029 153 1041 156
rect 1075 153 1087 187
rect 1029 147 1087 153
<< labels >>
rlabel locali s 765 265 805 475 6 D
port 1 nsew signal input
rlabel locali s 2892 165 2933 289 6 Q
port 2 nsew signal output
rlabel locali s 2883 289 2933 493 6 Q
port 2 nsew signal output
rlabel locali s 2883 51 2933 165 6 Q
port 2 nsew signal output
rlabel locali s 2532 143 2566 326 6 Q_N
port 3 nsew signal output
rlabel locali s 2516 326 2566 493 6 Q_N
port 3 nsew signal output
rlabel locali s 2516 51 2566 143 6 Q_N
port 3 nsew signal output
rlabel locali s 2318 219 2414 265 6 RESET_B
port 4 nsew signal input
rlabel locali s 283 205 339 337 6 SCD
port 5 nsew signal input
rlabel locali s 387 219 431 339 6 SCE
port 6 nsew signal input
rlabel locali s 387 153 467 219 6 SCE
port 6 nsew signal input
rlabel locali s 387 69 429 153 6 SCE
port 6 nsew signal input
rlabel locali s 1177 193 1243 213 6 SET_B
port 7 nsew signal input
rlabel locali s 1177 147 1259 193 6 SET_B
port 7 nsew signal input
rlabel locali s 1951 147 2026 213 6 SET_B
port 7 nsew signal input
rlabel metal1 s 1949 184 2007 193 6 SET_B
port 7 nsew signal input
rlabel metal1 s 1949 147 2007 156 6 SET_B
port 7 nsew signal input
rlabel metal1 s 1213 184 1271 193 6 SET_B
port 7 nsew signal input
rlabel metal1 s 1213 156 2007 184 6 SET_B
port 7 nsew signal input
rlabel metal1 s 1213 147 1271 156 6 SET_B
port 7 nsew signal input
rlabel locali s 17 195 87 325 6 CLK_N
port 8 nsew clock input
rlabel locali s 2967 17 3015 177 6 VGND
port 9 nsew ground bidirectional abutment
rlabel locali s 2790 17 2849 109 6 VGND
port 9 nsew ground bidirectional abutment
rlabel locali s 2600 17 2647 177 6 VGND
port 9 nsew ground bidirectional abutment
rlabel locali s 2416 17 2482 161 6 VGND
port 9 nsew ground bidirectional abutment
rlabel locali s 1912 17 1964 105 6 VGND
port 9 nsew ground bidirectional abutment
rlabel locali s 1529 17 1595 93 6 VGND
port 9 nsew ground bidirectional abutment
rlabel locali s 1177 17 1211 105 6 VGND
port 9 nsew ground bidirectional abutment
rlabel locali s 674 17 740 89 6 VGND
port 9 nsew ground bidirectional abutment
rlabel locali s 286 17 341 127 6 VGND
port 9 nsew ground bidirectional abutment
rlabel locali s 103 17 169 93 6 VGND
port 9 nsew ground bidirectional abutment
rlabel locali s 0 -17 3036 17 8 VGND
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 3036 48 8 VGND
port 9 nsew ground bidirectional abutment
rlabel locali s 2967 299 3015 527 6 VPWR
port 10 nsew power bidirectional abutment
rlabel locali s 2790 353 2849 527 6 VPWR
port 10 nsew power bidirectional abutment
rlabel locali s 2600 299 2647 527 6 VPWR
port 10 nsew power bidirectional abutment
rlabel locali s 2188 451 2482 527 6 VPWR
port 10 nsew power bidirectional abutment
rlabel locali s 1924 451 2000 527 6 VPWR
port 10 nsew power bidirectional abutment
rlabel locali s 1435 383 1501 527 6 VPWR
port 10 nsew power bidirectional abutment
rlabel locali s 1141 441 1217 527 6 VPWR
port 10 nsew power bidirectional abutment
rlabel locali s 659 443 728 527 6 VPWR
port 10 nsew power bidirectional abutment
rlabel locali s 286 377 357 527 6 VPWR
port 10 nsew power bidirectional abutment
rlabel locali s 103 427 169 527 6 VPWR
port 10 nsew power bidirectional abutment
rlabel locali s 0 527 3036 561 6 VPWR
port 10 nsew power bidirectional abutment
rlabel metal1 s 0 496 3036 592 6 VPWR
port 10 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 3036 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 264324
string GDS_START 240950
<< end >>
