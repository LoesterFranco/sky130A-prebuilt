magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1564 561
rect 103 427 169 527
rect 17 197 65 325
rect 103 17 169 93
rect 391 367 454 527
rect 751 427 918 527
rect 292 191 358 265
rect 1024 387 1178 527
rect 890 199 1087 265
rect 375 17 441 89
rect 747 17 814 106
rect 1024 17 1178 97
rect 1212 51 1282 493
rect 1402 367 1461 527
rect 1495 357 1547 493
rect 1513 119 1547 357
rect 1395 17 1461 93
rect 1495 51 1547 119
rect 0 -17 1564 17
<< obsli1 >>
rect 17 393 69 493
rect 17 359 156 393
rect 122 323 156 359
rect 122 280 156 289
rect 203 391 248 493
rect 203 357 214 391
rect 203 337 248 357
rect 122 214 168 280
rect 122 161 156 214
rect 17 127 156 161
rect 17 69 69 127
rect 203 69 237 337
rect 291 333 357 483
rect 549 451 717 485
rect 654 425 717 451
rect 661 415 717 425
rect 679 409 717 415
rect 679 403 721 409
rect 585 391 626 399
rect 683 398 721 403
rect 684 395 721 398
rect 686 392 721 395
rect 619 381 626 391
rect 619 357 653 381
rect 291 299 428 333
rect 394 219 428 299
rect 494 323 551 337
rect 528 289 551 323
rect 494 271 551 289
rect 585 315 653 357
rect 394 157 468 219
rect 585 207 619 315
rect 687 265 721 392
rect 956 373 990 487
rect 768 353 990 373
rect 768 307 1178 353
rect 687 233 840 265
rect 307 153 468 157
rect 520 153 619 207
rect 666 199 840 233
rect 307 123 428 153
rect 307 69 341 123
rect 666 107 700 199
rect 1131 165 1178 307
rect 554 73 700 107
rect 848 131 1178 165
rect 848 51 908 131
rect 1316 265 1366 493
rect 1316 199 1479 265
rect 1316 51 1361 199
<< obsli1c >>
rect 122 289 156 323
rect 214 357 248 391
rect 585 357 619 391
rect 494 289 528 323
<< metal1 >>
rect 0 496 1564 592
rect 0 -48 1564 48
<< obsm1 >>
rect 202 391 260 397
rect 202 357 214 391
rect 248 388 260 391
rect 573 391 631 397
rect 573 388 585 391
rect 248 360 585 388
rect 248 357 260 360
rect 202 351 260 357
rect 573 357 585 360
rect 619 357 631 391
rect 573 351 631 357
rect 110 323 168 329
rect 110 289 122 323
rect 156 320 168 323
rect 482 323 540 329
rect 482 320 494 323
rect 156 292 494 320
rect 156 289 168 292
rect 110 283 168 289
rect 482 289 494 292
rect 528 289 540 323
rect 482 283 540 289
<< labels >>
rlabel locali s 292 191 358 265 6 D
port 1 nsew signal input
rlabel locali s 1212 51 1282 493 6 Q
port 2 nsew signal output
rlabel locali s 1513 119 1547 357 6 Q_N
port 3 nsew signal output
rlabel locali s 1495 357 1547 493 6 Q_N
port 3 nsew signal output
rlabel locali s 1495 51 1547 119 6 Q_N
port 3 nsew signal output
rlabel locali s 890 199 1087 265 6 RESET_B
port 4 nsew signal input
rlabel locali s 17 197 65 325 6 GATE
port 5 nsew clock input
rlabel locali s 1395 17 1461 93 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1024 17 1178 97 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 747 17 814 106 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 375 17 441 89 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 103 17 169 93 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 1564 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1564 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1402 367 1461 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1024 387 1178 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 751 427 918 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 391 367 454 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 103 427 169 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 1564 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 1564 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1564 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2625894
string GDS_START 2612670
<< end >>
