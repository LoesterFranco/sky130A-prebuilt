magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 125 323 175 425
rect 313 323 363 425
rect 125 289 371 323
rect 789 289 1282 323
rect 331 255 371 289
rect 789 265 833 289
rect 18 215 287 255
rect 331 219 719 255
rect 331 181 371 219
rect 107 145 371 181
rect 107 51 183 145
rect 295 51 371 145
rect 675 164 719 219
rect 753 199 833 265
rect 867 199 1177 255
rect 1213 215 1282 289
rect 1317 289 1827 323
rect 1317 215 1393 289
rect 1793 255 1827 289
rect 1429 215 1751 255
rect 1793 215 2080 255
rect 1222 164 1426 181
rect 675 147 1717 164
rect 675 129 1256 147
rect 1392 129 1717 147
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 18 459 465 493
rect 18 289 81 459
rect 219 357 269 459
rect 415 323 465 459
rect 513 443 1331 493
rect 1365 443 1817 527
rect 513 359 563 443
rect 1281 409 1331 443
rect 1855 409 1889 493
rect 607 367 1237 409
rect 607 323 666 367
rect 1281 357 1905 409
rect 1949 359 1983 527
rect 1871 323 1905 357
rect 2035 323 2085 493
rect 415 289 666 323
rect 23 17 73 179
rect 227 17 261 111
rect 415 129 641 185
rect 1871 289 2085 323
rect 1761 145 1999 181
rect 415 17 449 129
rect 607 119 641 129
rect 487 85 572 95
rect 667 85 1237 95
rect 487 51 1237 85
rect 1291 17 1325 111
rect 1761 95 1811 145
rect 1359 51 1811 95
rect 1855 17 1889 111
rect 1923 51 1999 145
rect 2033 17 2067 181
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
<< metal1 >>
rect 0 561 2116 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 0 496 2116 527
rect 0 17 2116 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
rect 0 -48 2116 -17
<< labels >>
rlabel locali s 1429 215 1751 255 6 A1
port 1 nsew signal input
rlabel locali s 1793 255 1827 289 6 A2
port 2 nsew signal input
rlabel locali s 1793 215 2080 255 6 A2
port 2 nsew signal input
rlabel locali s 1317 289 1827 323 6 A2
port 2 nsew signal input
rlabel locali s 1317 215 1393 289 6 A2
port 2 nsew signal input
rlabel locali s 867 199 1177 255 6 B1
port 3 nsew signal input
rlabel locali s 1213 215 1282 289 6 B2
port 4 nsew signal input
rlabel locali s 789 289 1282 323 6 B2
port 4 nsew signal input
rlabel locali s 789 265 833 289 6 B2
port 4 nsew signal input
rlabel locali s 753 199 833 265 6 B2
port 4 nsew signal input
rlabel locali s 18 215 287 255 6 C1
port 5 nsew signal input
rlabel locali s 1392 129 1717 147 6 Y
port 6 nsew signal output
rlabel locali s 1222 164 1426 181 6 Y
port 6 nsew signal output
rlabel locali s 675 164 719 219 6 Y
port 6 nsew signal output
rlabel locali s 675 147 1717 164 6 Y
port 6 nsew signal output
rlabel locali s 675 129 1256 147 6 Y
port 6 nsew signal output
rlabel locali s 331 255 371 289 6 Y
port 6 nsew signal output
rlabel locali s 331 219 719 255 6 Y
port 6 nsew signal output
rlabel locali s 331 181 371 219 6 Y
port 6 nsew signal output
rlabel locali s 313 323 363 425 6 Y
port 6 nsew signal output
rlabel locali s 295 51 371 145 6 Y
port 6 nsew signal output
rlabel locali s 125 323 175 425 6 Y
port 6 nsew signal output
rlabel locali s 125 289 371 323 6 Y
port 6 nsew signal output
rlabel locali s 107 145 371 181 6 Y
port 6 nsew signal output
rlabel locali s 107 51 183 145 6 Y
port 6 nsew signal output
rlabel metal1 s 0 -48 2116 48 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 496 2116 592 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2116 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1245370
string GDS_START 1231422
<< end >>
