magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 127 424 180 596
rect 314 424 380 596
rect 566 424 632 596
rect 768 430 825 596
rect 768 424 935 430
rect 127 390 935 424
rect 25 270 218 356
rect 286 270 488 356
rect 536 270 743 356
rect 777 270 843 356
rect 889 236 935 390
rect 769 202 935 236
rect 769 129 835 202
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 23 390 90 649
rect 214 458 280 649
rect 416 458 530 649
rect 666 458 732 649
rect 859 464 925 649
rect 23 202 263 236
rect 23 70 89 202
rect 123 17 189 168
rect 229 85 263 202
rect 299 202 663 236
rect 299 119 365 202
rect 399 85 465 168
rect 229 51 465 85
rect 511 85 563 168
rect 597 129 663 202
rect 697 85 735 226
rect 869 85 935 168
rect 511 51 935 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
rlabel locali s 777 270 843 356 6 A
port 1 nsew signal input
rlabel locali s 536 270 743 356 6 B
port 2 nsew signal input
rlabel locali s 286 270 488 356 6 C
port 3 nsew signal input
rlabel locali s 25 270 218 356 6 D
port 4 nsew signal input
rlabel locali s 889 236 935 390 6 Y
port 5 nsew signal output
rlabel locali s 769 202 935 236 6 Y
port 5 nsew signal output
rlabel locali s 769 129 835 202 6 Y
port 5 nsew signal output
rlabel locali s 768 430 825 596 6 Y
port 5 nsew signal output
rlabel locali s 768 424 935 430 6 Y
port 5 nsew signal output
rlabel locali s 566 424 632 596 6 Y
port 5 nsew signal output
rlabel locali s 314 424 380 596 6 Y
port 5 nsew signal output
rlabel locali s 127 424 180 596 6 Y
port 5 nsew signal output
rlabel locali s 127 390 935 424 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -49 960 49 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 617 960 715 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1771812
string GDS_START 1762890
<< end >>
