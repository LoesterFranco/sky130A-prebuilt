magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 85 204 167 246
rect 217 238 333 369
rect 490 287 556 430
rect 658 270 737 356
rect 375 204 441 246
rect 85 170 441 204
rect 85 162 167 170
rect 2221 364 2287 596
rect 2243 210 2277 364
rect 2211 70 2277 210
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2400 683
rect 17 437 89 585
rect 123 471 189 649
rect 297 524 412 589
rect 537 558 627 649
rect 780 558 874 649
rect 1027 524 1077 596
rect 297 490 1077 524
rect 1111 504 1183 596
rect 1317 504 1367 649
rect 1401 581 1571 615
rect 297 471 624 490
rect 17 403 442 437
rect 17 294 183 403
rect 17 128 51 294
rect 376 355 442 403
rect 590 253 624 471
rect 668 390 829 456
rect 475 219 624 253
rect 771 260 829 390
rect 863 294 897 490
rect 931 364 1075 456
rect 1009 322 1075 364
rect 1111 360 1145 504
rect 1401 460 1435 581
rect 1179 426 1435 460
rect 1179 394 1245 426
rect 1369 360 1435 392
rect 1111 326 1435 360
rect 863 260 975 294
rect 771 236 805 260
rect 475 136 509 219
rect 661 202 805 236
rect 661 184 695 202
rect 17 78 98 128
rect 132 17 198 128
rect 296 70 509 136
rect 543 17 595 162
rect 629 66 695 184
rect 741 17 807 168
rect 841 85 907 226
rect 941 188 975 260
rect 941 119 1003 188
rect 1037 85 1071 322
rect 1111 188 1155 326
rect 1469 278 1503 522
rect 1537 386 1571 581
rect 1605 532 1655 584
rect 1605 498 1812 532
rect 1859 518 1985 649
rect 1657 398 1744 464
rect 1778 449 1812 498
rect 2019 483 2089 584
rect 1778 415 2021 449
rect 1537 320 1623 386
rect 1105 119 1155 188
rect 1189 178 1255 272
rect 1297 246 1503 278
rect 1657 272 1691 398
rect 1297 212 1578 246
rect 1189 144 1478 178
rect 1189 85 1223 144
rect 841 51 1223 85
rect 1344 17 1410 110
rect 1444 85 1478 144
rect 1512 119 1578 212
rect 1612 206 1691 272
rect 1612 85 1646 206
rect 1778 162 1812 415
rect 1846 248 1907 381
rect 1955 282 2021 415
rect 2055 310 2089 483
rect 2131 364 2181 649
rect 2327 364 2377 649
rect 2055 248 2209 310
rect 1846 244 2209 248
rect 1846 214 2089 244
rect 1444 51 1646 85
rect 1680 128 1812 162
rect 1680 70 1759 128
rect 1860 17 1926 162
rect 1960 70 2026 214
rect 2123 17 2177 210
rect 2311 17 2377 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2400 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
<< metal1 >>
rect 0 683 2400 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2400 683
rect 0 617 2400 649
rect 0 17 2400 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2400 17
rect 0 -49 2400 -17
<< labels >>
rlabel locali s 217 238 333 369 6 D
port 1 nsew signal input
rlabel locali s 2243 210 2277 364 6 Q
port 2 nsew signal output
rlabel locali s 2221 364 2287 596 6 Q
port 2 nsew signal output
rlabel locali s 2211 70 2277 210 6 Q
port 2 nsew signal output
rlabel locali s 490 287 556 430 6 SCD
port 3 nsew signal input
rlabel locali s 375 204 441 246 6 SCE
port 4 nsew signal input
rlabel locali s 85 204 167 246 6 SCE
port 4 nsew signal input
rlabel locali s 85 170 441 204 6 SCE
port 4 nsew signal input
rlabel locali s 85 162 167 170 6 SCE
port 4 nsew signal input
rlabel locali s 658 270 737 356 6 CLK
port 5 nsew clock input
rlabel metal1 s 0 -49 2400 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 2400 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2400 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 314198
string GDS_START 297156
<< end >>
