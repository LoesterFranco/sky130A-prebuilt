magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 25 290 182 356
rect 294 364 366 596
rect 332 226 366 364
rect 295 70 366 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 384 683
rect 94 424 160 596
rect 194 458 260 649
rect 94 390 260 424
rect 226 326 260 390
rect 226 260 298 326
rect 226 256 260 260
rect 23 222 260 256
rect 23 160 159 222
rect 195 17 261 188
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 384 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
<< metal1 >>
rect 0 683 384 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 384 683
rect 0 617 384 649
rect 0 17 384 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 384 17
rect 0 -49 384 -17
<< labels >>
rlabel locali s 25 290 182 356 6 A
port 1 nsew signal input
rlabel locali s 332 226 366 364 6 X
port 2 nsew signal output
rlabel locali s 295 70 366 226 6 X
port 2 nsew signal output
rlabel locali s 294 364 366 596 6 X
port 2 nsew signal output
rlabel metal1 s 0 -49 384 49 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 617 384 715 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 384 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3145768
string GDS_START 3141446
<< end >>
