magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 217 306 286 360
rect 880 272 1014 356
rect 1359 344 1425 596
rect 1549 356 1599 596
rect 1549 344 1703 356
rect 1359 310 1703 344
rect 1561 276 1603 310
rect 1367 242 1603 276
rect 1367 70 1433 242
rect 1553 70 1603 242
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 23 364 108 596
rect 157 462 232 649
rect 622 572 688 649
rect 287 504 497 570
rect 841 538 907 594
rect 661 504 907 538
rect 287 428 321 504
rect 661 470 695 504
rect 142 394 321 428
rect 355 410 695 470
rect 729 436 799 470
rect 23 204 73 364
rect 142 310 176 394
rect 107 272 176 310
rect 107 238 321 272
rect 23 170 253 204
rect 23 70 73 170
rect 110 17 185 136
rect 219 85 253 170
rect 287 196 321 238
rect 355 230 413 410
rect 661 392 695 410
rect 461 306 527 361
rect 661 340 731 392
rect 765 322 799 436
rect 841 418 907 504
rect 948 418 1014 649
rect 1048 398 1114 596
rect 1148 432 1325 649
rect 1048 364 1270 398
rect 765 306 831 322
rect 461 272 831 306
rect 1052 260 1161 326
rect 1052 238 1086 260
rect 563 204 1086 238
rect 1195 226 1270 364
rect 1459 378 1509 649
rect 1639 390 1705 649
rect 287 130 466 196
rect 563 85 629 204
rect 219 51 629 85
rect 663 17 729 170
rect 856 103 922 170
rect 763 51 922 103
rect 956 17 1022 170
rect 1120 134 1270 226
rect 1120 70 1195 134
rect 1232 17 1331 100
rect 1467 17 1517 208
rect 1639 17 1705 208
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
<< metal1 >>
rect 0 683 1728 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 0 617 1728 649
rect 0 17 1728 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
rect 0 -49 1728 -17
<< labels >>
rlabel locali s 217 306 286 360 6 GATE
port 1 nsew signal input
rlabel locali s 1561 276 1603 310 6 GCLK
port 2 nsew signal output
rlabel locali s 1553 70 1603 242 6 GCLK
port 2 nsew signal output
rlabel locali s 1549 356 1599 596 6 GCLK
port 2 nsew signal output
rlabel locali s 1549 344 1703 356 6 GCLK
port 2 nsew signal output
rlabel locali s 1367 242 1603 276 6 GCLK
port 2 nsew signal output
rlabel locali s 1367 70 1433 242 6 GCLK
port 2 nsew signal output
rlabel locali s 1359 344 1425 596 6 GCLK
port 2 nsew signal output
rlabel locali s 1359 310 1703 344 6 GCLK
port 2 nsew signal output
rlabel locali s 880 272 1014 356 6 CLK
port 3 nsew clock input
rlabel metal1 s 0 -49 1728 49 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 617 1728 715 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1728 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3043358
string GDS_START 3030404
<< end >>
