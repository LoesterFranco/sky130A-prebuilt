magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1472 561
rect 17 297 69 493
rect 103 430 153 527
rect 460 455 526 527
rect 648 451 714 527
rect 816 455 882 527
rect 1268 455 1334 527
rect 17 166 52 297
rect 260 289 340 376
rect 374 319 592 353
rect 182 255 216 265
rect 374 255 408 319
rect 182 199 248 255
rect 334 221 408 255
rect 446 206 524 272
rect 558 250 592 319
rect 640 287 712 353
rect 1031 337 1081 391
rect 757 303 1081 337
rect 757 250 791 303
rect 1127 289 1211 353
rect 1368 297 1448 493
rect 17 51 69 166
rect 558 193 791 250
rect 850 191 925 255
rect 1177 207 1265 255
rect 103 17 169 93
rect 460 17 526 89
rect 1382 162 1448 297
rect 648 17 714 98
rect 816 17 882 89
rect 1253 17 1319 89
rect 1368 51 1448 162
rect 0 -17 1472 17
<< obsli1 >>
rect 187 413 342 493
rect 392 421 426 493
rect 560 421 607 493
rect 187 389 221 413
rect 103 325 221 389
rect 392 387 607 421
rect 748 421 782 493
rect 916 421 950 493
rect 1017 425 1234 493
rect 748 387 950 421
rect 1200 421 1234 425
rect 103 265 137 325
rect 86 199 137 265
rect 1200 387 1333 421
rect 1299 265 1333 387
rect 103 161 137 199
rect 959 191 1092 225
rect 993 187 1092 191
rect 294 161 306 187
rect 103 153 306 161
rect 340 153 342 187
rect 103 127 342 153
rect 222 51 342 127
rect 392 123 594 157
rect 392 51 426 123
rect 560 51 594 123
rect 748 123 950 157
rect 993 153 1046 187
rect 1080 153 1092 187
rect 1299 199 1348 265
rect 1299 157 1333 199
rect 748 51 782 123
rect 916 51 950 123
rect 1185 123 1333 157
rect 1017 101 1051 119
rect 1185 101 1219 123
rect 1017 51 1219 101
<< obsli1c >>
rect 306 153 340 187
rect 1046 153 1080 187
<< metal1 >>
rect 0 496 1472 592
rect 294 320 352 329
rect 666 320 724 329
rect 1126 320 1184 329
rect 294 292 1184 320
rect 294 283 352 292
rect 666 283 724 292
rect 1126 283 1184 292
rect 202 252 260 261
rect 478 252 536 261
rect 850 252 908 261
rect 1218 252 1276 261
rect 202 224 1276 252
rect 202 215 260 224
rect 478 215 536 224
rect 850 215 908 224
rect 1218 215 1276 224
rect 0 -48 1472 48
<< obsm1 >>
rect 294 187 352 193
rect 294 153 306 187
rect 340 184 352 187
rect 1034 187 1092 193
rect 1034 184 1046 187
rect 340 156 1046 184
rect 340 153 352 156
rect 294 147 352 153
rect 1034 153 1046 156
rect 1080 153 1092 187
rect 1034 147 1092 153
<< labels >>
rlabel locali s 182 255 216 265 6 A
port 1 nsew signal input
rlabel locali s 182 199 248 255 6 A
port 1 nsew signal input
rlabel locali s 446 206 524 272 6 A
port 1 nsew signal input
rlabel locali s 850 191 925 255 6 A
port 1 nsew signal input
rlabel locali s 1177 207 1265 255 6 A
port 1 nsew signal input
rlabel metal1 s 1218 252 1276 261 6 A
port 1 nsew signal input
rlabel metal1 s 1218 215 1276 224 6 A
port 1 nsew signal input
rlabel metal1 s 850 252 908 261 6 A
port 1 nsew signal input
rlabel metal1 s 850 215 908 224 6 A
port 1 nsew signal input
rlabel metal1 s 478 252 536 261 6 A
port 1 nsew signal input
rlabel metal1 s 478 215 536 224 6 A
port 1 nsew signal input
rlabel metal1 s 202 252 260 261 6 A
port 1 nsew signal input
rlabel metal1 s 202 224 1276 252 6 A
port 1 nsew signal input
rlabel metal1 s 202 215 260 224 6 A
port 1 nsew signal input
rlabel locali s 260 289 340 376 6 B
port 2 nsew signal input
rlabel locali s 640 287 712 353 6 B
port 2 nsew signal input
rlabel locali s 1127 289 1211 353 6 B
port 2 nsew signal input
rlabel metal1 s 1126 320 1184 329 6 B
port 2 nsew signal input
rlabel metal1 s 1126 283 1184 292 6 B
port 2 nsew signal input
rlabel metal1 s 666 320 724 329 6 B
port 2 nsew signal input
rlabel metal1 s 666 283 724 292 6 B
port 2 nsew signal input
rlabel metal1 s 294 320 352 329 6 B
port 2 nsew signal input
rlabel metal1 s 294 292 1184 320 6 B
port 2 nsew signal input
rlabel metal1 s 294 283 352 292 6 B
port 2 nsew signal input
rlabel locali s 1031 337 1081 391 6 CIN
port 3 nsew signal input
rlabel locali s 757 303 1081 337 6 CIN
port 3 nsew signal input
rlabel locali s 757 250 791 303 6 CIN
port 3 nsew signal input
rlabel locali s 558 250 592 319 6 CIN
port 3 nsew signal input
rlabel locali s 558 193 791 250 6 CIN
port 3 nsew signal input
rlabel locali s 374 319 592 353 6 CIN
port 3 nsew signal input
rlabel locali s 374 255 408 319 6 CIN
port 3 nsew signal input
rlabel locali s 334 221 408 255 6 CIN
port 3 nsew signal input
rlabel locali s 17 297 69 493 6 COUT
port 4 nsew signal output
rlabel locali s 17 166 52 297 6 COUT
port 4 nsew signal output
rlabel locali s 17 51 69 166 6 COUT
port 4 nsew signal output
rlabel locali s 1382 162 1448 297 6 SUM
port 5 nsew signal output
rlabel locali s 1368 297 1448 493 6 SUM
port 5 nsew signal output
rlabel locali s 1368 51 1448 162 6 SUM
port 5 nsew signal output
rlabel locali s 1253 17 1319 89 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 816 17 882 89 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 648 17 714 98 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 460 17 526 89 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 103 17 169 93 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 1472 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1472 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1268 455 1334 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 816 455 882 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 648 451 714 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 460 455 526 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 103 430 153 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 1472 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 1472 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1472 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2019070
string GDS_START 2006120
<< end >>
