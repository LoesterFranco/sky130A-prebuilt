magic
tech sky130A
magscale 1 2
timestamp 1599588232
<< locali >>
rect 25 260 101 356
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2592 683
rect 23 424 89 596
rect 129 458 163 649
rect 23 390 169 424
rect 135 326 169 390
rect 203 394 269 596
rect 309 428 343 649
rect 383 394 449 596
rect 203 360 449 394
rect 498 364 548 649
rect 588 398 654 596
rect 694 432 728 649
rect 768 398 834 596
rect 874 432 908 649
rect 950 398 1016 596
rect 588 364 1016 398
rect 1056 385 1090 649
rect 1132 424 1198 596
rect 1132 390 1152 424
rect 1186 390 1198 424
rect 1132 384 1198 390
rect 1232 385 1282 649
rect 1322 424 1388 596
rect 1322 390 1335 424
rect 1369 390 1388 424
rect 1322 384 1388 390
rect 1428 385 1462 649
rect 1502 424 1568 596
rect 1502 390 1519 424
rect 1553 390 1568 424
rect 1502 384 1568 390
rect 1608 385 1642 649
rect 1682 424 1748 596
rect 1682 390 1697 424
rect 1731 390 1748 424
rect 1682 384 1748 390
rect 1788 385 1822 649
rect 1862 424 1928 596
rect 1862 390 1881 424
rect 1915 390 1928 424
rect 1862 384 1928 390
rect 1968 385 2002 649
rect 2042 424 2108 596
rect 2042 390 2059 424
rect 2093 390 2108 424
rect 2042 384 2108 390
rect 2148 385 2182 649
rect 2222 424 2288 596
rect 2222 390 2239 424
rect 2273 390 2288 424
rect 2222 384 2288 390
rect 2328 385 2378 649
rect 2412 424 2478 596
rect 2412 390 2423 424
rect 2457 404 2478 424
rect 2457 390 2469 404
rect 1132 380 1177 384
rect 409 330 449 360
rect 969 351 1016 364
rect 969 350 1081 351
rect 135 260 375 326
rect 409 264 896 330
rect 969 316 1036 350
rect 1070 316 1081 350
rect 969 264 1081 316
rect 135 226 169 260
rect 409 226 443 264
rect 969 230 1021 264
rect 26 192 169 226
rect 214 192 443 226
rect 26 70 76 192
rect 112 17 178 158
rect 214 70 248 192
rect 284 17 334 158
rect 371 70 443 192
rect 483 17 549 226
rect 583 196 1021 230
rect 583 70 633 196
rect 669 17 735 162
rect 769 70 819 196
rect 855 17 921 162
rect 955 70 1005 196
rect 1055 17 1091 226
rect 1127 70 1177 380
rect 1211 316 1225 350
rect 1259 316 1273 350
rect 1322 330 1356 384
rect 1211 264 1273 316
rect 1213 17 1263 226
rect 1307 70 1356 330
rect 1390 316 1400 350
rect 1434 316 1443 350
rect 1502 330 1536 384
rect 1390 264 1443 316
rect 1392 17 1435 226
rect 1477 70 1536 330
rect 1570 316 1580 350
rect 1614 316 1623 350
rect 1682 330 1716 384
rect 1570 264 1623 316
rect 1570 17 1623 226
rect 1657 70 1716 330
rect 1750 316 1764 350
rect 1798 316 1809 350
rect 1862 330 1896 384
rect 1750 264 1809 316
rect 1750 17 1809 226
rect 1843 70 1896 330
rect 1930 316 1946 350
rect 1980 316 1995 350
rect 2042 330 2079 384
rect 1930 264 1995 316
rect 1933 17 1995 226
rect 2029 70 2079 330
rect 2113 316 2135 350
rect 2169 316 2188 350
rect 2113 264 2188 316
rect 2115 17 2181 226
rect 2222 70 2265 384
rect 2299 316 2320 350
rect 2354 316 2378 350
rect 2299 264 2378 316
rect 2412 230 2469 390
rect 2518 364 2568 649
rect 2301 17 2367 226
rect 2403 70 2469 230
rect 2503 17 2569 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2592 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 1152 390 1186 424
rect 1335 390 1369 424
rect 1519 390 1553 424
rect 1697 390 1731 424
rect 1881 390 1915 424
rect 2059 390 2093 424
rect 2239 390 2273 424
rect 2423 390 2457 424
rect 1036 316 1070 350
rect 1225 316 1259 350
rect 1400 316 1434 350
rect 1580 316 1614 350
rect 1764 316 1798 350
rect 1946 316 1980 350
rect 2135 316 2169 350
rect 2320 316 2354 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
<< metal1 >>
rect 0 683 2592 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2592 683
rect 0 617 2592 649
rect 0 616 50 617
rect 1140 424 2476 430
rect 1140 390 1152 424
rect 1186 390 1335 424
rect 1369 390 1519 424
rect 1553 390 1697 424
rect 1731 390 1881 424
rect 1915 390 2059 424
rect 2093 390 2239 424
rect 2273 390 2423 424
rect 2457 390 2476 424
rect 1140 384 2476 390
rect 0 49 50 50
rect 0 17 2592 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2592 17
rect 0 -49 2592 -17
<< obsm1 >>
rect 1022 350 2366 356
rect 1022 316 1036 350
rect 1070 316 1225 350
rect 1259 316 1400 350
rect 1434 316 1580 350
rect 1614 316 1764 350
rect 1798 316 1946 350
rect 1980 316 2135 350
rect 2169 316 2320 350
rect 2354 316 2366 350
rect 1022 310 2366 316
<< labels >>
rlabel locali s 25 260 101 356 6 A
port 1 nsew signal input
rlabel metal1 s 1140 384 2476 430 6 X
port 2 nsew signal output
rlabel metal1 s 0 -49 2592 49 8 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 4 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 617 2592 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2592 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3449722
string GDS_START 3428542
<< end >>
