magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1196 561
rect 27 360 79 527
rect 113 326 161 487
rect 195 360 247 527
rect 281 326 329 487
rect 363 360 415 527
rect 449 326 499 487
rect 533 360 582 527
rect 616 326 665 487
rect 699 360 750 527
rect 784 326 835 487
rect 869 360 919 527
rect 953 326 1001 487
rect 1035 360 1086 527
rect 23 292 1088 326
rect 23 173 57 292
rect 91 207 973 258
rect 1034 173 1088 292
rect 23 139 1088 173
rect 207 17 273 105
rect 307 56 345 139
rect 379 17 445 105
rect 479 56 517 139
rect 551 17 617 105
rect 651 56 689 139
rect 723 17 789 105
rect 823 56 861 139
rect 895 17 961 105
rect 0 -17 1196 17
<< metal1 >>
rect 0 496 1196 592
rect 0 -48 1196 48
<< labels >>
rlabel locali s 91 207 973 258 6 A
port 1 nsew signal input
rlabel locali s 1034 173 1088 292 6 Y
port 2 nsew signal output
rlabel locali s 953 326 1001 487 6 Y
port 2 nsew signal output
rlabel locali s 823 56 861 139 6 Y
port 2 nsew signal output
rlabel locali s 784 326 835 487 6 Y
port 2 nsew signal output
rlabel locali s 651 56 689 139 6 Y
port 2 nsew signal output
rlabel locali s 616 326 665 487 6 Y
port 2 nsew signal output
rlabel locali s 479 56 517 139 6 Y
port 2 nsew signal output
rlabel locali s 449 326 499 487 6 Y
port 2 nsew signal output
rlabel locali s 307 56 345 139 6 Y
port 2 nsew signal output
rlabel locali s 281 326 329 487 6 Y
port 2 nsew signal output
rlabel locali s 113 326 161 487 6 Y
port 2 nsew signal output
rlabel locali s 23 292 1088 326 6 Y
port 2 nsew signal output
rlabel locali s 23 173 57 292 6 Y
port 2 nsew signal output
rlabel locali s 23 139 1088 173 6 Y
port 2 nsew signal output
rlabel locali s 895 17 961 105 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 723 17 789 105 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 551 17 617 105 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 379 17 445 105 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 207 17 273 105 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 0 -17 1196 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1196 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1035 360 1086 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 869 360 919 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 699 360 750 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 533 360 582 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 363 360 415 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 195 360 247 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 27 360 79 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 0 527 1196 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 496 1196 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3234598
string GDS_START 3225408
<< end >>
