magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 113 404 163 596
rect 303 404 359 600
rect 113 370 359 404
rect 1036 390 1319 424
rect 113 330 163 370
rect 25 296 163 330
rect 25 236 71 296
rect 501 290 567 356
rect 601 290 743 356
rect 25 186 380 236
rect 123 82 164 186
rect 314 86 380 186
rect 514 85 548 290
rect 1036 358 1070 390
rect 888 294 1070 358
rect 1127 290 1223 356
rect 1285 354 1319 390
rect 1285 288 1365 354
rect 1413 290 1607 356
rect 817 85 883 117
rect 514 51 883 85
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 23 364 73 649
rect 203 438 269 649
rect 393 458 459 649
rect 505 581 985 615
rect 505 458 571 581
rect 605 424 671 547
rect 705 458 771 581
rect 805 424 871 547
rect 403 390 871 424
rect 919 492 985 581
rect 1042 526 1123 649
rect 1157 492 1223 580
rect 1257 526 1329 649
rect 1363 492 1419 600
rect 919 458 1419 492
rect 1453 458 1509 649
rect 919 392 985 458
rect 1353 424 1419 458
rect 1543 424 1609 596
rect 1353 390 1609 424
rect 403 336 437 390
rect 197 270 437 336
rect 23 17 89 152
rect 198 17 280 152
rect 414 17 480 236
rect 777 256 811 390
rect 582 185 648 242
rect 684 222 1226 256
rect 684 219 750 222
rect 582 151 836 185
rect 870 151 951 188
rect 582 119 648 151
rect 917 17 951 151
rect 988 85 1038 188
rect 1074 153 1124 188
rect 1160 187 1226 222
rect 1262 153 1312 254
rect 1074 119 1312 153
rect 1348 220 1609 254
rect 1348 85 1398 220
rect 988 51 1398 85
rect 1438 17 1509 184
rect 1543 118 1609 220
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
rlabel locali s 1127 290 1223 356 6 A1
port 1 nsew signal input
rlabel locali s 1285 354 1319 390 6 A2
port 2 nsew signal input
rlabel locali s 1285 288 1365 354 6 A2
port 2 nsew signal input
rlabel locali s 1036 390 1319 424 6 A2
port 2 nsew signal input
rlabel locali s 1036 358 1070 390 6 A2
port 2 nsew signal input
rlabel locali s 888 294 1070 358 6 A2
port 2 nsew signal input
rlabel locali s 1413 290 1607 356 6 A3
port 3 nsew signal input
rlabel locali s 601 290 743 356 6 B1
port 4 nsew signal input
rlabel locali s 817 85 883 117 6 B2
port 5 nsew signal input
rlabel locali s 514 85 548 290 6 B2
port 5 nsew signal input
rlabel locali s 514 51 883 85 6 B2
port 5 nsew signal input
rlabel locali s 501 290 567 356 6 B2
port 5 nsew signal input
rlabel locali s 314 86 380 186 6 X
port 6 nsew signal output
rlabel locali s 303 404 359 600 6 X
port 6 nsew signal output
rlabel locali s 123 82 164 186 6 X
port 6 nsew signal output
rlabel locali s 113 404 163 596 6 X
port 6 nsew signal output
rlabel locali s 113 370 359 404 6 X
port 6 nsew signal output
rlabel locali s 113 330 163 370 6 X
port 6 nsew signal output
rlabel locali s 25 296 163 330 6 X
port 6 nsew signal output
rlabel locali s 25 236 71 296 6 X
port 6 nsew signal output
rlabel locali s 25 186 380 236 6 X
port 6 nsew signal output
rlabel metal1 s 0 -49 1632 49 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1632 715 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3712628
string GDS_START 3699320
<< end >>
