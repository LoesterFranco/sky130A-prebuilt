magic
tech sky130A
magscale 1 2
timestamp 1599588201
<< nwell >>
rect -38 261 1878 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 418 47 448 131
rect 513 47 543 119
rect 609 47 639 119
rect 775 47 805 131
rect 847 47 877 131
rect 979 47 1009 175
rect 1078 47 1108 119
rect 1187 47 1217 119
rect 1283 47 1313 131
rect 1432 47 1462 131
rect 1523 47 1553 131
rect 1731 47 1761 177
<< pmoshvt >>
rect 79 363 109 491
rect 163 363 193 491
rect 430 413 460 497
rect 522 413 552 497
rect 621 413 651 497
rect 761 413 791 497
rect 858 413 888 497
rect 1055 329 1085 497
rect 1154 413 1184 497
rect 1240 413 1270 497
rect 1324 413 1354 497
rect 1432 413 1462 497
rect 1516 413 1546 497
rect 1731 297 1761 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 313 89 418 131
rect 313 55 325 89
rect 359 55 418 89
rect 313 47 418 55
rect 448 119 498 131
rect 929 131 979 175
rect 657 119 775 131
rect 448 95 513 119
rect 448 61 458 95
rect 492 61 513 95
rect 448 47 513 61
rect 543 95 609 119
rect 543 61 565 95
rect 599 61 609 95
rect 543 47 609 61
rect 639 47 775 119
rect 805 47 847 131
rect 877 93 979 131
rect 877 59 911 93
rect 945 59 979 93
rect 877 47 979 59
rect 1009 119 1063 175
rect 1681 131 1731 177
rect 1233 119 1283 131
rect 1009 89 1078 119
rect 1009 55 1023 89
rect 1057 55 1078 89
rect 1009 47 1078 55
rect 1108 93 1187 119
rect 1108 59 1133 93
rect 1167 59 1187 93
rect 1108 47 1187 59
rect 1217 47 1283 119
rect 1313 89 1432 131
rect 1313 55 1345 89
rect 1379 55 1432 89
rect 1313 47 1432 55
rect 1462 47 1523 131
rect 1553 109 1605 131
rect 1553 75 1563 109
rect 1597 75 1605 109
rect 1553 47 1605 75
rect 1659 93 1731 131
rect 1659 59 1687 93
rect 1721 59 1731 93
rect 1659 47 1731 59
rect 1761 143 1813 177
rect 1761 109 1771 143
rect 1805 109 1813 143
rect 1761 47 1813 109
<< pdiff >>
rect 27 477 79 491
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 363 79 375
rect 109 461 163 491
rect 109 427 119 461
rect 153 427 163 461
rect 109 363 163 427
rect 193 477 245 491
rect 193 443 203 477
rect 237 443 245 477
rect 193 409 245 443
rect 378 485 430 497
rect 378 451 386 485
rect 420 451 430 485
rect 378 413 430 451
rect 460 477 522 497
rect 460 443 470 477
rect 504 443 522 477
rect 460 413 522 443
rect 552 483 621 497
rect 552 449 563 483
rect 597 449 621 483
rect 552 413 621 449
rect 651 459 761 497
rect 651 425 717 459
rect 751 425 761 459
rect 651 413 761 425
rect 791 475 858 497
rect 791 441 814 475
rect 848 441 858 475
rect 791 413 858 441
rect 888 459 940 497
rect 888 425 898 459
rect 932 425 940 459
rect 888 413 940 425
rect 1003 485 1055 497
rect 1003 451 1011 485
rect 1045 451 1055 485
rect 193 375 203 409
rect 237 375 245 409
rect 193 363 245 375
rect 1003 329 1055 451
rect 1085 477 1154 497
rect 1085 443 1099 477
rect 1133 443 1154 477
rect 1085 413 1154 443
rect 1184 484 1240 497
rect 1184 450 1196 484
rect 1230 450 1240 484
rect 1184 413 1240 450
rect 1270 413 1324 497
rect 1354 485 1432 497
rect 1354 451 1388 485
rect 1422 451 1432 485
rect 1354 413 1432 451
rect 1462 459 1516 497
rect 1462 425 1472 459
rect 1506 425 1516 459
rect 1462 413 1516 425
rect 1546 485 1600 497
rect 1546 451 1558 485
rect 1592 451 1600 485
rect 1546 413 1600 451
rect 1665 485 1731 497
rect 1665 451 1687 485
rect 1721 451 1731 485
rect 1665 417 1731 451
rect 1085 329 1139 413
rect 1665 383 1687 417
rect 1721 383 1731 417
rect 1665 369 1731 383
rect 1681 297 1731 369
rect 1761 449 1813 497
rect 1761 415 1771 449
rect 1805 415 1813 449
rect 1761 381 1813 415
rect 1761 347 1771 381
rect 1805 347 1813 381
rect 1761 297 1813 347
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 325 55 359 89
rect 458 61 492 95
rect 565 61 599 95
rect 911 59 945 93
rect 1023 55 1057 89
rect 1133 59 1167 93
rect 1345 55 1379 89
rect 1563 75 1597 109
rect 1687 59 1721 93
rect 1771 109 1805 143
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 427 153 461
rect 203 443 237 477
rect 386 451 420 485
rect 470 443 504 477
rect 563 449 597 483
rect 717 425 751 459
rect 814 441 848 475
rect 898 425 932 459
rect 1011 451 1045 485
rect 203 375 237 409
rect 1099 443 1133 477
rect 1196 450 1230 484
rect 1388 451 1422 485
rect 1472 425 1506 459
rect 1558 451 1592 485
rect 1687 451 1721 485
rect 1687 383 1721 417
rect 1771 415 1805 449
rect 1771 347 1805 381
<< poly >>
rect 79 491 109 517
rect 163 491 193 517
rect 430 497 460 523
rect 522 497 552 523
rect 621 497 651 523
rect 761 497 791 523
rect 858 497 888 523
rect 1055 497 1085 523
rect 1154 497 1184 523
rect 1240 497 1270 523
rect 1324 497 1354 523
rect 1432 497 1462 523
rect 1516 497 1546 523
rect 1731 497 1761 523
rect 79 348 109 363
rect 46 318 109 348
rect 46 265 76 318
rect 163 274 193 363
rect 430 326 460 413
rect 522 375 552 413
rect 22 249 76 265
rect 22 215 32 249
rect 66 215 76 249
rect 118 264 193 274
rect 118 230 134 264
rect 168 230 193 264
rect 331 310 460 326
rect 506 365 572 375
rect 506 331 522 365
rect 556 331 572 365
rect 506 321 572 331
rect 331 276 341 310
rect 375 296 460 310
rect 375 276 448 296
rect 621 279 651 413
rect 761 355 791 413
rect 761 339 816 355
rect 761 305 771 339
rect 805 305 816 339
rect 761 289 816 305
rect 331 260 448 276
rect 118 220 193 230
rect 22 199 76 215
rect 46 176 76 199
rect 46 146 109 176
rect 79 131 109 146
rect 163 131 193 220
rect 418 131 448 260
rect 513 249 651 279
rect 513 219 544 249
rect 490 203 544 219
rect 490 169 500 203
rect 534 169 544 203
rect 490 153 544 169
rect 586 197 652 207
rect 586 163 602 197
rect 636 163 652 197
rect 586 153 652 163
rect 513 119 543 153
rect 609 119 639 153
rect 775 131 805 289
rect 858 219 888 413
rect 1055 314 1085 329
rect 979 284 1085 314
rect 979 267 1009 284
rect 943 251 1009 267
rect 847 203 901 219
rect 847 169 857 203
rect 891 169 901 203
rect 943 217 953 251
rect 987 217 1009 251
rect 1154 279 1184 413
rect 1240 381 1270 413
rect 1226 365 1280 381
rect 1226 331 1236 365
rect 1270 331 1280 365
rect 1226 315 1280 331
rect 1154 267 1204 279
rect 1154 255 1217 267
rect 1154 249 1241 255
rect 1175 239 1241 249
rect 1175 237 1197 239
rect 943 201 1009 217
rect 979 175 1009 201
rect 1078 191 1145 207
rect 847 153 901 169
rect 847 131 877 153
rect 1078 157 1101 191
rect 1135 157 1145 191
rect 1078 141 1145 157
rect 1187 205 1197 237
rect 1231 205 1241 239
rect 1187 189 1241 205
rect 1324 229 1354 413
rect 1432 257 1462 413
rect 1516 365 1546 413
rect 1504 349 1558 365
rect 1504 315 1514 349
rect 1548 315 1558 349
rect 1504 299 1558 315
rect 1427 241 1481 257
rect 1324 213 1385 229
rect 1324 193 1341 213
rect 1078 119 1108 141
rect 1187 119 1217 189
rect 1283 179 1341 193
rect 1375 179 1385 213
rect 1427 207 1437 241
rect 1471 207 1481 241
rect 1427 191 1481 207
rect 1283 163 1385 179
rect 1283 131 1313 163
rect 1432 131 1462 191
rect 1523 131 1553 299
rect 1731 265 1761 297
rect 1702 249 1761 265
rect 1702 215 1712 249
rect 1746 215 1761 249
rect 1702 199 1761 215
rect 1731 177 1761 199
rect 79 21 109 47
rect 163 21 193 47
rect 418 21 448 47
rect 513 21 543 47
rect 609 21 639 47
rect 775 21 805 47
rect 847 21 877 47
rect 979 21 1009 47
rect 1078 21 1108 47
rect 1187 21 1217 47
rect 1283 21 1313 47
rect 1432 21 1462 47
rect 1523 21 1553 47
rect 1731 21 1761 47
<< polycont >>
rect 32 215 66 249
rect 134 230 168 264
rect 522 331 556 365
rect 341 276 375 310
rect 771 305 805 339
rect 500 169 534 203
rect 602 163 636 197
rect 857 169 891 203
rect 953 217 987 251
rect 1236 331 1270 365
rect 1101 157 1135 191
rect 1197 205 1231 239
rect 1514 315 1548 349
rect 1341 179 1375 213
rect 1437 207 1471 241
rect 1712 215 1746 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 18 477 69 493
rect 18 443 35 477
rect 18 409 69 443
rect 103 461 169 527
rect 103 427 119 461
rect 153 427 169 461
rect 203 477 237 493
rect 18 375 35 409
rect 203 409 237 443
rect 69 391 168 393
rect 69 375 131 391
rect 18 359 131 375
rect 122 357 131 359
rect 165 357 168 391
rect 18 249 88 325
rect 18 215 32 249
rect 66 215 88 249
rect 18 195 88 215
rect 122 264 168 357
rect 122 230 134 264
rect 122 161 168 230
rect 18 127 168 161
rect 203 255 237 375
rect 271 333 336 490
rect 370 485 420 527
rect 370 451 386 485
rect 370 435 420 451
rect 454 477 504 493
rect 454 443 470 477
rect 454 427 504 443
rect 547 483 683 493
rect 547 449 563 483
rect 597 449 683 483
rect 798 475 864 527
rect 991 485 1065 527
rect 547 427 683 449
rect 454 401 488 427
rect 409 367 488 401
rect 522 391 615 393
rect 18 119 69 127
rect 18 85 35 119
rect 203 119 237 221
rect 283 310 375 333
rect 283 276 341 310
rect 283 123 375 276
rect 18 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 409 95 443 367
rect 522 365 581 391
rect 556 357 581 365
rect 556 331 615 357
rect 522 315 615 331
rect 477 255 547 277
rect 477 221 489 255
rect 523 221 547 255
rect 477 203 547 221
rect 477 169 500 203
rect 534 169 547 203
rect 477 153 547 169
rect 581 197 615 315
rect 649 271 683 427
rect 717 459 751 475
rect 798 441 814 475
rect 848 441 864 475
rect 898 459 932 475
rect 717 407 751 425
rect 991 451 1011 485
rect 1045 451 1065 485
rect 991 435 1065 451
rect 1099 477 1133 493
rect 898 407 932 425
rect 717 373 932 407
rect 1099 401 1133 443
rect 1180 484 1354 493
rect 1180 450 1196 484
rect 1230 450 1354 484
rect 1180 425 1354 450
rect 1388 485 1438 527
rect 1422 451 1438 485
rect 1542 485 1608 527
rect 1388 435 1438 451
rect 1472 459 1506 475
rect 1021 367 1133 401
rect 1021 339 1055 367
rect 755 305 771 339
rect 805 305 1055 339
rect 1194 357 1205 391
rect 1239 365 1286 391
rect 1194 333 1236 357
rect 649 251 987 271
rect 649 237 953 251
rect 581 163 602 197
rect 636 163 652 197
rect 581 153 652 163
rect 686 95 720 237
rect 761 187 857 203
rect 795 153 833 187
rect 891 169 919 203
rect 953 201 987 217
rect 867 153 919 169
rect 1021 167 1055 305
rect 203 69 237 85
rect 103 17 169 59
rect 309 55 325 89
rect 359 55 375 89
rect 409 61 458 95
rect 492 61 508 95
rect 549 61 565 95
rect 599 61 720 95
rect 895 93 961 109
rect 309 17 375 55
rect 895 59 911 93
rect 945 59 961 93
rect 895 17 961 59
rect 1003 89 1055 167
rect 1093 331 1236 333
rect 1270 331 1286 365
rect 1320 349 1354 425
rect 1542 451 1558 485
rect 1592 451 1608 485
rect 1676 485 1737 527
rect 1676 451 1687 485
rect 1721 451 1737 485
rect 1472 417 1506 425
rect 1676 417 1737 451
rect 1472 383 1632 417
rect 1093 299 1228 331
rect 1320 315 1514 349
rect 1548 315 1564 349
rect 1093 191 1135 299
rect 1320 297 1354 315
rect 1093 157 1101 191
rect 1093 141 1135 157
rect 1169 255 1239 265
rect 1169 239 1205 255
rect 1169 205 1197 239
rect 1231 205 1239 221
rect 1169 141 1239 205
rect 1273 263 1354 297
rect 1273 107 1307 263
rect 1421 250 1529 281
rect 1598 265 1632 383
rect 1676 383 1687 417
rect 1721 383 1737 417
rect 1676 299 1737 383
rect 1771 449 1822 465
rect 1805 415 1822 449
rect 1771 381 1822 415
rect 1805 347 1822 381
rect 1771 289 1822 347
rect 1598 259 1746 265
rect 1455 241 1529 250
rect 1341 213 1385 229
rect 1375 179 1385 213
rect 1421 207 1437 216
rect 1471 207 1529 241
rect 1341 173 1385 179
rect 1481 187 1529 207
rect 1341 139 1447 173
rect 1117 93 1307 107
rect 1003 55 1023 89
rect 1057 55 1073 89
rect 1117 59 1133 93
rect 1167 59 1307 93
rect 1117 51 1307 59
rect 1341 89 1379 105
rect 1341 55 1345 89
rect 1413 93 1447 139
rect 1515 153 1529 187
rect 1481 127 1529 153
rect 1563 249 1746 259
rect 1563 215 1712 249
rect 1563 199 1746 215
rect 1563 164 1628 199
rect 1563 109 1627 164
rect 1780 159 1822 289
rect 1771 143 1822 159
rect 1805 109 1822 143
rect 1413 75 1563 93
rect 1597 75 1627 109
rect 1413 59 1627 75
rect 1676 93 1737 109
rect 1676 59 1687 93
rect 1721 59 1737 93
rect 1341 17 1379 55
rect 1676 17 1737 59
rect 1771 53 1822 109
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 131 357 165 391
rect 203 221 237 255
rect 581 357 615 391
rect 489 221 523 255
rect 1205 365 1239 391
rect 1205 357 1236 365
rect 1236 357 1239 365
rect 761 153 795 187
rect 833 169 857 187
rect 857 169 867 187
rect 833 153 867 169
rect 1205 239 1239 255
rect 1205 221 1231 239
rect 1231 221 1239 239
rect 1421 241 1455 250
rect 1421 216 1437 241
rect 1437 216 1455 241
rect 1481 153 1515 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
<< metal1 >>
rect 0 561 1840 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 0 496 1840 527
rect 119 391 177 397
rect 119 357 131 391
rect 165 388 177 391
rect 569 391 627 397
rect 569 388 581 391
rect 165 360 581 388
rect 165 357 177 360
rect 119 351 177 357
rect 569 357 581 360
rect 615 388 627 391
rect 1193 391 1251 397
rect 1193 388 1205 391
rect 615 360 1205 388
rect 615 357 627 360
rect 569 351 627 357
rect 1193 357 1205 360
rect 1239 357 1251 391
rect 1193 351 1251 357
rect 191 255 249 261
rect 191 221 203 255
rect 237 252 249 255
rect 477 255 535 261
rect 477 252 489 255
rect 237 224 489 252
rect 237 221 249 224
rect 191 215 249 221
rect 477 221 489 224
rect 523 252 535 255
rect 1193 255 1251 261
rect 1193 252 1205 255
rect 523 224 1205 252
rect 523 221 535 224
rect 477 215 535 221
rect 1193 221 1205 224
rect 1239 221 1251 255
rect 1193 215 1251 221
rect 1409 250 1467 256
rect 1409 216 1421 250
rect 1455 216 1467 250
rect 1409 193 1467 216
rect 749 187 879 193
rect 749 153 761 187
rect 795 153 833 187
rect 867 184 879 187
rect 1409 187 1527 193
rect 1409 184 1481 187
rect 867 156 1481 184
rect 867 153 879 156
rect 749 147 879 153
rect 1469 153 1481 156
rect 1515 153 1527 187
rect 1469 147 1527 153
rect 0 17 1840 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
rect 0 -48 1840 -17
<< labels >>
flabel corelocali s 30 220 66 252 0 FreeSans 200 0 0 0 CLK_N
port 1 nsew
flabel corelocali s 1776 425 1810 459 0 FreeSans 400 0 0 0 Q
port 8 nsew
flabel corelocali s 1776 357 1810 391 0 FreeSans 400 0 0 0 Q
port 8 nsew
flabel corelocali s 1776 289 1810 323 0 FreeSans 400 0 0 0 Q
port 8 nsew
flabel corelocali s 1776 85 1810 119 0 FreeSans 400 0 0 0 Q
port 8 nsew
flabel corelocali s 1481 153 1515 187 0 FreeSans 400 0 0 0 RESET_B
port 3 nsew
flabel corelocali s 305 289 339 323 0 FreeSans 400 0 0 0 D
port 2 nsew
flabel corelocali s 1481 221 1515 255 0 FreeSans 400 0 0 0 RESET_B
port 3 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
rlabel comment s 0 0 0 0 4 dfrtn_1
<< properties >>
string FIXED_BBOX 0 0 1840 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3369420
string GDS_START 3354318
string path 0.000 13.600 46.000 13.600 
<< end >>
