magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 346 383 431 493
rect 20 265 91 337
rect 20 215 133 265
rect 177 215 247 265
rect 372 109 431 383
rect 305 51 431 109
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 25 393 81 527
rect 125 349 185 459
rect 219 383 285 527
rect 125 315 315 349
rect 281 265 315 315
rect 281 199 332 265
rect 281 181 315 199
rect 25 143 315 181
rect 25 71 91 143
rect 221 17 271 109
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
rlabel locali s 20 265 91 337 6 A
port 1 nsew signal input
rlabel locali s 20 215 133 265 6 A
port 1 nsew signal input
rlabel locali s 177 215 247 265 6 B
port 2 nsew signal input
rlabel locali s 372 109 431 383 6 X
port 3 nsew signal output
rlabel locali s 346 383 431 493 6 X
port 3 nsew signal output
rlabel locali s 305 51 431 109 6 X
port 3 nsew signal output
rlabel metal1 s 0 -48 460 48 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 496 460 592 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 460 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1483452
string GDS_START 1478610
<< end >>
