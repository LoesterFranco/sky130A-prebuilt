magic
tech sky130A
magscale 1 2
timestamp 1599588238
<< locali >>
rect 210 300 455 360
rect 489 300 555 360
rect 25 88 168 134
rect 102 51 168 88
rect 319 98 359 134
rect 287 51 359 98
rect 401 98 449 134
rect 401 51 467 98
rect 772 74 839 596
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 72 428 138 596
rect 178 462 220 649
rect 260 428 326 596
rect 72 394 326 428
rect 506 428 572 596
rect 506 394 623 428
rect 72 388 138 394
rect 589 330 623 394
rect 682 364 732 649
rect 77 266 143 268
rect 589 266 738 330
rect 77 264 738 266
rect 77 232 623 264
rect 77 168 143 232
rect 219 132 285 198
rect 343 168 409 232
rect 219 17 253 132
rect 483 132 535 198
rect 569 132 623 232
rect 501 17 535 132
rect 687 17 737 230
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel locali s 102 51 168 88 6 A1
port 1 nsew signal input
rlabel locali s 25 88 168 134 6 A1
port 1 nsew signal input
rlabel locali s 210 300 455 360 6 A2
port 2 nsew signal input
rlabel locali s 319 98 359 134 6 B1
port 3 nsew signal input
rlabel locali s 287 51 359 98 6 B1
port 3 nsew signal input
rlabel locali s 401 98 449 134 6 C1
port 4 nsew signal input
rlabel locali s 401 51 467 98 6 C1
port 4 nsew signal input
rlabel locali s 489 300 555 360 6 D1
port 5 nsew signal input
rlabel locali s 772 74 839 596 6 X
port 6 nsew signal output
rlabel metal1 s 0 -49 864 49 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 617 864 715 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3884850
string GDS_START 3875986
<< end >>
