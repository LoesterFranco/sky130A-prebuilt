magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 89 53 119 137
rect 195 53 225 137
rect 289 53 319 137
rect 383 53 413 137
rect 481 47 511 177
rect 618 47 648 177
<< pmoshvt >>
rect 81 297 117 381
rect 187 297 223 381
rect 269 297 305 381
rect 375 297 411 381
rect 483 297 519 497
rect 610 297 646 497
<< ndiff >>
rect 428 137 481 177
rect 27 117 89 137
rect 27 83 35 117
rect 69 83 89 117
rect 27 53 89 83
rect 119 111 195 137
rect 119 77 135 111
rect 169 77 195 111
rect 119 53 195 77
rect 225 97 289 137
rect 225 63 235 97
rect 269 63 289 97
rect 225 53 289 63
rect 319 111 383 137
rect 319 77 329 111
rect 363 77 383 111
rect 319 53 383 77
rect 413 97 481 137
rect 413 63 433 97
rect 467 63 481 97
rect 413 53 481 63
rect 428 47 481 53
rect 511 135 618 177
rect 511 101 564 135
rect 598 101 618 135
rect 511 47 618 101
rect 648 165 709 177
rect 648 131 663 165
rect 697 131 709 165
rect 648 97 709 131
rect 648 63 663 97
rect 697 63 709 97
rect 648 47 709 63
<< pdiff >>
rect 428 485 483 497
rect 428 451 436 485
rect 470 451 483 485
rect 428 417 483 451
rect 428 383 436 417
rect 470 383 483 417
rect 428 381 483 383
rect 27 354 81 381
rect 27 320 35 354
rect 69 320 81 354
rect 27 297 81 320
rect 117 297 187 381
rect 223 297 269 381
rect 305 297 375 381
rect 411 297 483 381
rect 519 454 610 497
rect 519 420 564 454
rect 598 420 610 454
rect 519 386 610 420
rect 519 352 564 386
rect 598 352 610 386
rect 519 297 610 352
rect 646 485 709 497
rect 646 451 663 485
rect 697 451 709 485
rect 646 417 709 451
rect 646 383 663 417
rect 697 383 709 417
rect 646 349 709 383
rect 646 315 663 349
rect 697 315 709 349
rect 646 297 709 315
<< ndiffc >>
rect 35 83 69 117
rect 135 77 169 111
rect 235 63 269 97
rect 329 77 363 111
rect 433 63 467 97
rect 564 101 598 135
rect 663 131 697 165
rect 663 63 697 97
<< pdiffc >>
rect 436 451 470 485
rect 436 383 470 417
rect 35 320 69 354
rect 564 420 598 454
rect 564 352 598 386
rect 663 451 697 485
rect 663 383 697 417
rect 663 315 697 349
<< poly >>
rect 483 497 519 523
rect 610 497 646 523
rect 267 473 337 483
rect 267 439 287 473
rect 321 439 337 473
rect 267 429 337 439
rect 267 407 307 429
rect 81 381 117 407
rect 187 381 223 407
rect 269 381 305 407
rect 375 381 411 407
rect 81 282 117 297
rect 187 282 223 297
rect 269 282 305 297
rect 375 282 411 297
rect 483 282 519 297
rect 610 282 646 297
rect 79 265 119 282
rect 185 265 225 282
rect 25 249 119 265
rect 25 215 35 249
rect 69 215 119 249
rect 25 199 119 215
rect 161 249 225 265
rect 161 215 171 249
rect 205 215 225 249
rect 161 199 225 215
rect 89 137 119 199
rect 195 137 225 199
rect 267 182 307 282
rect 373 265 413 282
rect 481 265 521 282
rect 608 265 648 282
rect 358 249 422 265
rect 358 215 368 249
rect 402 215 422 249
rect 358 199 422 215
rect 481 249 648 265
rect 481 215 506 249
rect 540 215 648 249
rect 481 199 648 215
rect 267 152 319 182
rect 289 137 319 152
rect 383 137 413 199
rect 481 177 511 199
rect 618 177 648 199
rect 89 27 119 53
rect 195 27 225 53
rect 289 27 319 53
rect 383 27 413 53
rect 481 21 511 47
rect 618 21 648 47
<< polycont >>
rect 287 439 321 473
rect 35 215 69 249
rect 171 215 205 249
rect 368 215 402 249
rect 506 215 540 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 423 485 479 527
rect 17 473 379 483
rect 17 439 287 473
rect 321 439 379 473
rect 17 425 379 439
rect 423 451 436 485
rect 470 451 479 485
rect 423 417 479 451
rect 17 357 366 391
rect 423 383 436 417
rect 470 383 479 417
rect 423 367 479 383
rect 564 454 625 493
rect 598 420 625 454
rect 564 386 625 420
rect 17 354 82 357
rect 17 320 35 354
rect 69 320 82 354
rect 332 333 366 357
rect 598 352 625 386
rect 17 299 82 320
rect 17 249 87 265
rect 17 215 35 249
rect 69 215 87 249
rect 17 151 87 215
rect 121 249 261 323
rect 332 299 487 333
rect 564 299 625 352
rect 453 265 487 299
rect 121 215 171 249
rect 205 215 261 249
rect 121 199 261 215
rect 295 249 419 265
rect 295 215 368 249
rect 402 215 419 249
rect 295 199 419 215
rect 453 249 540 265
rect 453 215 506 249
rect 453 199 540 215
rect 453 165 487 199
rect 135 131 487 165
rect 578 152 625 299
rect 663 485 707 527
rect 697 451 707 485
rect 663 417 707 451
rect 697 383 707 417
rect 663 349 707 383
rect 697 315 707 349
rect 663 291 707 315
rect 564 135 625 152
rect 18 83 35 117
rect 69 83 85 117
rect 18 17 85 83
rect 135 111 169 131
rect 329 111 363 131
rect 135 61 169 77
rect 209 63 235 97
rect 269 63 285 97
rect 209 17 285 63
rect 598 101 625 135
rect 329 61 363 77
rect 397 63 433 97
rect 467 63 483 97
rect 564 83 625 101
rect 663 165 707 200
rect 697 131 707 165
rect 663 97 707 131
rect 397 17 483 63
rect 697 63 707 97
rect 663 17 707 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel corelocali s 303 425 337 459 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel corelocali s 215 221 249 255 0 FreeSans 400 0 0 0 C
port 3 nsew
flabel corelocali s 323 238 323 238 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 573 357 607 391 0 FreeSans 200 0 0 0 X
port 9 nsew
flabel corelocali s 125 221 159 255 0 FreeSans 400 0 0 0 C
port 3 nsew
flabel corelocali s 217 425 251 459 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel corelocali s 126 425 160 459 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel corelocali s 132 289 166 323 0 FreeSans 400 0 0 0 C
port 3 nsew
flabel corelocali s 30 425 64 459 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel corelocali s 221 289 255 323 0 FreeSans 400 0 0 0 C
port 3 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 400 0 0 0 D
port 4 nsew
flabel corelocali s 30 153 64 187 0 FreeSans 400 0 0 0 D
port 4 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
rlabel comment s 0 0 0 0 4 or4_2
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 505304
string GDS_START 498292
<< end >>
