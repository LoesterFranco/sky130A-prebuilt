magic
tech sky130A
magscale 1 2
timestamp 1601050058
<< locali >>
rect 17 215 96 257
rect 637 306 725 493
rect 669 128 725 306
rect 637 54 725 128
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 17 326 86 493
rect 120 360 186 527
rect 278 357 359 493
rect 17 291 254 326
rect 170 249 254 291
rect 325 249 359 357
rect 397 326 447 493
rect 537 360 603 527
rect 397 292 529 326
rect 759 360 811 527
rect 495 265 529 292
rect 153 215 287 249
rect 325 215 461 249
rect 170 181 254 215
rect 17 147 254 181
rect 325 180 359 215
rect 495 199 635 265
rect 495 181 529 199
rect 17 54 83 147
rect 117 17 183 113
rect 288 54 359 180
rect 397 147 529 181
rect 397 54 447 147
rect 537 17 603 113
rect 759 17 811 127
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
rlabel locali s 17 215 96 257 6 A
port 1 nsew signal input
rlabel locali s 669 128 725 306 6 X
port 2 nsew signal output
rlabel locali s 637 306 725 493 6 X
port 2 nsew signal output
rlabel locali s 637 54 725 128 6 X
port 2 nsew signal output
rlabel metal1 s 0 -48 828 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 828 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3198308
string GDS_START 3191708
<< end >>
