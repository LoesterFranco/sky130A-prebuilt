magic
tech sky130A
magscale 1 2
timestamp 1604502705
<< nwell >>
rect -38 335 2342 704
rect -38 332 278 335
rect 662 332 2342 335
rect 662 311 1386 332
<< pwell >>
rect 0 0 2304 49
<< scnmos >>
rect 87 78 117 162
rect 165 78 195 162
rect 382 119 412 267
rect 492 119 522 267
rect 693 138 723 222
rect 793 138 823 222
rect 871 138 901 222
rect 943 138 973 222
rect 1146 74 1176 222
rect 1241 74 1271 222
rect 1451 81 1481 165
rect 1529 81 1559 165
rect 1633 81 1663 165
rect 1711 81 1741 165
rect 1907 74 1937 222
rect 2105 74 2135 222
rect 2191 74 2221 222
<< pmoshvt >>
rect 84 508 114 592
rect 174 508 204 592
rect 366 390 396 590
rect 465 390 495 590
rect 667 463 697 547
rect 768 463 798 547
rect 840 463 870 547
rect 964 463 994 547
rect 1166 347 1196 547
rect 1267 362 1297 562
rect 1448 493 1478 577
rect 1532 493 1562 577
rect 1632 493 1662 577
rect 1774 493 1804 577
rect 1891 409 1921 577
rect 2098 368 2128 592
rect 2188 368 2218 592
<< ndiff >>
rect 323 210 382 267
rect 323 180 337 210
rect 313 176 337 180
rect 371 176 382 210
rect 30 137 87 162
rect 30 103 42 137
rect 76 103 87 137
rect 30 78 87 103
rect 117 78 165 162
rect 195 137 259 162
rect 195 103 213 137
rect 247 103 259 137
rect 195 78 259 103
rect 313 142 382 176
rect 313 108 325 142
rect 359 119 382 142
rect 412 160 492 267
rect 412 126 435 160
rect 469 126 492 160
rect 412 119 492 126
rect 522 225 572 267
rect 522 161 581 225
rect 522 127 535 161
rect 569 127 581 161
rect 636 193 693 222
rect 636 159 648 193
rect 682 159 693 193
rect 636 138 693 159
rect 723 189 793 222
rect 723 155 748 189
rect 782 155 793 189
rect 723 138 793 155
rect 823 138 871 222
rect 901 138 943 222
rect 973 138 1146 222
rect 522 119 581 127
rect 359 108 367 119
rect 313 96 367 108
rect 427 96 477 119
rect 988 74 1146 138
rect 1176 189 1241 222
rect 1176 155 1187 189
rect 1221 155 1241 189
rect 1176 74 1241 155
rect 1271 165 1321 222
rect 1851 194 1907 222
rect 1271 153 1451 165
rect 1271 119 1287 153
rect 1321 119 1373 153
rect 1407 119 1451 153
rect 1271 81 1451 119
rect 1481 81 1529 165
rect 1559 127 1633 165
rect 1559 93 1579 127
rect 1613 93 1633 127
rect 1559 81 1633 93
rect 1663 81 1711 165
rect 1741 140 1797 165
rect 1741 106 1752 140
rect 1786 106 1797 140
rect 1741 81 1797 106
rect 1851 160 1862 194
rect 1896 160 1907 194
rect 1851 120 1907 160
rect 1851 86 1862 120
rect 1896 86 1907 120
rect 1271 74 1321 81
rect 988 73 1065 74
rect 988 39 1009 73
rect 1043 39 1065 73
rect 1851 74 1907 86
rect 1937 209 1994 222
rect 1937 175 1948 209
rect 1982 175 1994 209
rect 1937 120 1994 175
rect 1937 86 1948 120
rect 1982 86 1994 120
rect 1937 74 1994 86
rect 2048 210 2105 222
rect 2048 176 2060 210
rect 2094 176 2105 210
rect 2048 120 2105 176
rect 2048 86 2060 120
rect 2094 86 2105 120
rect 2048 74 2105 86
rect 2135 210 2191 222
rect 2135 176 2146 210
rect 2180 176 2191 210
rect 2135 120 2191 176
rect 2135 86 2146 120
rect 2180 86 2191 120
rect 2135 74 2191 86
rect 2221 210 2277 222
rect 2221 176 2232 210
rect 2266 176 2277 210
rect 2221 120 2277 176
rect 2221 86 2232 120
rect 2266 86 2277 120
rect 2221 74 2277 86
rect 988 27 1065 39
<< pdiff >>
rect 27 567 84 592
rect 27 533 37 567
rect 71 533 84 567
rect 27 508 84 533
rect 114 567 174 592
rect 114 533 127 567
rect 161 533 174 567
rect 114 508 174 533
rect 204 580 261 592
rect 204 546 219 580
rect 253 546 261 580
rect 204 508 261 546
rect 315 482 366 590
rect 309 432 366 482
rect 309 398 321 432
rect 355 398 366 432
rect 309 390 366 398
rect 396 582 465 590
rect 396 548 407 582
rect 441 548 465 582
rect 396 390 465 548
rect 495 439 548 590
rect 495 405 506 439
rect 540 405 548 439
rect 495 390 548 405
rect 888 585 946 597
rect 888 551 900 585
rect 934 551 946 585
rect 2034 580 2098 592
rect 888 547 946 551
rect 1395 562 1448 577
rect 1214 547 1267 562
rect 614 516 667 547
rect 614 482 622 516
rect 656 482 667 516
rect 614 463 667 482
rect 697 539 768 547
rect 697 505 715 539
rect 749 505 768 539
rect 697 463 768 505
rect 798 463 840 547
rect 870 463 964 547
rect 994 512 1053 547
rect 994 478 1007 512
rect 1041 478 1053 512
rect 994 463 1053 478
rect 1107 535 1166 547
rect 1107 501 1119 535
rect 1153 501 1166 535
rect 1107 467 1166 501
rect 1107 433 1119 467
rect 1153 433 1166 467
rect 1107 399 1166 433
rect 1107 365 1119 399
rect 1153 365 1166 399
rect 1107 347 1166 365
rect 1196 535 1267 547
rect 1196 501 1219 535
rect 1253 501 1267 535
rect 1196 421 1267 501
rect 1196 387 1219 421
rect 1253 387 1267 421
rect 1196 362 1267 387
rect 1297 545 1448 562
rect 1297 511 1319 545
rect 1353 511 1401 545
rect 1435 511 1448 545
rect 1297 493 1448 511
rect 1478 493 1532 577
rect 1562 552 1632 577
rect 1562 518 1575 552
rect 1609 518 1632 552
rect 1562 493 1632 518
rect 1662 539 1774 577
rect 1662 505 1701 539
rect 1735 505 1774 539
rect 1662 493 1774 505
rect 1804 552 1891 577
rect 1804 518 1834 552
rect 1868 518 1891 552
rect 1804 493 1891 518
rect 1297 362 1350 493
rect 1196 347 1249 362
rect 1822 409 1891 493
rect 1921 565 1980 577
rect 1921 531 1934 565
rect 1968 531 1980 565
rect 1921 456 1980 531
rect 1921 422 1934 456
rect 1968 422 1980 456
rect 1921 409 1980 422
rect 2034 546 2046 580
rect 2080 546 2098 580
rect 2034 497 2098 546
rect 2034 463 2046 497
rect 2080 463 2098 497
rect 2034 414 2098 463
rect 2034 380 2046 414
rect 2080 380 2098 414
rect 2034 368 2098 380
rect 2128 580 2188 592
rect 2128 546 2141 580
rect 2175 546 2188 580
rect 2128 497 2188 546
rect 2128 463 2141 497
rect 2175 463 2188 497
rect 2128 414 2188 463
rect 2128 380 2141 414
rect 2175 380 2188 414
rect 2128 368 2188 380
rect 2218 580 2277 592
rect 2218 546 2231 580
rect 2265 546 2277 580
rect 2218 497 2277 546
rect 2218 463 2231 497
rect 2265 463 2277 497
rect 2218 414 2277 463
rect 2218 380 2231 414
rect 2265 380 2277 414
rect 2218 368 2277 380
<< ndiffc >>
rect 337 176 371 210
rect 42 103 76 137
rect 213 103 247 137
rect 325 108 359 142
rect 435 126 469 160
rect 535 127 569 161
rect 648 159 682 193
rect 748 155 782 189
rect 1187 155 1221 189
rect 1287 119 1321 153
rect 1373 119 1407 153
rect 1579 93 1613 127
rect 1752 106 1786 140
rect 1862 160 1896 194
rect 1862 86 1896 120
rect 1009 39 1043 73
rect 1948 175 1982 209
rect 1948 86 1982 120
rect 2060 176 2094 210
rect 2060 86 2094 120
rect 2146 176 2180 210
rect 2146 86 2180 120
rect 2232 176 2266 210
rect 2232 86 2266 120
<< pdiffc >>
rect 37 533 71 567
rect 127 533 161 567
rect 219 546 253 580
rect 321 398 355 432
rect 407 548 441 582
rect 506 405 540 439
rect 900 551 934 585
rect 622 482 656 516
rect 715 505 749 539
rect 1007 478 1041 512
rect 1119 501 1153 535
rect 1119 433 1153 467
rect 1119 365 1153 399
rect 1219 501 1253 535
rect 1219 387 1253 421
rect 1319 511 1353 545
rect 1401 511 1435 545
rect 1575 518 1609 552
rect 1701 505 1735 539
rect 1834 518 1868 552
rect 1934 531 1968 565
rect 1934 422 1968 456
rect 2046 546 2080 580
rect 2046 463 2080 497
rect 2046 380 2080 414
rect 2141 546 2175 580
rect 2141 463 2175 497
rect 2141 380 2175 414
rect 2231 546 2265 580
rect 2231 463 2265 497
rect 2231 380 2265 414
<< poly >>
rect 84 592 114 618
rect 174 592 204 618
rect 366 590 396 616
rect 465 590 495 616
rect 563 615 1300 645
rect 84 493 114 508
rect 174 493 204 508
rect 81 402 117 493
rect 171 430 214 493
rect 44 386 117 402
rect 44 352 60 386
rect 94 352 117 386
rect 44 318 117 352
rect 44 284 60 318
rect 94 284 117 318
rect 44 250 117 284
rect 44 216 60 250
rect 94 216 117 250
rect 44 200 117 216
rect 87 162 117 200
rect 165 414 271 430
rect 165 380 207 414
rect 241 380 271 414
rect 165 346 271 380
rect 366 355 396 390
rect 465 375 495 390
rect 563 375 593 615
rect 667 547 697 573
rect 768 547 798 615
rect 840 547 870 573
rect 1264 577 1300 615
rect 1448 577 1478 603
rect 1532 577 1562 603
rect 1632 577 1662 603
rect 1774 577 1804 603
rect 1891 577 1921 603
rect 2098 592 2128 618
rect 2188 592 2218 618
rect 964 547 994 573
rect 1166 547 1196 573
rect 1267 562 1297 577
rect 667 398 697 463
rect 768 437 798 463
rect 840 442 870 463
rect 964 442 994 463
rect 840 425 873 442
rect 961 425 997 442
rect 839 409 911 425
rect 667 397 701 398
rect 465 364 593 375
rect 165 312 207 346
rect 241 312 271 346
rect 165 278 271 312
rect 356 351 421 355
rect 356 339 425 351
rect 356 305 375 339
rect 409 305 425 339
rect 356 287 425 305
rect 467 339 593 364
rect 467 305 503 339
rect 537 312 593 339
rect 635 381 701 397
rect 635 347 651 381
rect 685 361 701 381
rect 839 375 855 409
rect 889 375 911 409
rect 685 347 795 361
rect 839 359 911 375
rect 961 409 1057 425
rect 961 375 1007 409
rect 1041 375 1057 409
rect 961 359 1057 375
rect 635 337 795 347
rect 637 335 795 337
rect 639 333 795 335
rect 641 331 795 333
rect 537 307 598 312
rect 765 311 795 331
rect 537 305 601 307
rect 467 304 601 305
rect 467 301 604 304
rect 467 298 607 301
rect 467 296 609 298
rect 467 293 612 296
rect 467 290 615 293
rect 165 244 207 278
rect 241 244 271 278
rect 382 267 412 287
rect 467 282 617 290
rect 492 267 522 282
rect 580 280 617 282
rect 765 281 823 311
rect 581 279 617 280
rect 583 278 617 279
rect 584 276 617 278
rect 585 275 617 276
rect 587 270 617 275
rect 165 228 271 244
rect 165 162 195 228
rect 587 240 723 270
rect 693 222 723 240
rect 793 222 823 281
rect 871 222 901 359
rect 961 267 991 359
rect 1448 478 1478 493
rect 1532 478 1562 493
rect 1632 478 1662 493
rect 1774 478 1804 493
rect 1445 461 1481 478
rect 1391 445 1481 461
rect 1391 411 1407 445
rect 1441 411 1481 445
rect 1391 395 1481 411
rect 1529 395 1565 478
rect 1629 455 1665 478
rect 1613 439 1679 455
rect 1613 405 1629 439
rect 1663 405 1679 439
rect 1267 347 1297 362
rect 1166 332 1196 347
rect 1163 315 1199 332
rect 1264 317 1481 347
rect 943 237 991 267
rect 1071 299 1199 315
rect 1071 265 1087 299
rect 1121 285 1199 299
rect 1121 265 1176 285
rect 1071 249 1176 265
rect 943 222 973 237
rect 1146 222 1176 249
rect 1241 253 1409 269
rect 1241 239 1359 253
rect 1241 222 1271 239
rect 382 93 412 119
rect 492 93 522 119
rect 693 112 723 138
rect 793 112 823 138
rect 871 112 901 138
rect 87 52 117 78
rect 165 51 195 78
rect 943 51 973 138
rect 165 21 973 51
rect 1343 219 1359 239
rect 1393 219 1409 253
rect 1343 203 1409 219
rect 1451 165 1481 317
rect 1529 278 1559 395
rect 1613 389 1679 405
rect 1525 262 1591 278
rect 1525 228 1541 262
rect 1575 228 1591 262
rect 1525 212 1591 228
rect 1529 165 1559 212
rect 1633 165 1663 389
rect 1771 378 1807 478
rect 1891 394 1921 409
rect 1741 362 1807 378
rect 1741 341 1757 362
rect 1711 328 1757 341
rect 1791 341 1807 362
rect 1888 341 1924 394
rect 2098 353 2128 368
rect 2188 353 2218 368
rect 1791 328 1937 341
rect 1711 311 1937 328
rect 1711 165 1741 311
rect 1907 222 1937 311
rect 1985 310 2051 326
rect 1985 276 2001 310
rect 2035 290 2051 310
rect 2095 290 2131 353
rect 2185 290 2221 353
rect 2035 276 2221 290
rect 1985 260 2221 276
rect 2105 222 2135 260
rect 2191 222 2221 260
rect 1146 48 1176 74
rect 1241 48 1271 74
rect 1451 55 1481 81
rect 1529 55 1559 81
rect 1633 55 1663 81
rect 1711 55 1741 81
rect 1907 48 1937 74
rect 2105 48 2135 74
rect 2191 48 2221 74
<< polycont >>
rect 60 352 94 386
rect 60 284 94 318
rect 60 216 94 250
rect 207 380 241 414
rect 207 312 241 346
rect 375 305 409 339
rect 503 305 537 339
rect 651 347 685 381
rect 855 375 889 409
rect 1007 375 1041 409
rect 207 244 241 278
rect 1407 411 1441 445
rect 1629 405 1663 439
rect 1087 265 1121 299
rect 1359 219 1393 253
rect 1541 228 1575 262
rect 1757 328 1791 362
rect 2001 276 2035 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2304 683
rect 21 567 87 649
rect 21 533 37 567
rect 71 533 87 567
rect 21 504 87 533
rect 127 567 167 596
rect 161 533 167 567
rect 203 580 269 649
rect 203 546 219 580
rect 253 546 269 580
rect 391 582 457 649
rect 391 548 407 582
rect 441 548 457 582
rect 884 585 950 649
rect 884 551 900 585
rect 934 551 950 585
rect 127 526 167 533
rect 127 521 174 526
rect 609 523 665 545
rect 481 521 665 523
rect 127 512 178 521
rect 478 519 665 521
rect 475 518 665 519
rect 473 517 665 518
rect 471 516 665 517
rect 469 515 622 516
rect 466 514 622 515
rect 281 512 622 514
rect 127 504 622 512
rect 133 489 622 504
rect 133 488 497 489
rect 133 487 494 488
rect 133 486 492 487
rect 133 484 488 486
rect 133 481 484 484
rect 589 482 622 489
rect 656 482 665 516
rect 699 539 850 550
rect 884 548 950 551
rect 699 505 715 539
rect 749 514 850 539
rect 1103 535 1169 649
rect 749 512 1057 514
rect 749 505 1007 512
rect 133 479 481 481
rect 589 480 665 482
rect 787 480 1007 505
rect 133 476 477 479
rect 133 471 472 476
rect 589 475 674 480
rect 622 471 674 475
rect 133 466 468 471
rect 25 386 99 434
rect 25 352 60 386
rect 94 352 99 386
rect 25 318 99 352
rect 25 284 60 318
rect 94 284 99 318
rect 25 250 99 284
rect 25 216 60 250
rect 94 216 99 250
rect 25 200 99 216
rect 133 166 167 466
rect 506 446 555 455
rect 622 446 753 471
rect 503 441 555 446
rect 503 439 588 441
rect 201 424 257 430
rect 201 414 223 424
rect 201 380 207 414
rect 241 380 257 390
rect 201 346 257 380
rect 201 312 207 346
rect 241 312 257 346
rect 201 278 257 312
rect 201 244 207 278
rect 241 244 257 278
rect 201 228 257 244
rect 291 398 321 432
rect 355 398 373 432
rect 291 380 373 398
rect 503 405 506 439
rect 540 416 588 439
rect 640 437 753 446
rect 540 407 602 416
rect 540 405 619 407
rect 503 397 619 405
rect 503 389 685 397
rect 562 381 685 389
rect 562 380 651 381
rect 291 230 325 380
rect 409 346 455 356
rect 359 339 455 346
rect 359 305 375 339
rect 409 305 455 339
rect 503 339 537 355
rect 359 264 455 305
rect 489 305 503 310
rect 489 230 537 305
rect 291 210 537 230
rect 291 176 337 210
rect 371 195 537 210
rect 573 347 651 380
rect 573 325 685 347
rect 371 194 508 195
rect 371 176 375 194
rect 26 137 167 166
rect 26 103 42 137
rect 76 132 167 137
rect 201 137 257 166
rect 76 103 92 132
rect 26 74 92 103
rect 201 103 213 137
rect 247 103 257 137
rect 201 17 257 103
rect 291 142 375 176
rect 573 161 614 325
rect 719 278 753 437
rect 664 244 753 278
rect 664 209 698 244
rect 787 210 821 480
rect 923 478 1007 480
rect 1041 478 1057 512
rect 923 464 1057 478
rect 1103 501 1119 535
rect 1153 501 1169 535
rect 1103 467 1169 501
rect 291 108 325 142
rect 359 108 375 142
rect 291 70 375 108
rect 419 126 435 160
rect 469 126 485 160
rect 419 17 485 126
rect 519 127 535 161
rect 569 127 614 161
rect 648 193 698 209
rect 682 159 698 193
rect 648 134 698 159
rect 732 189 821 210
rect 855 409 889 425
rect 855 225 889 375
rect 923 315 957 464
rect 1103 433 1119 467
rect 1153 433 1169 467
rect 991 424 1057 430
rect 1025 409 1057 424
rect 991 375 1007 390
rect 1041 375 1057 409
rect 991 359 1057 375
rect 1103 399 1169 433
rect 1103 365 1119 399
rect 1153 365 1169 399
rect 1103 349 1169 365
rect 1203 535 1269 551
rect 1203 501 1219 535
rect 1253 501 1269 535
rect 1203 421 1269 501
rect 1203 387 1219 421
rect 1253 387 1269 421
rect 1203 371 1269 387
rect 1303 545 1525 561
rect 1303 511 1319 545
rect 1353 511 1401 545
rect 1435 511 1525 545
rect 1303 495 1525 511
rect 923 299 1137 315
rect 923 265 1087 299
rect 1121 265 1137 299
rect 923 259 1137 265
rect 1203 226 1237 371
rect 1303 337 1337 495
rect 1171 225 1237 226
rect 855 191 1237 225
rect 732 155 748 189
rect 782 155 821 189
rect 1171 189 1237 191
rect 732 134 821 155
rect 519 100 614 127
rect 861 123 1137 157
rect 861 100 895 123
rect 519 66 895 100
rect 984 73 1069 89
rect 984 39 1009 73
rect 1043 39 1069 73
rect 1103 85 1137 123
rect 1171 155 1187 189
rect 1221 155 1237 189
rect 1171 119 1237 155
rect 1271 303 1337 337
rect 1391 445 1457 461
rect 1391 411 1407 445
rect 1441 411 1457 445
rect 1271 169 1305 303
rect 1391 269 1457 411
rect 1491 346 1525 495
rect 1559 552 1625 649
rect 1559 518 1575 552
rect 1609 518 1625 552
rect 1559 489 1625 518
rect 1659 539 1777 555
rect 1659 505 1701 539
rect 1735 505 1777 539
rect 1659 489 1777 505
rect 1818 552 1884 649
rect 1818 518 1834 552
rect 1868 518 1884 552
rect 1818 489 1884 518
rect 1918 565 1984 581
rect 1918 531 1934 565
rect 1968 531 1984 565
rect 1743 455 1777 489
rect 1918 456 1984 531
rect 1561 439 1679 455
rect 1561 424 1629 439
rect 1561 390 1567 424
rect 1601 405 1629 424
rect 1663 405 1679 439
rect 1743 421 1875 455
rect 1601 390 1679 405
rect 1561 384 1679 390
rect 1741 362 1807 378
rect 1741 346 1757 362
rect 1491 328 1757 346
rect 1791 328 1807 362
rect 1491 312 1807 328
rect 1841 278 1875 421
rect 1918 422 1934 456
rect 1968 422 1984 456
rect 1918 406 1984 422
rect 1345 253 1491 269
rect 1345 219 1359 253
rect 1393 219 1491 253
rect 1345 203 1491 219
rect 1525 262 1875 278
rect 1525 228 1541 262
rect 1575 244 1875 262
rect 1932 326 1984 406
rect 2030 580 2096 649
rect 2030 546 2046 580
rect 2080 546 2096 580
rect 2030 497 2096 546
rect 2030 463 2046 497
rect 2080 463 2096 497
rect 2030 414 2096 463
rect 2030 380 2046 414
rect 2080 380 2096 414
rect 2030 364 2096 380
rect 2130 580 2196 596
rect 2130 546 2141 580
rect 2175 546 2196 580
rect 2130 497 2196 546
rect 2130 463 2141 497
rect 2175 463 2196 497
rect 2130 414 2196 463
rect 2130 380 2141 414
rect 2175 380 2196 414
rect 1932 310 2038 326
rect 1932 276 2001 310
rect 2035 276 2038 310
rect 1932 260 2038 276
rect 1575 228 1591 244
rect 1525 212 1591 228
rect 1271 153 1423 169
rect 1271 119 1287 153
rect 1321 119 1373 153
rect 1407 119 1423 153
rect 1457 85 1491 203
rect 1103 51 1491 85
rect 1554 127 1638 143
rect 1554 93 1579 127
rect 1613 93 1638 127
rect 984 17 1069 39
rect 1554 17 1638 93
rect 1736 140 1802 244
rect 1736 106 1752 140
rect 1786 106 1802 140
rect 1736 77 1802 106
rect 1846 194 1896 210
rect 1846 160 1862 194
rect 1846 120 1896 160
rect 1846 86 1862 120
rect 1846 17 1896 86
rect 1932 209 1998 260
rect 1932 175 1948 209
rect 1982 175 1998 209
rect 1932 120 1998 175
rect 1932 86 1948 120
rect 1982 86 1998 120
rect 1932 70 1998 86
rect 2044 210 2094 226
rect 2044 176 2060 210
rect 2044 120 2094 176
rect 2044 86 2060 120
rect 2044 17 2094 86
rect 2130 210 2196 380
rect 2231 580 2281 649
rect 2265 546 2281 580
rect 2231 497 2281 546
rect 2265 463 2281 497
rect 2231 414 2281 463
rect 2265 380 2281 414
rect 2231 364 2281 380
rect 2130 176 2146 210
rect 2180 176 2196 210
rect 2130 120 2196 176
rect 2130 86 2146 120
rect 2180 86 2196 120
rect 2130 70 2196 86
rect 2232 210 2282 226
rect 2266 176 2282 210
rect 2232 120 2282 176
rect 2266 86 2282 120
rect 2232 17 2282 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2304 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 223 414 257 424
rect 223 390 241 414
rect 241 390 257 414
rect 991 409 1025 424
rect 991 390 1007 409
rect 1007 390 1025 409
rect 1567 390 1601 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
<< metal1 >>
rect 0 683 2304 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2304 683
rect 0 617 2304 649
rect 211 424 269 430
rect 211 390 223 424
rect 257 421 269 424
rect 979 424 1037 430
rect 979 421 991 424
rect 257 393 991 421
rect 257 390 269 393
rect 211 384 269 390
rect 979 390 991 393
rect 1025 421 1037 424
rect 1555 424 1613 430
rect 1555 421 1567 424
rect 1025 393 1567 421
rect 1025 390 1037 393
rect 979 384 1037 390
rect 1555 390 1567 393
rect 1601 390 1613 424
rect 1555 384 1613 390
rect 0 17 2304 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2304 17
rect 0 -49 2304 -17
<< labels >>
flabel comment s 926 630 926 630 0 FreeSans 300 0 0 0 no_jumper_check
flabel comment s 587 36 587 36 0 FreeSans 300 0 0 0 no_jumper_check
rlabel comment s 0 0 0 0 4 dfrtp_2
flabel pwell s 0 0 2304 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 2304 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 223 390 257 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew
flabel metal1 s 0 617 2304 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 2304 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 31 390 65 424 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 2143 94 2177 128 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 2143 168 2177 202 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 2143 242 2177 276 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 2143 316 2177 350 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 2143 390 2177 424 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 2143 464 2177 498 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 2143 538 2177 572 0 FreeSans 340 0 0 0 Q
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 2304 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2623918
string GDS_START 2605032
<< end >>
