magic
tech sky130A
magscale 1 2
timestamp 1604502697
<< nwell >>
rect -38 261 2522 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 466 47 496 131
rect 562 47 592 131
rect 658 47 688 131
rect 754 47 784 131
rect 850 47 880 131
rect 946 47 976 131
rect 1049 47 1079 131
rect 1176 47 1206 131
rect 1272 47 1302 131
rect 1368 47 1398 131
rect 1464 47 1494 131
rect 1560 47 1590 131
rect 1656 47 1686 131
rect 1752 47 1782 131
rect 1848 47 1878 131
rect 1944 47 1974 131
<< pmoshvt >>
rect 84 297 120 497
rect 180 297 216 497
rect 276 297 312 497
rect 372 297 408 497
rect 468 297 504 497
rect 564 297 600 497
rect 660 297 696 497
rect 756 297 792 497
rect 852 297 888 497
rect 948 297 984 497
rect 1051 297 1087 497
rect 1178 297 1214 497
rect 1274 297 1310 497
rect 1370 297 1406 497
rect 1466 297 1502 497
rect 1562 297 1598 497
rect 1658 297 1694 497
rect 1754 297 1790 497
rect 1850 297 1886 497
rect 1946 297 1982 497
rect 2042 297 2078 497
rect 2138 297 2174 497
rect 2234 297 2270 497
rect 2330 297 2366 497
<< ndiff >>
rect 413 106 466 131
rect 413 72 421 106
rect 455 72 466 106
rect 413 47 466 72
rect 496 106 562 131
rect 496 72 517 106
rect 551 72 562 106
rect 496 47 562 72
rect 592 106 658 131
rect 592 72 613 106
rect 647 72 658 106
rect 592 47 658 72
rect 688 106 754 131
rect 688 72 709 106
rect 743 72 754 106
rect 688 47 754 72
rect 784 106 850 131
rect 784 72 805 106
rect 839 72 850 106
rect 784 47 850 72
rect 880 106 946 131
rect 880 72 901 106
rect 935 72 946 106
rect 880 47 946 72
rect 976 106 1049 131
rect 976 72 1002 106
rect 1036 72 1049 106
rect 976 47 1049 72
rect 1079 106 1176 131
rect 1079 72 1106 106
rect 1140 72 1176 106
rect 1079 47 1176 72
rect 1206 106 1272 131
rect 1206 72 1227 106
rect 1261 72 1272 106
rect 1206 47 1272 72
rect 1302 106 1368 131
rect 1302 72 1323 106
rect 1357 72 1368 106
rect 1302 47 1368 72
rect 1398 106 1464 131
rect 1398 72 1419 106
rect 1453 72 1464 106
rect 1398 47 1464 72
rect 1494 106 1560 131
rect 1494 72 1515 106
rect 1549 72 1560 106
rect 1494 47 1560 72
rect 1590 106 1656 131
rect 1590 72 1611 106
rect 1645 72 1656 106
rect 1590 47 1656 72
rect 1686 106 1752 131
rect 1686 72 1707 106
rect 1741 72 1752 106
rect 1686 47 1752 72
rect 1782 106 1848 131
rect 1782 72 1803 106
rect 1837 72 1848 106
rect 1782 47 1848 72
rect 1878 106 1944 131
rect 1878 72 1899 106
rect 1933 72 1944 106
rect 1878 47 1944 72
rect 1974 106 2037 131
rect 1974 72 1995 106
rect 2029 72 2037 106
rect 1974 47 2037 72
<< pdiff >>
rect 27 485 84 497
rect 27 451 38 485
rect 72 451 84 485
rect 27 417 84 451
rect 27 383 38 417
rect 72 383 84 417
rect 27 349 84 383
rect 27 315 38 349
rect 72 315 84 349
rect 27 297 84 315
rect 120 477 180 497
rect 120 443 133 477
rect 167 443 180 477
rect 120 409 180 443
rect 120 375 133 409
rect 167 375 180 409
rect 120 341 180 375
rect 120 307 133 341
rect 167 307 180 341
rect 120 297 180 307
rect 216 485 276 497
rect 216 451 229 485
rect 263 451 276 485
rect 216 417 276 451
rect 216 383 229 417
rect 263 383 276 417
rect 216 297 276 383
rect 312 474 372 497
rect 312 440 325 474
rect 359 440 372 474
rect 312 341 372 440
rect 312 307 325 341
rect 359 307 372 341
rect 312 297 372 307
rect 408 485 468 497
rect 408 451 421 485
rect 455 451 468 485
rect 408 417 468 451
rect 408 383 421 417
rect 455 383 468 417
rect 408 297 468 383
rect 504 474 564 497
rect 504 440 517 474
rect 551 440 564 474
rect 504 341 564 440
rect 504 307 517 341
rect 551 307 564 341
rect 504 297 564 307
rect 600 485 660 497
rect 600 451 613 485
rect 647 451 660 485
rect 600 417 660 451
rect 600 383 613 417
rect 647 383 660 417
rect 600 297 660 383
rect 696 474 756 497
rect 696 440 709 474
rect 743 440 756 474
rect 696 341 756 440
rect 696 307 709 341
rect 743 307 756 341
rect 696 297 756 307
rect 792 485 852 497
rect 792 451 805 485
rect 839 451 852 485
rect 792 417 852 451
rect 792 383 805 417
rect 839 383 852 417
rect 792 297 852 383
rect 888 474 948 497
rect 888 440 901 474
rect 935 440 948 474
rect 888 341 948 440
rect 888 307 901 341
rect 935 307 948 341
rect 888 297 948 307
rect 984 485 1051 497
rect 984 451 1001 485
rect 1035 451 1051 485
rect 984 417 1051 451
rect 984 383 1001 417
rect 1035 383 1051 417
rect 984 297 1051 383
rect 1087 474 1178 497
rect 1087 440 1126 474
rect 1160 440 1178 474
rect 1087 341 1178 440
rect 1087 307 1126 341
rect 1160 307 1178 341
rect 1087 297 1178 307
rect 1214 485 1274 497
rect 1214 451 1226 485
rect 1260 451 1274 485
rect 1214 417 1274 451
rect 1214 383 1226 417
rect 1260 383 1274 417
rect 1214 297 1274 383
rect 1310 474 1370 497
rect 1310 440 1323 474
rect 1357 440 1370 474
rect 1310 341 1370 440
rect 1310 307 1323 341
rect 1357 307 1370 341
rect 1310 297 1370 307
rect 1406 485 1466 497
rect 1406 451 1419 485
rect 1453 451 1466 485
rect 1406 417 1466 451
rect 1406 383 1419 417
rect 1453 383 1466 417
rect 1406 297 1466 383
rect 1502 474 1562 497
rect 1502 440 1515 474
rect 1549 440 1562 474
rect 1502 341 1562 440
rect 1502 307 1515 341
rect 1549 307 1562 341
rect 1502 297 1562 307
rect 1598 485 1658 497
rect 1598 451 1611 485
rect 1645 451 1658 485
rect 1598 417 1658 451
rect 1598 383 1611 417
rect 1645 383 1658 417
rect 1598 297 1658 383
rect 1694 474 1754 497
rect 1694 440 1707 474
rect 1741 440 1754 474
rect 1694 341 1754 440
rect 1694 307 1707 341
rect 1741 307 1754 341
rect 1694 297 1754 307
rect 1790 485 1850 497
rect 1790 451 1803 485
rect 1837 451 1850 485
rect 1790 417 1850 451
rect 1790 383 1803 417
rect 1837 383 1850 417
rect 1790 297 1850 383
rect 1886 474 1946 497
rect 1886 440 1899 474
rect 1933 440 1946 474
rect 1886 341 1946 440
rect 1886 307 1899 341
rect 1933 307 1946 341
rect 1886 297 1946 307
rect 1982 485 2042 497
rect 1982 451 1995 485
rect 2029 451 2042 485
rect 1982 417 2042 451
rect 1982 383 1995 417
rect 2029 383 2042 417
rect 1982 297 2042 383
rect 2078 474 2138 497
rect 2078 440 2091 474
rect 2125 440 2138 474
rect 2078 341 2138 440
rect 2078 307 2091 341
rect 2125 307 2138 341
rect 2078 297 2138 307
rect 2174 485 2234 497
rect 2174 451 2187 485
rect 2221 451 2234 485
rect 2174 417 2234 451
rect 2174 383 2187 417
rect 2221 383 2234 417
rect 2174 297 2234 383
rect 2270 474 2330 497
rect 2270 440 2283 474
rect 2317 440 2330 474
rect 2270 341 2330 440
rect 2270 307 2283 341
rect 2317 307 2330 341
rect 2270 297 2330 307
rect 2366 485 2421 497
rect 2366 451 2378 485
rect 2412 451 2421 485
rect 2366 417 2421 451
rect 2366 383 2378 417
rect 2412 383 2421 417
rect 2366 297 2421 383
<< ndiffc >>
rect 421 72 455 106
rect 517 72 551 106
rect 613 72 647 106
rect 709 72 743 106
rect 805 72 839 106
rect 901 72 935 106
rect 1002 72 1036 106
rect 1106 72 1140 106
rect 1227 72 1261 106
rect 1323 72 1357 106
rect 1419 72 1453 106
rect 1515 72 1549 106
rect 1611 72 1645 106
rect 1707 72 1741 106
rect 1803 72 1837 106
rect 1899 72 1933 106
rect 1995 72 2029 106
<< pdiffc >>
rect 38 451 72 485
rect 38 383 72 417
rect 38 315 72 349
rect 133 443 167 477
rect 133 375 167 409
rect 133 307 167 341
rect 229 451 263 485
rect 229 383 263 417
rect 325 440 359 474
rect 325 307 359 341
rect 421 451 455 485
rect 421 383 455 417
rect 517 440 551 474
rect 517 307 551 341
rect 613 451 647 485
rect 613 383 647 417
rect 709 440 743 474
rect 709 307 743 341
rect 805 451 839 485
rect 805 383 839 417
rect 901 440 935 474
rect 901 307 935 341
rect 1001 451 1035 485
rect 1001 383 1035 417
rect 1126 440 1160 474
rect 1126 307 1160 341
rect 1226 451 1260 485
rect 1226 383 1260 417
rect 1323 440 1357 474
rect 1323 307 1357 341
rect 1419 451 1453 485
rect 1419 383 1453 417
rect 1515 440 1549 474
rect 1515 307 1549 341
rect 1611 451 1645 485
rect 1611 383 1645 417
rect 1707 440 1741 474
rect 1707 307 1741 341
rect 1803 451 1837 485
rect 1803 383 1837 417
rect 1899 440 1933 474
rect 1899 307 1933 341
rect 1995 451 2029 485
rect 1995 383 2029 417
rect 2091 440 2125 474
rect 2091 307 2125 341
rect 2187 451 2221 485
rect 2187 383 2221 417
rect 2283 440 2317 474
rect 2283 307 2317 341
rect 2378 451 2412 485
rect 2378 383 2412 417
<< poly >>
rect 84 497 120 523
rect 180 497 216 523
rect 276 497 312 523
rect 372 497 408 523
rect 468 497 504 523
rect 564 497 600 523
rect 660 497 696 523
rect 756 497 792 523
rect 852 497 888 523
rect 948 497 984 523
rect 1051 497 1087 523
rect 1178 497 1214 523
rect 1274 497 1310 523
rect 1370 497 1406 523
rect 1466 497 1502 523
rect 1562 497 1598 523
rect 1658 497 1694 523
rect 1754 497 1790 523
rect 1850 497 1886 523
rect 1946 497 1982 523
rect 2042 497 2078 523
rect 2138 497 2174 523
rect 2234 497 2270 523
rect 2330 497 2366 523
rect 84 282 120 297
rect 180 282 216 297
rect 276 282 312 297
rect 372 282 408 297
rect 468 282 504 297
rect 564 282 600 297
rect 660 282 696 297
rect 756 282 792 297
rect 852 282 888 297
rect 948 282 984 297
rect 1051 282 1087 297
rect 1178 282 1214 297
rect 1274 282 1310 297
rect 1370 282 1406 297
rect 1466 282 1502 297
rect 1562 282 1598 297
rect 1658 282 1694 297
rect 1754 282 1790 297
rect 1850 282 1886 297
rect 1946 282 1982 297
rect 2042 282 2078 297
rect 2138 282 2174 297
rect 2234 282 2270 297
rect 2330 282 2366 297
rect 82 270 122 282
rect 178 270 218 282
rect 274 270 314 282
rect 370 270 410 282
rect 466 270 506 282
rect 562 270 602 282
rect 658 270 698 282
rect 754 270 794 282
rect 850 270 890 282
rect 946 270 986 282
rect 1049 270 1089 282
rect 1176 270 1216 282
rect 1272 270 1312 282
rect 1368 270 1408 282
rect 1464 270 1504 282
rect 1560 270 1600 282
rect 1656 270 1696 282
rect 1752 270 1792 282
rect 1848 270 1888 282
rect 1944 270 1984 282
rect 2040 270 2080 282
rect 2136 270 2176 282
rect 2232 270 2272 282
rect 2328 270 2368 282
rect 82 249 2368 270
rect 82 215 101 249
rect 135 215 179 249
rect 213 215 257 249
rect 291 215 335 249
rect 369 215 413 249
rect 447 215 2003 249
rect 2037 215 2081 249
rect 2115 215 2149 249
rect 2183 215 2227 249
rect 2261 215 2305 249
rect 2339 215 2368 249
rect 82 198 2368 215
rect 466 131 496 198
rect 562 131 592 198
rect 658 131 688 198
rect 754 131 784 198
rect 850 131 880 198
rect 946 131 976 198
rect 1049 131 1079 198
rect 1176 131 1206 198
rect 1272 131 1302 198
rect 1368 131 1398 198
rect 1464 131 1494 198
rect 1560 131 1590 198
rect 1656 131 1686 198
rect 1752 131 1782 198
rect 1848 131 1878 198
rect 1944 131 1974 198
rect 466 21 496 47
rect 562 21 592 47
rect 658 21 688 47
rect 754 21 784 47
rect 850 21 880 47
rect 946 21 976 47
rect 1049 21 1079 47
rect 1176 21 1206 47
rect 1272 21 1302 47
rect 1368 21 1398 47
rect 1464 21 1494 47
rect 1560 21 1590 47
rect 1656 21 1686 47
rect 1752 21 1782 47
rect 1848 21 1878 47
rect 1944 21 1974 47
<< polycont >>
rect 101 215 135 249
rect 179 215 213 249
rect 257 215 291 249
rect 335 215 369 249
rect 413 215 447 249
rect 2003 215 2037 249
rect 2081 215 2115 249
rect 2149 215 2183 249
rect 2227 215 2261 249
rect 2305 215 2339 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2484 561
rect 28 485 81 527
rect 28 451 38 485
rect 72 451 81 485
rect 28 417 81 451
rect 28 383 38 417
rect 72 383 81 417
rect 28 349 81 383
rect 28 315 38 349
rect 72 315 81 349
rect 28 299 81 315
rect 125 477 176 493
rect 125 443 133 477
rect 167 443 176 477
rect 125 409 176 443
rect 125 375 133 409
rect 167 375 176 409
rect 125 341 176 375
rect 220 485 272 527
rect 220 451 229 485
rect 263 451 272 485
rect 220 417 272 451
rect 220 383 229 417
rect 263 383 272 417
rect 220 367 272 383
rect 317 474 368 490
rect 317 440 325 474
rect 359 440 368 474
rect 125 307 133 341
rect 167 333 176 341
rect 317 341 368 440
rect 413 485 464 527
rect 413 451 421 485
rect 455 451 464 485
rect 413 417 464 451
rect 413 383 421 417
rect 455 383 464 417
rect 413 367 464 383
rect 515 474 560 493
rect 515 440 517 474
rect 551 440 560 474
rect 317 333 325 341
rect 167 307 325 333
rect 359 333 368 341
rect 515 341 560 440
rect 604 485 656 527
rect 604 451 613 485
rect 647 451 656 485
rect 604 417 656 451
rect 604 383 613 417
rect 647 383 656 417
rect 604 367 656 383
rect 701 474 752 490
rect 701 440 709 474
rect 743 440 752 474
rect 515 333 517 341
rect 359 307 517 333
rect 551 333 560 341
rect 701 341 752 440
rect 797 485 848 527
rect 797 451 805 485
rect 839 451 848 485
rect 797 417 848 451
rect 797 383 805 417
rect 839 383 848 417
rect 797 367 848 383
rect 893 474 941 490
rect 893 440 901 474
rect 935 440 941 474
rect 701 333 709 341
rect 551 307 709 333
rect 743 333 752 341
rect 893 341 941 440
rect 993 485 1044 527
rect 993 451 1001 485
rect 1035 451 1044 485
rect 993 417 1044 451
rect 993 383 1001 417
rect 1035 383 1044 417
rect 993 367 1044 383
rect 1091 474 1166 490
rect 1091 440 1126 474
rect 1160 440 1166 474
rect 893 333 901 341
rect 743 307 901 333
rect 935 333 941 341
rect 1091 341 1166 440
rect 1218 485 1270 527
rect 1218 451 1226 485
rect 1260 451 1270 485
rect 1218 424 1270 451
rect 1315 474 1365 490
rect 1315 440 1323 474
rect 1357 440 1365 474
rect 1218 417 1269 424
rect 1218 383 1226 417
rect 1260 383 1269 417
rect 1218 367 1269 383
rect 1091 333 1126 341
rect 935 307 1126 333
rect 1160 333 1166 341
rect 1315 341 1365 440
rect 1411 485 1462 527
rect 1411 451 1419 485
rect 1453 451 1462 485
rect 1411 417 1462 451
rect 1411 383 1419 417
rect 1453 383 1462 417
rect 1411 367 1462 383
rect 1507 474 1557 490
rect 1507 440 1515 474
rect 1549 440 1557 474
rect 1315 333 1323 341
rect 1160 307 1323 333
rect 1357 333 1365 341
rect 1507 341 1557 440
rect 1603 485 1654 527
rect 1603 451 1611 485
rect 1645 451 1654 485
rect 1603 417 1654 451
rect 1603 383 1611 417
rect 1645 383 1654 417
rect 1603 367 1654 383
rect 1699 474 1749 490
rect 1699 440 1707 474
rect 1741 440 1749 474
rect 1507 333 1515 341
rect 1357 307 1515 333
rect 1549 333 1557 341
rect 1699 341 1749 440
rect 1795 485 1846 527
rect 1795 451 1803 485
rect 1837 451 1846 485
rect 1795 417 1846 451
rect 1795 383 1803 417
rect 1837 383 1846 417
rect 1795 367 1846 383
rect 1891 474 1941 490
rect 1891 440 1899 474
rect 1933 440 1941 474
rect 1699 333 1707 341
rect 1549 307 1707 333
rect 1741 333 1749 341
rect 1891 341 1941 440
rect 1987 485 2038 527
rect 1987 451 1995 485
rect 2029 451 2038 485
rect 1987 417 2038 451
rect 1987 383 1995 417
rect 2029 383 2038 417
rect 1987 367 2038 383
rect 2083 474 2131 490
rect 2083 440 2091 474
rect 2125 440 2131 474
rect 1891 333 1899 341
rect 1741 307 1899 333
rect 1933 333 1941 341
rect 2083 341 2131 440
rect 2179 485 2230 527
rect 2179 451 2187 485
rect 2221 451 2230 485
rect 2179 417 2230 451
rect 2179 383 2187 417
rect 2221 383 2230 417
rect 2179 367 2230 383
rect 2275 474 2326 490
rect 2275 440 2283 474
rect 2317 440 2326 474
rect 2083 333 2091 341
rect 1933 307 2091 333
rect 2125 333 2131 341
rect 2275 341 2326 440
rect 2370 485 2422 527
rect 2370 451 2378 485
rect 2412 451 2422 485
rect 2370 417 2422 451
rect 2370 383 2378 417
rect 2412 383 2422 417
rect 2370 367 2422 383
rect 2275 333 2283 341
rect 2125 307 2283 333
rect 2317 307 2326 341
rect 125 291 2326 307
rect 515 283 1941 291
rect 69 249 335 255
rect 369 249 437 255
rect 69 215 101 249
rect 135 215 179 249
rect 213 215 257 249
rect 291 215 335 249
rect 369 215 413 249
rect 447 215 471 221
rect 69 179 471 215
rect 411 106 465 122
rect 411 72 421 106
rect 455 72 465 106
rect 411 17 465 72
rect 515 106 560 283
rect 515 72 517 106
rect 551 72 560 106
rect 515 56 560 72
rect 604 106 657 122
rect 604 72 613 106
rect 647 72 657 106
rect 604 17 657 72
rect 701 106 752 283
rect 701 72 709 106
rect 743 72 752 106
rect 701 56 752 72
rect 796 106 849 122
rect 796 72 805 106
rect 839 72 849 106
rect 796 17 849 72
rect 893 106 941 283
rect 893 72 901 106
rect 935 72 941 106
rect 893 56 941 72
rect 993 106 1046 122
rect 993 72 1002 106
rect 1036 72 1046 106
rect 993 17 1046 72
rect 1091 106 1161 283
rect 1091 72 1106 106
rect 1140 72 1161 106
rect 1091 56 1161 72
rect 1218 106 1271 122
rect 1218 72 1227 106
rect 1261 72 1271 106
rect 1218 17 1271 72
rect 1315 106 1365 283
rect 1315 72 1323 106
rect 1357 72 1365 106
rect 1315 56 1365 72
rect 1410 106 1455 122
rect 1410 72 1419 106
rect 1453 72 1455 106
rect 1410 17 1455 72
rect 1507 106 1557 283
rect 1507 72 1515 106
rect 1549 72 1557 106
rect 1507 56 1557 72
rect 1602 106 1655 122
rect 1602 72 1611 106
rect 1645 72 1655 106
rect 1602 17 1655 72
rect 1699 106 1749 283
rect 1699 72 1707 106
rect 1741 72 1749 106
rect 1699 56 1749 72
rect 1794 106 1847 122
rect 1794 72 1803 106
rect 1837 72 1847 106
rect 1794 17 1847 72
rect 1891 106 1941 283
rect 1986 249 2079 255
rect 2113 249 2181 255
rect 2215 249 2382 255
rect 1986 215 2003 249
rect 2037 221 2079 249
rect 2037 215 2081 221
rect 2115 215 2149 249
rect 2215 221 2227 249
rect 2183 215 2227 221
rect 2261 215 2305 249
rect 2339 215 2382 249
rect 1986 179 2382 215
rect 1891 72 1899 106
rect 1933 72 1941 106
rect 1891 56 1941 72
rect 1986 106 2039 122
rect 1986 72 1995 106
rect 2029 72 2039 106
rect 1986 17 2039 72
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2484 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 335 249 369 255
rect 437 249 471 255
rect 335 221 369 249
rect 437 221 447 249
rect 447 221 471 249
rect 2079 249 2113 255
rect 2181 249 2215 255
rect 2079 221 2081 249
rect 2081 221 2113 249
rect 2181 221 2183 249
rect 2183 221 2215 249
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
<< metal1 >>
rect 0 561 2484 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2484 561
rect 0 496 2484 527
rect 323 255 483 261
rect 323 221 335 255
rect 369 221 437 255
rect 471 252 483 255
rect 2057 255 2227 261
rect 2057 252 2079 255
rect 471 224 2079 252
rect 471 221 483 224
rect 323 215 483 221
rect 2057 221 2079 224
rect 2113 221 2181 255
rect 2215 221 2227 255
rect 2057 215 2227 221
rect 0 17 2484 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2484 17
rect 0 -48 2484 -17
<< labels >>
flabel corelocali s 1058 306 1058 306 0 FreeSans 400 0 0 0 Y
port 6 nsew
flabel corelocali s 397 221 431 255 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew
rlabel comment s 0 0 0 0 4 clkinv_16
<< properties >>
string FIXED_BBOX 0 0 2484 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1797500
string GDS_START 1783280
<< end >>
