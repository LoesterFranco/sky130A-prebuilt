magic
tech sky130A
magscale 1 2
timestamp 1601050088
<< locali >>
rect 127 364 193 596
rect 127 226 161 364
rect 309 286 375 356
rect 409 286 500 356
rect 542 286 647 356
rect 681 260 747 356
rect 107 164 173 226
rect 107 70 158 164
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 27 364 93 649
rect 227 458 358 649
rect 470 424 536 588
rect 227 390 536 424
rect 680 390 746 649
rect 227 326 261 390
rect 195 260 261 326
rect 227 226 261 260
rect 21 17 73 226
rect 227 176 459 226
rect 401 160 459 176
rect 493 192 745 226
rect 193 17 259 128
rect 301 104 367 142
rect 493 104 559 192
rect 301 70 559 104
rect 593 17 659 158
rect 695 70 745 192
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel locali s 681 260 747 356 6 A1
port 1 nsew signal input
rlabel locali s 542 286 647 356 6 A2
port 2 nsew signal input
rlabel locali s 309 286 375 356 6 B1
port 3 nsew signal input
rlabel locali s 409 286 500 356 6 B2
port 4 nsew signal input
rlabel locali s 127 364 193 596 6 X
port 5 nsew signal output
rlabel locali s 127 226 161 364 6 X
port 5 nsew signal output
rlabel locali s 107 164 173 226 6 X
port 5 nsew signal output
rlabel locali s 107 70 158 164 6 X
port 5 nsew signal output
rlabel metal1 s 0 -49 768 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 768 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1282800
string GDS_START 1275870
<< end >>
