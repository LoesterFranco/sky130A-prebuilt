magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 136 333 212 493
rect 324 333 400 493
rect 512 333 588 493
rect 700 333 776 493
rect 17 299 901 333
rect 17 181 86 299
rect 136 215 777 265
rect 837 181 901 299
rect 17 143 901 181
rect 136 51 212 143
rect 324 51 400 143
rect 512 51 588 143
rect 700 51 776 143
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 51 367 102 527
rect 256 367 290 527
rect 444 367 478 527
rect 632 367 666 527
rect 820 367 880 527
rect 51 17 102 109
rect 256 17 290 109
rect 444 17 478 109
rect 632 17 666 109
rect 820 17 881 109
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
rlabel locali s 136 215 777 265 6 A
port 1 nsew signal input
rlabel locali s 837 181 901 299 6 Y
port 2 nsew signal output
rlabel locali s 700 333 776 493 6 Y
port 2 nsew signal output
rlabel locali s 700 51 776 143 6 Y
port 2 nsew signal output
rlabel locali s 512 333 588 493 6 Y
port 2 nsew signal output
rlabel locali s 512 51 588 143 6 Y
port 2 nsew signal output
rlabel locali s 324 333 400 493 6 Y
port 2 nsew signal output
rlabel locali s 324 51 400 143 6 Y
port 2 nsew signal output
rlabel locali s 136 333 212 493 6 Y
port 2 nsew signal output
rlabel locali s 136 51 212 143 6 Y
port 2 nsew signal output
rlabel locali s 17 299 901 333 6 Y
port 2 nsew signal output
rlabel locali s 17 181 86 299 6 Y
port 2 nsew signal output
rlabel locali s 17 143 901 181 6 Y
port 2 nsew signal output
rlabel metal1 s 0 -48 920 48 8 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 496 920 592 6 VPWR
port 4 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 920 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2121748
string GDS_START 2113832
<< end >>
