magic
tech sky130A
magscale 1 2
timestamp 1604502697
<< nwell >>
rect -38 261 1786 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 80 47 110 177
rect 176 47 206 177
rect 282 47 312 177
rect 368 47 398 177
rect 464 47 494 177
rect 560 47 590 177
rect 666 47 696 177
rect 764 47 794 177
rect 856 47 886 177
rect 952 47 982 177
rect 1058 47 1088 177
rect 1142 47 1172 177
rect 1236 47 1266 177
rect 1330 47 1360 177
rect 1434 47 1464 177
rect 1540 47 1570 177
<< pmoshvt >>
rect 82 297 118 497
rect 178 297 214 497
rect 274 297 310 497
rect 370 297 406 497
rect 466 297 502 497
rect 562 297 598 497
rect 658 297 694 497
rect 754 297 790 497
rect 858 297 894 497
rect 954 297 990 497
rect 1050 297 1086 497
rect 1144 297 1180 497
rect 1238 297 1274 497
rect 1332 297 1368 497
rect 1426 297 1462 497
rect 1520 297 1556 497
<< ndiff >>
rect 27 157 80 177
rect 27 123 35 157
rect 69 123 80 157
rect 27 47 80 123
rect 110 89 176 177
rect 110 55 131 89
rect 165 55 176 89
rect 110 47 176 55
rect 206 159 282 177
rect 206 125 227 159
rect 261 125 282 159
rect 206 47 282 125
rect 312 89 368 177
rect 312 55 323 89
rect 357 55 368 89
rect 312 47 368 55
rect 398 159 464 177
rect 398 125 419 159
rect 453 125 464 159
rect 398 47 464 125
rect 494 89 560 177
rect 494 55 515 89
rect 549 55 560 89
rect 494 47 560 55
rect 590 159 666 177
rect 590 125 611 159
rect 645 125 666 159
rect 590 47 666 125
rect 696 89 764 177
rect 696 55 707 89
rect 741 55 764 89
rect 696 47 764 55
rect 794 116 856 177
rect 794 82 807 116
rect 841 82 856 116
rect 794 47 856 82
rect 886 163 952 177
rect 886 129 907 163
rect 941 129 952 163
rect 886 47 952 129
rect 982 90 1058 177
rect 982 56 1003 90
rect 1037 56 1058 90
rect 982 47 1058 56
rect 1088 47 1142 177
rect 1172 90 1236 177
rect 1172 56 1192 90
rect 1226 56 1236 90
rect 1172 47 1236 56
rect 1266 162 1330 177
rect 1266 128 1286 162
rect 1320 128 1330 162
rect 1266 47 1330 128
rect 1360 90 1434 177
rect 1360 56 1380 90
rect 1414 56 1434 90
rect 1360 47 1434 56
rect 1464 47 1540 177
rect 1570 96 1649 177
rect 1570 62 1581 96
rect 1615 62 1649 96
rect 1570 47 1649 62
<< pdiff >>
rect 27 485 82 497
rect 27 451 35 485
rect 69 451 82 485
rect 27 383 82 451
rect 27 349 35 383
rect 69 349 82 383
rect 27 297 82 349
rect 118 422 178 497
rect 118 388 131 422
rect 165 388 178 422
rect 118 297 178 388
rect 214 489 274 497
rect 214 455 227 489
rect 261 455 274 489
rect 214 297 274 455
rect 310 449 370 497
rect 310 415 323 449
rect 357 415 370 449
rect 310 297 370 415
rect 406 405 466 497
rect 406 371 419 405
rect 453 371 466 405
rect 406 297 466 371
rect 502 489 562 497
rect 502 455 515 489
rect 549 455 562 489
rect 502 297 562 455
rect 598 405 658 497
rect 598 371 611 405
rect 645 371 658 405
rect 598 297 658 371
rect 694 489 754 497
rect 694 455 707 489
rect 741 455 754 489
rect 694 297 754 455
rect 790 489 858 497
rect 790 455 807 489
rect 841 455 858 489
rect 790 297 858 455
rect 894 405 954 497
rect 894 371 907 405
rect 941 371 954 405
rect 894 297 954 371
rect 990 489 1050 497
rect 990 455 1003 489
rect 1037 455 1050 489
rect 990 297 1050 455
rect 1086 405 1144 497
rect 1086 371 1098 405
rect 1132 371 1144 405
rect 1086 297 1144 371
rect 1180 489 1238 497
rect 1180 455 1192 489
rect 1226 455 1238 489
rect 1180 297 1238 455
rect 1274 405 1332 497
rect 1274 371 1286 405
rect 1320 371 1332 405
rect 1274 297 1332 371
rect 1368 489 1426 497
rect 1368 455 1380 489
rect 1414 455 1426 489
rect 1368 297 1426 455
rect 1462 405 1520 497
rect 1462 371 1474 405
rect 1508 371 1520 405
rect 1462 297 1520 371
rect 1556 489 1693 497
rect 1556 455 1647 489
rect 1681 455 1693 489
rect 1556 297 1693 455
<< ndiffc >>
rect 35 123 69 157
rect 131 55 165 89
rect 227 125 261 159
rect 323 55 357 89
rect 419 125 453 159
rect 515 55 549 89
rect 611 125 645 159
rect 707 55 741 89
rect 807 82 841 116
rect 907 129 941 163
rect 1003 56 1037 90
rect 1192 56 1226 90
rect 1286 128 1320 162
rect 1380 56 1414 90
rect 1581 62 1615 96
<< pdiffc >>
rect 35 451 69 485
rect 35 349 69 383
rect 131 388 165 422
rect 227 455 261 489
rect 323 415 357 449
rect 419 371 453 405
rect 515 455 549 489
rect 611 371 645 405
rect 707 455 741 489
rect 807 455 841 489
rect 907 371 941 405
rect 1003 455 1037 489
rect 1098 371 1132 405
rect 1192 455 1226 489
rect 1286 371 1320 405
rect 1380 455 1414 489
rect 1474 371 1508 405
rect 1647 455 1681 489
<< poly >>
rect 82 497 118 523
rect 178 497 214 523
rect 274 497 310 523
rect 370 497 406 523
rect 466 497 502 523
rect 562 497 598 523
rect 658 497 694 523
rect 754 497 790 523
rect 858 497 894 523
rect 954 497 990 523
rect 1050 497 1086 523
rect 1144 497 1180 523
rect 1238 497 1274 523
rect 1332 497 1368 523
rect 1426 497 1462 523
rect 1520 497 1556 523
rect 82 282 118 297
rect 178 282 214 297
rect 274 282 310 297
rect 370 282 406 297
rect 466 282 502 297
rect 562 282 598 297
rect 658 282 694 297
rect 754 282 790 297
rect 858 282 894 297
rect 954 282 990 297
rect 1050 282 1086 297
rect 1144 282 1180 297
rect 1238 282 1274 297
rect 1332 282 1368 297
rect 1426 282 1462 297
rect 1520 282 1556 297
rect 80 265 120 282
rect 176 265 216 282
rect 272 265 312 282
rect 80 249 312 265
rect 80 215 96 249
rect 130 215 174 249
rect 208 215 252 249
rect 286 215 312 249
rect 80 199 312 215
rect 80 177 110 199
rect 176 177 206 199
rect 282 177 312 199
rect 368 275 408 282
rect 464 275 504 282
rect 560 275 600 282
rect 656 275 696 282
rect 368 249 696 275
rect 752 265 792 282
rect 856 265 896 282
rect 952 265 992 282
rect 1048 265 1088 282
rect 368 215 387 249
rect 421 215 465 249
rect 499 215 543 249
rect 577 215 621 249
rect 655 215 696 249
rect 368 199 696 215
rect 738 249 814 265
rect 738 215 754 249
rect 788 215 814 249
rect 738 199 814 215
rect 856 249 1088 265
rect 856 215 872 249
rect 906 215 950 249
rect 984 215 1028 249
rect 1062 215 1088 249
rect 856 199 1088 215
rect 368 177 398 199
rect 464 177 494 199
rect 560 177 590 199
rect 666 177 696 199
rect 764 177 794 199
rect 856 177 886 199
rect 952 177 982 199
rect 1058 177 1088 199
rect 1142 265 1182 282
rect 1236 265 1276 282
rect 1330 265 1370 282
rect 1424 265 1464 282
rect 1518 265 1558 282
rect 1142 249 1464 265
rect 1142 215 1222 249
rect 1256 215 1300 249
rect 1334 215 1378 249
rect 1412 215 1464 249
rect 1142 199 1464 215
rect 1506 249 1570 265
rect 1506 215 1516 249
rect 1550 215 1570 249
rect 1506 199 1570 215
rect 1142 177 1172 199
rect 1236 177 1266 199
rect 1330 177 1360 199
rect 1434 177 1464 199
rect 1540 177 1570 199
rect 80 21 110 47
rect 176 21 206 47
rect 282 21 312 47
rect 368 21 398 47
rect 464 21 494 47
rect 560 21 590 47
rect 666 21 696 47
rect 764 21 794 47
rect 856 21 886 47
rect 952 21 982 47
rect 1058 21 1088 47
rect 1142 21 1172 47
rect 1236 21 1266 47
rect 1330 21 1360 47
rect 1434 21 1464 47
rect 1540 21 1570 47
<< polycont >>
rect 96 215 130 249
rect 174 215 208 249
rect 252 215 286 249
rect 387 215 421 249
rect 465 215 499 249
rect 543 215 577 249
rect 621 215 655 249
rect 754 215 788 249
rect 872 215 906 249
rect 950 215 984 249
rect 1028 215 1062 249
rect 1222 215 1256 249
rect 1300 215 1334 249
rect 1378 215 1412 249
rect 1516 215 1550 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 18 485 77 527
rect 18 451 35 485
rect 69 451 77 485
rect 201 489 277 527
rect 201 455 227 489
rect 261 455 277 489
rect 321 489 757 493
rect 321 455 515 489
rect 549 455 707 489
rect 741 455 757 489
rect 803 489 857 527
rect 803 455 807 489
rect 841 455 857 489
rect 977 489 1053 527
rect 977 455 1003 489
rect 1037 455 1053 489
rect 1166 489 1242 527
rect 1166 455 1192 489
rect 1226 455 1242 489
rect 1354 489 1431 527
rect 1354 455 1380 489
rect 1414 455 1431 489
rect 1631 489 1697 527
rect 1631 455 1647 489
rect 1681 455 1697 489
rect 18 383 77 451
rect 321 449 357 455
rect 18 349 35 383
rect 69 349 77 383
rect 121 422 165 438
rect 121 388 131 422
rect 321 421 323 449
rect 165 415 323 421
rect 803 439 857 455
rect 165 388 357 415
rect 121 387 357 388
rect 391 405 764 421
rect 899 405 1696 421
rect 121 372 165 387
rect 391 371 419 405
rect 453 371 611 405
rect 645 371 907 405
rect 941 371 1098 405
rect 1132 371 1286 405
rect 1320 371 1474 405
rect 1508 371 1696 405
rect 18 333 77 349
rect 203 303 806 337
rect 203 266 312 303
rect 80 249 312 266
rect 80 215 96 249
rect 130 215 174 249
rect 208 215 252 249
rect 286 215 312 249
rect 371 249 706 269
rect 371 215 387 249
rect 421 215 465 249
rect 499 215 543 249
rect 577 215 621 249
rect 655 215 706 249
rect 740 249 806 303
rect 942 303 1560 337
rect 942 282 1105 303
rect 740 215 754 249
rect 788 215 806 249
rect 740 199 806 215
rect 840 249 1105 282
rect 840 215 872 249
rect 906 215 950 249
rect 984 215 1028 249
rect 1062 215 1105 249
rect 1194 249 1428 269
rect 1194 215 1222 249
rect 1256 215 1300 249
rect 1334 215 1378 249
rect 1412 215 1428 249
rect 1516 249 1560 303
rect 1550 215 1560 249
rect 840 199 1105 215
rect 1516 199 1560 215
rect 1596 268 1696 371
rect 31 159 696 181
rect 1596 165 1632 268
rect 31 157 227 159
rect 31 123 35 157
rect 69 125 227 157
rect 261 125 419 159
rect 453 125 611 159
rect 645 125 847 159
rect 881 129 907 163
rect 941 162 1374 163
rect 941 129 1286 162
rect 881 128 1286 129
rect 1320 128 1374 162
rect 881 127 1374 128
rect 1453 131 1632 165
rect 69 123 71 125
rect 31 107 71 123
rect 225 119 268 125
rect 105 55 131 89
rect 165 55 181 89
rect 225 85 234 119
rect 801 116 847 125
rect 307 89 373 91
rect 105 17 181 55
rect 307 55 323 89
rect 357 55 373 89
rect 307 17 373 55
rect 489 55 515 89
rect 549 55 565 89
rect 489 17 565 55
rect 681 55 707 89
rect 741 55 757 89
rect 681 17 757 55
rect 801 82 807 116
rect 841 91 847 116
rect 841 90 1094 91
rect 1453 90 1497 131
rect 841 82 1003 90
rect 801 56 1003 82
rect 1037 56 1094 90
rect 801 51 1094 56
rect 1166 56 1192 90
rect 1226 56 1380 90
rect 1414 56 1497 90
rect 1546 62 1581 96
rect 1615 85 1664 96
rect 1615 62 1698 85
rect 1166 54 1497 56
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 234 85 268 119
rect 1664 85 1698 119
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
<< metal1 >>
rect 0 561 1748 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 0 496 1748 527
rect 222 119 280 125
rect 222 85 234 119
rect 268 116 280 119
rect 1652 119 1710 125
rect 1652 116 1664 119
rect 268 88 1664 116
rect 268 85 280 88
rect 222 79 280 85
rect 1652 85 1664 88
rect 1698 85 1710 119
rect 1652 79 1710 85
rect 0 17 1748 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
rect 0 -48 1748 -17
<< labels >>
flabel corelocali s 215 289 249 323 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 967 306 967 306 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 415 238 415 238 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 1243 238 1243 238 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 1599 357 1633 391 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
rlabel comment s 0 0 0 0 4 o211ai_4
<< properties >>
string FIXED_BBOX 0 0 1748 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 979962
string GDS_START 969190
<< end >>
