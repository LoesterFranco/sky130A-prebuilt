magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 86 199 166 339
rect 200 199 268 265
rect 541 425 679 491
rect 831 299 891 493
rect 568 199 719 265
rect 852 152 891 299
rect 831 83 891 152
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 17 407 69 491
rect 103 441 179 527
rect 327 441 486 475
rect 17 373 408 407
rect 17 165 52 373
rect 209 305 340 339
rect 302 249 340 305
rect 374 317 408 373
rect 452 391 486 441
rect 452 357 679 391
rect 723 367 779 527
rect 645 333 679 357
rect 374 283 514 317
rect 645 299 787 333
rect 302 215 391 249
rect 302 165 340 215
rect 480 199 514 283
rect 753 265 787 299
rect 753 199 808 265
rect 753 165 787 199
rect 17 90 81 165
rect 142 17 176 165
rect 236 131 340 165
rect 438 131 787 165
rect 930 288 964 527
rect 236 90 270 131
rect 319 17 394 97
rect 438 61 472 131
rect 509 17 585 97
rect 629 61 663 131
rect 697 17 783 97
rect 930 17 964 183
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
rlabel locali s 568 199 719 265 6 A
port 1 nsew signal input
rlabel locali s 541 425 679 491 6 B
port 2 nsew signal input
rlabel locali s 86 199 166 339 6 C_N
port 3 nsew signal input
rlabel locali s 200 199 268 265 6 D_N
port 4 nsew signal input
rlabel locali s 852 152 891 299 6 X
port 5 nsew signal output
rlabel locali s 831 299 891 493 6 X
port 5 nsew signal output
rlabel locali s 831 83 891 152 6 X
port 5 nsew signal output
rlabel metal1 s 0 -48 1012 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 1012 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1012 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 8094
string GDS_START 134
<< end >>
