magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 644 561
rect 17 425 77 527
rect 211 425 337 527
rect 453 425 529 459
rect 563 425 623 527
rect 495 391 529 425
rect 85 289 393 323
rect 85 199 134 289
rect 186 215 325 255
rect 359 249 393 289
rect 495 351 627 391
rect 359 215 479 249
rect 211 17 245 181
rect 593 165 627 351
rect 379 17 449 95
rect 563 69 627 165
rect 0 -17 644 17
<< obsli1 >>
rect 111 391 177 493
rect 17 357 461 391
rect 17 165 51 357
rect 427 317 461 357
rect 427 283 559 317
rect 525 199 559 283
rect 17 56 110 165
rect 279 165 461 181
rect 279 147 529 165
rect 279 51 345 147
rect 427 131 529 147
rect 483 51 529 131
<< metal1 >>
rect 0 496 644 592
rect 0 -48 644 48
<< labels >>
rlabel locali s 186 215 325 255 6 A
port 1 nsew signal input
rlabel locali s 359 249 393 289 6 B
port 2 nsew signal input
rlabel locali s 359 215 479 249 6 B
port 2 nsew signal input
rlabel locali s 85 289 393 323 6 B
port 2 nsew signal input
rlabel locali s 85 199 134 289 6 B
port 2 nsew signal input
rlabel locali s 593 165 627 351 6 Y
port 3 nsew signal output
rlabel locali s 563 69 627 165 6 Y
port 3 nsew signal output
rlabel locali s 495 391 529 425 6 Y
port 3 nsew signal output
rlabel locali s 495 351 627 391 6 Y
port 3 nsew signal output
rlabel locali s 453 425 529 459 6 Y
port 3 nsew signal output
rlabel locali s 379 17 449 95 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 211 17 245 181 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 644 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 644 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 563 425 623 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 211 425 337 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 17 425 77 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 644 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 644 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 632352
string GDS_START 627048
<< end >>
