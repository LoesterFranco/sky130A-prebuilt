magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1196 561
rect 103 333 169 419
rect 287 435 321 527
rect 555 333 621 417
rect 103 299 621 333
rect 924 367 965 527
rect 1099 299 1143 527
rect 18 215 169 265
rect 203 215 341 265
rect 375 221 434 299
rect 375 181 409 221
rect 481 215 613 265
rect 674 215 896 265
rect 950 215 1173 265
rect 103 131 409 181
rect 524 17 590 109
rect 727 17 761 109
rect 981 17 1047 109
rect 0 -17 1196 17
<< obsli1 >>
rect 18 459 253 493
rect 18 299 69 459
rect 203 401 253 459
rect 355 401 421 491
rect 203 367 421 401
rect 467 451 877 489
rect 467 367 517 451
rect 655 299 689 451
rect 723 333 789 417
rect 827 367 877 451
rect 999 333 1065 492
rect 723 299 1065 333
rect 18 97 69 181
rect 447 143 1151 181
rect 447 97 481 143
rect 18 51 481 97
rect 627 51 693 143
rect 811 51 945 143
rect 1085 51 1151 143
<< metal1 >>
rect 0 496 1196 592
rect 0 -48 1196 48
<< labels >>
rlabel locali s 950 215 1173 265 6 A1
port 1 nsew signal input
rlabel locali s 674 215 896 265 6 A2
port 2 nsew signal input
rlabel locali s 481 215 613 265 6 A3
port 3 nsew signal input
rlabel locali s 203 215 341 265 6 B1
port 4 nsew signal input
rlabel locali s 18 215 169 265 6 B2
port 5 nsew signal input
rlabel locali s 555 333 621 417 6 Y
port 6 nsew signal output
rlabel locali s 375 221 434 299 6 Y
port 6 nsew signal output
rlabel locali s 375 181 409 221 6 Y
port 6 nsew signal output
rlabel locali s 103 333 169 419 6 Y
port 6 nsew signal output
rlabel locali s 103 299 621 333 6 Y
port 6 nsew signal output
rlabel locali s 103 131 409 181 6 Y
port 6 nsew signal output
rlabel locali s 981 17 1047 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 727 17 761 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 524 17 590 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 1196 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1196 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1099 299 1143 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 924 367 965 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 287 435 321 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 1196 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 1196 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 905868
string GDS_START 895942
<< end >>
