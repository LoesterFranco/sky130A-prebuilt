magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 364 424 430 596
rect 564 424 686 596
rect 934 424 1056 596
rect 1464 424 1602 596
rect 364 390 1703 424
rect 25 270 455 356
rect 505 270 839 356
rect 889 270 1232 356
rect 1347 270 1617 356
rect 1657 226 1703 390
rect 1349 176 1703 226
rect 1363 160 1401 176
rect 1551 160 1589 176
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 23 390 330 649
rect 464 458 530 649
rect 720 458 900 649
rect 1090 458 1428 649
rect 1638 458 1704 649
rect 23 202 515 236
rect 23 70 89 202
rect 123 17 189 168
rect 223 70 289 202
rect 323 17 389 168
rect 449 136 515 202
rect 549 176 1243 226
rect 549 170 787 176
rect 1019 160 1057 176
rect 1191 160 1229 176
rect 449 70 873 136
rect 919 104 985 142
rect 1091 104 1157 142
rect 1263 104 1329 142
rect 1435 104 1501 142
rect 1639 104 1705 142
rect 919 70 1705 104
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
<< metal1 >>
rect 0 683 1728 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 0 617 1728 649
rect 0 17 1728 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
rect 0 -49 1728 -17
<< labels >>
rlabel locali s 1347 270 1617 356 6 A
port 1 nsew signal input
rlabel locali s 889 270 1232 356 6 B
port 2 nsew signal input
rlabel locali s 505 270 839 356 6 C
port 3 nsew signal input
rlabel locali s 25 270 455 356 6 D
port 4 nsew signal input
rlabel locali s 1657 226 1703 390 6 Y
port 5 nsew signal output
rlabel locali s 1551 160 1589 176 6 Y
port 5 nsew signal output
rlabel locali s 1464 424 1602 596 6 Y
port 5 nsew signal output
rlabel locali s 1363 160 1401 176 6 Y
port 5 nsew signal output
rlabel locali s 1349 176 1703 226 6 Y
port 5 nsew signal output
rlabel locali s 934 424 1056 596 6 Y
port 5 nsew signal output
rlabel locali s 564 424 686 596 6 Y
port 5 nsew signal output
rlabel locali s 364 424 430 596 6 Y
port 5 nsew signal output
rlabel locali s 364 390 1703 424 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -49 1728 49 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1728 715 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1728 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1762834
string GDS_START 1748584
<< end >>
