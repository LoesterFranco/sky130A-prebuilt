magic
tech sky130A
magscale 1 2
timestamp 1604502710
<< nwell >>
rect -38 332 998 704
<< pwell >>
rect 0 0 960 49
<< scpmos >>
rect 113 392 149 592
rect 203 392 239 592
rect 293 392 329 592
rect 513 378 549 578
rect 591 378 627 578
rect 693 368 729 592
rect 783 368 819 592
<< nmoslvt >>
rect 119 74 149 222
rect 191 74 221 222
rect 299 74 329 222
rect 499 74 529 184
rect 585 74 615 184
rect 693 74 723 222
rect 779 74 809 222
<< ndiff >>
rect 62 196 119 222
rect 62 162 74 196
rect 108 162 119 196
rect 62 120 119 162
rect 62 86 74 120
rect 108 86 119 120
rect 62 74 119 86
rect 149 74 191 222
rect 221 199 299 222
rect 221 165 243 199
rect 277 165 299 199
rect 221 116 299 165
rect 221 82 243 116
rect 277 82 299 116
rect 221 74 299 82
rect 329 184 379 222
rect 643 184 693 222
rect 329 127 499 184
rect 329 93 346 127
rect 380 93 454 127
rect 488 93 499 127
rect 329 74 499 93
rect 529 146 585 184
rect 529 112 540 146
rect 574 112 585 146
rect 529 74 585 112
rect 615 146 693 184
rect 615 112 627 146
rect 661 112 693 146
rect 615 74 693 112
rect 723 210 779 222
rect 723 176 734 210
rect 768 176 779 210
rect 723 120 779 176
rect 723 86 734 120
rect 768 86 779 120
rect 723 74 779 86
rect 809 210 862 222
rect 809 176 820 210
rect 854 176 862 210
rect 809 120 862 176
rect 809 86 820 120
rect 854 86 862 120
rect 809 74 862 86
<< pdiff >>
rect 61 580 113 592
rect 61 546 69 580
rect 103 546 113 580
rect 61 509 113 546
rect 61 475 69 509
rect 103 475 113 509
rect 61 438 113 475
rect 61 404 69 438
rect 103 404 113 438
rect 61 392 113 404
rect 149 580 203 592
rect 149 546 159 580
rect 193 546 203 580
rect 149 462 203 546
rect 149 428 159 462
rect 193 428 203 462
rect 149 392 203 428
rect 239 580 293 592
rect 239 546 249 580
rect 283 546 293 580
rect 239 509 293 546
rect 239 475 249 509
rect 283 475 293 509
rect 239 438 293 475
rect 239 404 249 438
rect 283 404 293 438
rect 239 392 293 404
rect 329 580 381 592
rect 329 546 339 580
rect 373 546 381 580
rect 643 578 693 592
rect 329 509 381 546
rect 329 475 339 509
rect 373 475 381 509
rect 329 438 381 475
rect 329 404 339 438
rect 373 404 381 438
rect 329 392 381 404
rect 461 512 513 578
rect 461 478 469 512
rect 503 478 513 512
rect 461 427 513 478
rect 461 393 469 427
rect 503 393 513 427
rect 461 378 513 393
rect 549 378 591 578
rect 627 566 693 578
rect 627 532 643 566
rect 677 532 693 566
rect 627 378 693 532
rect 643 368 693 378
rect 729 414 783 592
rect 729 380 739 414
rect 773 380 783 414
rect 729 368 783 380
rect 819 573 871 592
rect 819 539 829 573
rect 863 539 871 573
rect 819 368 871 539
<< ndiffc >>
rect 74 162 108 196
rect 74 86 108 120
rect 243 165 277 199
rect 243 82 277 116
rect 346 93 380 127
rect 454 93 488 127
rect 540 112 574 146
rect 627 112 661 146
rect 734 176 768 210
rect 734 86 768 120
rect 820 176 854 210
rect 820 86 854 120
<< pdiffc >>
rect 69 546 103 580
rect 69 475 103 509
rect 69 404 103 438
rect 159 546 193 580
rect 159 428 193 462
rect 249 546 283 580
rect 249 475 283 509
rect 249 404 283 438
rect 339 546 373 580
rect 339 475 373 509
rect 339 404 373 438
rect 469 478 503 512
rect 469 393 503 427
rect 643 532 677 566
rect 739 380 773 414
rect 829 539 863 573
<< poly >>
rect 113 592 149 618
rect 203 592 239 618
rect 293 592 329 618
rect 513 578 549 604
rect 591 578 627 604
rect 693 592 729 618
rect 783 592 819 618
rect 113 310 149 392
rect 203 310 239 392
rect 293 333 329 392
rect 299 310 329 333
rect 513 332 549 378
rect 21 294 149 310
rect 21 260 37 294
rect 71 260 149 294
rect 21 244 149 260
rect 119 222 149 244
rect 191 294 257 310
rect 191 260 207 294
rect 241 260 257 294
rect 191 244 257 260
rect 299 294 435 310
rect 513 302 543 332
rect 591 310 627 378
rect 693 336 729 368
rect 783 336 819 368
rect 693 320 884 336
rect 299 260 385 294
rect 419 260 435 294
rect 299 244 435 260
rect 477 286 543 302
rect 477 252 493 286
rect 527 252 543 286
rect 191 222 221 244
rect 299 222 329 244
rect 477 236 543 252
rect 585 294 651 310
rect 585 260 601 294
rect 635 260 651 294
rect 585 244 651 260
rect 693 306 834 320
rect 499 184 529 236
rect 585 184 615 244
rect 693 222 723 306
rect 779 286 834 306
rect 868 286 884 320
rect 779 270 884 286
rect 779 222 809 270
rect 119 48 149 74
rect 191 48 221 74
rect 299 48 329 74
rect 499 48 529 74
rect 585 48 615 74
rect 693 48 723 74
rect 779 48 809 74
<< polycont >>
rect 37 260 71 294
rect 207 260 241 294
rect 385 260 419 294
rect 493 252 527 286
rect 601 260 635 294
rect 834 286 868 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 53 580 103 596
rect 53 546 69 580
rect 53 509 103 546
rect 53 475 69 509
rect 53 438 103 475
rect 53 404 69 438
rect 143 580 209 649
rect 143 546 159 580
rect 193 546 209 580
rect 143 462 209 546
rect 143 428 159 462
rect 193 428 209 462
rect 143 412 209 428
rect 249 580 283 596
rect 249 509 283 546
rect 249 438 283 475
rect 53 378 103 404
rect 249 378 283 404
rect 53 344 283 378
rect 317 580 584 596
rect 317 546 339 580
rect 373 562 584 580
rect 373 546 389 562
rect 317 509 389 546
rect 317 475 339 509
rect 373 475 389 509
rect 317 438 389 475
rect 317 404 339 438
rect 373 404 389 438
rect 453 512 516 528
rect 453 478 469 512
rect 503 478 516 512
rect 453 427 516 478
rect 550 498 584 562
rect 621 566 699 649
rect 621 532 643 566
rect 677 532 699 566
rect 813 573 879 649
rect 813 539 829 573
rect 863 539 879 573
rect 813 532 879 539
rect 550 464 894 498
rect 317 310 351 404
rect 453 393 469 427
rect 503 393 516 427
rect 453 370 516 393
rect 21 294 87 310
rect 21 260 37 294
rect 71 260 87 294
rect 21 236 87 260
rect 121 294 263 310
rect 121 260 207 294
rect 241 260 263 294
rect 121 236 263 260
rect 297 276 351 310
rect 385 336 516 370
rect 385 294 435 336
rect 297 202 331 276
rect 58 196 124 202
rect 58 162 74 196
rect 108 162 124 196
rect 58 120 124 162
rect 58 86 74 120
rect 108 86 124 120
rect 58 17 124 86
rect 216 199 331 202
rect 216 165 243 199
rect 277 168 331 199
rect 419 260 435 294
rect 385 202 435 260
rect 477 286 551 302
rect 477 252 493 286
rect 527 252 551 286
rect 477 236 551 252
rect 585 294 651 430
rect 585 260 601 294
rect 635 260 651 294
rect 585 236 651 260
rect 697 414 784 430
rect 697 380 739 414
rect 773 380 784 414
rect 697 210 784 380
rect 818 320 894 464
rect 818 286 834 320
rect 868 286 894 320
rect 818 270 894 286
rect 385 168 574 202
rect 277 165 296 168
rect 216 116 296 165
rect 538 146 574 168
rect 216 82 243 116
rect 277 82 296 116
rect 216 70 296 82
rect 330 127 504 134
rect 330 93 346 127
rect 380 93 454 127
rect 488 93 504 127
rect 330 17 504 93
rect 538 112 540 146
rect 538 70 574 112
rect 610 146 663 188
rect 610 112 627 146
rect 661 112 663 146
rect 610 17 663 112
rect 697 176 734 210
rect 768 176 784 210
rect 697 120 784 176
rect 697 86 734 120
rect 768 86 784 120
rect 697 70 784 86
rect 820 210 870 226
rect 854 176 870 210
rect 820 120 870 176
rect 854 86 870 120
rect 820 17 870 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
rlabel comment s 0 0 0 0 4 a2bb2o_2
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 127 242 161 276 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 223 242 257 276 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 511 242 545 276 0 FreeSans 340 0 0 0 A2_N
port 2 nsew
flabel corelocali s 703 94 737 128 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 703 168 737 202 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 703 242 737 276 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 703 390 737 424 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 607 242 641 276 0 FreeSans 340 0 0 0 A1_N
port 1 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 A1_N
port 1 nsew
flabel corelocali s 607 390 641 424 0 FreeSans 340 0 0 0 A1_N
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 960 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3540562
string GDS_START 3532212
<< end >>
