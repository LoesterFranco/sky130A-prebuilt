magic
tech sky130A
magscale 1 2
timestamp 1601050082
<< locali >>
rect 25 241 110 375
rect 161 241 263 375
rect 297 296 363 362
rect 694 270 760 356
rect 2978 364 3055 596
rect 2815 238 2876 310
rect 3021 226 3055 364
rect 2983 70 3055 226
rect 3271 364 3343 596
rect 3309 210 3343 364
rect 3267 70 3343 210
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3360 683
rect 23 443 79 596
rect 113 477 179 649
rect 213 581 449 615
rect 213 443 247 581
rect 293 460 343 547
rect 383 464 449 581
rect 494 460 544 649
rect 578 460 650 596
rect 23 409 247 443
rect 309 430 343 460
rect 309 396 431 430
rect 397 262 431 396
rect 578 362 612 460
rect 696 424 746 596
rect 786 458 836 649
rect 696 390 828 424
rect 502 296 612 362
rect 297 228 512 262
rect 297 207 331 228
rect 28 17 94 207
rect 192 173 331 207
rect 192 115 258 173
rect 378 17 444 194
rect 478 85 512 228
rect 546 119 612 296
rect 794 334 828 390
rect 876 368 956 596
rect 1004 493 1054 649
rect 1088 581 1501 615
rect 1088 459 1122 581
rect 1385 564 1501 581
rect 990 425 1122 459
rect 1173 449 1239 547
rect 1273 496 1339 547
rect 1385 530 1586 564
rect 1625 530 1659 649
rect 1552 496 1586 530
rect 1699 496 1766 596
rect 1273 462 1518 496
rect 1205 428 1239 449
rect 990 393 1043 425
rect 1205 394 1450 428
rect 922 344 956 368
rect 1081 360 1151 381
rect 1081 344 1342 360
rect 794 268 888 334
rect 922 310 1342 344
rect 794 234 828 268
rect 922 234 958 310
rect 1276 294 1342 310
rect 658 184 828 234
rect 862 184 958 234
rect 992 241 1194 275
rect 1384 260 1450 394
rect 992 150 1026 241
rect 646 116 1026 150
rect 646 85 680 116
rect 478 51 680 85
rect 760 17 826 82
rect 1060 17 1126 207
rect 1160 85 1194 241
rect 1234 226 1450 260
rect 1234 119 1284 226
rect 1484 192 1518 462
rect 1319 158 1518 192
rect 1552 462 1766 496
rect 1810 494 1876 649
rect 1552 216 1586 462
rect 1732 460 1766 462
rect 1657 424 1698 428
rect 1732 426 1906 460
rect 1657 390 1663 424
rect 1697 392 1698 424
rect 1697 390 1798 392
rect 1657 358 1798 390
rect 1732 326 1798 358
rect 1840 326 1906 426
rect 1978 456 2044 596
rect 2180 594 2246 649
rect 2292 560 2358 596
rect 2399 594 2465 649
rect 2590 560 2656 596
rect 2133 526 2656 560
rect 1978 422 2082 456
rect 1620 292 1686 324
rect 1945 311 2014 388
rect 2048 379 2082 422
rect 2133 413 2199 526
rect 2234 458 2556 492
rect 2234 379 2268 458
rect 2048 345 2268 379
rect 1620 258 1911 292
rect 1319 85 1385 158
rect 1160 51 1385 85
rect 1430 85 1496 124
rect 1552 119 1618 216
rect 1652 85 1718 216
rect 1430 51 1718 85
rect 1759 17 1825 216
rect 1877 107 1911 258
rect 1945 252 2200 311
rect 2234 218 2268 345
rect 2326 390 2335 424
rect 2369 390 2392 424
rect 2326 294 2392 390
rect 2522 378 2556 458
rect 2590 476 2656 526
rect 2800 510 2938 649
rect 2590 442 2944 476
rect 2590 412 2656 442
rect 2522 344 2688 378
rect 2440 260 2506 310
rect 2554 294 2688 344
rect 2722 358 2826 408
rect 2722 260 2756 358
rect 2910 326 2944 442
rect 1949 184 2268 218
rect 2302 226 2781 260
rect 2910 260 2987 326
rect 1949 141 2116 184
rect 2302 150 2336 226
rect 2150 116 2336 150
rect 2150 107 2184 116
rect 1877 73 2184 107
rect 2387 85 2453 192
rect 2493 158 2713 192
rect 2493 119 2559 158
rect 2595 85 2645 124
rect 2283 17 2351 82
rect 2387 51 2645 85
rect 2679 100 2713 158
rect 2747 134 2781 226
rect 2910 204 2944 260
rect 2815 170 2944 204
rect 2815 100 2849 170
rect 2679 66 2849 100
rect 2883 17 2947 136
rect 3090 310 3140 556
rect 3181 380 3231 649
rect 3090 244 3275 310
rect 3090 70 3145 244
rect 3181 17 3231 210
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3360 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 3199 649 3233 683
rect 3295 649 3329 683
rect 1663 390 1697 424
rect 2335 390 2369 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
<< metal1 >>
rect 0 683 3360 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3360 683
rect 0 617 3360 649
rect 1651 424 1709 430
rect 1651 390 1663 424
rect 1697 421 1709 424
rect 2323 424 2381 430
rect 2323 421 2335 424
rect 1697 393 2335 421
rect 1697 390 1709 393
rect 1651 384 1709 390
rect 2323 390 2335 393
rect 2369 390 2381 424
rect 2323 384 2381 390
rect 0 17 3360 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3360 17
rect 0 -49 3360 -17
<< obsm1 >>
rect 1075 347 1133 356
rect 1939 347 1997 356
rect 1075 319 1997 347
rect 1075 310 1133 319
rect 1939 310 1997 319
<< labels >>
rlabel locali s 297 296 363 362 6 D
port 1 nsew signal input
rlabel locali s 3309 210 3343 364 6 Q
port 2 nsew signal output
rlabel locali s 3271 364 3343 596 6 Q
port 2 nsew signal output
rlabel locali s 3267 70 3343 210 6 Q
port 2 nsew signal output
rlabel locali s 3021 226 3055 364 6 Q_N
port 3 nsew signal output
rlabel locali s 2983 70 3055 226 6 Q_N
port 3 nsew signal output
rlabel locali s 2978 364 3055 596 6 Q_N
port 3 nsew signal output
rlabel locali s 2815 238 2876 310 6 RESET_B
port 4 nsew signal input
rlabel locali s 25 241 110 375 6 SCD
port 5 nsew signal input
rlabel locali s 161 241 263 375 6 SCE
port 6 nsew signal input
rlabel metal1 s 2323 421 2381 430 6 SET_B
port 7 nsew signal input
rlabel metal1 s 2323 384 2381 393 6 SET_B
port 7 nsew signal input
rlabel metal1 s 1651 421 1709 430 6 SET_B
port 7 nsew signal input
rlabel metal1 s 1651 393 2381 421 6 SET_B
port 7 nsew signal input
rlabel metal1 s 1651 384 1709 393 6 SET_B
port 7 nsew signal input
rlabel locali s 694 270 760 356 6 CLK_N
port 8 nsew clock input
rlabel metal1 s 0 -49 3360 49 8 VGND
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 617 3360 715 6 VPWR
port 10 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 3360 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 24514
string GDS_START 132
<< end >>
