magic
tech sky130A
magscale 1 2
timestamp 1604502741
<< locali >>
rect 25 260 91 356
rect 697 378 763 547
rect 877 378 943 547
rect 697 344 943 378
rect 697 310 763 344
rect 723 226 763 310
rect 807 236 1031 310
rect 723 202 773 226
rect 723 154 931 202
rect 897 119 931 154
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 35 390 85 649
rect 125 262 191 596
rect 237 330 287 596
rect 327 364 377 649
rect 417 330 467 596
rect 507 364 573 649
rect 607 581 1033 615
rect 607 330 657 581
rect 237 296 657 330
rect 803 412 837 581
rect 983 364 1033 581
rect 125 226 259 262
rect 23 17 73 226
rect 109 60 259 226
rect 293 228 687 262
rect 293 70 327 228
rect 363 17 429 194
rect 465 70 499 228
rect 535 17 601 194
rect 637 120 687 228
rect 637 85 861 120
rect 967 85 1033 202
rect 637 51 1033 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 683 1056 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 0 617 1056 649
rect 0 17 1056 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -49 1056 -17
<< labels >>
rlabel locali s 807 236 1031 310 6 A
port 1 nsew signal input
rlabel locali s 25 260 91 356 6 TE_B
port 2 nsew signal input
rlabel locali s 897 119 931 154 6 Z
port 3 nsew signal output
rlabel locali s 877 378 943 547 6 Z
port 3 nsew signal output
rlabel locali s 723 226 763 310 6 Z
port 3 nsew signal output
rlabel locali s 723 202 773 226 6 Z
port 3 nsew signal output
rlabel locali s 723 154 931 202 6 Z
port 3 nsew signal output
rlabel locali s 697 378 763 547 6 Z
port 3 nsew signal output
rlabel locali s 697 344 943 378 6 Z
port 3 nsew signal output
rlabel locali s 697 310 763 344 6 Z
port 3 nsew signal output
rlabel metal1 s 0 -49 1056 49 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 617 1056 715 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1056 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 2280866
string GDS_START 2271994
<< end >>
