magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 422 704
<< pwell >>
rect 0 0 384 49
<< scnmos >>
rect 79 47 305 202
<< scpmos >>
rect 79 368 305 619
<< ndiff >>
rect 27 190 79 202
rect 27 156 35 190
rect 69 156 79 190
rect 27 93 79 156
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 305 190 357 202
rect 305 156 315 190
rect 349 156 357 190
rect 305 93 357 156
rect 305 59 315 93
rect 349 59 357 93
rect 305 47 357 59
<< pdiff >>
rect 27 607 79 619
rect 27 573 35 607
rect 69 573 79 607
rect 27 510 79 573
rect 27 476 35 510
rect 69 476 79 510
rect 27 414 79 476
rect 27 380 35 414
rect 69 380 79 414
rect 27 368 79 380
rect 305 607 357 619
rect 305 573 315 607
rect 349 573 357 607
rect 305 510 357 573
rect 305 476 315 510
rect 349 476 357 510
rect 305 414 357 476
rect 305 380 315 414
rect 349 380 357 414
rect 305 368 357 380
<< ndiffc >>
rect 35 156 69 190
rect 35 59 69 93
rect 315 156 349 190
rect 315 59 349 93
<< pdiffc >>
rect 35 573 69 607
rect 35 476 69 510
rect 35 380 69 414
rect 315 573 349 607
rect 315 476 349 510
rect 315 380 349 414
<< poly >>
rect 79 619 305 645
rect 79 342 305 368
rect 79 320 148 342
rect 79 286 98 320
rect 132 286 148 320
rect 79 270 148 286
rect 238 284 305 300
rect 238 250 254 284
rect 288 250 305 284
rect 238 228 305 250
rect 79 202 305 228
rect 79 21 305 47
<< polycont >>
rect 98 286 132 320
rect 254 250 288 284
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 384 683
rect 17 607 367 649
rect 17 573 35 607
rect 69 573 315 607
rect 349 573 367 607
rect 17 510 367 573
rect 17 476 35 510
rect 69 476 315 510
rect 349 476 367 510
rect 17 414 367 476
rect 17 380 35 414
rect 69 380 315 414
rect 349 380 367 414
rect 17 354 367 380
rect 17 286 98 320
rect 132 286 178 320
rect 17 216 178 286
rect 212 284 367 354
rect 212 250 254 284
rect 288 250 367 284
rect 17 190 367 216
rect 17 156 35 190
rect 69 156 315 190
rect 349 156 367 190
rect 17 93 367 156
rect 17 59 35 93
rect 69 59 315 93
rect 349 59 367 93
rect 17 17 367 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 384 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
<< metal1 >>
rect 0 683 384 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 384 683
rect 0 617 384 649
rect 0 17 384 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 384 17
rect 0 -49 384 -17
<< labels >>
flabel metal1 s 0 617 384 666 0 FreeSans 340 0 0 0 VPWR
port 4 nsew
flabel metal1 s 0 0 384 49 0 FreeSans 340 0 0 0 VGND
port 1 nsew
rlabel comment s 0 0 0 0 4 decaphe_4
flabel nwell s 0 617 384 666 0 FreeSans 200 0 0 0 VPB
port 3 nsew
flabel pwell s 0 0 384 49 0 FreeSans 200 0 0 0 VNB
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 384 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2458340
string GDS_START 2455412
<< end >>
