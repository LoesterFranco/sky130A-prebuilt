magic
tech sky130A
magscale 1 2
timestamp 1604502693
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 84 47 114 177
rect 170 47 200 177
rect 256 47 286 177
rect 342 47 372 177
rect 535 47 565 177
rect 619 47 649 177
rect 711 47 741 177
rect 787 47 817 177
rect 871 47 901 177
rect 955 47 985 177
<< pmoshvt >>
rect 84 297 114 497
rect 170 297 200 497
rect 256 297 286 497
rect 342 297 372 497
rect 535 297 565 497
rect 619 297 649 497
rect 703 297 733 497
rect 787 297 817 497
rect 871 297 901 497
rect 955 297 985 497
<< ndiff >>
rect 27 89 84 177
rect 27 55 39 89
rect 73 55 84 89
rect 27 47 84 55
rect 114 157 170 177
rect 114 123 125 157
rect 159 123 170 157
rect 114 47 170 123
rect 200 89 256 177
rect 200 55 211 89
rect 245 55 256 89
rect 200 47 256 55
rect 286 157 342 177
rect 286 123 297 157
rect 331 123 342 157
rect 286 47 342 123
rect 372 89 535 177
rect 372 55 405 89
rect 439 55 487 89
rect 521 55 535 89
rect 372 47 535 55
rect 565 169 619 177
rect 565 135 575 169
rect 609 135 619 169
rect 565 101 619 135
rect 565 67 575 101
rect 609 67 619 101
rect 565 47 619 67
rect 649 89 711 177
rect 649 55 667 89
rect 701 55 711 89
rect 649 47 711 55
rect 741 47 787 177
rect 817 131 871 177
rect 817 97 827 131
rect 861 97 871 131
rect 817 47 871 97
rect 901 47 955 177
rect 985 161 1037 177
rect 985 127 995 161
rect 1029 127 1037 161
rect 985 93 1037 127
rect 985 59 995 93
rect 1029 59 1037 93
rect 985 47 1037 59
<< pdiff >>
rect 27 489 84 497
rect 27 455 39 489
rect 73 455 84 489
rect 27 421 84 455
rect 27 387 39 421
rect 73 387 84 421
rect 27 297 84 387
rect 114 421 170 497
rect 114 387 125 421
rect 159 387 170 421
rect 114 351 170 387
rect 114 317 125 351
rect 159 317 170 351
rect 114 297 170 317
rect 200 489 256 497
rect 200 455 211 489
rect 245 455 256 489
rect 200 421 256 455
rect 200 387 211 421
rect 245 387 256 421
rect 200 297 256 387
rect 286 421 342 497
rect 286 387 297 421
rect 331 387 342 421
rect 286 351 342 387
rect 286 317 297 351
rect 331 317 342 351
rect 286 297 342 317
rect 372 489 429 497
rect 372 455 383 489
rect 417 455 429 489
rect 372 421 429 455
rect 372 387 383 421
rect 417 387 429 421
rect 372 353 429 387
rect 372 319 383 353
rect 417 319 429 353
rect 372 297 429 319
rect 483 459 535 497
rect 483 425 491 459
rect 525 425 535 459
rect 483 389 535 425
rect 483 355 491 389
rect 525 355 535 389
rect 483 297 535 355
rect 565 409 619 497
rect 565 375 575 409
rect 609 375 619 409
rect 565 341 619 375
rect 565 307 575 341
rect 609 307 619 341
rect 565 297 619 307
rect 649 428 703 497
rect 649 394 659 428
rect 693 394 703 428
rect 649 339 703 394
rect 649 305 659 339
rect 693 305 703 339
rect 649 297 703 305
rect 733 489 787 497
rect 733 455 743 489
rect 777 455 787 489
rect 733 297 787 455
rect 817 477 871 497
rect 817 443 827 477
rect 861 443 871 477
rect 817 404 871 443
rect 817 370 827 404
rect 861 370 871 404
rect 817 297 871 370
rect 901 489 955 497
rect 901 455 911 489
rect 945 455 955 489
rect 901 297 955 455
rect 985 479 1064 497
rect 985 445 1022 479
rect 1056 445 1064 479
rect 985 411 1064 445
rect 985 377 1022 411
rect 1056 377 1064 411
rect 985 343 1064 377
rect 985 309 1022 343
rect 1056 309 1064 343
rect 985 297 1064 309
<< ndiffc >>
rect 39 55 73 89
rect 125 123 159 157
rect 211 55 245 89
rect 297 123 331 157
rect 405 55 439 89
rect 487 55 521 89
rect 575 135 609 169
rect 575 67 609 101
rect 667 55 701 89
rect 827 97 861 131
rect 995 127 1029 161
rect 995 59 1029 93
<< pdiffc >>
rect 39 455 73 489
rect 39 387 73 421
rect 125 387 159 421
rect 125 317 159 351
rect 211 455 245 489
rect 211 387 245 421
rect 297 387 331 421
rect 297 317 331 351
rect 383 455 417 489
rect 383 387 417 421
rect 383 319 417 353
rect 491 425 525 459
rect 491 355 525 389
rect 575 375 609 409
rect 575 307 609 341
rect 659 394 693 428
rect 659 305 693 339
rect 743 455 777 489
rect 827 443 861 477
rect 827 370 861 404
rect 911 455 945 489
rect 1022 445 1056 479
rect 1022 377 1056 411
rect 1022 309 1056 343
<< poly >>
rect 84 497 114 523
rect 170 497 200 523
rect 256 497 286 523
rect 342 497 372 523
rect 535 497 565 523
rect 619 497 649 523
rect 703 497 733 523
rect 787 497 817 523
rect 871 497 901 523
rect 955 497 985 523
rect 84 265 114 297
rect 170 265 200 297
rect 256 265 286 297
rect 342 265 372 297
rect 535 265 565 297
rect 619 265 649 297
rect 703 265 733 297
rect 787 265 817 297
rect 871 265 901 297
rect 84 249 395 265
rect 84 215 215 249
rect 249 215 283 249
rect 317 215 351 249
rect 385 215 395 249
rect 84 199 395 215
rect 497 249 649 265
rect 497 215 507 249
rect 541 215 649 249
rect 497 199 649 215
rect 691 249 745 265
rect 691 215 701 249
rect 735 215 745 249
rect 691 199 745 215
rect 787 249 901 265
rect 787 215 821 249
rect 855 215 901 249
rect 787 199 901 215
rect 84 177 114 199
rect 170 177 200 199
rect 256 177 286 199
rect 342 177 372 199
rect 535 177 565 199
rect 619 177 649 199
rect 711 177 741 199
rect 787 177 817 199
rect 871 177 901 199
rect 955 265 985 297
rect 955 249 1009 265
rect 955 215 965 249
rect 999 215 1009 249
rect 955 199 1009 215
rect 955 177 985 199
rect 84 21 114 47
rect 170 21 200 47
rect 256 21 286 47
rect 342 21 372 47
rect 535 21 565 47
rect 619 21 649 47
rect 711 21 741 47
rect 787 21 817 47
rect 871 21 901 47
rect 955 21 985 47
<< polycont >>
rect 215 215 249 249
rect 283 215 317 249
rect 351 215 385 249
rect 507 215 541 249
rect 701 215 735 249
rect 821 215 855 249
rect 965 215 999 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 23 489 89 527
rect 23 455 39 489
rect 73 455 89 489
rect 23 421 89 455
rect 195 489 261 527
rect 195 455 211 489
rect 245 455 261 489
rect 23 387 39 421
rect 73 387 89 421
rect 125 421 159 437
rect 195 421 261 455
rect 383 489 433 527
rect 417 455 433 489
rect 195 387 211 421
rect 245 387 261 421
rect 297 421 347 437
rect 331 387 347 421
rect 125 351 159 387
rect 297 351 347 387
rect 29 317 125 351
rect 159 317 297 351
rect 331 317 347 351
rect 383 421 433 455
rect 417 387 433 421
rect 383 353 433 387
rect 417 319 433 353
rect 491 459 693 493
rect 657 428 693 459
rect 727 489 793 527
rect 727 455 743 489
rect 777 455 793 489
rect 827 477 861 493
rect 491 389 525 425
rect 491 339 525 355
rect 575 409 609 425
rect 575 341 609 375
rect 29 157 126 317
rect 383 303 433 319
rect 160 249 441 265
rect 160 215 215 249
rect 249 215 283 249
rect 317 215 351 249
rect 385 215 441 249
rect 160 199 441 215
rect 479 249 541 305
rect 479 215 507 249
rect 479 199 541 215
rect 407 157 441 199
rect 575 169 609 307
rect 657 394 659 428
rect 895 489 961 527
rect 895 455 911 489
rect 945 455 961 489
rect 827 404 861 443
rect 1006 445 1022 479
rect 1056 445 1072 479
rect 1006 411 1072 445
rect 1006 404 1022 411
rect 693 394 827 404
rect 657 370 827 394
rect 861 377 1022 404
rect 1056 377 1072 411
rect 861 370 1072 377
rect 657 339 693 370
rect 657 305 659 339
rect 1021 343 1072 370
rect 657 289 693 305
rect 729 302 987 336
rect 729 255 764 302
rect 937 258 987 302
rect 1021 309 1022 343
rect 1056 309 1072 343
rect 1021 292 1072 309
rect 685 249 764 255
rect 685 215 701 249
rect 735 215 764 249
rect 685 202 764 215
rect 798 249 903 255
rect 798 215 821 249
rect 855 215 903 249
rect 798 202 903 215
rect 937 249 1020 258
rect 937 215 965 249
rect 999 215 1020 249
rect 937 211 1020 215
rect 29 123 125 157
rect 159 123 297 157
rect 331 123 347 157
rect 407 135 575 157
rect 609 135 873 168
rect 407 134 873 135
rect 407 123 609 134
rect 575 101 609 123
rect 21 55 39 89
rect 73 55 89 89
rect 21 17 89 55
rect 195 55 211 89
rect 245 55 261 89
rect 195 17 261 55
rect 382 55 405 89
rect 439 55 487 89
rect 521 55 537 89
rect 382 17 537 55
rect 817 131 873 134
rect 817 97 827 131
rect 861 97 873 131
rect 575 51 609 67
rect 651 55 667 89
rect 701 55 717 89
rect 817 81 873 97
rect 989 161 1045 177
rect 989 127 995 161
rect 1029 127 1045 161
rect 989 93 1045 127
rect 651 17 717 55
rect 989 59 995 93
rect 1029 59 1045 93
rect 989 17 1045 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
flabel corelocali s 953 289 987 323 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 861 221 895 255 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 29 289 63 323 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 493 221 527 255 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
rlabel comment s 0 0 0 0 4 a21o_4
<< properties >>
string FIXED_BBOX 0 0 1104 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 4028982
string GDS_START 4020818
string path 0.000 0.000 27.600 0.000 
<< end >>
