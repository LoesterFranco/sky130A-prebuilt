magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 552 561
rect 18 425 349 483
rect 383 367 439 527
rect 18 151 88 265
rect 122 199 264 323
rect 481 299 535 493
rect 298 199 379 265
rect 501 152 535 299
rect 19 17 85 117
rect 199 17 265 97
rect 367 17 443 97
rect 481 83 535 152
rect 0 -17 552 17
<< obsli1 >>
rect 18 357 336 391
rect 18 299 82 357
rect 302 333 336 357
rect 302 299 447 333
rect 413 265 447 299
rect 413 199 467 265
rect 413 165 447 199
rect 125 131 447 165
rect 125 61 159 131
rect 299 61 333 131
<< metal1 >>
rect 0 496 552 592
rect 0 -48 552 48
<< labels >>
rlabel locali s 298 199 379 265 6 A
port 1 nsew signal input
rlabel locali s 18 425 349 483 6 B
port 2 nsew signal input
rlabel locali s 122 199 264 323 6 C
port 3 nsew signal input
rlabel locali s 18 151 88 265 6 D
port 4 nsew signal input
rlabel locali s 501 152 535 299 6 X
port 5 nsew signal output
rlabel locali s 481 299 535 493 6 X
port 5 nsew signal output
rlabel locali s 481 83 535 152 6 X
port 5 nsew signal output
rlabel locali s 367 17 443 97 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 199 17 265 97 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 19 17 85 117 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 552 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 552 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 383 367 439 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 552 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 552 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 552 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1069060
string GDS_START 1063038
<< end >>
