magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 828 561
rect 103 369 190 527
rect 396 455 462 527
rect 659 353 725 425
rect 98 153 156 335
rect 381 325 725 353
rect 381 289 811 325
rect 190 153 256 255
rect 765 171 811 289
rect 103 17 170 119
rect 468 17 534 97
rect 659 127 811 171
rect 0 -17 828 17
<< obsli1 >>
rect 17 369 69 493
rect 17 255 64 369
rect 224 353 282 493
rect 320 421 362 493
rect 496 459 811 493
rect 496 421 625 459
rect 320 387 625 421
rect 759 359 811 459
rect 17 221 30 255
rect 17 123 64 221
rect 224 289 347 353
rect 290 255 347 289
rect 290 205 593 255
rect 649 221 676 255
rect 710 221 731 255
rect 649 205 731 221
rect 17 56 69 123
rect 290 119 346 205
rect 204 51 346 119
rect 380 131 625 171
rect 380 51 434 131
rect 568 93 625 131
rect 568 55 810 93
<< obsli1c >>
rect 30 221 64 255
rect 676 221 710 255
<< metal1 >>
rect 0 496 828 592
rect 0 -48 828 48
<< obsm1 >>
rect 17 255 76 261
rect 17 221 30 255
rect 64 252 76 255
rect 664 255 722 261
rect 664 252 676 255
rect 64 224 676 252
rect 64 221 76 224
rect 17 215 76 221
rect 664 221 676 224
rect 710 221 722 255
rect 664 215 722 221
<< labels >>
rlabel locali s 98 153 156 335 6 A
port 1 nsew signal input
rlabel locali s 190 153 256 255 6 TE_B
port 2 nsew signal input
rlabel locali s 765 171 811 289 6 Z
port 3 nsew signal output
rlabel locali s 659 353 725 425 6 Z
port 3 nsew signal output
rlabel locali s 659 127 811 171 6 Z
port 3 nsew signal output
rlabel locali s 381 325 725 353 6 Z
port 3 nsew signal output
rlabel locali s 381 289 811 325 6 Z
port 3 nsew signal output
rlabel locali s 468 17 534 97 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 103 17 170 119 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 828 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 828 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 396 455 462 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 103 369 190 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 828 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 828 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2860906
string GDS_START 2853710
<< end >>
