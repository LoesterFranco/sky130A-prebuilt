magic
tech sky130A
magscale 1 2
timestamp 1601050088
<< locali >>
rect 217 291 326 357
rect 476 310 545 430
rect 85 191 410 257
rect 313 162 410 191
rect 647 236 737 310
rect 2130 364 2183 596
rect 2149 226 2183 364
rect 2100 70 2183 226
rect 2409 364 2475 596
rect 2431 210 2475 364
rect 2407 70 2475 210
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2496 683
rect 17 371 106 596
rect 140 460 206 649
rect 314 512 380 596
rect 512 546 630 649
rect 766 546 867 649
rect 997 526 1047 584
rect 901 512 1047 526
rect 314 492 1047 512
rect 1082 492 1153 584
rect 1290 572 1356 649
rect 1187 504 1547 538
rect 314 478 935 492
rect 314 460 380 478
rect 149 391 434 425
rect 149 371 183 391
rect 17 305 183 371
rect 368 359 434 391
rect 17 157 51 305
rect 579 270 613 478
rect 654 398 720 444
rect 654 364 805 398
rect 444 236 613 270
rect 17 70 93 157
rect 127 17 193 146
rect 444 128 478 236
rect 771 202 805 364
rect 839 330 873 478
rect 982 444 1048 456
rect 907 364 1048 444
rect 839 296 980 330
rect 607 168 805 202
rect 291 78 478 128
rect 523 17 573 162
rect 607 70 673 168
rect 719 17 787 134
rect 839 85 889 226
rect 930 119 980 296
rect 1014 85 1048 364
rect 1082 340 1116 492
rect 1187 440 1221 504
rect 1150 374 1221 440
rect 1397 420 1479 470
rect 1338 340 1404 386
rect 1082 306 1404 340
rect 1082 119 1116 306
rect 1438 272 1472 420
rect 1513 392 1547 504
rect 1581 426 1647 596
rect 1772 530 1886 649
rect 1920 470 1990 596
rect 1513 326 1576 392
rect 1613 390 1647 426
rect 1742 424 1990 470
rect 1613 356 1804 390
rect 1920 388 1990 424
rect 1610 284 1736 322
rect 1150 172 1207 272
rect 1249 206 1472 272
rect 1506 271 1736 284
rect 1506 250 1644 271
rect 1770 254 1804 356
rect 1856 254 1922 354
rect 1506 218 1572 250
rect 1770 230 1922 254
rect 1438 184 1472 206
rect 1150 138 1404 172
rect 1150 85 1207 138
rect 839 51 1207 85
rect 1286 17 1336 104
rect 1370 85 1404 138
rect 1438 119 1504 184
rect 1538 85 1572 218
rect 1678 220 1922 230
rect 1956 330 1990 388
rect 2024 364 2090 649
rect 1956 264 2115 330
rect 1678 196 1804 220
rect 1678 162 1712 196
rect 1956 186 1990 264
rect 1370 51 1572 85
rect 1606 70 1712 162
rect 1748 17 1882 162
rect 1918 70 1990 186
rect 2030 17 2064 226
rect 2218 310 2268 575
rect 2308 399 2374 649
rect 2218 244 2397 310
rect 2218 108 2262 244
rect 2298 17 2373 204
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2496 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
<< metal1 >>
rect 0 683 2496 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2496 683
rect 0 617 2496 649
rect 0 17 2496 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2496 17
rect 0 -49 2496 -17
<< labels >>
rlabel locali s 217 291 326 357 6 D
port 1 nsew signal input
rlabel locali s 2149 226 2183 364 6 Q
port 2 nsew signal output
rlabel locali s 2130 364 2183 596 6 Q
port 2 nsew signal output
rlabel locali s 2100 70 2183 226 6 Q
port 2 nsew signal output
rlabel locali s 2431 210 2475 364 6 Q_N
port 3 nsew signal output
rlabel locali s 2409 364 2475 596 6 Q_N
port 3 nsew signal output
rlabel locali s 2407 70 2475 210 6 Q_N
port 3 nsew signal output
rlabel locali s 476 310 545 430 6 SCD
port 4 nsew signal input
rlabel locali s 313 162 410 191 6 SCE
port 5 nsew signal input
rlabel locali s 85 191 410 257 6 SCE
port 5 nsew signal input
rlabel locali s 647 236 737 310 6 CLK
port 6 nsew clock input
rlabel metal1 s 0 -49 2496 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 617 2496 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2496 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 59618
string GDS_START 41090
<< end >>
