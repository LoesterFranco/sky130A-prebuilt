magic
tech sky130A
magscale 1 2
timestamp 1604502710
<< nwell >>
rect -38 332 1574 704
<< pwell >>
rect 0 0 1536 49
<< scpmos >>
rect 161 368 197 536
rect 251 368 287 536
rect 507 368 543 592
rect 597 368 633 592
rect 720 368 756 592
rect 886 368 922 592
rect 1074 368 1110 592
rect 1164 368 1200 592
<< nmoslvt >>
rect 146 82 176 230
rect 267 82 297 230
rect 353 82 383 230
rect 503 82 533 230
rect 603 82 633 230
rect 801 74 831 222
rect 892 74 922 222
rect 978 74 1008 222
rect 1064 74 1094 222
rect 1164 74 1194 222
rect 1250 74 1280 222
rect 1336 74 1366 222
rect 1422 74 1452 222
<< ndiff >>
rect 89 218 146 230
rect 89 184 101 218
rect 135 184 146 218
rect 89 172 146 184
rect 96 82 146 172
rect 176 82 267 230
rect 297 140 353 230
rect 297 106 308 140
rect 342 106 353 140
rect 297 82 353 106
rect 383 84 503 230
rect 383 82 426 84
rect 191 48 204 82
rect 238 48 252 82
rect 191 36 252 48
rect 398 50 426 82
rect 460 82 503 84
rect 533 140 603 230
rect 533 106 544 140
rect 578 106 603 140
rect 533 82 603 106
rect 633 164 683 230
rect 633 140 690 164
rect 633 106 644 140
rect 678 106 690 140
rect 751 138 801 222
rect 633 82 690 106
rect 744 123 801 138
rect 744 89 756 123
rect 790 89 801 123
rect 460 50 488 82
rect 744 74 801 89
rect 831 210 892 222
rect 831 176 844 210
rect 878 176 892 210
rect 831 74 892 176
rect 922 120 978 222
rect 922 86 933 120
rect 967 86 978 120
rect 922 74 978 86
rect 1008 199 1064 222
rect 1008 165 1019 199
rect 1053 165 1064 199
rect 1008 74 1064 165
rect 1094 127 1164 222
rect 1094 93 1119 127
rect 1153 93 1164 127
rect 1094 74 1164 93
rect 1194 202 1250 222
rect 1194 168 1205 202
rect 1239 168 1250 202
rect 1194 74 1250 168
rect 1280 127 1336 222
rect 1280 93 1291 127
rect 1325 93 1336 127
rect 1280 74 1336 93
rect 1366 202 1422 222
rect 1366 168 1377 202
rect 1411 168 1422 202
rect 1366 74 1422 168
rect 1452 146 1502 222
rect 1452 127 1509 146
rect 1452 93 1463 127
rect 1497 93 1509 127
rect 1452 74 1509 93
rect 398 38 488 50
<< pdiff >>
rect 302 580 507 592
rect 302 546 314 580
rect 348 546 388 580
rect 422 546 463 580
rect 497 546 507 580
rect 302 536 507 546
rect 27 516 161 536
rect 27 482 39 516
rect 73 482 161 516
rect 27 368 161 482
rect 197 426 251 536
rect 197 392 207 426
rect 241 392 251 426
rect 197 368 251 392
rect 287 368 507 536
rect 543 426 597 592
rect 543 392 553 426
rect 587 392 597 426
rect 543 368 597 392
rect 633 580 720 592
rect 633 546 659 580
rect 693 546 720 580
rect 633 368 720 546
rect 756 414 886 592
rect 756 380 766 414
rect 800 380 842 414
rect 876 380 886 414
rect 756 368 886 380
rect 922 580 1074 592
rect 922 546 932 580
rect 966 546 1030 580
rect 1064 546 1074 580
rect 922 368 1074 546
rect 1110 421 1164 592
rect 1110 387 1120 421
rect 1154 387 1164 421
rect 1110 368 1164 387
rect 1200 580 1509 592
rect 1200 546 1210 580
rect 1244 546 1294 580
rect 1328 546 1379 580
rect 1413 546 1463 580
rect 1497 546 1509 580
rect 1200 482 1509 546
rect 1200 448 1294 482
rect 1328 448 1379 482
rect 1413 448 1463 482
rect 1497 448 1509 482
rect 1200 368 1509 448
<< ndiffc >>
rect 101 184 135 218
rect 308 106 342 140
rect 204 48 238 82
rect 426 50 460 84
rect 544 106 578 140
rect 644 106 678 140
rect 756 89 790 123
rect 844 176 878 210
rect 933 86 967 120
rect 1019 165 1053 199
rect 1119 93 1153 127
rect 1205 168 1239 202
rect 1291 93 1325 127
rect 1377 168 1411 202
rect 1463 93 1497 127
<< pdiffc >>
rect 314 546 348 580
rect 388 546 422 580
rect 463 546 497 580
rect 39 482 73 516
rect 207 392 241 426
rect 553 392 587 426
rect 659 546 693 580
rect 766 380 800 414
rect 842 380 876 414
rect 932 546 966 580
rect 1030 546 1064 580
rect 1120 387 1154 421
rect 1210 546 1244 580
rect 1294 546 1328 580
rect 1379 546 1413 580
rect 1463 546 1497 580
rect 1294 448 1328 482
rect 1379 448 1413 482
rect 1463 448 1497 482
<< poly >>
rect 507 592 543 618
rect 597 592 633 618
rect 720 592 756 618
rect 886 592 922 618
rect 1074 592 1110 618
rect 1164 592 1200 618
rect 161 536 197 562
rect 251 536 287 562
rect 161 353 197 368
rect 251 353 287 368
rect 85 323 287 353
rect 507 336 543 368
rect 597 336 633 368
rect 85 320 219 323
rect 85 286 101 320
rect 135 286 169 320
rect 203 286 219 320
rect 85 270 219 286
rect 353 320 633 336
rect 353 286 369 320
rect 403 286 437 320
rect 471 286 505 320
rect 539 286 573 320
rect 607 286 633 320
rect 353 275 633 286
rect 146 230 176 270
rect 267 245 633 275
rect 267 230 297 245
rect 353 230 383 245
rect 503 230 533 245
rect 603 230 633 245
rect 720 326 756 368
rect 886 326 922 368
rect 720 310 922 326
rect 1074 345 1110 368
rect 1164 345 1200 368
rect 1074 315 1431 345
rect 720 276 736 310
rect 770 276 804 310
rect 838 276 872 310
rect 906 276 922 310
rect 720 267 922 276
rect 1148 314 1431 315
rect 1148 280 1172 314
rect 1206 280 1240 314
rect 1274 280 1308 314
rect 1342 280 1376 314
rect 1410 294 1431 314
rect 1410 280 1452 294
rect 720 237 1094 267
rect 1148 264 1452 280
rect 146 56 176 82
rect 267 56 297 82
rect 353 56 383 82
rect 801 222 831 237
rect 892 222 922 237
rect 978 222 1008 237
rect 1064 222 1094 237
rect 1164 222 1194 264
rect 1250 222 1280 264
rect 1336 222 1366 264
rect 1422 222 1452 264
rect 503 56 533 82
rect 603 56 633 82
rect 801 48 831 74
rect 892 48 922 74
rect 978 48 1008 74
rect 1064 48 1094 74
rect 1164 48 1194 74
rect 1250 48 1280 74
rect 1336 48 1366 74
rect 1422 48 1452 74
<< polycont >>
rect 101 286 135 320
rect 169 286 203 320
rect 369 286 403 320
rect 437 286 471 320
rect 505 286 539 320
rect 573 286 607 320
rect 736 276 770 310
rect 804 276 838 310
rect 872 276 906 310
rect 1172 280 1206 314
rect 1240 280 1274 314
rect 1308 280 1342 314
rect 1376 280 1410 314
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 23 516 89 649
rect 298 580 513 649
rect 298 546 314 580
rect 348 546 388 580
rect 422 546 463 580
rect 497 546 513 580
rect 298 530 513 546
rect 627 580 726 649
rect 627 546 659 580
rect 693 546 726 580
rect 627 530 726 546
rect 916 580 1080 649
rect 916 546 932 580
rect 966 546 1030 580
rect 1064 546 1080 580
rect 916 530 1080 546
rect 1194 580 1513 649
rect 1194 546 1210 580
rect 1244 546 1294 580
rect 1328 546 1379 580
rect 1413 546 1463 580
rect 1497 546 1513 580
rect 1194 530 1513 546
rect 23 482 39 516
rect 73 482 89 516
rect 23 458 89 482
rect 123 462 1246 496
rect 123 424 157 462
rect 17 390 157 424
rect 191 426 287 428
rect 191 392 207 426
rect 241 392 287 426
rect 191 390 287 392
rect 537 426 1170 428
rect 537 392 553 426
rect 587 421 1170 426
rect 587 414 1120 421
rect 587 392 766 414
rect 537 390 766 392
rect 17 150 51 390
rect 85 320 219 356
rect 85 286 101 320
rect 135 286 169 320
rect 203 286 219 320
rect 85 270 219 286
rect 253 236 287 390
rect 750 380 766 390
rect 800 380 842 414
rect 876 387 1120 414
rect 1154 387 1170 421
rect 876 380 1170 387
rect 750 364 1170 380
rect 1212 398 1246 462
rect 1280 482 1513 530
rect 1280 448 1294 482
rect 1328 448 1379 482
rect 1413 448 1463 482
rect 1497 448 1513 482
rect 1280 432 1513 448
rect 1212 364 1483 398
rect 353 320 647 356
rect 353 286 369 320
rect 403 286 437 320
rect 471 286 505 320
rect 539 286 573 320
rect 607 286 647 320
rect 353 270 647 286
rect 720 310 922 326
rect 720 276 736 310
rect 770 276 804 310
rect 838 276 872 310
rect 906 276 922 310
rect 720 260 922 276
rect 720 236 754 260
rect 85 218 754 236
rect 985 226 1031 364
rect 1164 314 1415 330
rect 1164 280 1172 314
rect 1206 280 1240 314
rect 1274 280 1308 314
rect 1342 280 1376 314
rect 1410 280 1415 314
rect 1164 236 1415 280
rect 85 184 101 218
rect 135 202 754 218
rect 826 210 1069 226
rect 135 184 151 202
rect 826 176 844 210
rect 878 199 1069 210
rect 1449 202 1483 364
rect 878 176 1019 199
rect 292 150 594 168
rect 17 140 594 150
rect 17 116 308 140
rect 292 106 308 116
rect 342 134 544 140
rect 342 106 358 134
rect 187 48 204 82
rect 238 48 256 82
rect 292 78 358 106
rect 528 106 544 134
rect 578 106 594 140
rect 394 84 492 100
rect 187 17 256 48
rect 394 50 426 84
rect 460 50 492 84
rect 528 78 594 106
rect 628 140 694 168
rect 826 165 1019 176
rect 1053 165 1069 199
rect 1189 168 1205 202
rect 1239 168 1377 202
rect 1411 168 1483 202
rect 826 160 1069 165
rect 985 154 1069 160
rect 628 106 644 140
rect 678 106 694 140
rect 1103 127 1513 134
rect 394 17 492 50
rect 628 17 694 106
rect 740 123 806 126
rect 740 89 756 123
rect 790 120 806 123
rect 1103 120 1119 127
rect 790 89 933 120
rect 740 86 933 89
rect 967 93 1119 120
rect 1153 93 1291 127
rect 1325 93 1463 127
rect 1497 93 1513 127
rect 967 86 1513 93
rect 740 70 1513 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
flabel pwell s 0 0 1536 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 1536 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
rlabel comment s 0 0 0 0 4 nand3b_4
flabel metal1 s 0 617 1536 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 1536 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 1183 242 1217 276 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 1279 242 1313 276 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 1375 242 1409 276 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 991 168 1025 202 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 991 242 1025 276 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 Y
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 1536 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 2066032
string GDS_START 2055924
<< end >>
