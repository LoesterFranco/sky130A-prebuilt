magic
tech sky130A
magscale 1 2
timestamp 1599588244
<< locali >>
rect 25 464 424 504
rect 25 326 59 464
rect 25 260 110 326
rect 212 290 278 356
rect 358 290 424 464
rect 793 364 935 434
rect 973 364 1039 434
rect 901 210 935 364
rect 795 176 935 210
rect 977 226 1011 364
rect 977 70 1043 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 23 538 89 649
rect 203 538 280 649
rect 616 536 769 649
rect 883 536 949 649
rect 1063 536 1129 649
rect 113 396 179 430
rect 144 256 178 396
rect 458 468 1111 502
rect 458 322 492 468
rect 526 384 698 434
rect 458 256 607 322
rect 664 310 698 384
rect 144 226 492 256
rect 23 222 492 226
rect 664 244 866 310
rect 664 222 698 244
rect 23 192 178 222
rect 23 70 89 192
rect 527 188 698 222
rect 273 154 493 188
rect 187 17 253 120
rect 359 17 425 120
rect 459 85 493 154
rect 527 119 561 188
rect 1077 326 1111 468
rect 1045 260 1111 326
rect 597 85 663 154
rect 459 51 663 85
rect 709 17 775 142
rect 891 17 941 142
rect 1079 17 1129 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
rlabel locali s 212 290 278 356 6 A
port 1 nsew signal input
rlabel locali s 358 290 424 464 6 B
port 2 nsew signal input
rlabel locali s 25 464 424 504 6 B
port 2 nsew signal input
rlabel locali s 25 326 59 464 6 B
port 2 nsew signal input
rlabel locali s 25 260 110 326 6 B
port 2 nsew signal input
rlabel locali s 977 226 1011 364 6 COUT
port 3 nsew signal output
rlabel locali s 977 70 1043 226 6 COUT
port 3 nsew signal output
rlabel locali s 973 364 1039 434 6 COUT
port 3 nsew signal output
rlabel locali s 901 210 935 364 6 SUM
port 4 nsew signal output
rlabel locali s 795 176 935 210 6 SUM
port 4 nsew signal output
rlabel locali s 793 364 935 434 6 SUM
port 4 nsew signal output
rlabel metal1 s 0 -49 1152 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 6 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 617 1152 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1785718
string GDS_START 1776966
<< end >>
