magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1104 561
rect 180 370 428 421
rect 738 455 804 527
rect 914 455 980 527
rect 25 289 360 336
rect 394 325 428 370
rect 394 289 651 325
rect 25 209 91 289
rect 323 255 360 289
rect 151 215 285 255
rect 323 206 395 255
rect 437 206 571 255
rect 605 169 651 289
rect 693 289 1058 335
rect 693 197 743 289
rect 794 203 945 255
rect 979 199 1058 289
rect 24 161 651 169
rect 24 123 1071 161
rect 24 51 76 123
rect 110 17 176 89
rect 210 51 259 123
rect 293 17 359 89
rect 393 51 459 123
rect 493 17 559 89
rect 593 55 659 123
rect 825 17 891 89
rect 1004 59 1071 123
rect 0 -17 1104 17
<< obsli1 >>
rect 20 459 597 493
rect 20 455 437 459
rect 20 374 92 455
rect 563 427 597 459
rect 631 419 704 493
rect 838 421 880 493
rect 1014 421 1080 493
rect 838 419 1080 421
rect 462 393 528 412
rect 631 393 1080 419
rect 462 369 1080 393
rect 462 359 667 369
<< metal1 >>
rect 0 496 1104 592
rect 0 -48 1104 48
<< labels >>
rlabel locali s 979 199 1058 289 6 A1
port 1 nsew signal input
rlabel locali s 693 289 1058 335 6 A1
port 1 nsew signal input
rlabel locali s 693 197 743 289 6 A1
port 1 nsew signal input
rlabel locali s 794 203 945 255 6 A2
port 2 nsew signal input
rlabel locali s 437 206 571 255 6 B1
port 3 nsew signal input
rlabel locali s 323 255 360 289 6 C1
port 4 nsew signal input
rlabel locali s 323 206 395 255 6 C1
port 4 nsew signal input
rlabel locali s 25 289 360 336 6 C1
port 4 nsew signal input
rlabel locali s 25 209 91 289 6 C1
port 4 nsew signal input
rlabel locali s 151 215 285 255 6 D1
port 5 nsew signal input
rlabel locali s 1004 59 1071 123 6 Y
port 6 nsew signal output
rlabel locali s 605 169 651 289 6 Y
port 6 nsew signal output
rlabel locali s 593 55 659 123 6 Y
port 6 nsew signal output
rlabel locali s 394 325 428 370 6 Y
port 6 nsew signal output
rlabel locali s 394 289 651 325 6 Y
port 6 nsew signal output
rlabel locali s 393 51 459 123 6 Y
port 6 nsew signal output
rlabel locali s 210 51 259 123 6 Y
port 6 nsew signal output
rlabel locali s 180 370 428 421 6 Y
port 6 nsew signal output
rlabel locali s 24 161 651 169 6 Y
port 6 nsew signal output
rlabel locali s 24 123 1071 161 6 Y
port 6 nsew signal output
rlabel locali s 24 51 76 123 6 Y
port 6 nsew signal output
rlabel locali s 825 17 891 89 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 493 17 559 89 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 293 17 359 89 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 110 17 176 89 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 1104 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1104 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 914 455 980 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 738 455 804 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 1104 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 1104 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1104 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3912856
string GDS_START 3904628
<< end >>
