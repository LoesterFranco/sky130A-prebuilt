magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 998 704
rect 375 311 765 332
<< pwell >>
rect 0 0 960 49
<< scnmos >>
rect 88 74 118 222
rect 174 74 204 222
rect 383 74 413 222
rect 461 74 491 222
rect 547 74 577 222
rect 643 74 673 222
rect 763 74 793 222
rect 841 74 871 222
<< pmoshvt >>
rect 90 368 120 592
rect 180 368 210 592
rect 363 368 393 568
rect 464 347 494 547
rect 554 347 584 547
rect 646 347 676 547
rect 760 368 790 568
rect 844 368 874 568
<< ndiff >>
rect 31 210 88 222
rect 31 176 43 210
rect 77 176 88 210
rect 31 120 88 176
rect 31 86 43 120
rect 77 86 88 120
rect 31 74 88 86
rect 118 210 174 222
rect 118 176 129 210
rect 163 176 174 210
rect 118 120 174 176
rect 118 86 129 120
rect 163 86 174 120
rect 118 74 174 86
rect 204 186 383 222
rect 204 152 215 186
rect 249 152 325 186
rect 359 152 383 186
rect 204 118 383 152
rect 204 84 215 118
rect 249 84 325 118
rect 359 84 383 118
rect 204 74 383 84
rect 413 74 461 222
rect 491 199 547 222
rect 491 165 502 199
rect 536 165 547 199
rect 491 120 547 165
rect 491 86 502 120
rect 536 86 547 120
rect 491 74 547 86
rect 577 74 643 222
rect 673 130 763 222
rect 673 96 701 130
rect 735 96 763 130
rect 673 74 763 96
rect 793 74 841 222
rect 871 210 928 222
rect 871 176 882 210
rect 916 176 928 210
rect 871 120 928 176
rect 871 86 882 120
rect 916 86 928 120
rect 871 74 928 86
<< pdiff >>
rect 31 580 90 592
rect 31 546 43 580
rect 77 546 90 580
rect 31 497 90 546
rect 31 463 43 497
rect 77 463 90 497
rect 31 414 90 463
rect 31 380 43 414
rect 77 380 90 414
rect 31 368 90 380
rect 120 580 180 592
rect 120 546 133 580
rect 167 546 180 580
rect 120 497 180 546
rect 120 463 133 497
rect 167 463 180 497
rect 120 414 180 463
rect 120 380 133 414
rect 167 380 180 414
rect 120 368 180 380
rect 210 579 279 592
rect 210 545 224 579
rect 258 568 279 579
rect 258 560 363 568
rect 258 545 315 560
rect 210 526 315 545
rect 349 526 363 560
rect 210 474 363 526
rect 210 440 224 474
rect 258 440 315 474
rect 349 440 363 474
rect 210 368 363 440
rect 393 547 446 568
rect 697 560 760 568
rect 697 547 713 560
rect 393 368 464 547
rect 411 347 464 368
rect 494 535 554 547
rect 494 501 507 535
rect 541 501 554 535
rect 494 440 554 501
rect 494 406 507 440
rect 541 406 554 440
rect 494 347 554 406
rect 584 347 646 547
rect 676 526 713 547
rect 747 526 760 560
rect 676 492 760 526
rect 676 458 713 492
rect 747 458 760 492
rect 676 368 760 458
rect 790 368 844 568
rect 874 556 933 568
rect 874 522 887 556
rect 921 522 933 556
rect 874 485 933 522
rect 874 451 887 485
rect 921 451 933 485
rect 874 414 933 451
rect 874 380 887 414
rect 921 380 933 414
rect 874 368 933 380
rect 676 347 729 368
<< ndiffc >>
rect 43 176 77 210
rect 43 86 77 120
rect 129 176 163 210
rect 129 86 163 120
rect 215 152 249 186
rect 325 152 359 186
rect 215 84 249 118
rect 325 84 359 118
rect 502 165 536 199
rect 502 86 536 120
rect 701 96 735 130
rect 882 176 916 210
rect 882 86 916 120
<< pdiffc >>
rect 43 546 77 580
rect 43 463 77 497
rect 43 380 77 414
rect 133 546 167 580
rect 133 463 167 497
rect 133 380 167 414
rect 224 545 258 579
rect 315 526 349 560
rect 224 440 258 474
rect 315 440 349 474
rect 507 501 541 535
rect 507 406 541 440
rect 713 526 747 560
rect 713 458 747 492
rect 887 522 921 556
rect 887 451 921 485
rect 887 380 921 414
<< poly >>
rect 90 592 120 618
rect 180 592 210 618
rect 360 615 793 645
rect 360 583 396 615
rect 757 583 793 615
rect 363 568 393 583
rect 464 547 494 573
rect 554 547 584 573
rect 646 547 676 573
rect 760 568 790 583
rect 844 568 874 594
rect 90 353 120 368
rect 180 353 210 368
rect 363 353 393 368
rect 87 330 123 353
rect 177 330 213 353
rect 87 314 245 330
rect 87 280 195 314
rect 229 280 245 314
rect 360 310 396 353
rect 760 353 790 368
rect 844 353 874 368
rect 464 332 494 347
rect 554 332 584 347
rect 646 332 676 347
rect 461 315 497 332
rect 551 315 587 332
rect 643 315 679 332
rect 757 323 793 353
rect 87 264 245 280
rect 293 294 413 310
rect 88 222 118 264
rect 174 222 204 264
rect 293 260 309 294
rect 343 260 413 294
rect 293 244 413 260
rect 383 222 413 244
rect 461 299 595 315
rect 461 265 477 299
rect 511 265 545 299
rect 579 265 595 299
rect 461 249 595 265
rect 643 299 709 315
rect 643 265 659 299
rect 693 265 709 299
rect 643 249 709 265
rect 461 222 491 249
rect 547 222 577 249
rect 643 222 673 249
rect 763 222 793 323
rect 841 326 877 353
rect 841 310 907 326
rect 841 276 857 310
rect 891 276 907 310
rect 841 260 907 276
rect 841 222 871 260
rect 88 48 118 74
rect 174 48 204 74
rect 383 48 413 74
rect 461 48 491 74
rect 547 48 577 74
rect 643 48 673 74
rect 763 48 793 74
rect 841 48 871 74
<< polycont >>
rect 195 280 229 314
rect 309 260 343 294
rect 477 265 511 299
rect 545 265 579 299
rect 659 265 693 299
rect 857 276 891 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 27 580 77 649
rect 27 546 43 580
rect 27 497 77 546
rect 27 463 43 497
rect 27 414 77 463
rect 27 380 43 414
rect 27 364 77 380
rect 111 580 183 596
rect 111 546 133 580
rect 167 546 183 580
rect 111 497 183 546
rect 111 463 133 497
rect 167 463 183 497
rect 111 414 183 463
rect 217 579 356 649
rect 217 545 224 579
rect 258 560 356 579
rect 258 545 315 560
rect 217 526 315 545
rect 349 526 356 560
rect 697 560 763 649
rect 217 474 356 526
rect 217 440 224 474
rect 258 440 315 474
rect 349 440 356 474
rect 217 424 356 440
rect 393 535 557 551
rect 393 501 507 535
rect 541 501 557 535
rect 393 440 557 501
rect 697 526 713 560
rect 747 526 763 560
rect 697 492 763 526
rect 697 458 713 492
rect 747 458 763 492
rect 871 556 937 572
rect 871 522 887 556
rect 921 522 937 556
rect 871 485 937 522
rect 111 380 133 414
rect 167 380 183 414
rect 393 406 507 440
rect 541 424 557 440
rect 871 451 887 485
rect 921 451 937 485
rect 871 424 937 451
rect 541 414 937 424
rect 541 406 887 414
rect 393 390 887 406
rect 111 364 183 380
rect 111 226 145 364
rect 217 356 427 390
rect 871 380 887 390
rect 921 380 937 414
rect 871 364 937 380
rect 217 330 251 356
rect 179 314 251 330
rect 179 280 195 314
rect 229 280 251 314
rect 179 264 251 280
rect 293 294 359 310
rect 293 260 309 294
rect 343 260 359 294
rect 293 236 359 260
rect 27 210 77 226
rect 27 176 43 210
rect 27 120 77 176
rect 27 86 43 120
rect 27 17 77 86
rect 111 210 179 226
rect 111 176 129 210
rect 163 176 179 210
rect 393 215 427 356
rect 461 299 595 356
rect 461 265 477 299
rect 511 265 545 299
rect 579 265 595 299
rect 461 249 595 265
rect 643 326 743 356
rect 643 310 907 326
rect 643 299 857 310
rect 643 265 659 299
rect 693 276 857 299
rect 891 276 907 310
rect 693 265 907 276
rect 643 260 907 265
rect 643 249 743 260
rect 866 215 932 226
rect 393 210 932 215
rect 111 120 179 176
rect 111 86 129 120
rect 163 86 179 120
rect 111 70 179 86
rect 215 186 359 202
rect 249 152 325 186
rect 215 118 359 152
rect 249 84 325 118
rect 215 17 359 84
rect 393 199 882 210
rect 393 165 502 199
rect 536 181 882 199
rect 536 165 552 181
rect 393 120 552 165
rect 866 176 882 181
rect 916 176 932 210
rect 393 86 502 120
rect 536 86 552 120
rect 393 70 552 86
rect 668 130 768 136
rect 668 96 701 130
rect 735 96 768 130
rect 668 17 768 96
rect 866 120 932 176
rect 866 86 882 120
rect 916 86 932 120
rect 866 70 932 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
rlabel comment s 0 0 0 0 4 maj3_2
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 127 390 161 424 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 127 464 161 498 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 127 538 161 572 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 319 242 353 276 0 FreeSans 340 0 0 0 A
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 960 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2428082
string GDS_START 2420226
<< end >>
