magic
tech sky130A
magscale 1 2
timestamp 1599588232
<< locali >>
rect 115 236 167 596
rect 115 202 196 236
rect 162 70 196 202
rect 309 252 375 356
rect 409 252 507 356
rect 549 252 647 356
rect 681 290 747 356
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 25 364 75 649
rect 205 458 271 649
rect 309 492 375 596
rect 415 526 473 649
rect 507 492 573 596
rect 309 458 573 492
rect 681 424 747 596
rect 233 390 747 424
rect 233 336 267 390
rect 201 270 267 336
rect 60 17 126 168
rect 233 218 267 270
rect 698 218 748 226
rect 233 184 748 218
rect 232 70 374 150
rect 466 70 540 184
rect 574 70 662 150
rect 698 70 748 184
rect 232 17 266 70
rect 574 17 608 70
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel locali s 409 252 507 356 6 A1
port 1 nsew signal input
rlabel locali s 309 252 375 356 6 A2
port 2 nsew signal input
rlabel locali s 549 252 647 356 6 B1
port 3 nsew signal input
rlabel locali s 681 290 747 356 6 C1
port 4 nsew signal input
rlabel locali s 162 70 196 202 6 X
port 5 nsew signal output
rlabel locali s 115 236 167 596 6 X
port 5 nsew signal output
rlabel locali s 115 202 196 236 6 X
port 5 nsew signal output
rlabel metal1 s 0 -49 768 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 7 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 617 768 715 6 VPWR
port 9 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3982222
string GDS_START 3974818
<< end >>
