magic
tech sky130A
magscale 1 2
timestamp 1599588232
<< locali >>
rect 217 410 505 444
rect 85 270 167 356
rect 217 236 290 410
rect 224 150 290 236
rect 675 270 743 356
rect 1273 290 1415 356
rect 1505 236 1707 310
rect 224 116 555 150
rect 224 70 290 116
rect 428 84 555 116
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 17 512 89 572
rect 130 546 199 649
rect 313 546 398 649
rect 568 546 634 649
rect 967 596 1223 615
rect 787 581 1223 596
rect 787 526 1033 581
rect 17 478 573 512
rect 17 390 89 478
rect 17 226 51 390
rect 539 376 573 478
rect 17 90 89 226
rect 123 17 183 226
rect 324 342 573 376
rect 607 458 943 492
rect 324 218 358 342
rect 607 308 641 458
rect 675 390 811 424
rect 392 252 641 308
rect 777 318 811 390
rect 877 386 943 458
rect 1067 454 1133 547
rect 1173 488 1223 581
rect 1269 581 1515 615
rect 1269 488 1335 581
rect 1375 454 1409 547
rect 1067 420 1409 454
rect 1315 390 1409 420
rect 1449 448 1515 581
rect 1549 482 1615 649
rect 1650 448 1705 598
rect 1449 390 1705 448
rect 1639 388 1705 390
rect 877 352 1229 386
rect 777 284 1161 318
rect 889 252 1161 284
rect 1195 252 1229 352
rect 789 218 855 250
rect 324 184 855 218
rect 889 150 923 252
rect 1195 218 1471 252
rect 326 17 392 82
rect 589 17 655 150
rect 691 116 923 150
rect 691 90 757 116
rect 803 17 921 82
rect 957 70 1256 218
rect 1290 17 1356 184
rect 1405 70 1471 218
rect 1528 17 1662 197
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
<< metal1 >>
rect 0 683 1728 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 0 617 1728 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 1728 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
rect 0 -49 1728 -17
<< labels >>
rlabel locali s 1505 236 1707 310 6 A
port 1 nsew signal input
rlabel locali s 1273 290 1415 356 6 B
port 2 nsew signal input
rlabel locali s 675 270 743 356 6 C_N
port 3 nsew signal input
rlabel locali s 85 270 167 356 6 D_N
port 4 nsew signal input
rlabel locali s 428 84 555 116 6 X
port 5 nsew signal output
rlabel locali s 224 150 290 236 6 X
port 5 nsew signal output
rlabel locali s 224 116 555 150 6 X
port 5 nsew signal output
rlabel locali s 224 70 290 116 6 X
port 5 nsew signal output
rlabel locali s 217 410 505 444 6 X
port 5 nsew signal output
rlabel locali s 217 236 290 410 6 X
port 5 nsew signal output
rlabel metal1 s 0 -49 1728 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 7 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 617 1728 715 6 VPWR
port 9 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1728 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 940304
string GDS_START 927488
<< end >>
