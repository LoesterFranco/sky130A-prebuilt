magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1840 561
rect 19 365 78 527
rect 198 365 250 527
rect 370 526 1625 527
rect 370 367 422 526
rect 456 347 508 492
rect 542 381 594 526
rect 628 347 680 492
rect 714 381 766 526
rect 800 347 852 492
rect 886 381 938 526
rect 972 347 1024 492
rect 1058 381 1107 526
rect 1141 347 1193 492
rect 1230 381 1279 526
rect 1313 347 1365 492
rect 1402 381 1451 526
rect 1485 347 1537 492
rect 1574 381 1625 526
rect 456 344 1537 347
rect 1659 344 1717 492
rect 1751 378 1805 527
rect 456 299 1805 344
rect 17 153 80 265
rect 17 17 78 119
rect 198 17 250 122
rect 1572 181 1805 299
rect 456 147 1805 181
rect 370 17 422 129
rect 456 56 508 147
rect 542 17 594 113
rect 628 56 680 147
rect 714 17 766 113
rect 800 56 852 147
rect 886 17 935 113
rect 969 56 1024 147
rect 1058 17 1107 113
rect 1141 56 1193 147
rect 1229 17 1279 113
rect 1313 56 1365 147
rect 1401 17 1451 113
rect 1485 56 1537 147
rect 1573 17 1625 113
rect 1659 56 1711 147
rect 1745 17 1805 113
rect 0 -17 1840 17
<< obsli1 >>
rect 114 265 163 493
rect 286 265 336 492
rect 114 215 1538 265
rect 114 53 164 215
rect 286 53 336 215
<< metal1 >>
rect 0 496 1840 592
rect 0 -48 1840 48
<< labels >>
rlabel locali s 17 153 80 265 6 A
port 1 nsew signal input
rlabel locali s 1659 344 1717 492 6 X
port 2 nsew signal output
rlabel locali s 1659 56 1711 147 6 X
port 2 nsew signal output
rlabel locali s 1572 181 1805 299 6 X
port 2 nsew signal output
rlabel locali s 1485 347 1537 492 6 X
port 2 nsew signal output
rlabel locali s 1485 56 1537 147 6 X
port 2 nsew signal output
rlabel locali s 1313 347 1365 492 6 X
port 2 nsew signal output
rlabel locali s 1313 56 1365 147 6 X
port 2 nsew signal output
rlabel locali s 1141 347 1193 492 6 X
port 2 nsew signal output
rlabel locali s 1141 56 1193 147 6 X
port 2 nsew signal output
rlabel locali s 972 347 1024 492 6 X
port 2 nsew signal output
rlabel locali s 969 56 1024 147 6 X
port 2 nsew signal output
rlabel locali s 800 347 852 492 6 X
port 2 nsew signal output
rlabel locali s 800 56 852 147 6 X
port 2 nsew signal output
rlabel locali s 628 347 680 492 6 X
port 2 nsew signal output
rlabel locali s 628 56 680 147 6 X
port 2 nsew signal output
rlabel locali s 456 347 508 492 6 X
port 2 nsew signal output
rlabel locali s 456 344 1537 347 6 X
port 2 nsew signal output
rlabel locali s 456 299 1805 344 6 X
port 2 nsew signal output
rlabel locali s 456 147 1805 181 6 X
port 2 nsew signal output
rlabel locali s 456 56 508 147 6 X
port 2 nsew signal output
rlabel locali s 1745 17 1805 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1573 17 1625 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1401 17 1451 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1229 17 1279 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1058 17 1107 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 886 17 935 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 714 17 766 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 542 17 594 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 370 17 422 129 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 198 17 250 122 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 17 17 78 119 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 0 -17 1840 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1840 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1751 378 1805 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1574 381 1625 526 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1402 381 1451 526 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1230 381 1279 526 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1058 381 1107 526 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 886 381 938 526 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 714 381 766 526 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 542 381 594 526 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 370 526 1625 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 370 367 422 526 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 198 365 250 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 19 365 78 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 0 527 1840 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 496 1840 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1840 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3185428
string GDS_START 3172756
<< end >>
