magic
tech sky130A
magscale 1 2
timestamp 1599588218
<< nwell >>
rect -38 332 806 704
<< pwell >>
rect 0 0 768 49
<< scpmos >>
rect 83 368 119 592
rect 209 413 245 581
rect 309 413 345 581
rect 460 413 496 581
rect 567 381 603 581
rect 651 381 687 581
<< nmoslvt >>
rect 82 74 112 222
rect 291 74 321 222
rect 363 74 393 222
rect 441 74 471 222
rect 543 74 573 222
rect 651 74 681 222
<< ndiff >>
rect 27 192 82 222
rect 27 158 37 192
rect 71 158 82 192
rect 27 120 82 158
rect 27 86 37 120
rect 71 86 82 120
rect 27 74 82 86
rect 112 192 167 222
rect 112 158 123 192
rect 157 158 167 192
rect 112 120 167 158
rect 112 86 123 120
rect 157 86 167 120
rect 112 74 167 86
rect 221 210 291 222
rect 221 176 232 210
rect 266 176 291 210
rect 221 120 291 176
rect 221 86 232 120
rect 266 86 291 120
rect 221 74 291 86
rect 321 74 363 222
rect 393 74 441 222
rect 471 210 543 222
rect 471 176 492 210
rect 526 176 543 210
rect 471 120 543 176
rect 471 86 492 120
rect 526 86 543 120
rect 471 74 543 86
rect 573 131 651 222
rect 573 97 592 131
rect 626 97 651 131
rect 573 74 651 97
rect 681 210 738 222
rect 681 176 692 210
rect 726 176 738 210
rect 681 120 738 176
rect 681 86 692 120
rect 726 86 738 120
rect 681 74 738 86
<< pdiff >>
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 497 83 546
rect 27 463 39 497
rect 73 463 83 497
rect 27 414 83 463
rect 27 380 39 414
rect 73 380 83 414
rect 27 368 83 380
rect 119 584 190 592
rect 119 550 139 584
rect 173 581 190 584
rect 173 550 209 581
rect 119 516 209 550
rect 119 482 139 516
rect 173 482 209 516
rect 119 413 209 482
rect 245 569 309 581
rect 245 535 255 569
rect 289 535 309 569
rect 245 465 309 535
rect 245 431 255 465
rect 289 431 309 465
rect 245 413 309 431
rect 345 541 460 581
rect 345 507 386 541
rect 420 507 460 541
rect 345 413 460 507
rect 496 569 567 581
rect 496 535 523 569
rect 557 535 567 569
rect 496 459 567 535
rect 496 425 523 459
rect 557 425 567 459
rect 496 413 567 425
rect 119 368 169 413
rect 511 381 567 413
rect 603 381 651 581
rect 687 569 741 581
rect 687 535 697 569
rect 731 535 741 569
rect 687 501 741 535
rect 687 467 697 501
rect 731 467 741 501
rect 687 433 741 467
rect 687 399 697 433
rect 731 399 741 433
rect 687 381 741 399
<< ndiffc >>
rect 37 158 71 192
rect 37 86 71 120
rect 123 158 157 192
rect 123 86 157 120
rect 232 176 266 210
rect 232 86 266 120
rect 492 176 526 210
rect 492 86 526 120
rect 592 97 626 131
rect 692 176 726 210
rect 692 86 726 120
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 139 550 173 584
rect 139 482 173 516
rect 255 535 289 569
rect 255 431 289 465
rect 386 507 420 541
rect 523 535 557 569
rect 523 425 557 459
rect 697 535 731 569
rect 697 467 731 501
rect 697 399 731 433
<< poly >>
rect 83 592 119 618
rect 209 581 245 607
rect 309 581 345 607
rect 460 581 496 607
rect 567 581 603 607
rect 651 581 687 607
rect 209 376 245 413
rect 309 380 345 413
rect 83 310 119 368
rect 201 360 267 376
rect 201 326 217 360
rect 251 326 267 360
rect 201 310 267 326
rect 309 364 393 380
rect 309 330 325 364
rect 359 330 393 364
rect 460 349 496 413
rect 567 349 603 381
rect 309 314 393 330
rect 82 294 153 310
rect 82 260 103 294
rect 137 260 153 294
rect 82 244 153 260
rect 237 267 267 310
rect 82 222 112 244
rect 237 237 321 267
rect 291 222 321 237
rect 363 222 393 314
rect 435 333 501 349
rect 435 299 451 333
rect 485 299 501 333
rect 435 283 501 299
rect 543 333 609 349
rect 543 299 559 333
rect 593 299 609 333
rect 543 283 609 299
rect 651 326 687 381
rect 651 310 747 326
rect 441 222 471 283
rect 543 222 573 283
rect 651 276 697 310
rect 731 276 747 310
rect 651 260 747 276
rect 651 222 681 260
rect 82 48 112 74
rect 291 48 321 74
rect 363 48 393 74
rect 441 48 471 74
rect 543 48 573 74
rect 651 48 681 74
<< polycont >>
rect 217 326 251 360
rect 325 330 359 364
rect 103 260 137 294
rect 451 299 485 333
rect 559 299 593 333
rect 697 276 731 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 19 580 89 596
rect 19 546 39 580
rect 73 546 89 580
rect 19 497 89 546
rect 19 463 39 497
rect 73 463 89 497
rect 123 584 189 649
rect 123 550 139 584
rect 173 550 189 584
rect 123 516 189 550
rect 123 482 139 516
rect 173 482 189 516
rect 239 569 305 585
rect 239 535 255 569
rect 289 535 305 569
rect 19 414 89 463
rect 239 465 305 535
rect 348 541 458 649
rect 348 507 386 541
rect 420 507 458 541
rect 348 491 458 507
rect 507 569 573 585
rect 507 535 523 569
rect 557 535 573 569
rect 239 448 255 465
rect 19 380 39 414
rect 73 380 89 414
rect 19 364 89 380
rect 123 431 255 448
rect 289 449 305 465
rect 507 459 573 535
rect 507 449 523 459
rect 289 431 523 449
rect 123 425 523 431
rect 557 425 573 459
rect 123 414 573 425
rect 19 208 53 364
rect 123 310 157 414
rect 507 409 573 414
rect 681 569 747 649
rect 681 535 697 569
rect 731 535 747 569
rect 681 501 747 535
rect 681 467 697 501
rect 731 467 747 501
rect 681 433 747 467
rect 681 399 697 433
rect 731 399 747 433
rect 681 390 747 399
rect 201 360 267 376
rect 201 326 217 360
rect 251 326 267 360
rect 201 310 267 326
rect 309 364 375 380
rect 309 330 325 364
rect 359 330 375 364
rect 87 294 157 310
rect 87 260 103 294
rect 137 276 157 294
rect 137 260 266 276
rect 87 242 266 260
rect 216 210 266 242
rect 19 192 71 208
rect 19 158 37 192
rect 19 120 71 158
rect 19 86 37 120
rect 19 70 71 86
rect 107 192 173 208
rect 107 158 123 192
rect 157 158 173 192
rect 107 120 173 158
rect 107 86 123 120
rect 157 86 173 120
rect 107 17 173 86
rect 216 176 232 210
rect 216 120 266 176
rect 216 86 232 120
rect 309 88 375 330
rect 409 333 501 356
rect 409 299 451 333
rect 485 299 501 333
rect 409 283 501 299
rect 543 333 647 356
rect 543 299 559 333
rect 593 299 647 333
rect 543 283 647 299
rect 681 310 747 356
rect 681 276 697 310
rect 731 276 747 310
rect 681 260 747 276
rect 476 210 742 226
rect 476 176 492 210
rect 526 192 692 210
rect 526 176 542 192
rect 476 120 542 176
rect 676 176 692 192
rect 726 176 742 210
rect 216 70 266 86
rect 476 86 492 120
rect 526 86 542 120
rect 476 70 542 86
rect 576 131 642 158
rect 576 97 592 131
rect 626 97 642 131
rect 576 17 642 97
rect 676 120 742 176
rect 676 86 692 120
rect 726 86 742 120
rect 676 70 742 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
rlabel comment s 0 0 0 0 4 o2111a_1
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 319 94 353 128 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 319 168 353 202 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 319 242 353 276 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 D1
port 5 nsew
flabel corelocali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 10 nsew
flabel corelocali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 10 nsew
flabel corelocali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 768 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1667120
string GDS_START 1659512
<< end >>
