magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 2534 704
<< pwell >>
rect 0 0 2496 49
<< scnmos >>
rect 88 74 118 158
rect 188 74 218 158
rect 266 74 296 158
rect 404 74 434 158
rect 482 74 512 158
rect 582 74 612 222
rect 798 74 828 222
rect 991 100 1021 184
rect 1127 100 1157 184
rect 1249 100 1279 184
rect 1412 74 1442 184
rect 1499 74 1529 184
rect 1651 74 1681 158
rect 1723 74 1753 158
rect 1877 74 1907 184
rect 2075 74 2105 222
rect 2273 112 2303 222
rect 2382 74 2412 222
<< pmoshvt >>
rect 103 464 133 592
rect 203 464 233 592
rect 287 464 317 592
rect 377 464 407 592
rect 485 464 515 592
rect 627 368 657 592
rect 864 368 894 592
rect 1060 496 1090 580
rect 1150 496 1180 580
rect 1246 496 1276 580
rect 1370 424 1400 592
rect 1554 424 1584 592
rect 1661 508 1691 592
rect 1745 508 1775 592
rect 1893 392 1923 592
rect 2087 368 2117 592
rect 2281 403 2311 571
rect 2382 368 2412 592
<< ndiff >>
rect 532 158 582 222
rect 31 130 88 158
rect 31 96 43 130
rect 77 96 88 130
rect 31 74 88 96
rect 118 133 188 158
rect 118 99 143 133
rect 177 99 188 133
rect 118 74 188 99
rect 218 74 266 158
rect 296 128 404 158
rect 296 94 333 128
rect 367 94 404 128
rect 296 74 404 94
rect 434 74 482 158
rect 512 133 582 158
rect 512 99 531 133
rect 565 99 582 133
rect 512 74 582 99
rect 612 202 669 222
rect 612 168 623 202
rect 657 168 669 202
rect 612 120 669 168
rect 612 86 623 120
rect 657 86 669 120
rect 612 74 669 86
rect 723 118 798 222
rect 723 84 736 118
rect 770 84 798 118
rect 723 74 798 84
rect 828 210 882 222
rect 828 176 839 210
rect 873 176 882 210
rect 828 120 882 176
rect 828 86 839 120
rect 873 86 882 120
rect 936 170 991 184
rect 936 136 946 170
rect 980 136 991 170
rect 936 100 991 136
rect 1021 170 1127 184
rect 1021 136 1082 170
rect 1116 136 1127 170
rect 1021 100 1127 136
rect 1157 100 1249 184
rect 1279 100 1412 184
rect 828 74 882 86
rect 1294 88 1412 100
rect 723 72 783 74
rect 1294 54 1302 88
rect 1336 74 1412 88
rect 1442 160 1499 184
rect 1442 126 1454 160
rect 1488 126 1499 160
rect 1442 74 1499 126
rect 1529 158 1579 184
rect 2018 210 2075 222
rect 1820 158 1877 184
rect 1529 133 1651 158
rect 1529 99 1606 133
rect 1640 99 1651 133
rect 1529 74 1651 99
rect 1681 74 1723 158
rect 1753 133 1877 158
rect 1753 99 1764 133
rect 1798 99 1832 133
rect 1866 99 1877 133
rect 1753 74 1877 99
rect 1907 145 1964 184
rect 1907 111 1918 145
rect 1952 111 1964 145
rect 1907 74 1964 111
rect 2018 176 2030 210
rect 2064 176 2075 210
rect 2018 120 2075 176
rect 2018 86 2030 120
rect 2064 86 2075 120
rect 2018 74 2075 86
rect 2105 210 2162 222
rect 2105 176 2116 210
rect 2150 176 2162 210
rect 2105 120 2162 176
rect 2105 86 2116 120
rect 2150 86 2162 120
rect 2216 184 2273 222
rect 2216 150 2228 184
rect 2262 150 2273 184
rect 2216 112 2273 150
rect 2303 200 2382 222
rect 2303 166 2318 200
rect 2352 166 2382 200
rect 2303 120 2382 166
rect 2303 112 2333 120
rect 2318 86 2333 112
rect 2367 86 2382 120
rect 2105 74 2162 86
rect 2318 74 2382 86
rect 2412 194 2469 222
rect 2412 160 2423 194
rect 2457 160 2469 194
rect 2412 120 2469 160
rect 2412 86 2423 120
rect 2457 86 2469 120
rect 2412 74 2469 86
rect 1336 54 1348 74
rect 1294 42 1348 54
<< pdiff >>
rect 1294 622 1352 634
rect 44 580 103 592
rect 44 546 56 580
rect 90 546 103 580
rect 44 510 103 546
rect 44 476 56 510
rect 90 476 103 510
rect 44 464 103 476
rect 133 580 203 592
rect 133 546 156 580
rect 190 546 203 580
rect 133 510 203 546
rect 133 476 156 510
rect 190 476 203 510
rect 133 464 203 476
rect 233 464 287 592
rect 317 580 377 592
rect 317 546 330 580
rect 364 546 377 580
rect 317 510 377 546
rect 317 476 330 510
rect 364 476 377 510
rect 317 464 377 476
rect 407 464 485 592
rect 515 580 627 592
rect 515 546 554 580
rect 588 546 627 580
rect 515 464 627 546
rect 574 368 627 464
rect 657 421 716 592
rect 657 387 670 421
rect 704 387 716 421
rect 657 368 716 387
rect 770 580 864 592
rect 770 546 799 580
rect 833 546 864 580
rect 770 368 864 546
rect 894 421 950 592
rect 1294 588 1306 622
rect 1340 592 1352 622
rect 1340 588 1370 592
rect 1294 580 1370 588
rect 1004 555 1060 580
rect 1004 521 1013 555
rect 1047 521 1060 555
rect 1004 496 1060 521
rect 1090 555 1150 580
rect 1090 521 1103 555
rect 1137 521 1150 555
rect 1090 496 1150 521
rect 1180 496 1246 580
rect 1276 496 1370 580
rect 894 387 907 421
rect 941 387 950 421
rect 894 368 950 387
rect 1317 424 1370 496
rect 1400 470 1554 592
rect 1400 436 1421 470
rect 1455 436 1554 470
rect 1400 424 1554 436
rect 1584 580 1661 592
rect 1584 546 1597 580
rect 1631 546 1661 580
rect 1584 508 1661 546
rect 1691 508 1745 592
rect 1775 580 1893 592
rect 1775 546 1815 580
rect 1849 546 1893 580
rect 1775 508 1893 546
rect 1584 476 1643 508
rect 1584 442 1597 476
rect 1631 442 1643 476
rect 1584 424 1643 442
rect 1840 392 1893 508
rect 1923 580 1978 592
rect 1923 546 1936 580
rect 1970 546 1978 580
rect 1923 509 1978 546
rect 1923 475 1936 509
rect 1970 475 1978 509
rect 1923 438 1978 475
rect 1923 404 1936 438
rect 1970 404 1978 438
rect 1923 392 1978 404
rect 2032 580 2087 592
rect 2032 546 2040 580
rect 2074 546 2087 580
rect 2032 497 2087 546
rect 2032 463 2040 497
rect 2074 463 2087 497
rect 2032 414 2087 463
rect 2032 380 2040 414
rect 2074 380 2087 414
rect 2032 368 2087 380
rect 2117 580 2172 592
rect 2117 546 2130 580
rect 2164 546 2172 580
rect 2329 571 2382 592
rect 2117 497 2172 546
rect 2117 463 2130 497
rect 2164 463 2172 497
rect 2117 414 2172 463
rect 2117 380 2130 414
rect 2164 380 2172 414
rect 2226 559 2281 571
rect 2226 525 2234 559
rect 2268 525 2281 559
rect 2226 449 2281 525
rect 2226 415 2234 449
rect 2268 415 2281 449
rect 2226 403 2281 415
rect 2311 559 2382 571
rect 2311 525 2324 559
rect 2358 525 2382 559
rect 2311 449 2382 525
rect 2311 415 2324 449
rect 2358 415 2382 449
rect 2311 403 2382 415
rect 2117 368 2172 380
rect 2329 368 2382 403
rect 2412 580 2469 592
rect 2412 546 2425 580
rect 2459 546 2469 580
rect 2412 497 2469 546
rect 2412 463 2425 497
rect 2459 463 2469 497
rect 2412 414 2469 463
rect 2412 380 2425 414
rect 2459 380 2469 414
rect 2412 368 2469 380
<< ndiffc >>
rect 43 96 77 130
rect 143 99 177 133
rect 333 94 367 128
rect 531 99 565 133
rect 623 168 657 202
rect 623 86 657 120
rect 736 84 770 118
rect 839 176 873 210
rect 839 86 873 120
rect 946 136 980 170
rect 1082 136 1116 170
rect 1302 54 1336 88
rect 1454 126 1488 160
rect 1606 99 1640 133
rect 1764 99 1798 133
rect 1832 99 1866 133
rect 1918 111 1952 145
rect 2030 176 2064 210
rect 2030 86 2064 120
rect 2116 176 2150 210
rect 2116 86 2150 120
rect 2228 150 2262 184
rect 2318 166 2352 200
rect 2333 86 2367 120
rect 2423 160 2457 194
rect 2423 86 2457 120
<< pdiffc >>
rect 56 546 90 580
rect 56 476 90 510
rect 156 546 190 580
rect 156 476 190 510
rect 330 546 364 580
rect 330 476 364 510
rect 554 546 588 580
rect 670 387 704 421
rect 799 546 833 580
rect 1306 588 1340 622
rect 1013 521 1047 555
rect 1103 521 1137 555
rect 907 387 941 421
rect 1421 436 1455 470
rect 1597 546 1631 580
rect 1815 546 1849 580
rect 1597 442 1631 476
rect 1936 546 1970 580
rect 1936 475 1970 509
rect 1936 404 1970 438
rect 2040 546 2074 580
rect 2040 463 2074 497
rect 2040 380 2074 414
rect 2130 546 2164 580
rect 2130 463 2164 497
rect 2130 380 2164 414
rect 2234 525 2268 559
rect 2234 415 2268 449
rect 2324 525 2358 559
rect 2324 415 2358 449
rect 2425 546 2459 580
rect 2425 463 2459 497
rect 2425 380 2459 414
<< poly >>
rect 103 592 133 618
rect 203 592 233 618
rect 287 592 317 618
rect 377 592 407 618
rect 485 592 515 618
rect 627 592 657 618
rect 864 592 894 618
rect 103 449 133 464
rect 203 449 233 464
rect 287 449 317 464
rect 377 449 407 464
rect 485 449 515 464
rect 39 419 236 449
rect 39 257 69 419
rect 117 355 218 371
rect 284 357 320 449
rect 374 425 410 449
rect 368 409 434 425
rect 368 375 384 409
rect 418 375 434 409
rect 482 388 518 449
rect 368 359 434 375
rect 476 372 542 388
rect 117 321 133 355
rect 167 321 218 355
rect 117 305 218 321
rect 39 241 146 257
rect 39 227 96 241
rect 80 207 96 227
rect 130 207 146 241
rect 80 191 146 207
rect 88 158 118 191
rect 188 158 218 305
rect 260 341 326 357
rect 260 307 276 341
rect 310 307 326 341
rect 476 338 492 372
rect 526 338 542 372
rect 1060 580 1090 606
rect 1150 580 1180 606
rect 1246 580 1276 606
rect 1370 592 1400 618
rect 1554 592 1584 618
rect 1661 592 1691 618
rect 1745 592 1775 618
rect 1893 592 1923 618
rect 2087 592 2117 618
rect 1060 481 1090 496
rect 1150 481 1180 496
rect 1246 481 1276 496
rect 1057 464 1093 481
rect 982 448 1093 464
rect 982 414 998 448
rect 1032 434 1093 448
rect 1147 440 1183 481
rect 1032 414 1048 434
rect 982 398 1048 414
rect 1135 424 1201 440
rect 1135 390 1151 424
rect 1185 390 1201 424
rect 1243 398 1279 481
rect 1661 493 1691 508
rect 1745 493 1775 508
rect 1658 434 1694 493
rect 1742 476 1778 493
rect 1742 460 1808 476
rect 1370 409 1400 424
rect 1554 409 1584 424
rect 627 353 657 368
rect 864 353 894 368
rect 476 322 542 338
rect 260 291 326 307
rect 266 158 296 291
rect 344 230 434 246
rect 344 196 360 230
rect 394 196 434 230
rect 344 180 434 196
rect 404 158 434 180
rect 482 158 512 322
rect 624 310 660 353
rect 861 350 897 353
rect 1135 350 1201 390
rect 755 320 1201 350
rect 624 294 713 310
rect 624 274 663 294
rect 582 260 663 274
rect 697 260 713 294
rect 755 286 771 320
rect 805 286 828 320
rect 755 270 828 286
rect 582 244 713 260
rect 582 222 612 244
rect 798 222 828 270
rect 991 184 1021 320
rect 1249 272 1279 398
rect 1367 386 1403 409
rect 1551 392 1587 409
rect 1658 404 1700 434
rect 1742 426 1758 460
rect 1792 426 1808 460
rect 1742 410 1808 426
rect 1338 370 1442 386
rect 1338 336 1354 370
rect 1388 336 1442 370
rect 1338 320 1442 336
rect 1511 376 1587 392
rect 1511 342 1527 376
rect 1561 356 1587 376
rect 1561 342 1628 356
rect 1511 326 1628 342
rect 1127 256 1207 272
rect 1127 222 1157 256
rect 1191 222 1207 256
rect 1127 206 1207 222
rect 1249 256 1315 272
rect 1249 222 1265 256
rect 1299 222 1315 256
rect 1249 206 1315 222
rect 1127 184 1157 206
rect 1249 184 1279 206
rect 1412 184 1442 320
rect 1490 268 1556 284
rect 1490 234 1506 268
rect 1540 234 1556 268
rect 1490 218 1556 234
rect 1598 223 1628 326
rect 1670 337 1700 404
rect 1670 321 1736 337
rect 1670 287 1686 321
rect 1720 287 1736 321
rect 1670 271 1736 287
rect 1778 229 1808 410
rect 1893 377 1923 392
rect 1890 354 1926 377
rect 2281 571 2311 597
rect 2382 592 2412 618
rect 2281 388 2311 403
rect 1499 184 1529 218
rect 1598 193 1681 223
rect 991 74 1021 100
rect 1127 74 1157 100
rect 1249 74 1279 100
rect 88 48 118 74
rect 188 48 218 74
rect 266 48 296 74
rect 404 48 434 74
rect 482 48 512 74
rect 582 48 612 74
rect 798 48 828 74
rect 1651 158 1681 193
rect 1723 199 1808 229
rect 1856 338 1926 354
rect 2087 353 2117 368
rect 2273 358 2314 388
rect 1856 304 1872 338
rect 1906 304 1926 338
rect 2084 330 2120 353
rect 1856 270 1926 304
rect 1856 236 1872 270
rect 1906 236 1926 270
rect 1981 318 2120 330
rect 2273 318 2303 358
rect 2382 353 2412 368
rect 1981 314 2303 318
rect 1981 280 1997 314
rect 2031 280 2065 314
rect 2099 280 2303 314
rect 2379 310 2415 353
rect 1981 264 2303 280
rect 1856 220 1926 236
rect 2075 222 2105 264
rect 2273 222 2303 264
rect 2345 294 2412 310
rect 2345 260 2361 294
rect 2395 260 2412 294
rect 2345 244 2412 260
rect 2382 222 2412 244
rect 1723 158 1753 199
rect 1877 184 1907 220
rect 2273 86 2303 112
rect 1412 48 1442 74
rect 1499 48 1529 74
rect 1651 48 1681 74
rect 1723 48 1753 74
rect 1877 48 1907 74
rect 2075 48 2105 74
rect 2382 48 2412 74
<< polycont >>
rect 384 375 418 409
rect 133 321 167 355
rect 96 207 130 241
rect 276 307 310 341
rect 492 338 526 372
rect 998 414 1032 448
rect 1151 390 1185 424
rect 360 196 394 230
rect 663 260 697 294
rect 771 286 805 320
rect 1758 426 1792 460
rect 1354 336 1388 370
rect 1527 342 1561 376
rect 1157 222 1191 256
rect 1265 222 1299 256
rect 1506 234 1540 268
rect 1686 287 1720 321
rect 1872 304 1906 338
rect 1872 236 1906 270
rect 1997 280 2031 314
rect 2065 280 2099 314
rect 2361 260 2395 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2496 683
rect 17 580 106 596
rect 17 546 56 580
rect 90 546 106 580
rect 17 510 106 546
rect 17 476 56 510
rect 90 476 106 510
rect 17 371 106 476
rect 140 580 206 649
rect 140 546 156 580
rect 190 546 206 580
rect 140 510 206 546
rect 140 476 156 510
rect 190 476 206 510
rect 140 460 206 476
rect 314 580 380 596
rect 314 546 330 580
rect 364 546 380 580
rect 512 580 630 649
rect 512 546 554 580
rect 588 546 630 580
rect 766 580 867 649
rect 1290 622 1356 649
rect 1290 588 1306 622
rect 1340 588 1356 622
rect 766 546 799 580
rect 833 546 867 580
rect 997 555 1047 584
rect 314 512 380 546
rect 997 526 1013 555
rect 901 521 1013 526
rect 901 512 1047 521
rect 314 510 1047 512
rect 314 476 330 510
rect 364 492 1047 510
rect 1082 555 1153 584
rect 1290 572 1356 588
rect 1581 580 1647 596
rect 1082 521 1103 555
rect 1137 521 1153 555
rect 1581 546 1597 580
rect 1631 546 1647 580
rect 1082 492 1153 521
rect 1187 504 1547 538
rect 364 478 935 492
rect 364 476 380 478
rect 314 460 380 476
rect 149 409 434 425
rect 149 391 384 409
rect 149 371 183 391
rect 17 355 183 371
rect 368 375 384 391
rect 418 375 434 409
rect 368 359 434 375
rect 476 372 545 430
rect 17 321 133 355
rect 167 321 183 355
rect 17 305 183 321
rect 217 341 326 357
rect 217 307 276 341
rect 310 307 326 341
rect 476 338 492 372
rect 526 338 545 372
rect 476 310 545 338
rect 17 157 51 305
rect 217 291 326 307
rect 579 270 613 478
rect 654 421 720 444
rect 654 387 670 421
rect 704 398 720 421
rect 704 387 805 398
rect 654 364 805 387
rect 771 320 805 364
rect 85 241 410 257
rect 85 207 96 241
rect 130 230 410 241
rect 130 207 360 230
rect 85 196 360 207
rect 394 196 410 230
rect 85 191 410 196
rect 313 162 410 191
rect 444 236 613 270
rect 647 294 737 310
rect 647 260 663 294
rect 697 260 737 294
rect 647 236 737 260
rect 839 330 873 478
rect 982 448 1048 456
rect 982 444 998 448
rect 907 421 998 444
rect 941 414 998 421
rect 1032 414 1048 448
rect 941 387 1048 414
rect 907 364 1048 387
rect 839 296 980 330
rect 17 130 93 157
rect 17 96 43 130
rect 77 96 93 130
rect 17 70 93 96
rect 127 133 193 146
rect 127 99 143 133
rect 177 99 193 133
rect 444 128 478 236
rect 771 202 805 286
rect 607 168 623 202
rect 657 168 805 202
rect 839 210 889 226
rect 873 176 889 210
rect 127 17 193 99
rect 291 94 333 128
rect 367 94 478 128
rect 291 78 478 94
rect 523 133 573 162
rect 523 99 531 133
rect 565 99 573 133
rect 523 17 573 99
rect 607 120 673 168
rect 607 86 623 120
rect 657 86 673 120
rect 607 70 673 86
rect 719 118 787 134
rect 719 84 736 118
rect 770 84 787 118
rect 719 17 787 84
rect 839 120 889 176
rect 873 86 889 120
rect 930 170 980 296
rect 930 136 946 170
rect 930 119 980 136
rect 839 85 889 86
rect 1014 85 1048 364
rect 1082 340 1116 492
rect 1187 440 1221 504
rect 1150 424 1221 440
rect 1150 390 1151 424
rect 1185 390 1221 424
rect 1397 436 1421 470
rect 1455 436 1479 470
rect 1397 420 1479 436
rect 1150 374 1221 390
rect 1338 370 1404 386
rect 1338 340 1354 370
rect 1082 336 1354 340
rect 1388 336 1404 370
rect 1082 306 1404 336
rect 1082 170 1116 306
rect 1438 272 1472 420
rect 1513 392 1547 504
rect 1581 476 1647 546
rect 1772 580 1886 649
rect 1772 546 1815 580
rect 1849 546 1886 580
rect 1772 530 1886 546
rect 1920 580 1990 596
rect 1920 546 1936 580
rect 1970 546 1990 580
rect 1581 442 1597 476
rect 1631 442 1647 476
rect 1920 509 1990 546
rect 1920 475 1936 509
rect 1970 475 1990 509
rect 1920 470 1990 475
rect 1581 426 1647 442
rect 1513 376 1576 392
rect 1513 342 1527 376
rect 1561 342 1576 376
rect 1613 390 1647 426
rect 1742 460 1990 470
rect 1742 426 1758 460
rect 1792 438 1990 460
rect 1792 426 1936 438
rect 1742 424 1936 426
rect 1920 404 1936 424
rect 1970 404 1990 438
rect 1613 356 1804 390
rect 1920 388 1990 404
rect 1513 326 1576 342
rect 1610 321 1736 322
rect 1610 287 1686 321
rect 1720 287 1736 321
rect 1610 284 1736 287
rect 1082 119 1116 136
rect 1150 256 1207 272
rect 1150 222 1157 256
rect 1191 222 1207 256
rect 1150 172 1207 222
rect 1249 256 1472 272
rect 1249 222 1265 256
rect 1299 222 1472 256
rect 1249 206 1472 222
rect 1506 271 1736 284
rect 1506 268 1644 271
rect 1540 250 1644 268
rect 1770 254 1804 356
rect 1856 338 1922 354
rect 1856 304 1872 338
rect 1906 304 1922 338
rect 1856 270 1922 304
rect 1856 254 1872 270
rect 1540 234 1572 250
rect 1506 218 1572 234
rect 1770 236 1872 254
rect 1906 236 1922 270
rect 1770 230 1922 236
rect 1438 184 1472 206
rect 1150 138 1404 172
rect 1150 85 1207 138
rect 839 51 1207 85
rect 1286 88 1336 104
rect 1286 54 1302 88
rect 1286 17 1336 54
rect 1370 85 1404 138
rect 1438 160 1504 184
rect 1438 126 1454 160
rect 1488 126 1504 160
rect 1438 119 1504 126
rect 1538 85 1572 218
rect 1678 220 1922 230
rect 1956 330 1990 388
rect 2024 580 2090 649
rect 2024 546 2040 580
rect 2074 546 2090 580
rect 2024 497 2090 546
rect 2024 463 2040 497
rect 2074 463 2090 497
rect 2024 414 2090 463
rect 2024 380 2040 414
rect 2074 380 2090 414
rect 2024 364 2090 380
rect 2130 580 2183 596
rect 2164 546 2183 580
rect 2130 497 2183 546
rect 2164 463 2183 497
rect 2130 414 2183 463
rect 2164 380 2183 414
rect 2130 364 2183 380
rect 1956 314 2115 330
rect 1956 280 1997 314
rect 2031 280 2065 314
rect 2099 280 2115 314
rect 1956 264 2115 280
rect 1678 196 1804 220
rect 1678 162 1712 196
rect 1956 186 1990 264
rect 2149 226 2183 364
rect 1370 51 1572 85
rect 1606 133 1712 162
rect 1640 99 1712 133
rect 1606 70 1712 99
rect 1748 133 1882 162
rect 1748 99 1764 133
rect 1798 99 1832 133
rect 1866 99 1882 133
rect 1748 17 1882 99
rect 1918 145 1990 186
rect 1952 111 1990 145
rect 1918 70 1990 111
rect 2030 210 2064 226
rect 2030 120 2064 176
rect 2030 17 2064 86
rect 2100 210 2183 226
rect 2100 176 2116 210
rect 2150 176 2183 210
rect 2100 120 2183 176
rect 2100 86 2116 120
rect 2150 86 2183 120
rect 2218 559 2268 575
rect 2218 525 2234 559
rect 2218 449 2268 525
rect 2218 415 2234 449
rect 2218 310 2268 415
rect 2308 559 2374 649
rect 2308 525 2324 559
rect 2358 525 2374 559
rect 2308 449 2374 525
rect 2308 415 2324 449
rect 2358 415 2374 449
rect 2308 399 2374 415
rect 2409 580 2475 596
rect 2409 546 2425 580
rect 2459 546 2475 580
rect 2409 497 2475 546
rect 2409 463 2425 497
rect 2459 463 2475 497
rect 2409 414 2475 463
rect 2409 380 2425 414
rect 2459 380 2475 414
rect 2409 364 2475 380
rect 2218 294 2397 310
rect 2218 260 2361 294
rect 2395 260 2397 294
rect 2218 244 2397 260
rect 2218 184 2262 244
rect 2431 210 2475 364
rect 2218 150 2228 184
rect 2218 108 2262 150
rect 2298 200 2373 204
rect 2298 166 2318 200
rect 2352 166 2373 200
rect 2298 120 2373 166
rect 2100 70 2183 86
rect 2298 86 2333 120
rect 2367 86 2373 120
rect 2298 17 2373 86
rect 2407 194 2475 210
rect 2407 160 2423 194
rect 2457 160 2475 194
rect 2407 120 2475 160
rect 2407 86 2423 120
rect 2457 86 2475 120
rect 2407 70 2475 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2496 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
<< metal1 >>
rect 0 683 2496 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2496 683
rect 0 617 2496 649
rect 0 17 2496 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2496 17
rect 0 -49 2496 -17
<< labels >>
rlabel comment s 0 0 0 0 4 sdfxbp_1
flabel comment s 969 337 969 337 0 FreeSans 200 0 0 0 no_jumper_check
flabel pwell s 0 0 2496 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 2496 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 2496 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 2496 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 2431 94 2465 128 0 FreeSans 340 0 0 0 Q_N
port 10 nsew
flabel corelocali s 2431 168 2465 202 0 FreeSans 340 0 0 0 Q_N
port 10 nsew
flabel corelocali s 2431 242 2465 276 0 FreeSans 340 0 0 0 Q_N
port 10 nsew
flabel corelocali s 2431 316 2465 350 0 FreeSans 340 0 0 0 Q_N
port 10 nsew
flabel corelocali s 2431 390 2465 424 0 FreeSans 340 0 0 0 Q_N
port 10 nsew
flabel corelocali s 2431 464 2465 498 0 FreeSans 340 0 0 0 Q_N
port 10 nsew
flabel corelocali s 2431 538 2465 572 0 FreeSans 340 0 0 0 Q_N
port 10 nsew
flabel corelocali s 2143 94 2177 128 0 FreeSans 340 0 0 0 Q
port 9 nsew
flabel corelocali s 2143 168 2177 202 0 FreeSans 340 0 0 0 Q
port 9 nsew
flabel corelocali s 703 242 737 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 319 168 353 202 0 FreeSans 340 0 0 0 SCE
port 4 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 SCD
port 3 nsew
flabel corelocali s 511 390 545 424 0 FreeSans 340 0 0 0 SCD
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 2496 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 296864
string GDS_START 277900
<< end >>
