magic
tech sky130A
magscale 1 2
timestamp 1604502705
<< nwell >>
rect -38 332 3494 704
<< pwell >>
rect 0 0 3456 49
<< scnmos >>
rect 111 74 141 158
rect 189 74 219 158
rect 397 113 427 197
rect 497 113 527 197
rect 575 113 605 197
rect 661 113 691 197
rect 953 125 983 209
rect 1061 125 1091 209
rect 1139 125 1169 209
rect 1358 74 1388 222
rect 1556 74 1586 222
rect 1754 97 1784 181
rect 1890 97 1920 181
rect 2013 97 2043 181
rect 2165 74 2195 202
rect 2387 74 2417 202
rect 2459 74 2489 202
rect 2561 74 2591 158
rect 2639 74 2669 158
rect 2876 74 2906 222
rect 3074 74 3104 222
rect 3160 74 3190 222
rect 3246 74 3276 222
rect 3332 74 3362 222
<< pmoshvt >>
rect 102 464 132 592
rect 186 464 216 592
rect 412 462 442 590
rect 548 462 578 590
rect 626 462 656 590
rect 716 462 746 590
rect 920 453 950 581
rect 1058 453 1088 581
rect 1142 453 1172 581
rect 1344 368 1374 592
rect 1622 368 1652 592
rect 1824 508 1854 592
rect 1914 508 1944 592
rect 2016 508 2046 592
rect 2125 398 2155 566
rect 2344 392 2374 592
rect 2535 392 2565 592
rect 2642 508 2672 592
rect 2726 508 2756 592
rect 2868 368 2898 592
rect 3070 368 3100 592
rect 3160 368 3190 592
rect 3250 368 3280 592
rect 3340 368 3370 592
<< ndiff >>
rect 340 172 397 197
rect 32 134 111 158
rect 32 100 66 134
rect 100 100 111 134
rect 32 74 111 100
rect 141 74 189 158
rect 219 133 276 158
rect 219 99 230 133
rect 264 99 276 133
rect 340 138 352 172
rect 386 138 397 172
rect 340 113 397 138
rect 427 172 497 197
rect 427 138 452 172
rect 486 138 497 172
rect 427 113 497 138
rect 527 113 575 197
rect 605 172 661 197
rect 605 138 616 172
rect 650 138 661 172
rect 605 113 661 138
rect 691 172 762 197
rect 691 138 716 172
rect 750 138 762 172
rect 691 113 762 138
rect 896 178 953 209
rect 896 144 908 178
rect 942 144 953 178
rect 896 125 953 144
rect 983 178 1061 209
rect 983 144 1008 178
rect 1042 144 1061 178
rect 983 125 1061 144
rect 1091 125 1139 209
rect 1169 184 1226 209
rect 1169 150 1180 184
rect 1214 150 1226 184
rect 1169 125 1226 150
rect 1287 184 1358 222
rect 1287 150 1299 184
rect 1333 150 1358 184
rect 219 74 276 99
rect 1287 116 1358 150
rect 1287 82 1299 116
rect 1333 82 1358 116
rect 1287 74 1358 82
rect 1388 202 1445 222
rect 1388 168 1399 202
rect 1433 168 1445 202
rect 1388 120 1445 168
rect 1388 86 1399 120
rect 1433 86 1445 120
rect 1388 74 1445 86
rect 1499 210 1556 222
rect 1499 176 1511 210
rect 1545 176 1556 210
rect 1499 120 1556 176
rect 1499 86 1511 120
rect 1545 86 1556 120
rect 1499 74 1556 86
rect 1586 210 1643 222
rect 1586 176 1597 210
rect 1631 176 1643 210
rect 2115 181 2165 202
rect 1586 120 1643 176
rect 1586 86 1597 120
rect 1631 86 1643 120
rect 1697 169 1754 181
rect 1697 135 1709 169
rect 1743 135 1754 169
rect 1697 97 1754 135
rect 1784 169 1890 181
rect 1784 135 1845 169
rect 1879 135 1890 169
rect 1784 97 1890 135
rect 1920 97 2013 181
rect 2043 120 2165 181
rect 2043 97 2070 120
rect 1586 74 1643 86
rect 2058 86 2070 97
rect 2104 86 2165 120
rect 2058 74 2165 86
rect 2195 178 2252 202
rect 2195 144 2206 178
rect 2240 144 2252 178
rect 2195 74 2252 144
rect 2330 120 2387 202
rect 2330 86 2342 120
rect 2376 86 2387 120
rect 2330 74 2387 86
rect 2417 74 2459 202
rect 2489 188 2546 202
rect 2489 154 2500 188
rect 2534 158 2546 188
rect 2803 208 2876 222
rect 2803 174 2831 208
rect 2865 174 2876 208
rect 2803 158 2876 174
rect 2534 154 2561 158
rect 2489 120 2561 154
rect 2489 86 2500 120
rect 2534 86 2561 120
rect 2489 74 2561 86
rect 2591 74 2639 158
rect 2669 120 2876 158
rect 2669 86 2680 120
rect 2714 86 2752 120
rect 2786 86 2831 120
rect 2865 86 2876 120
rect 2669 74 2876 86
rect 2906 210 2963 222
rect 2906 176 2917 210
rect 2951 176 2963 210
rect 2906 120 2963 176
rect 2906 86 2917 120
rect 2951 86 2963 120
rect 2906 74 2963 86
rect 3017 210 3074 222
rect 3017 176 3029 210
rect 3063 176 3074 210
rect 3017 120 3074 176
rect 3017 86 3029 120
rect 3063 86 3074 120
rect 3017 74 3074 86
rect 3104 210 3160 222
rect 3104 176 3115 210
rect 3149 176 3160 210
rect 3104 120 3160 176
rect 3104 86 3115 120
rect 3149 86 3160 120
rect 3104 74 3160 86
rect 3190 210 3246 222
rect 3190 176 3201 210
rect 3235 176 3246 210
rect 3190 120 3246 176
rect 3190 86 3201 120
rect 3235 86 3246 120
rect 3190 74 3246 86
rect 3276 210 3332 222
rect 3276 176 3287 210
rect 3321 176 3332 210
rect 3276 120 3332 176
rect 3276 86 3287 120
rect 3321 86 3332 120
rect 3276 74 3332 86
rect 3362 142 3419 222
rect 3362 108 3373 142
rect 3407 108 3419 142
rect 3362 74 3419 108
<< pdiff >>
rect 43 580 102 592
rect 43 546 55 580
rect 89 546 102 580
rect 43 510 102 546
rect 43 476 55 510
rect 89 476 102 510
rect 43 464 102 476
rect 132 464 186 592
rect 216 578 275 592
rect 216 544 229 578
rect 263 544 275 578
rect 216 464 275 544
rect 353 519 412 590
rect 353 485 365 519
rect 399 485 412 519
rect 353 462 412 485
rect 442 577 548 590
rect 442 543 501 577
rect 535 543 548 577
rect 442 462 548 543
rect 578 462 626 590
rect 656 578 716 590
rect 656 544 669 578
rect 703 544 716 578
rect 656 508 716 544
rect 656 474 669 508
rect 703 474 716 508
rect 656 462 716 474
rect 746 578 805 590
rect 2268 596 2326 608
rect 746 544 759 578
rect 793 544 805 578
rect 746 508 805 544
rect 746 474 759 508
rect 793 474 805 508
rect 746 462 805 474
rect 859 515 920 581
rect 859 481 871 515
rect 905 481 920 515
rect 859 453 920 481
rect 950 569 1058 581
rect 950 535 1009 569
rect 1043 535 1058 569
rect 950 453 1058 535
rect 1088 453 1142 581
rect 1172 569 1231 581
rect 1172 535 1185 569
rect 1219 535 1231 569
rect 1172 501 1231 535
rect 1172 467 1185 501
rect 1219 467 1231 501
rect 1172 453 1231 467
rect 1285 580 1344 592
rect 1285 546 1297 580
rect 1331 546 1344 580
rect 1285 368 1344 546
rect 1374 421 1433 592
rect 1563 580 1622 592
rect 1563 546 1575 580
rect 1609 546 1622 580
rect 1374 387 1387 421
rect 1421 387 1433 421
rect 1374 368 1433 387
rect 1563 368 1622 546
rect 1652 421 1711 592
rect 1765 567 1824 592
rect 1765 533 1777 567
rect 1811 533 1824 567
rect 1765 508 1824 533
rect 1854 568 1914 592
rect 1854 534 1867 568
rect 1901 534 1914 568
rect 1854 508 1914 534
rect 1944 508 2016 592
rect 2046 580 2107 592
rect 2046 546 2061 580
rect 2095 566 2107 580
rect 2095 546 2125 566
rect 2046 508 2125 546
rect 1652 387 1665 421
rect 1699 387 1711 421
rect 1652 368 1711 387
rect 2072 398 2125 508
rect 2155 444 2214 566
rect 2155 410 2168 444
rect 2202 410 2214 444
rect 2155 398 2214 410
rect 2268 562 2280 596
rect 2314 592 2326 596
rect 2314 562 2344 592
rect 2268 392 2344 562
rect 2374 392 2535 592
rect 2565 567 2642 592
rect 2565 533 2578 567
rect 2612 533 2642 567
rect 2565 508 2642 533
rect 2672 508 2726 592
rect 2756 580 2868 592
rect 2756 546 2790 580
rect 2824 546 2868 580
rect 2756 508 2868 546
rect 2565 392 2624 508
rect 2815 368 2868 508
rect 2898 580 2957 592
rect 2898 546 2911 580
rect 2945 546 2957 580
rect 2898 497 2957 546
rect 2898 463 2911 497
rect 2945 463 2957 497
rect 2898 414 2957 463
rect 2898 380 2911 414
rect 2945 380 2957 414
rect 2898 368 2957 380
rect 3011 573 3070 592
rect 3011 539 3023 573
rect 3057 539 3070 573
rect 3011 368 3070 539
rect 3100 414 3160 592
rect 3100 380 3113 414
rect 3147 380 3160 414
rect 3100 368 3160 380
rect 3190 573 3250 592
rect 3190 539 3203 573
rect 3237 539 3250 573
rect 3190 368 3250 539
rect 3280 414 3340 592
rect 3280 380 3293 414
rect 3327 380 3340 414
rect 3280 368 3340 380
rect 3370 573 3429 592
rect 3370 539 3383 573
rect 3417 539 3429 573
rect 3370 467 3429 539
rect 3370 433 3383 467
rect 3417 433 3429 467
rect 3370 368 3429 433
<< ndiffc >>
rect 66 100 100 134
rect 230 99 264 133
rect 352 138 386 172
rect 452 138 486 172
rect 616 138 650 172
rect 716 138 750 172
rect 908 144 942 178
rect 1008 144 1042 178
rect 1180 150 1214 184
rect 1299 150 1333 184
rect 1299 82 1333 116
rect 1399 168 1433 202
rect 1399 86 1433 120
rect 1511 176 1545 210
rect 1511 86 1545 120
rect 1597 176 1631 210
rect 1597 86 1631 120
rect 1709 135 1743 169
rect 1845 135 1879 169
rect 2070 86 2104 120
rect 2206 144 2240 178
rect 2342 86 2376 120
rect 2500 154 2534 188
rect 2831 174 2865 208
rect 2500 86 2534 120
rect 2680 86 2714 120
rect 2752 86 2786 120
rect 2831 86 2865 120
rect 2917 176 2951 210
rect 2917 86 2951 120
rect 3029 176 3063 210
rect 3029 86 3063 120
rect 3115 176 3149 210
rect 3115 86 3149 120
rect 3201 176 3235 210
rect 3201 86 3235 120
rect 3287 176 3321 210
rect 3287 86 3321 120
rect 3373 108 3407 142
<< pdiffc >>
rect 55 546 89 580
rect 55 476 89 510
rect 229 544 263 578
rect 365 485 399 519
rect 501 543 535 577
rect 669 544 703 578
rect 669 474 703 508
rect 759 544 793 578
rect 759 474 793 508
rect 871 481 905 515
rect 1009 535 1043 569
rect 1185 535 1219 569
rect 1185 467 1219 501
rect 1297 546 1331 580
rect 1575 546 1609 580
rect 1387 387 1421 421
rect 1777 533 1811 567
rect 1867 534 1901 568
rect 2061 546 2095 580
rect 1665 387 1699 421
rect 2168 410 2202 444
rect 2280 562 2314 596
rect 2578 533 2612 567
rect 2790 546 2824 580
rect 2911 546 2945 580
rect 2911 463 2945 497
rect 2911 380 2945 414
rect 3023 539 3057 573
rect 3113 380 3147 414
rect 3203 539 3237 573
rect 3293 380 3327 414
rect 3383 539 3417 573
rect 3383 433 3417 467
<< poly >>
rect 102 592 132 618
rect 186 592 216 618
rect 412 590 442 616
rect 548 590 578 616
rect 626 590 656 616
rect 713 605 953 635
rect 716 590 746 605
rect 917 596 953 605
rect 102 449 132 464
rect 186 449 216 464
rect 920 581 950 596
rect 1058 581 1088 607
rect 1142 581 1172 607
rect 1344 592 1374 618
rect 1622 592 1652 618
rect 1824 592 1854 618
rect 1914 592 1944 618
rect 2016 592 2046 618
rect 99 398 135 449
rect 183 424 219 449
rect 412 447 442 462
rect 548 447 578 462
rect 626 447 656 462
rect 183 408 267 424
rect 75 382 141 398
rect 75 348 91 382
rect 125 348 141 382
rect 75 314 141 348
rect 75 280 91 314
rect 125 280 141 314
rect 183 374 217 408
rect 251 374 267 408
rect 183 340 267 374
rect 351 417 581 447
rect 351 356 381 417
rect 623 369 659 447
rect 716 436 746 462
rect 920 438 950 453
rect 1058 438 1088 453
rect 1142 438 1172 453
rect 183 306 217 340
rect 251 306 267 340
rect 183 290 267 306
rect 315 340 381 356
rect 315 306 331 340
rect 365 306 381 340
rect 315 290 381 306
rect 461 353 527 369
rect 461 319 477 353
rect 511 319 527 353
rect 461 303 527 319
rect 75 246 141 280
rect 75 212 91 246
rect 125 212 141 246
rect 315 242 345 290
rect 75 196 141 212
rect 111 158 141 196
rect 189 212 427 242
rect 189 158 219 212
rect 397 197 427 212
rect 497 197 527 303
rect 575 353 659 369
rect 575 319 591 353
rect 625 319 659 353
rect 575 303 659 319
rect 803 395 869 411
rect 803 361 819 395
rect 853 361 869 395
rect 803 327 869 361
rect 575 197 605 303
rect 803 293 819 327
rect 853 293 869 327
rect 803 259 869 293
rect 803 242 819 259
rect 661 225 819 242
rect 853 225 869 259
rect 917 302 953 438
rect 1055 302 1091 438
rect 917 286 983 302
rect 917 252 933 286
rect 967 252 983 286
rect 917 236 983 252
rect 1025 286 1091 302
rect 1025 252 1041 286
rect 1075 252 1091 286
rect 1139 417 1175 438
rect 1139 401 1227 417
rect 1139 367 1177 401
rect 1211 367 1227 401
rect 1465 412 1531 428
rect 1465 378 1481 412
rect 1515 378 1531 412
rect 1139 333 1227 367
rect 1344 353 1374 368
rect 1139 299 1177 333
rect 1211 299 1227 333
rect 1139 283 1227 299
rect 1341 310 1377 353
rect 1465 347 1531 378
rect 2125 566 2155 592
rect 1824 493 1854 508
rect 1914 493 1944 508
rect 2016 493 2046 508
rect 1821 461 1857 493
rect 1911 472 1947 493
rect 1745 445 1857 461
rect 1745 411 1761 445
rect 1795 431 1857 445
rect 1905 456 1971 472
rect 1795 411 1811 431
rect 1745 395 1811 411
rect 1905 422 1921 456
rect 1955 422 1971 456
rect 1905 406 1971 422
rect 1622 353 1652 368
rect 1619 347 1655 353
rect 1905 347 1935 406
rect 1465 344 1935 347
rect 1465 310 1481 344
rect 1515 317 1935 344
rect 1515 310 1586 317
rect 1341 294 1407 310
rect 1465 294 1586 310
rect 1025 236 1091 252
rect 1341 260 1357 294
rect 1391 260 1407 294
rect 1341 244 1407 260
rect 661 212 869 225
rect 661 197 691 212
rect 803 191 869 212
rect 953 209 983 236
rect 1061 209 1091 236
rect 1139 209 1169 235
rect 1358 222 1388 244
rect 1556 222 1586 294
rect 803 157 819 191
rect 853 157 869 191
rect 803 123 869 157
rect 397 87 427 113
rect 497 87 527 113
rect 575 87 605 113
rect 661 87 691 113
rect 803 89 819 123
rect 853 89 869 123
rect 111 48 141 74
rect 189 48 219 74
rect 803 73 869 89
rect 953 51 983 125
rect 1061 99 1091 125
rect 1139 51 1169 125
rect 1754 181 1784 317
rect 2013 304 2049 493
rect 2344 592 2374 618
rect 2535 592 2565 618
rect 2642 592 2672 618
rect 2726 592 2756 618
rect 2868 592 2898 618
rect 3070 592 3100 618
rect 3160 592 3190 618
rect 3250 592 3280 618
rect 3340 592 3370 618
rect 2125 383 2155 398
rect 2642 493 2672 508
rect 2726 493 2756 508
rect 2122 366 2158 383
rect 2344 377 2374 392
rect 2535 377 2565 392
rect 2122 350 2195 366
rect 2122 316 2138 350
rect 2172 316 2195 350
rect 2013 288 2079 304
rect 2122 300 2195 316
rect 2341 304 2377 377
rect 2532 360 2568 377
rect 1890 253 1971 269
rect 1890 219 1921 253
rect 1955 219 1971 253
rect 1890 203 1971 219
rect 2013 254 2029 288
rect 2063 254 2079 288
rect 2013 238 2079 254
rect 1890 181 1920 203
rect 2013 181 2043 238
rect 2165 202 2195 300
rect 2243 288 2377 304
rect 2419 344 2489 360
rect 2419 310 2435 344
rect 2469 310 2489 344
rect 2419 294 2489 310
rect 2531 344 2597 360
rect 2531 310 2547 344
rect 2581 310 2597 344
rect 2531 294 2597 310
rect 2639 311 2675 493
rect 2723 476 2759 493
rect 2717 460 2783 476
rect 2717 426 2733 460
rect 2767 426 2783 460
rect 2717 410 2783 426
rect 2639 295 2705 311
rect 2243 254 2259 288
rect 2293 254 2327 288
rect 2361 254 2377 288
rect 2243 252 2377 254
rect 2243 222 2417 252
rect 2387 202 2417 222
rect 2459 202 2489 294
rect 953 21 1169 51
rect 1358 48 1388 74
rect 1556 48 1586 74
rect 1754 71 1784 97
rect 1890 71 1920 97
rect 2013 71 2043 97
rect 2561 158 2591 294
rect 2639 261 2655 295
rect 2689 261 2705 295
rect 2639 245 2705 261
rect 2753 203 2783 410
rect 2868 353 2898 368
rect 3070 353 3100 368
rect 3160 353 3190 368
rect 3250 353 3280 368
rect 3340 353 3370 368
rect 2865 326 2901 353
rect 3067 326 3103 353
rect 3157 326 3193 353
rect 3247 327 3283 353
rect 2833 310 3193 326
rect 2833 276 2849 310
rect 2883 276 3193 310
rect 2833 260 3193 276
rect 3246 326 3283 327
rect 3337 326 3373 353
rect 3246 310 3373 326
rect 3246 276 3262 310
rect 3296 276 3373 310
rect 3246 260 3373 276
rect 2876 222 2906 260
rect 3074 222 3104 260
rect 3160 222 3190 260
rect 3246 222 3276 260
rect 3332 222 3362 260
rect 2639 173 2783 203
rect 2639 158 2669 173
rect 2165 48 2195 74
rect 2387 48 2417 74
rect 2459 48 2489 74
rect 2561 48 2591 74
rect 2639 48 2669 74
rect 2876 48 2906 74
rect 3074 48 3104 74
rect 3160 48 3190 74
rect 3246 48 3276 74
rect 3332 48 3362 74
<< polycont >>
rect 91 348 125 382
rect 91 280 125 314
rect 217 374 251 408
rect 217 306 251 340
rect 331 306 365 340
rect 477 319 511 353
rect 91 212 125 246
rect 591 319 625 353
rect 819 361 853 395
rect 819 293 853 327
rect 819 225 853 259
rect 933 252 967 286
rect 1041 252 1075 286
rect 1177 367 1211 401
rect 1481 378 1515 412
rect 1177 299 1211 333
rect 1761 411 1795 445
rect 1921 422 1955 456
rect 1481 310 1515 344
rect 1357 260 1391 294
rect 819 157 853 191
rect 819 89 853 123
rect 2138 316 2172 350
rect 1921 219 1955 253
rect 2029 254 2063 288
rect 2435 310 2469 344
rect 2547 310 2581 344
rect 2733 426 2767 460
rect 2259 254 2293 288
rect 2327 254 2361 288
rect 2655 261 2689 295
rect 2849 276 2883 310
rect 3262 276 3296 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3391 683
rect 3425 649 3456 683
rect 17 580 105 596
rect 17 546 55 580
rect 89 546 105 580
rect 17 510 105 546
rect 213 578 263 649
rect 213 544 229 578
rect 213 526 263 544
rect 297 581 467 615
rect 17 476 55 510
rect 89 492 105 510
rect 297 492 331 581
rect 89 476 331 492
rect 17 458 331 476
rect 365 519 399 547
rect 17 146 51 458
rect 365 424 399 485
rect 433 492 467 581
rect 501 577 551 649
rect 535 543 551 577
rect 501 526 551 543
rect 653 578 709 594
rect 653 544 669 578
rect 703 544 709 578
rect 653 508 709 544
rect 653 492 669 508
rect 433 474 669 492
rect 703 474 709 508
rect 433 458 709 474
rect 201 408 527 424
rect 85 382 167 398
rect 85 348 91 382
rect 125 348 167 382
rect 85 314 167 348
rect 85 280 91 314
rect 125 280 167 314
rect 85 246 167 280
rect 85 212 91 246
rect 125 212 167 246
rect 201 374 217 408
rect 251 390 527 408
rect 251 374 267 390
rect 201 340 267 374
rect 201 306 217 340
rect 251 306 267 340
rect 201 256 267 306
rect 313 340 381 356
rect 313 306 331 340
rect 365 306 381 340
rect 313 290 381 306
rect 461 353 527 390
rect 461 319 477 353
rect 511 319 527 353
rect 461 303 527 319
rect 575 353 641 369
rect 575 319 591 353
rect 625 350 641 353
rect 575 316 607 319
rect 575 303 641 316
rect 675 269 709 458
rect 201 222 402 256
rect 85 196 167 212
rect 336 172 402 222
rect 600 235 709 269
rect 743 581 973 615
rect 743 578 793 581
rect 743 544 759 578
rect 743 508 793 544
rect 743 474 759 508
rect 743 458 793 474
rect 827 515 905 547
rect 827 481 871 515
rect 17 134 116 146
rect 17 100 66 134
rect 100 100 116 134
rect 17 84 116 100
rect 214 133 280 162
rect 214 99 230 133
rect 264 99 280 133
rect 336 138 352 172
rect 386 138 402 172
rect 336 109 402 138
rect 436 172 502 201
rect 436 138 452 172
rect 486 138 502 172
rect 214 17 280 99
rect 436 17 502 138
rect 600 172 666 235
rect 743 201 777 458
rect 827 449 905 481
rect 939 485 973 581
rect 1007 569 1061 649
rect 1007 535 1009 569
rect 1043 535 1061 569
rect 1007 519 1061 535
rect 1169 569 1261 585
rect 1169 535 1185 569
rect 1219 535 1261 569
rect 1169 501 1261 535
rect 1297 580 1347 649
rect 1331 546 1347 580
rect 1297 530 1347 546
rect 1559 580 1625 649
rect 1559 546 1575 580
rect 1609 546 1625 580
rect 1559 530 1625 546
rect 1761 567 1811 596
rect 1761 533 1777 567
rect 1761 530 1811 533
rect 1169 485 1185 501
rect 939 467 1185 485
rect 1219 496 1261 501
rect 1659 496 1811 530
rect 1845 568 1917 596
rect 1845 534 1867 568
rect 1901 534 1917 568
rect 2045 580 2111 649
rect 2045 546 2061 580
rect 2095 546 2111 580
rect 2264 596 2330 649
rect 2264 562 2280 596
rect 2314 562 2330 596
rect 2264 546 2330 562
rect 2578 567 2665 596
rect 1845 506 1917 534
rect 2612 533 2665 567
rect 1219 467 1693 496
rect 939 462 1693 467
rect 939 451 1295 462
rect 827 411 861 449
rect 600 138 616 172
rect 650 138 666 172
rect 600 109 666 138
rect 700 172 777 201
rect 700 138 716 172
rect 750 138 777 172
rect 700 109 777 138
rect 811 395 861 411
rect 811 361 819 395
rect 853 370 861 395
rect 1161 401 1227 417
rect 1161 370 1177 401
rect 853 367 1177 370
rect 1211 367 1227 401
rect 853 361 1227 367
rect 811 336 1227 361
rect 811 327 861 336
rect 811 293 819 327
rect 853 293 861 327
rect 1161 333 1227 336
rect 811 259 861 293
rect 811 225 819 259
rect 853 225 861 259
rect 895 286 983 302
rect 895 252 933 286
rect 967 252 983 286
rect 895 236 983 252
rect 1025 286 1127 302
rect 1161 299 1177 333
rect 1211 299 1227 333
rect 1161 286 1227 299
rect 1025 252 1041 286
rect 1075 252 1127 286
rect 1261 252 1295 451
rect 1371 421 1531 428
rect 1371 387 1387 421
rect 1421 412 1531 421
rect 1421 387 1481 412
rect 1371 378 1481 387
rect 1515 378 1531 412
rect 1371 364 1531 378
rect 1443 344 1531 364
rect 1443 310 1481 344
rect 1515 310 1531 344
rect 1025 236 1127 252
rect 811 202 861 225
rect 1164 218 1295 252
rect 1341 294 1409 310
rect 1341 260 1357 294
rect 1391 260 1409 294
rect 1341 236 1409 260
rect 1443 294 1531 310
rect 1581 330 1615 462
rect 1745 445 1811 461
rect 1745 428 1761 445
rect 1649 421 1761 428
rect 1649 387 1665 421
rect 1699 411 1761 421
rect 1795 411 1811 445
rect 1699 387 1811 411
rect 1649 364 1811 387
rect 1581 296 1743 330
rect 811 191 958 202
rect 811 157 819 191
rect 853 178 958 191
rect 853 157 908 178
rect 811 144 908 157
rect 942 144 958 178
rect 811 123 958 144
rect 811 89 819 123
rect 853 121 958 123
rect 992 178 1058 202
rect 992 144 1008 178
rect 1042 144 1058 178
rect 853 89 861 121
rect 811 73 861 89
rect 992 17 1058 144
rect 1164 184 1230 218
rect 1443 202 1477 294
rect 1164 150 1180 184
rect 1214 150 1230 184
rect 1164 121 1230 150
rect 1283 150 1299 184
rect 1333 150 1349 184
rect 1283 116 1349 150
rect 1283 82 1299 116
rect 1333 82 1349 116
rect 1283 17 1349 82
rect 1383 168 1399 202
rect 1433 168 1477 202
rect 1383 120 1477 168
rect 1383 86 1399 120
rect 1433 86 1477 120
rect 1383 70 1477 86
rect 1511 210 1545 226
rect 1511 120 1545 176
rect 1511 17 1545 86
rect 1581 210 1647 226
rect 1581 176 1597 210
rect 1631 176 1647 210
rect 1581 120 1647 176
rect 1581 86 1597 120
rect 1631 86 1647 120
rect 1693 169 1743 296
rect 1693 135 1709 169
rect 1693 119 1743 135
rect 1581 85 1647 86
rect 1777 85 1811 364
rect 1845 372 1879 506
rect 1951 478 2544 512
rect 2578 504 2665 533
rect 2753 580 2861 649
rect 2753 546 2790 580
rect 2824 546 2861 580
rect 2753 530 2861 546
rect 2895 580 2967 596
rect 2895 546 2911 580
rect 2945 546 2967 580
rect 1951 472 1985 478
rect 1913 456 1985 472
rect 1913 422 1921 456
rect 1955 422 1985 456
rect 1913 406 1985 422
rect 2152 410 2168 444
rect 2202 410 2277 444
rect 1845 350 2188 372
rect 1845 338 2138 350
rect 1845 169 1879 338
rect 2122 316 2138 338
rect 2172 316 2188 350
rect 2122 306 2188 316
rect 2243 304 2277 410
rect 2510 360 2544 478
rect 2631 377 2665 504
rect 2895 498 2967 546
rect 3007 573 3073 649
rect 3007 539 3023 573
rect 3057 539 3073 573
rect 3007 532 3073 539
rect 3187 573 3253 649
rect 3187 539 3203 573
rect 3237 539 3253 573
rect 3187 532 3253 539
rect 2895 497 3237 498
rect 2895 476 2911 497
rect 2717 463 2911 476
rect 2945 464 3237 497
rect 2945 463 3047 464
rect 2717 460 3047 463
rect 2717 426 2733 460
rect 2767 426 3047 460
rect 2717 414 3047 426
rect 2717 411 2911 414
rect 2895 380 2911 411
rect 2945 380 3047 414
rect 2416 344 2476 360
rect 2416 310 2435 344
rect 2469 310 2476 344
rect 2013 288 2079 304
rect 1845 119 1879 135
rect 1913 253 1971 269
rect 1913 219 1921 253
rect 1955 219 1971 253
rect 2013 254 2029 288
rect 2063 272 2079 288
rect 2243 288 2377 304
rect 2243 272 2259 288
rect 2063 254 2259 272
rect 2293 254 2327 288
rect 2361 254 2377 288
rect 2013 238 2377 254
rect 2416 260 2476 310
rect 2510 344 2597 360
rect 2510 310 2547 344
rect 2581 310 2597 344
rect 2631 343 2773 377
rect 2895 360 3047 380
rect 2510 294 2597 310
rect 2739 326 2773 343
rect 2933 350 3047 360
rect 2739 310 2899 326
rect 2639 295 2705 309
rect 2639 261 2655 295
rect 2689 261 2705 295
rect 2639 260 2705 261
rect 1913 204 1971 219
rect 1913 170 2172 204
rect 1913 85 1947 170
rect 1581 51 1947 85
rect 2054 120 2104 136
rect 2054 86 2070 120
rect 2054 17 2104 86
rect 2138 85 2172 170
rect 2206 178 2240 238
rect 2416 226 2705 260
rect 2739 276 2849 310
rect 2883 276 2899 310
rect 2739 260 2899 276
rect 2933 316 3007 350
rect 3041 316 3047 350
rect 2933 310 3047 316
rect 3097 414 3165 430
rect 3097 380 3113 414
rect 3147 380 3165 414
rect 2416 204 2450 226
rect 2206 119 2240 144
rect 2274 170 2450 204
rect 2739 188 2773 260
rect 2933 226 2967 310
rect 2274 85 2308 170
rect 2484 154 2500 188
rect 2534 154 2773 188
rect 2813 208 2867 224
rect 2813 174 2831 208
rect 2865 174 2867 208
rect 2138 51 2308 85
rect 2342 120 2392 136
rect 2376 86 2392 120
rect 2342 17 2392 86
rect 2484 120 2550 154
rect 2813 120 2867 174
rect 2484 86 2500 120
rect 2534 86 2550 120
rect 2484 70 2550 86
rect 2664 86 2680 120
rect 2714 86 2752 120
rect 2786 86 2831 120
rect 2865 86 2867 120
rect 2664 17 2867 86
rect 2901 210 2967 226
rect 2901 176 2917 210
rect 2951 176 2967 210
rect 2901 120 2967 176
rect 2901 86 2917 120
rect 2951 86 2967 120
rect 2901 70 2967 86
rect 3013 210 3063 226
rect 3013 176 3029 210
rect 3013 120 3063 176
rect 3013 86 3029 120
rect 3013 17 3063 86
rect 3097 210 3165 380
rect 3199 327 3237 464
rect 3287 414 3333 602
rect 3367 573 3433 649
rect 3367 539 3383 573
rect 3417 539 3433 573
rect 3367 467 3433 539
rect 3367 433 3383 467
rect 3417 433 3433 467
rect 3367 429 3433 433
rect 3287 380 3293 414
rect 3327 395 3333 414
rect 3327 380 3433 395
rect 3287 361 3433 380
rect 3199 310 3302 327
rect 3199 276 3262 310
rect 3296 276 3302 310
rect 3199 260 3302 276
rect 3340 226 3433 361
rect 3097 176 3115 210
rect 3149 176 3165 210
rect 3097 120 3165 176
rect 3097 86 3115 120
rect 3149 86 3165 120
rect 3097 70 3165 86
rect 3201 210 3235 226
rect 3201 120 3235 176
rect 3201 17 3235 86
rect 3271 210 3433 226
rect 3271 176 3287 210
rect 3321 192 3433 210
rect 3321 176 3337 192
rect 3271 120 3337 176
rect 3271 86 3287 120
rect 3321 86 3337 120
rect 3271 70 3337 86
rect 3371 142 3423 158
rect 3371 108 3373 142
rect 3407 108 3423 142
rect 3371 17 3423 108
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3456 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 3199 649 3233 683
rect 3295 649 3329 683
rect 3391 649 3425 683
rect 607 319 625 350
rect 625 319 641 350
rect 607 316 641 319
rect 3007 316 3041 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
<< metal1 >>
rect 0 683 3456 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3391 683
rect 3425 649 3456 683
rect 0 617 3456 649
rect 595 350 653 356
rect 595 316 607 350
rect 641 347 653 350
rect 2995 350 3053 356
rect 2995 347 3007 350
rect 641 319 3007 347
rect 641 316 653 319
rect 595 310 653 316
rect 2995 316 3007 319
rect 3041 316 3053 350
rect 2995 310 3053 316
rect 0 17 3456 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3456 17
rect 0 -49 3456 -17
<< labels >>
rlabel comment s 0 0 0 0 4 sedfxbp_2
flabel comment s 1687 337 1687 337 0 FreeSans 200 0 0 0 no_jumper_check
flabel pwell s 0 0 3456 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 0 617 3456 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 0 617 3456 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 3456 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 3103 94 3137 128 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 3103 168 3137 202 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 3103 242 3137 276 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 3103 316 3137 350 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 3103 390 3137 424 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 3295 94 3329 128 0 FreeSans 340 0 0 0 Q_N
port 11 nsew
flabel corelocali s 3295 168 3329 202 0 FreeSans 340 0 0 0 Q_N
port 11 nsew
flabel corelocali s 3295 390 3329 424 0 FreeSans 340 0 0 0 Q_N
port 11 nsew
flabel corelocali s 3295 464 3329 498 0 FreeSans 340 0 0 0 Q_N
port 11 nsew
flabel corelocali s 3295 538 3329 572 0 FreeSans 340 0 0 0 Q_N
port 11 nsew
flabel corelocali s 127 242 161 276 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 1375 242 1409 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 1087 242 1121 276 0 FreeSans 340 0 0 0 SCD
port 4 nsew
flabel corelocali s 895 242 929 276 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 DE
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 3456 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 500578
string GDS_START 476390
<< end >>
