magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 18 195 88 325
rect 291 333 354 401
rect 291 123 381 333
rect 1848 325 1906 493
rect 1848 291 2002 325
rect 1925 181 2002 291
rect 1830 147 2002 181
rect 1830 51 1906 147
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 18 393 69 493
rect 103 427 179 527
rect 18 359 178 393
rect 132 255 178 359
rect 166 221 178 255
rect 132 161 178 221
rect 18 127 178 161
rect 223 391 257 493
rect 354 435 388 527
rect 434 427 484 493
rect 537 427 673 493
rect 434 401 468 427
rect 18 69 69 127
rect 103 17 179 93
rect 223 69 257 357
rect 415 367 468 401
rect 502 391 605 393
rect 415 95 449 367
rect 502 357 545 391
rect 579 357 605 391
rect 502 315 605 357
rect 485 255 537 277
rect 485 221 496 255
rect 530 221 537 255
rect 485 153 537 221
rect 571 197 605 315
rect 639 271 673 427
rect 707 407 741 475
rect 798 441 864 527
rect 908 407 942 475
rect 1001 435 1085 527
rect 707 373 942 407
rect 1129 401 1163 493
rect 1210 425 1401 493
rect 1468 435 1518 527
rect 1031 367 1163 401
rect 1031 339 1065 367
rect 745 305 1065 339
rect 1229 357 1294 391
rect 1328 357 1332 391
rect 1229 333 1332 357
rect 639 237 997 271
rect 571 153 642 197
rect 686 95 720 237
rect 761 187 929 203
rect 963 201 997 237
rect 761 153 821 187
rect 855 153 893 187
rect 927 153 929 187
rect 1031 167 1065 305
rect 315 17 381 89
rect 415 61 499 95
rect 539 61 720 95
rect 905 17 971 109
rect 1013 89 1065 167
rect 1121 331 1332 333
rect 1367 349 1401 425
rect 1562 417 1596 475
rect 1632 451 1708 527
rect 1562 383 1722 417
rect 1121 299 1263 331
rect 1367 315 1654 349
rect 1121 141 1155 299
rect 1367 297 1411 315
rect 1189 255 1263 265
rect 1189 221 1204 255
rect 1238 221 1263 255
rect 1189 141 1263 221
rect 1297 263 1411 297
rect 1297 107 1331 263
rect 1391 173 1445 229
rect 1501 187 1581 281
rect 1688 259 1722 383
rect 1762 315 1796 527
rect 1950 359 1984 527
rect 1391 139 1467 173
rect 1013 55 1093 89
rect 1147 51 1331 107
rect 1365 17 1399 105
rect 1433 93 1467 139
rect 1501 153 1527 187
rect 1561 153 1581 187
rect 1501 127 1581 153
rect 1658 257 1722 259
rect 1658 215 1867 257
rect 1658 93 1727 215
rect 1433 59 1727 93
rect 1762 17 1796 179
rect 1950 17 1984 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 132 221 166 255
rect 223 357 257 391
rect 545 357 579 391
rect 496 221 530 255
rect 1294 357 1328 391
rect 821 153 855 187
rect 893 153 927 187
rect 1204 221 1238 255
rect 1527 153 1561 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
<< metal1 >>
rect 0 561 2024 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 0 496 2024 527
rect 799 187 949 193
rect 799 153 821 187
rect 855 153 893 187
rect 927 184 949 187
rect 1515 187 1573 193
rect 1515 184 1527 187
rect 927 156 1527 184
rect 927 153 949 156
rect 799 147 949 153
rect 1515 153 1527 156
rect 1561 153 1573 187
rect 1515 147 1573 153
rect 0 17 2024 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
rect 0 -48 2024 -17
<< obsm1 >>
rect 201 391 269 397
rect 201 357 223 391
rect 257 388 269 391
rect 533 391 591 397
rect 533 388 545 391
rect 257 360 545 388
rect 257 357 269 360
rect 201 351 269 357
rect 533 357 545 360
rect 579 388 591 391
rect 1282 391 1340 397
rect 1282 388 1294 391
rect 579 360 1294 388
rect 579 357 591 360
rect 533 351 591 357
rect 1282 357 1294 360
rect 1328 357 1340 391
rect 1282 351 1340 357
rect 120 255 178 261
rect 120 221 132 255
rect 166 252 178 255
rect 484 255 542 261
rect 484 252 496 255
rect 166 224 496 252
rect 166 221 178 224
rect 120 215 178 221
rect 484 221 496 224
rect 530 252 542 255
rect 1192 255 1250 261
rect 1192 252 1204 255
rect 530 224 1204 252
rect 530 221 542 224
rect 484 215 542 221
rect 1192 221 1204 224
rect 1238 221 1250 255
rect 1192 215 1250 221
<< labels >>
rlabel locali s 18 195 88 325 6 CLK
port 1 nsew signal input
rlabel locali s 291 333 354 401 6 D
port 2 nsew signal input
rlabel locali s 291 123 381 333 6 D
port 2 nsew signal input
rlabel locali s 1925 181 2002 291 6 Q
port 3 nsew signal output
rlabel locali s 1848 325 1906 493 6 Q
port 3 nsew signal output
rlabel locali s 1848 291 2002 325 6 Q
port 3 nsew signal output
rlabel locali s 1830 147 2002 181 6 Q
port 3 nsew signal output
rlabel locali s 1830 51 1906 147 6 Q
port 3 nsew signal output
rlabel metal1 s 1515 184 1573 193 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 1515 147 1573 156 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 799 184 949 193 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 799 156 1573 184 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 799 147 949 156 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 0 -48 2024 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 2024 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2024 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1860434
string GDS_START 1845400
<< end >>
