magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 17 199 75 394
rect 109 342 171 493
rect 325 342 363 493
rect 605 342 681 425
rect 109 308 681 342
rect 109 134 185 308
rect 243 215 442 273
rect 534 215 727 271
rect 761 215 983 259
rect 893 153 983 215
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 23 435 75 527
rect 205 383 281 527
rect 397 383 473 527
rect 519 459 763 493
rect 519 420 571 459
rect 725 339 763 459
rect 797 373 873 527
rect 917 339 969 493
rect 725 305 969 339
rect 229 93 267 178
rect 301 127 859 169
rect 821 103 859 127
rect 229 89 473 93
rect 19 51 473 89
rect 519 17 585 89
rect 705 17 781 89
rect 893 17 974 89
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
rlabel locali s 893 153 983 215 6 A1
port 1 nsew signal input
rlabel locali s 761 215 983 259 6 A1
port 1 nsew signal input
rlabel locali s 534 215 727 271 6 A2
port 2 nsew signal input
rlabel locali s 243 215 442 273 6 B1
port 3 nsew signal input
rlabel locali s 17 199 75 394 6 C1
port 4 nsew signal input
rlabel locali s 605 342 681 425 6 Y
port 5 nsew signal output
rlabel locali s 325 342 363 493 6 Y
port 5 nsew signal output
rlabel locali s 109 342 171 493 6 Y
port 5 nsew signal output
rlabel locali s 109 308 681 342 6 Y
port 5 nsew signal output
rlabel locali s 109 134 185 308 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -48 1012 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 1012 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1012 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 987786
string GDS_START 980022
<< end >>
