magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 2430 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 89 47 119 131
rect 183 47 213 131
rect 381 47 411 175
rect 476 47 506 119
rect 606 47 636 119
rect 702 47 732 131
rect 836 47 866 131
rect 908 47 938 131
rect 1126 47 1156 131
rect 1208 47 1238 131
rect 1314 47 1344 131
rect 1386 47 1416 131
rect 1458 47 1488 131
rect 1602 47 1632 155
rect 1800 47 1830 131
rect 1895 47 1925 177
rect 1989 47 2019 177
rect 2083 47 2113 177
rect 2177 47 2207 177
rect 2281 47 2311 177
<< pmoshvt >>
rect 81 363 117 491
rect 175 363 211 491
rect 373 329 409 497
rect 480 413 516 497
rect 574 413 610 497
rect 704 413 740 497
rect 820 413 856 497
rect 914 413 950 497
rect 1008 413 1044 497
rect 1090 413 1126 497
rect 1208 413 1244 497
rect 1290 413 1326 497
rect 1488 413 1524 497
rect 1594 329 1630 497
rect 1792 369 1828 497
rect 1897 297 1933 497
rect 1991 297 2027 497
rect 2085 297 2121 497
rect 2179 297 2215 497
rect 2273 297 2309 497
<< ndiff >>
rect 27 119 89 131
rect 27 85 35 119
rect 69 85 89 119
rect 27 47 89 85
rect 119 93 183 131
rect 119 59 129 93
rect 163 59 183 93
rect 119 47 183 59
rect 213 119 265 131
rect 213 85 223 119
rect 257 85 265 119
rect 213 47 265 85
rect 319 93 381 175
rect 319 59 327 93
rect 361 59 381 93
rect 319 47 381 59
rect 411 119 461 175
rect 1542 131 1602 155
rect 651 119 702 131
rect 411 111 476 119
rect 411 77 421 111
rect 455 77 476 111
rect 411 47 476 77
rect 506 93 606 119
rect 506 59 541 93
rect 575 59 606 93
rect 506 47 606 59
rect 636 47 702 119
rect 732 89 836 131
rect 732 55 782 89
rect 816 55 836 89
rect 732 47 836 55
rect 866 47 908 131
rect 938 109 1000 131
rect 938 75 958 109
rect 992 75 1000 109
rect 938 47 1000 75
rect 1064 93 1126 131
rect 1064 59 1072 93
rect 1106 59 1126 93
rect 1064 47 1126 59
rect 1156 47 1208 131
rect 1238 95 1314 131
rect 1238 61 1254 95
rect 1288 61 1314 95
rect 1238 47 1314 61
rect 1344 47 1386 131
rect 1416 47 1458 131
rect 1488 113 1602 131
rect 1488 79 1528 113
rect 1562 79 1602 113
rect 1488 47 1602 79
rect 1632 120 1684 155
rect 1845 131 1895 177
rect 1632 86 1642 120
rect 1676 86 1684 120
rect 1632 47 1684 86
rect 1738 119 1800 131
rect 1738 85 1746 119
rect 1780 85 1800 119
rect 1738 47 1800 85
rect 1830 93 1895 131
rect 1830 59 1851 93
rect 1885 59 1895 93
rect 1830 47 1895 59
rect 1925 143 1989 177
rect 1925 109 1945 143
rect 1979 109 1989 143
rect 1925 47 1989 109
rect 2019 93 2083 177
rect 2019 59 2039 93
rect 2073 59 2083 93
rect 2019 47 2083 59
rect 2113 143 2177 177
rect 2113 109 2133 143
rect 2167 109 2177 143
rect 2113 47 2177 109
rect 2207 93 2281 177
rect 2207 59 2227 93
rect 2261 59 2281 93
rect 2207 47 2281 59
rect 2311 143 2363 177
rect 2311 109 2321 143
rect 2355 109 2363 143
rect 2311 47 2363 109
<< pdiff >>
rect 27 477 81 491
rect 27 443 35 477
rect 69 443 81 477
rect 27 409 81 443
rect 27 375 35 409
rect 69 375 81 409
rect 27 363 81 375
rect 117 461 175 491
rect 117 427 129 461
rect 163 427 175 461
rect 117 363 175 427
rect 211 477 265 491
rect 211 443 223 477
rect 257 443 265 477
rect 211 409 265 443
rect 211 375 223 409
rect 257 375 265 409
rect 211 363 265 375
rect 319 461 373 497
rect 319 427 327 461
rect 361 427 373 461
rect 319 329 373 427
rect 409 477 480 497
rect 409 443 421 477
rect 455 443 480 477
rect 409 413 480 443
rect 516 484 574 497
rect 516 450 528 484
rect 562 450 574 484
rect 516 413 574 450
rect 610 413 704 497
rect 740 485 820 497
rect 740 451 762 485
rect 796 451 820 485
rect 740 413 820 451
rect 856 459 914 497
rect 856 425 868 459
rect 902 425 914 459
rect 856 413 914 425
rect 950 485 1008 497
rect 950 451 962 485
rect 996 451 1008 485
rect 950 413 1008 451
rect 1044 413 1090 497
rect 1126 483 1208 497
rect 1126 449 1138 483
rect 1172 449 1208 483
rect 1126 413 1208 449
rect 1244 413 1290 497
rect 1326 485 1380 497
rect 1326 451 1338 485
rect 1372 451 1380 485
rect 1326 413 1380 451
rect 1434 459 1488 497
rect 1434 425 1442 459
rect 1476 425 1488 459
rect 1434 413 1488 425
rect 1524 459 1594 497
rect 1524 425 1548 459
rect 1582 425 1594 459
rect 1524 413 1594 425
rect 409 409 463 413
rect 409 375 421 409
rect 455 375 463 409
rect 409 329 463 375
rect 1541 329 1594 413
rect 1630 459 1684 497
rect 1630 425 1642 459
rect 1676 425 1684 459
rect 1630 391 1684 425
rect 1630 357 1642 391
rect 1676 357 1684 391
rect 1738 485 1792 497
rect 1738 451 1746 485
rect 1780 451 1792 485
rect 1738 417 1792 451
rect 1738 383 1746 417
rect 1780 383 1792 417
rect 1738 369 1792 383
rect 1828 485 1897 497
rect 1828 451 1851 485
rect 1885 451 1897 485
rect 1828 417 1897 451
rect 1828 383 1851 417
rect 1885 383 1897 417
rect 1828 369 1897 383
rect 1630 329 1684 357
rect 1845 297 1897 369
rect 1933 449 1991 497
rect 1933 415 1945 449
rect 1979 415 1991 449
rect 1933 381 1991 415
rect 1933 347 1945 381
rect 1979 347 1991 381
rect 1933 297 1991 347
rect 2027 449 2085 497
rect 2027 415 2039 449
rect 2073 415 2085 449
rect 2027 297 2085 415
rect 2121 449 2179 497
rect 2121 415 2133 449
rect 2167 415 2179 449
rect 2121 381 2179 415
rect 2121 347 2133 381
rect 2167 347 2179 381
rect 2121 297 2179 347
rect 2215 489 2273 497
rect 2215 455 2227 489
rect 2261 455 2273 489
rect 2215 421 2273 455
rect 2215 387 2227 421
rect 2261 387 2273 421
rect 2215 297 2273 387
rect 2309 449 2363 497
rect 2309 415 2321 449
rect 2355 415 2363 449
rect 2309 381 2363 415
rect 2309 347 2321 381
rect 2355 347 2363 381
rect 2309 297 2363 347
<< ndiffc >>
rect 35 85 69 119
rect 129 59 163 93
rect 223 85 257 119
rect 327 59 361 93
rect 421 77 455 111
rect 541 59 575 93
rect 782 55 816 89
rect 958 75 992 109
rect 1072 59 1106 93
rect 1254 61 1288 95
rect 1528 79 1562 113
rect 1642 86 1676 120
rect 1746 85 1780 119
rect 1851 59 1885 93
rect 1945 109 1979 143
rect 2039 59 2073 93
rect 2133 109 2167 143
rect 2227 59 2261 93
rect 2321 109 2355 143
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 129 427 163 461
rect 223 443 257 477
rect 223 375 257 409
rect 327 427 361 461
rect 421 443 455 477
rect 528 450 562 484
rect 762 451 796 485
rect 868 425 902 459
rect 962 451 996 485
rect 1138 449 1172 483
rect 1338 451 1372 485
rect 1442 425 1476 459
rect 1548 425 1582 459
rect 421 375 455 409
rect 1642 425 1676 459
rect 1642 357 1676 391
rect 1746 451 1780 485
rect 1746 383 1780 417
rect 1851 451 1885 485
rect 1851 383 1885 417
rect 1945 415 1979 449
rect 1945 347 1979 381
rect 2039 415 2073 449
rect 2133 415 2167 449
rect 2133 347 2167 381
rect 2227 455 2261 489
rect 2227 387 2261 421
rect 2321 415 2355 449
rect 2321 347 2355 381
<< poly >>
rect 81 491 117 517
rect 175 491 211 517
rect 373 497 409 523
rect 480 497 516 523
rect 574 497 610 523
rect 704 497 740 523
rect 820 497 856 523
rect 914 497 950 523
rect 1008 497 1044 523
rect 1090 497 1126 523
rect 1208 497 1244 523
rect 1290 497 1326 523
rect 1488 497 1524 523
rect 1594 497 1630 523
rect 1792 497 1828 523
rect 1897 497 1933 523
rect 1991 497 2027 523
rect 2085 497 2121 523
rect 2179 497 2215 523
rect 2273 497 2309 523
rect 81 348 117 363
rect 175 348 211 363
rect 46 318 119 348
rect 46 280 76 318
rect 22 264 76 280
rect 173 274 213 348
rect 480 398 516 413
rect 574 398 610 413
rect 704 398 740 413
rect 820 398 856 413
rect 914 398 950 413
rect 1008 398 1044 413
rect 1090 398 1126 413
rect 1208 398 1244 413
rect 1290 398 1326 413
rect 1488 398 1524 413
rect 373 314 409 329
rect 22 230 32 264
rect 66 230 76 264
rect 22 214 76 230
rect 128 264 213 274
rect 371 267 411 314
rect 478 279 518 398
rect 572 375 612 398
rect 702 381 742 398
rect 560 365 636 375
rect 560 331 576 365
rect 610 331 636 365
rect 560 321 636 331
rect 702 365 776 381
rect 702 331 722 365
rect 756 331 776 365
rect 702 315 776 331
rect 128 230 144 264
rect 178 230 213 264
rect 128 220 213 230
rect 46 176 76 214
rect 46 146 119 176
rect 89 131 119 146
rect 183 131 213 220
rect 364 251 428 267
rect 364 217 374 251
rect 408 217 428 251
rect 478 249 636 279
rect 364 201 428 217
rect 606 219 636 249
rect 381 175 411 201
rect 476 191 554 207
rect 476 157 500 191
rect 534 157 554 191
rect 476 141 554 157
rect 606 203 660 219
rect 606 169 616 203
rect 650 169 660 203
rect 606 153 660 169
rect 476 119 506 141
rect 606 119 636 153
rect 702 131 732 315
rect 818 229 858 398
rect 912 313 952 398
rect 1006 313 1046 398
rect 1088 375 1128 398
rect 1088 365 1164 375
rect 1088 331 1104 365
rect 1138 331 1164 365
rect 1088 321 1164 331
rect 900 297 1046 313
rect 900 263 910 297
rect 944 263 1046 297
rect 1206 291 1246 398
rect 1194 279 1246 291
rect 900 247 1046 263
rect 1130 269 1246 279
rect 788 213 858 229
rect 788 179 798 213
rect 832 193 858 213
rect 832 179 866 193
rect 788 163 866 179
rect 836 131 866 163
rect 908 183 948 247
rect 1130 235 1146 269
rect 1180 261 1246 269
rect 1288 365 1328 398
rect 1288 349 1362 365
rect 1288 315 1308 349
rect 1342 315 1362 349
rect 1486 337 1526 398
rect 1288 291 1362 315
rect 1482 307 1526 337
rect 1792 354 1828 369
rect 1594 314 1630 329
rect 1288 261 1416 291
rect 1180 235 1238 261
rect 1130 225 1238 235
rect 908 147 1156 183
rect 908 131 938 147
rect 1126 131 1156 147
rect 1208 131 1238 225
rect 1280 203 1344 219
rect 1280 169 1290 203
rect 1324 169 1344 203
rect 1280 153 1344 169
rect 1314 131 1344 153
rect 1386 131 1416 261
rect 1482 229 1522 307
rect 1592 285 1632 314
rect 1790 285 1830 354
rect 1458 213 1522 229
rect 1564 269 1830 285
rect 1897 282 1933 297
rect 1991 282 2027 297
rect 2085 282 2121 297
rect 2179 282 2215 297
rect 2273 282 2309 297
rect 1564 235 1574 269
rect 1608 235 1830 269
rect 1564 219 1830 235
rect 1458 179 1468 213
rect 1502 179 1522 213
rect 1458 163 1522 179
rect 1458 131 1488 163
rect 1602 155 1632 219
rect 1800 131 1830 219
rect 1895 259 1935 282
rect 1989 259 2029 282
rect 2083 259 2123 282
rect 2177 259 2217 282
rect 2271 259 2311 282
rect 1895 249 2311 259
rect 1895 215 1911 249
rect 1945 215 1989 249
rect 2023 215 2067 249
rect 2101 215 2145 249
rect 2179 215 2223 249
rect 2257 215 2311 249
rect 1895 205 2311 215
rect 1895 177 1925 205
rect 1989 177 2019 205
rect 2083 177 2113 205
rect 2177 177 2207 205
rect 2281 177 2311 205
rect 89 21 119 47
rect 183 21 213 47
rect 381 21 411 47
rect 476 21 506 47
rect 606 21 636 47
rect 702 21 732 47
rect 836 21 866 47
rect 908 21 938 47
rect 1126 21 1156 47
rect 1208 21 1238 47
rect 1314 21 1344 47
rect 1386 21 1416 47
rect 1458 21 1488 47
rect 1602 21 1632 47
rect 1800 21 1830 47
rect 1895 21 1925 47
rect 1989 21 2019 47
rect 2083 21 2113 47
rect 2177 21 2207 47
rect 2281 21 2311 47
<< polycont >>
rect 32 230 66 264
rect 576 331 610 365
rect 722 331 756 365
rect 144 230 178 264
rect 374 217 408 251
rect 500 157 534 191
rect 616 169 650 203
rect 1104 331 1138 365
rect 910 263 944 297
rect 798 179 832 213
rect 1146 235 1180 269
rect 1308 315 1342 349
rect 1290 169 1324 203
rect 1574 235 1608 269
rect 1468 179 1502 213
rect 1911 215 1945 249
rect 1989 215 2023 249
rect 2067 215 2101 249
rect 2145 215 2179 249
rect 2223 215 2257 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2392 561
rect 35 477 69 493
rect 35 409 69 443
rect 103 461 179 527
rect 103 427 129 461
rect 163 427 179 461
rect 223 477 268 493
rect 257 443 268 477
rect 223 409 268 443
rect 311 461 377 527
rect 311 427 327 461
rect 361 427 377 461
rect 421 477 455 493
rect 746 485 822 527
rect 502 450 528 484
rect 562 450 688 484
rect 746 451 762 485
rect 796 451 822 485
rect 936 485 1012 527
rect 868 459 902 475
rect 69 382 178 393
rect 69 375 133 382
rect 35 359 133 375
rect 132 348 133 359
rect 167 348 178 382
rect 18 264 88 325
rect 18 230 32 264
rect 66 230 88 264
rect 18 195 88 230
rect 132 264 178 348
rect 132 230 144 264
rect 132 161 178 230
rect 35 127 178 161
rect 257 375 268 409
rect 421 409 455 443
rect 223 178 268 375
rect 223 144 233 178
rect 267 144 268 178
rect 35 119 69 127
rect 223 119 268 144
rect 306 375 421 393
rect 306 359 455 375
rect 500 382 620 391
rect 306 165 340 359
rect 500 348 529 382
rect 563 365 620 382
rect 563 348 576 365
rect 500 331 576 348
rect 610 331 620 365
rect 374 251 466 325
rect 408 217 466 251
rect 374 201 466 217
rect 500 315 620 331
rect 500 191 554 315
rect 654 281 688 450
rect 936 451 962 485
rect 996 451 1012 485
rect 1294 485 1388 527
rect 1112 449 1138 483
rect 1172 449 1258 483
rect 1294 451 1338 485
rect 1372 451 1388 485
rect 1428 459 1476 475
rect 1112 433 1258 449
rect 868 417 902 425
rect 1214 417 1258 433
rect 1428 425 1442 459
rect 1428 417 1476 425
rect 722 367 1022 417
rect 722 365 782 367
rect 756 331 782 365
rect 722 315 782 331
rect 894 297 954 313
rect 894 281 910 297
rect 654 263 910 281
rect 944 263 954 297
rect 654 247 954 263
rect 654 246 748 247
rect 306 127 455 165
rect 534 157 554 191
rect 500 141 554 157
rect 590 169 616 203
rect 650 178 670 203
rect 590 144 631 169
rect 665 144 670 178
rect 590 129 670 144
rect 35 69 69 85
rect 103 59 129 93
rect 163 59 179 93
rect 257 85 268 119
rect 421 111 455 127
rect 223 69 268 85
rect 103 17 179 59
rect 311 59 327 93
rect 361 59 377 93
rect 704 93 748 246
rect 988 213 1022 367
rect 782 179 798 213
rect 832 187 902 213
rect 832 179 856 187
rect 782 153 856 179
rect 890 153 902 187
rect 782 147 902 153
rect 958 145 1022 213
rect 1066 382 1180 393
rect 1066 365 1141 382
rect 1066 331 1104 365
rect 1138 348 1141 365
rect 1175 348 1180 382
rect 1138 331 1180 348
rect 1214 383 1476 417
rect 1542 459 1608 527
rect 1838 485 1909 527
rect 1542 425 1548 459
rect 1582 425 1608 459
rect 1542 389 1608 425
rect 1642 459 1676 475
rect 1642 391 1676 425
rect 1066 179 1100 331
rect 1144 269 1180 295
rect 1144 256 1146 269
rect 1144 222 1145 256
rect 1214 281 1258 383
rect 1730 451 1746 485
rect 1780 451 1796 485
rect 1730 417 1796 451
rect 1730 383 1746 417
rect 1780 383 1796 417
rect 1642 353 1676 357
rect 1642 349 1710 353
rect 1292 315 1308 349
rect 1342 315 1710 349
rect 1214 269 1634 281
rect 1214 247 1574 269
rect 1179 222 1180 235
rect 1144 213 1180 222
rect 1274 179 1290 203
rect 1066 169 1290 179
rect 1324 169 1350 203
rect 1066 145 1350 169
rect 958 109 992 145
rect 421 61 455 77
rect 311 17 377 59
rect 525 59 541 93
rect 575 59 748 93
rect 525 53 748 59
rect 782 89 874 105
rect 816 55 874 89
rect 958 59 992 75
rect 1028 93 1106 109
rect 1384 95 1418 247
rect 1558 235 1574 247
rect 1608 235 1634 269
rect 1452 179 1468 213
rect 1502 201 1528 213
rect 1502 187 1556 201
rect 1452 153 1501 179
rect 1535 153 1556 187
rect 1452 147 1556 153
rect 1668 136 1710 315
rect 1642 120 1710 136
rect 1028 59 1072 93
rect 1238 61 1254 95
rect 1288 61 1418 95
rect 1464 79 1528 113
rect 1562 79 1606 113
rect 782 17 874 55
rect 1028 17 1106 59
rect 1464 17 1606 79
rect 1676 86 1710 120
rect 1642 70 1710 86
rect 1746 255 1796 383
rect 1838 451 1851 485
rect 1885 451 1909 485
rect 1838 417 1909 451
rect 1838 383 1851 417
rect 1885 383 1909 417
rect 1838 367 1909 383
rect 1945 449 1999 493
rect 1979 415 1999 449
rect 1945 381 1999 415
rect 1979 347 1999 381
rect 2033 449 2084 527
rect 2033 415 2039 449
rect 2073 415 2084 449
rect 2033 362 2084 415
rect 2133 449 2167 493
rect 2133 381 2167 415
rect 1945 328 1999 347
rect 2211 489 2287 527
rect 2211 455 2227 489
rect 2261 455 2287 489
rect 2211 421 2287 455
rect 2211 387 2227 421
rect 2261 387 2287 421
rect 2211 362 2287 387
rect 2321 449 2372 493
rect 2355 415 2372 449
rect 2321 381 2372 415
rect 2133 328 2167 347
rect 2355 347 2372 381
rect 2321 328 2372 347
rect 1945 294 2372 328
rect 1746 249 2288 255
rect 1746 215 1911 249
rect 1945 215 1989 249
rect 2023 215 2067 249
rect 2101 215 2145 249
rect 2179 215 2223 249
rect 2257 215 2288 249
rect 1746 211 2288 215
rect 1746 119 1796 211
rect 2322 177 2372 294
rect 1780 85 1796 119
rect 1945 143 2372 177
rect 1979 109 2005 143
rect 2355 109 2372 143
rect 1746 69 1796 85
rect 1838 93 1895 109
rect 1838 59 1851 93
rect 1885 59 1895 93
rect 1838 17 1895 59
rect 1945 53 2005 109
rect 2039 93 2099 109
rect 2073 59 2099 93
rect 2039 17 2099 59
rect 2133 53 2167 109
rect 2211 93 2287 109
rect 2211 59 2227 93
rect 2261 59 2287 93
rect 2211 17 2287 59
rect 2321 53 2372 109
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2392 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 133 348 167 382
rect 233 144 267 178
rect 529 348 563 382
rect 631 169 650 178
rect 650 169 665 178
rect 631 144 665 169
rect 856 153 890 187
rect 1141 348 1175 382
rect 1145 235 1146 256
rect 1146 235 1179 256
rect 1145 222 1179 235
rect 1501 179 1502 187
rect 1502 179 1535 187
rect 1501 153 1535 179
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
<< metal1 >>
rect 0 561 2392 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2392 561
rect 0 496 2392 527
rect 121 382 1187 388
rect 121 348 133 382
rect 167 360 529 382
rect 167 348 179 360
rect 121 342 179 348
rect 517 348 529 360
rect 563 360 1141 382
rect 563 348 575 360
rect 517 342 575 348
rect 1129 348 1141 360
rect 1175 348 1187 382
rect 1129 342 1187 348
rect 1133 256 1191 262
rect 1133 252 1145 256
rect 634 224 1145 252
rect 634 184 677 224
rect 1133 222 1145 224
rect 1179 222 1191 256
rect 1133 216 1191 222
rect 221 178 677 184
rect 221 144 233 178
rect 267 156 631 178
rect 267 144 279 156
rect 221 138 279 144
rect 619 144 631 156
rect 665 144 677 178
rect 844 187 902 193
rect 844 153 856 187
rect 890 184 902 187
rect 1489 187 1547 193
rect 1489 184 1501 187
rect 890 156 1501 184
rect 890 153 902 156
rect 844 147 902 153
rect 1489 153 1501 156
rect 1535 153 1547 187
rect 1489 147 1547 153
rect 619 138 677 144
rect 0 17 2392 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2392 17
rect 0 -48 2392 -17
<< labels >>
flabel corelocali s 2329 357 2363 391 0 FreeSans 400 0 0 0 Q
port 8 nsew
flabel corelocali s 2329 425 2363 459 0 FreeSans 400 0 0 0 Q
port 8 nsew
flabel corelocali s 2329 153 2363 187 0 FreeSans 400 0 0 0 Q
port 8 nsew
flabel corelocali s 2329 85 2363 119 0 FreeSans 400 0 0 0 Q
port 8 nsew
flabel corelocali s 2329 289 2363 323 0 FreeSans 400 0 0 0 Q
port 8 nsew
flabel corelocali s 2329 221 2363 255 0 FreeSans 400 0 0 0 Q
port 8 nsew
flabel corelocali s 397 289 431 323 0 FreeSans 200 0 0 0 D
port 2 nsew
flabel corelocali s 397 221 431 255 0 FreeSans 200 0 0 0 D
port 2 nsew
flabel corelocali s 29 527 63 561 3 FreeSans 400 0 0 0 VPWR
port 7 nsew
flabel corelocali s 1960 425 1994 459 0 FreeSans 400 0 0 0 Q
port 8 nsew
flabel corelocali s 1960 357 1994 391 0 FreeSans 400 0 0 0 Q
port 8 nsew
flabel corelocali s 1960 85 1994 119 0 FreeSans 400 0 0 0 Q
port 8 nsew
flabel corelocali s 29 289 63 323 0 FreeSans 400 0 0 0 CLK
port 1 nsew
flabel corelocali s 29 221 63 255 0 FreeSans 400 0 0 0 CLK
port 1 nsew
flabel corelocali s 29 -17 63 17 3 FreeSans 400 0 0 0 VGND
port 4 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel nbase s 46 544 46 544 3 FreeSans 400 0 0 0 VPB
port 6 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel pwell s 46 0 46 0 3 FreeSans 400 0 0 0 VNB
port 5 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 857 153 891 187 0 FreeSans 400 0 0 0 SET_B
port 3 nsew
rlabel comment s 0 0 0 0 4 dfstp_4
<< properties >>
string FIXED_BBOX 0 0 2392 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1928260
string GDS_START 1909802
<< end >>
