magic
tech sky130A
magscale 1 2
timestamp 1604502741
<< locali >>
rect 763 378 829 547
rect 25 236 96 310
rect 217 286 455 356
rect 505 344 829 378
rect 505 252 551 344
rect 130 218 551 252
rect 601 236 743 310
rect 793 236 935 310
rect 130 127 166 218
rect 517 202 551 218
rect 517 168 718 202
rect 592 66 718 168
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 21 364 71 649
rect 111 424 161 596
rect 201 458 267 649
rect 307 446 341 596
rect 381 480 447 649
rect 493 581 919 615
rect 493 480 559 581
rect 593 446 649 547
rect 307 424 649 446
rect 111 412 649 424
rect 689 412 723 581
rect 111 390 471 412
rect 111 364 161 390
rect 869 364 919 581
rect 30 85 96 202
rect 202 150 448 184
rect 202 85 252 150
rect 30 51 252 85
rect 288 66 362 116
rect 398 66 448 150
rect 288 17 322 66
rect 492 17 558 134
rect 752 17 818 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
rlabel locali s 25 236 96 310 6 A1
port 1 nsew signal input
rlabel locali s 217 286 455 356 6 A2
port 2 nsew signal input
rlabel locali s 601 236 743 310 6 B1
port 3 nsew signal input
rlabel locali s 793 236 935 310 6 C1
port 4 nsew signal input
rlabel locali s 763 378 829 547 6 Y
port 5 nsew signal output
rlabel locali s 592 66 718 168 6 Y
port 5 nsew signal output
rlabel locali s 517 202 551 218 6 Y
port 5 nsew signal output
rlabel locali s 517 168 718 202 6 Y
port 5 nsew signal output
rlabel locali s 505 344 829 378 6 Y
port 5 nsew signal output
rlabel locali s 505 252 551 344 6 Y
port 5 nsew signal output
rlabel locali s 130 218 551 252 6 Y
port 5 nsew signal output
rlabel locali s 130 127 166 218 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -49 960 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 960 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3814888
string GDS_START 3806206
<< end >>
