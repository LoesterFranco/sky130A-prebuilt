magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 131 47 161 131
rect 299 47 329 177
rect 393 47 423 177
rect 499 47 529 177
rect 571 47 601 177
rect 667 47 697 177
rect 763 47 793 177
<< pmoshvt >>
rect 82 378 118 462
rect 291 297 327 497
rect 385 297 421 497
rect 479 297 515 497
rect 573 297 609 497
rect 669 297 705 497
rect 765 297 801 497
<< ndiff >>
rect 186 161 299 177
rect 186 131 224 161
rect 61 106 131 131
rect 61 72 69 106
rect 103 72 131 106
rect 61 47 131 72
rect 161 127 224 131
rect 258 127 299 161
rect 161 93 299 127
rect 161 59 224 93
rect 258 59 299 93
rect 161 47 299 59
rect 329 169 393 177
rect 329 135 339 169
rect 373 135 393 169
rect 329 101 393 135
rect 329 67 339 101
rect 373 67 393 101
rect 329 47 393 67
rect 423 89 499 177
rect 423 55 444 89
rect 478 55 499 89
rect 423 47 499 55
rect 529 47 571 177
rect 601 157 667 177
rect 601 123 622 157
rect 656 123 667 157
rect 601 89 667 123
rect 601 55 622 89
rect 656 55 667 89
rect 601 47 667 55
rect 697 47 763 177
rect 793 157 860 177
rect 793 123 814 157
rect 848 123 860 157
rect 793 89 860 123
rect 793 55 814 89
rect 848 55 860 89
rect 793 47 860 55
<< pdiff >>
rect 228 477 291 497
rect 27 450 82 462
rect 27 416 35 450
rect 69 416 82 450
rect 27 378 82 416
rect 118 437 173 462
rect 118 403 131 437
rect 165 403 173 437
rect 118 378 173 403
rect 228 443 236 477
rect 270 443 291 477
rect 228 409 291 443
rect 228 375 236 409
rect 270 375 291 409
rect 228 297 291 375
rect 327 407 385 497
rect 327 373 339 407
rect 373 373 385 407
rect 327 339 385 373
rect 327 305 339 339
rect 373 305 385 339
rect 327 297 385 305
rect 421 489 479 497
rect 421 455 433 489
rect 467 455 479 489
rect 421 421 479 455
rect 421 387 433 421
rect 467 387 479 421
rect 421 297 479 387
rect 515 489 573 497
rect 515 455 527 489
rect 561 455 573 489
rect 515 297 573 455
rect 609 477 669 497
rect 609 443 622 477
rect 656 443 669 477
rect 609 405 669 443
rect 609 371 622 405
rect 656 371 669 405
rect 609 297 669 371
rect 705 489 765 497
rect 705 455 718 489
rect 752 455 765 489
rect 705 297 765 455
rect 801 477 860 497
rect 801 443 814 477
rect 848 443 860 477
rect 801 409 860 443
rect 801 375 814 409
rect 848 375 860 409
rect 801 297 860 375
<< ndiffc >>
rect 69 72 103 106
rect 224 127 258 161
rect 224 59 258 93
rect 339 135 373 169
rect 339 67 373 101
rect 444 55 478 89
rect 622 123 656 157
rect 622 55 656 89
rect 814 123 848 157
rect 814 55 848 89
<< pdiffc >>
rect 35 416 69 450
rect 131 403 165 437
rect 236 443 270 477
rect 236 375 270 409
rect 339 373 373 407
rect 339 305 373 339
rect 433 455 467 489
rect 433 387 467 421
rect 527 455 561 489
rect 622 443 656 477
rect 622 371 656 405
rect 718 455 752 489
rect 814 443 848 477
rect 814 375 848 409
<< poly >>
rect 291 497 327 523
rect 385 497 421 523
rect 479 497 515 523
rect 573 497 609 523
rect 669 497 705 523
rect 765 497 801 523
rect 82 462 118 488
rect 82 363 118 378
rect 80 287 120 363
rect 35 271 120 287
rect 291 282 327 297
rect 385 282 421 297
rect 479 282 515 297
rect 573 282 609 297
rect 669 282 705 297
rect 765 282 801 297
rect 35 237 51 271
rect 85 237 120 271
rect 289 265 329 282
rect 35 203 120 237
rect 35 169 51 203
rect 85 176 120 203
rect 211 261 329 265
rect 383 261 423 282
rect 477 265 517 282
rect 571 265 611 282
rect 667 265 707 282
rect 763 265 803 282
rect 211 249 423 261
rect 211 215 221 249
rect 255 215 423 249
rect 211 203 423 215
rect 211 199 329 203
rect 299 177 329 199
rect 393 177 423 203
rect 465 249 529 265
rect 465 215 475 249
rect 509 215 529 249
rect 465 199 529 215
rect 499 177 529 199
rect 571 249 713 265
rect 571 215 581 249
rect 615 215 659 249
rect 693 215 713 249
rect 571 199 713 215
rect 763 249 817 265
rect 763 215 773 249
rect 807 215 817 249
rect 763 199 817 215
rect 571 177 601 199
rect 667 177 697 199
rect 763 177 793 199
rect 85 169 161 176
rect 35 146 161 169
rect 131 131 161 146
rect 131 21 161 47
rect 299 21 329 47
rect 393 21 423 47
rect 499 21 529 47
rect 571 21 601 47
rect 667 21 697 47
rect 763 21 793 47
<< polycont >>
rect 51 237 85 271
rect 51 169 85 203
rect 221 215 255 249
rect 475 215 509 249
rect 581 215 615 249
rect 659 215 693 249
rect 773 215 807 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 19 450 85 527
rect 220 489 483 493
rect 220 477 433 489
rect 19 416 35 450
rect 69 416 85 450
rect 129 437 165 453
rect 129 403 131 437
rect 24 271 85 361
rect 24 237 51 271
rect 24 203 85 237
rect 24 169 51 203
rect 24 153 85 169
rect 129 257 165 403
rect 220 443 236 477
rect 270 457 433 477
rect 220 409 270 443
rect 407 455 433 457
rect 467 455 483 489
rect 220 375 236 409
rect 220 359 270 375
rect 305 407 373 423
rect 305 373 339 407
rect 305 339 373 373
rect 407 421 483 455
rect 527 489 561 527
rect 527 439 561 455
rect 622 477 656 493
rect 692 489 768 527
rect 692 455 718 489
rect 752 455 768 489
rect 812 477 864 493
rect 407 387 433 421
rect 467 405 483 421
rect 622 421 656 443
rect 812 443 814 477
rect 848 443 864 477
rect 812 421 864 443
rect 622 409 864 421
rect 622 405 814 409
rect 467 387 622 405
rect 407 371 622 387
rect 656 375 814 405
rect 848 375 864 409
rect 656 371 864 375
rect 305 305 339 339
rect 129 249 271 257
rect 129 215 221 249
rect 255 215 271 249
rect 129 214 271 215
rect 129 106 165 214
rect 53 72 69 106
rect 103 72 165 106
rect 217 161 265 177
rect 217 127 224 161
rect 258 127 265 161
rect 217 93 265 127
rect 217 59 224 93
rect 258 59 265 93
rect 217 17 265 59
rect 305 169 373 305
rect 460 299 817 335
rect 460 249 535 299
rect 459 215 475 249
rect 509 215 535 249
rect 571 249 713 265
rect 571 215 581 249
rect 615 215 659 249
rect 693 215 713 249
rect 571 199 713 215
rect 747 249 817 299
rect 747 215 773 249
rect 807 215 817 249
rect 747 199 817 215
rect 305 135 339 169
rect 373 135 622 157
rect 305 123 622 135
rect 656 123 672 157
rect 305 101 374 123
rect 305 67 339 101
rect 373 67 374 101
rect 596 89 672 123
rect 305 51 374 67
rect 428 55 444 89
rect 478 55 494 89
rect 428 17 494 55
rect 596 55 622 89
rect 656 55 672 89
rect 596 51 672 55
rect 798 123 814 157
rect 848 123 866 157
rect 798 89 866 123
rect 798 55 814 89
rect 848 55 866 89
rect 798 17 866 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel corelocali s 30 153 64 187 0 FreeSans 340 0 0 0 B1_N
port 3 nsew
flabel corelocali s 785 306 785 306 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 603 238 603 238 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 327 102 327 102 0 FreeSans 340 0 0 0 Y
port 8 nsew
rlabel comment s 0 0 0 0 4 a21boi_2
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1163918
string GDS_START 1156918
<< end >>
