magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1196 561
rect 103 448 169 527
rect 85 199 156 339
rect 190 199 247 265
rect 580 289 799 341
rect 1032 359 1074 527
rect 715 181 799 289
rect 833 215 992 255
rect 1026 215 1179 255
rect 127 17 161 165
rect 412 145 1090 181
rect 312 17 378 96
rect 412 51 478 145
rect 512 17 546 111
rect 580 51 646 145
rect 680 17 822 111
rect 856 51 922 145
rect 956 17 990 111
rect 1024 51 1090 145
rect 1124 17 1179 181
rect 0 -17 1196 17
<< obsli1 >>
rect 17 411 69 491
rect 328 459 730 493
rect 328 445 394 459
rect 496 443 730 459
rect 772 443 998 493
rect 17 377 383 411
rect 17 165 51 377
rect 199 305 315 343
rect 281 249 315 305
rect 349 317 383 377
rect 428 409 462 425
rect 428 375 922 409
rect 428 359 462 375
rect 349 283 546 317
rect 864 291 922 375
rect 956 325 998 443
rect 1108 325 1174 493
rect 956 291 1174 325
rect 512 255 546 283
rect 281 215 478 249
rect 512 215 681 255
rect 281 165 315 215
rect 17 90 93 165
rect 211 131 315 165
rect 211 90 250 131
<< metal1 >>
rect 0 496 1196 592
rect 0 -48 1196 48
<< labels >>
rlabel locali s 1026 215 1179 255 6 A
port 1 nsew signal input
rlabel locali s 833 215 992 255 6 B
port 2 nsew signal input
rlabel locali s 190 199 247 265 6 C_N
port 3 nsew signal input
rlabel locali s 85 199 156 339 6 D_N
port 4 nsew signal input
rlabel locali s 1024 51 1090 145 6 Y
port 5 nsew signal output
rlabel locali s 856 51 922 145 6 Y
port 5 nsew signal output
rlabel locali s 715 181 799 289 6 Y
port 5 nsew signal output
rlabel locali s 580 289 799 341 6 Y
port 5 nsew signal output
rlabel locali s 580 51 646 145 6 Y
port 5 nsew signal output
rlabel locali s 412 145 1090 181 6 Y
port 5 nsew signal output
rlabel locali s 412 51 478 145 6 Y
port 5 nsew signal output
rlabel locali s 1124 17 1179 181 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 956 17 990 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 680 17 822 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 512 17 546 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 312 17 378 96 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 127 17 161 165 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 1196 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1196 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1032 359 1074 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 103 448 169 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 1196 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 1196 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1206872
string GDS_START 1197548
<< end >>
