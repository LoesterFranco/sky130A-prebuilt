magic
tech sky130A
magscale 1 2
timestamp 1599588218
<< nwell >>
rect -38 332 1670 704
<< pwell >>
rect 0 0 1632 49
<< scpmos >>
rect 83 368 119 592
rect 173 368 209 592
rect 273 368 309 592
rect 363 368 399 592
rect 463 368 499 592
rect 553 368 589 592
rect 653 368 689 592
rect 743 368 779 592
rect 833 368 869 592
rect 923 368 959 592
rect 1017 368 1053 592
rect 1113 368 1149 592
rect 1223 368 1259 592
rect 1313 368 1349 592
rect 1423 368 1459 592
rect 1513 368 1549 592
<< nmoslvt >>
rect 98 74 128 222
rect 184 74 214 222
rect 284 74 314 222
rect 370 74 400 222
rect 470 74 500 222
rect 556 74 586 222
rect 656 74 686 222
rect 742 74 772 222
rect 828 74 858 222
rect 914 74 944 222
rect 1014 74 1044 222
rect 1100 74 1130 222
rect 1214 74 1244 222
rect 1300 74 1330 222
rect 1418 74 1448 222
rect 1504 74 1534 222
<< ndiff >>
rect 45 210 98 222
rect 45 176 53 210
rect 87 176 98 210
rect 45 120 98 176
rect 45 86 53 120
rect 87 86 98 120
rect 45 74 98 86
rect 128 210 184 222
rect 128 176 139 210
rect 173 176 184 210
rect 128 120 184 176
rect 128 86 139 120
rect 173 86 184 120
rect 128 74 184 86
rect 214 210 284 222
rect 214 176 239 210
rect 273 176 284 210
rect 214 120 284 176
rect 214 86 239 120
rect 273 86 284 120
rect 214 74 284 86
rect 314 210 370 222
rect 314 176 325 210
rect 359 176 370 210
rect 314 120 370 176
rect 314 86 325 120
rect 359 86 370 120
rect 314 74 370 86
rect 400 210 470 222
rect 400 176 411 210
rect 445 176 470 210
rect 400 120 470 176
rect 400 86 411 120
rect 445 86 470 120
rect 400 74 470 86
rect 500 210 556 222
rect 500 176 511 210
rect 545 176 556 210
rect 500 120 556 176
rect 500 86 511 120
rect 545 86 556 120
rect 500 74 556 86
rect 586 210 656 222
rect 586 176 607 210
rect 641 176 656 210
rect 586 120 656 176
rect 586 86 607 120
rect 641 86 656 120
rect 586 74 656 86
rect 686 210 742 222
rect 686 176 697 210
rect 731 176 742 210
rect 686 120 742 176
rect 686 86 697 120
rect 731 86 742 120
rect 686 74 742 86
rect 772 210 828 222
rect 772 176 783 210
rect 817 176 828 210
rect 772 120 828 176
rect 772 86 783 120
rect 817 86 828 120
rect 772 74 828 86
rect 858 210 914 222
rect 858 176 869 210
rect 903 176 914 210
rect 858 120 914 176
rect 858 86 869 120
rect 903 86 914 120
rect 858 74 914 86
rect 944 210 1014 222
rect 944 176 962 210
rect 996 176 1014 210
rect 944 123 1014 176
rect 944 89 962 123
rect 996 89 1014 123
rect 944 74 1014 89
rect 1044 210 1100 222
rect 1044 176 1055 210
rect 1089 176 1100 210
rect 1044 120 1100 176
rect 1044 86 1055 120
rect 1089 86 1100 120
rect 1044 74 1100 86
rect 1130 210 1214 222
rect 1130 176 1155 210
rect 1189 176 1214 210
rect 1130 123 1214 176
rect 1130 89 1155 123
rect 1189 89 1214 123
rect 1130 74 1214 89
rect 1244 210 1300 222
rect 1244 176 1255 210
rect 1289 176 1300 210
rect 1244 120 1300 176
rect 1244 86 1255 120
rect 1289 86 1300 120
rect 1244 74 1300 86
rect 1330 210 1418 222
rect 1330 176 1357 210
rect 1391 176 1418 210
rect 1330 123 1418 176
rect 1330 89 1357 123
rect 1391 89 1418 123
rect 1330 74 1418 89
rect 1448 210 1504 222
rect 1448 176 1459 210
rect 1493 176 1504 210
rect 1448 120 1504 176
rect 1448 86 1459 120
rect 1493 86 1504 120
rect 1448 74 1504 86
rect 1534 210 1587 222
rect 1534 176 1545 210
rect 1579 176 1587 210
rect 1534 120 1587 176
rect 1534 86 1545 120
rect 1579 86 1587 120
rect 1534 74 1587 86
<< pdiff >>
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 497 83 546
rect 27 463 39 497
rect 73 463 83 497
rect 27 414 83 463
rect 27 380 39 414
rect 73 380 83 414
rect 27 368 83 380
rect 119 580 173 592
rect 119 546 129 580
rect 163 546 173 580
rect 119 497 173 546
rect 119 463 129 497
rect 163 463 173 497
rect 119 414 173 463
rect 119 380 129 414
rect 163 380 173 414
rect 119 368 173 380
rect 209 580 273 592
rect 209 546 219 580
rect 253 546 273 580
rect 209 506 273 546
rect 209 472 219 506
rect 253 472 273 506
rect 209 438 273 472
rect 209 404 219 438
rect 253 404 273 438
rect 209 368 273 404
rect 309 580 363 592
rect 309 546 319 580
rect 353 546 363 580
rect 309 501 363 546
rect 309 467 319 501
rect 353 467 363 501
rect 309 422 363 467
rect 309 388 319 422
rect 353 388 363 422
rect 309 368 363 388
rect 399 580 463 592
rect 399 546 409 580
rect 443 546 463 580
rect 399 506 463 546
rect 399 472 409 506
rect 443 472 463 506
rect 399 438 463 472
rect 399 404 409 438
rect 443 404 463 438
rect 399 368 463 404
rect 499 580 553 592
rect 499 546 509 580
rect 543 546 553 580
rect 499 497 553 546
rect 499 463 509 497
rect 543 463 553 497
rect 499 414 553 463
rect 499 380 509 414
rect 543 380 553 414
rect 499 368 553 380
rect 589 580 653 592
rect 589 546 599 580
rect 633 546 653 580
rect 589 506 653 546
rect 589 472 599 506
rect 633 472 653 506
rect 589 438 653 472
rect 589 404 599 438
rect 633 404 653 438
rect 589 368 653 404
rect 689 580 743 592
rect 689 546 699 580
rect 733 546 743 580
rect 689 497 743 546
rect 689 463 699 497
rect 733 463 743 497
rect 689 414 743 463
rect 689 380 699 414
rect 733 380 743 414
rect 689 368 743 380
rect 779 580 833 592
rect 779 546 789 580
rect 823 546 833 580
rect 779 506 833 546
rect 779 472 789 506
rect 823 472 833 506
rect 779 438 833 472
rect 779 404 789 438
rect 823 404 833 438
rect 779 368 833 404
rect 869 580 923 592
rect 869 546 879 580
rect 913 546 923 580
rect 869 497 923 546
rect 869 463 879 497
rect 913 463 923 497
rect 869 414 923 463
rect 869 380 879 414
rect 913 380 923 414
rect 869 368 923 380
rect 959 580 1017 592
rect 959 546 969 580
rect 1003 546 1017 580
rect 959 506 1017 546
rect 959 472 969 506
rect 1003 472 1017 506
rect 959 438 1017 472
rect 959 404 969 438
rect 1003 404 1017 438
rect 959 368 1017 404
rect 1053 580 1113 592
rect 1053 546 1069 580
rect 1103 546 1113 580
rect 1053 497 1113 546
rect 1053 463 1069 497
rect 1103 463 1113 497
rect 1053 414 1113 463
rect 1053 380 1069 414
rect 1103 380 1113 414
rect 1053 368 1113 380
rect 1149 580 1223 592
rect 1149 546 1169 580
rect 1203 546 1223 580
rect 1149 506 1223 546
rect 1149 472 1169 506
rect 1203 472 1223 506
rect 1149 438 1223 472
rect 1149 404 1169 438
rect 1203 404 1223 438
rect 1149 368 1223 404
rect 1259 580 1313 592
rect 1259 546 1269 580
rect 1303 546 1313 580
rect 1259 497 1313 546
rect 1259 463 1269 497
rect 1303 463 1313 497
rect 1259 414 1313 463
rect 1259 380 1269 414
rect 1303 380 1313 414
rect 1259 368 1313 380
rect 1349 580 1423 592
rect 1349 546 1369 580
rect 1403 546 1423 580
rect 1349 506 1423 546
rect 1349 472 1369 506
rect 1403 472 1423 506
rect 1349 438 1423 472
rect 1349 404 1369 438
rect 1403 404 1423 438
rect 1349 368 1423 404
rect 1459 580 1513 592
rect 1459 546 1469 580
rect 1503 546 1513 580
rect 1459 497 1513 546
rect 1459 463 1469 497
rect 1503 463 1513 497
rect 1459 414 1513 463
rect 1459 380 1469 414
rect 1503 380 1513 414
rect 1459 368 1513 380
rect 1549 580 1605 592
rect 1549 546 1559 580
rect 1593 546 1605 580
rect 1549 497 1605 546
rect 1549 463 1559 497
rect 1593 463 1605 497
rect 1549 414 1605 463
rect 1549 380 1559 414
rect 1593 380 1605 414
rect 1549 368 1605 380
<< ndiffc >>
rect 53 176 87 210
rect 53 86 87 120
rect 139 176 173 210
rect 139 86 173 120
rect 239 176 273 210
rect 239 86 273 120
rect 325 176 359 210
rect 325 86 359 120
rect 411 176 445 210
rect 411 86 445 120
rect 511 176 545 210
rect 511 86 545 120
rect 607 176 641 210
rect 607 86 641 120
rect 697 176 731 210
rect 697 86 731 120
rect 783 176 817 210
rect 783 86 817 120
rect 869 176 903 210
rect 869 86 903 120
rect 962 176 996 210
rect 962 89 996 123
rect 1055 176 1089 210
rect 1055 86 1089 120
rect 1155 176 1189 210
rect 1155 89 1189 123
rect 1255 176 1289 210
rect 1255 86 1289 120
rect 1357 176 1391 210
rect 1357 89 1391 123
rect 1459 176 1493 210
rect 1459 86 1493 120
rect 1545 176 1579 210
rect 1545 86 1579 120
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 129 546 163 580
rect 129 463 163 497
rect 129 380 163 414
rect 219 546 253 580
rect 219 472 253 506
rect 219 404 253 438
rect 319 546 353 580
rect 319 467 353 501
rect 319 388 353 422
rect 409 546 443 580
rect 409 472 443 506
rect 409 404 443 438
rect 509 546 543 580
rect 509 463 543 497
rect 509 380 543 414
rect 599 546 633 580
rect 599 472 633 506
rect 599 404 633 438
rect 699 546 733 580
rect 699 463 733 497
rect 699 380 733 414
rect 789 546 823 580
rect 789 472 823 506
rect 789 404 823 438
rect 879 546 913 580
rect 879 463 913 497
rect 879 380 913 414
rect 969 546 1003 580
rect 969 472 1003 506
rect 969 404 1003 438
rect 1069 546 1103 580
rect 1069 463 1103 497
rect 1069 380 1103 414
rect 1169 546 1203 580
rect 1169 472 1203 506
rect 1169 404 1203 438
rect 1269 546 1303 580
rect 1269 463 1303 497
rect 1269 380 1303 414
rect 1369 546 1403 580
rect 1369 472 1403 506
rect 1369 404 1403 438
rect 1469 546 1503 580
rect 1469 463 1503 497
rect 1469 380 1503 414
rect 1559 546 1593 580
rect 1559 463 1593 497
rect 1559 380 1593 414
<< poly >>
rect 83 592 119 618
rect 173 592 209 618
rect 273 592 309 618
rect 363 592 399 618
rect 463 592 499 618
rect 553 592 589 618
rect 653 592 689 618
rect 743 592 779 618
rect 833 592 869 618
rect 923 592 959 618
rect 1017 592 1053 618
rect 1113 592 1149 618
rect 1223 592 1259 618
rect 1313 592 1349 618
rect 1423 592 1459 618
rect 1513 592 1549 618
rect 83 336 119 368
rect 173 336 209 368
rect 273 336 309 368
rect 363 336 399 368
rect 463 336 499 368
rect 553 336 589 368
rect 653 336 689 368
rect 743 336 779 368
rect 833 336 869 368
rect 923 336 959 368
rect 1017 336 1053 368
rect 1113 336 1149 368
rect 1223 336 1259 368
rect 1313 336 1349 368
rect 1423 336 1459 368
rect 1513 336 1549 368
rect 83 320 1549 336
rect 83 286 229 320
rect 263 286 417 320
rect 451 286 605 320
rect 639 286 788 320
rect 822 286 970 320
rect 1004 286 1169 320
rect 1203 286 1368 320
rect 1402 286 1549 320
rect 83 270 1549 286
rect 98 222 128 270
rect 184 222 214 270
rect 284 222 314 270
rect 370 222 400 270
rect 470 222 500 270
rect 556 222 586 270
rect 656 222 686 270
rect 742 222 772 270
rect 828 222 858 270
rect 914 222 944 270
rect 1014 222 1044 270
rect 1100 222 1130 270
rect 1214 222 1244 270
rect 1300 222 1330 270
rect 1418 222 1448 270
rect 1504 222 1534 270
rect 98 48 128 74
rect 184 48 214 74
rect 284 48 314 74
rect 370 48 400 74
rect 470 48 500 74
rect 556 48 586 74
rect 656 48 686 74
rect 742 48 772 74
rect 828 48 858 74
rect 914 48 944 74
rect 1014 48 1044 74
rect 1100 48 1130 74
rect 1214 48 1244 74
rect 1300 48 1330 74
rect 1418 48 1448 74
rect 1504 48 1534 74
<< polycont >>
rect 229 286 263 320
rect 417 286 451 320
rect 605 286 639 320
rect 788 286 822 320
rect 970 286 1004 320
rect 1169 286 1203 320
rect 1368 286 1402 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 23 580 73 649
rect 23 546 39 580
rect 23 497 73 546
rect 23 463 39 497
rect 23 414 73 463
rect 23 380 39 414
rect 23 364 73 380
rect 113 580 177 599
rect 113 546 129 580
rect 163 546 177 580
rect 113 497 177 546
rect 113 463 129 497
rect 163 463 177 497
rect 113 424 177 463
rect 113 380 129 424
rect 163 380 177 424
rect 211 580 269 649
rect 211 546 219 580
rect 253 546 269 580
rect 211 506 269 546
rect 211 472 219 506
rect 253 472 269 506
rect 211 438 269 472
rect 211 404 219 438
rect 253 404 269 438
rect 211 388 269 404
rect 303 580 369 596
rect 303 546 319 580
rect 353 546 369 580
rect 303 501 369 546
rect 303 467 319 501
rect 353 467 369 501
rect 303 424 369 467
rect 303 388 319 424
rect 353 388 369 424
rect 409 580 459 649
rect 443 546 459 580
rect 409 506 459 546
rect 443 472 459 506
rect 409 438 459 472
rect 443 404 459 438
rect 409 388 459 404
rect 493 580 559 596
rect 493 546 509 580
rect 543 546 559 580
rect 493 497 559 546
rect 493 463 509 497
rect 543 463 559 497
rect 493 424 559 463
rect 493 388 509 424
rect 113 266 177 380
rect 214 350 276 354
rect 214 286 229 350
rect 263 286 276 350
rect 214 270 276 286
rect 123 226 177 266
rect 37 210 89 226
rect 37 176 53 210
rect 87 176 89 210
rect 37 120 89 176
rect 37 86 53 120
rect 87 86 89 120
rect 37 17 89 86
rect 123 210 189 226
rect 123 176 139 210
rect 173 176 189 210
rect 123 120 189 176
rect 123 86 139 120
rect 173 86 189 120
rect 123 70 189 86
rect 223 210 275 226
rect 223 176 239 210
rect 273 176 275 210
rect 223 120 275 176
rect 223 86 239 120
rect 273 86 275 120
rect 223 17 275 86
rect 311 210 369 388
rect 497 380 509 388
rect 543 380 559 424
rect 599 580 649 649
rect 633 546 649 580
rect 599 506 649 546
rect 633 472 649 506
rect 599 438 649 472
rect 633 404 649 438
rect 599 388 649 404
rect 683 580 742 596
rect 683 546 699 580
rect 733 546 742 580
rect 683 497 742 546
rect 683 463 699 497
rect 733 463 742 497
rect 683 424 742 463
rect 404 350 462 354
rect 404 286 417 350
rect 451 286 462 350
rect 404 270 462 286
rect 311 176 325 210
rect 359 176 369 210
rect 311 120 369 176
rect 311 86 325 120
rect 359 86 369 120
rect 311 70 369 86
rect 405 210 461 226
rect 405 176 411 210
rect 445 176 461 210
rect 405 120 461 176
rect 405 86 411 120
rect 445 86 461 120
rect 405 17 461 86
rect 497 210 559 380
rect 683 380 699 424
rect 733 380 742 424
rect 783 580 830 649
rect 783 546 789 580
rect 823 546 830 580
rect 783 506 830 546
rect 783 472 789 506
rect 823 472 830 506
rect 783 438 830 472
rect 783 404 789 438
rect 823 404 830 438
rect 783 388 830 404
rect 868 580 926 596
rect 868 546 879 580
rect 913 546 926 580
rect 868 497 926 546
rect 868 463 879 497
rect 913 463 926 497
rect 868 424 926 463
rect 594 350 649 354
rect 594 286 605 350
rect 639 286 649 350
rect 594 270 649 286
rect 497 176 511 210
rect 545 176 559 210
rect 497 120 559 176
rect 497 86 511 120
rect 545 86 559 120
rect 497 70 559 86
rect 595 210 649 226
rect 595 176 607 210
rect 641 176 649 210
rect 595 120 649 176
rect 595 86 607 120
rect 641 86 649 120
rect 595 17 649 86
rect 683 210 742 380
rect 868 380 879 424
rect 913 388 926 424
rect 962 580 1019 649
rect 962 546 969 580
rect 1003 546 1019 580
rect 962 506 1019 546
rect 962 472 969 506
rect 1003 472 1019 506
rect 962 438 1019 472
rect 962 404 969 438
rect 1003 404 1019 438
rect 962 388 1019 404
rect 1053 580 1116 596
rect 1053 546 1069 580
rect 1103 546 1116 580
rect 1053 497 1116 546
rect 1053 463 1069 497
rect 1103 463 1116 497
rect 1053 424 1116 463
rect 913 380 919 388
rect 777 350 833 354
rect 777 286 788 350
rect 822 286 833 350
rect 777 270 833 286
rect 683 176 697 210
rect 731 176 742 210
rect 683 120 742 176
rect 683 86 697 120
rect 731 86 742 120
rect 683 70 742 86
rect 778 210 830 226
rect 778 176 783 210
rect 817 176 830 210
rect 778 120 830 176
rect 778 86 783 120
rect 817 86 830 120
rect 778 17 830 86
rect 868 210 919 380
rect 1053 380 1069 424
rect 1103 380 1116 424
rect 1153 580 1219 649
rect 1153 546 1169 580
rect 1203 546 1219 580
rect 1153 506 1219 546
rect 1153 472 1169 506
rect 1203 472 1219 506
rect 1153 438 1219 472
rect 1153 404 1169 438
rect 1203 404 1219 438
rect 1153 388 1219 404
rect 1253 580 1319 596
rect 1253 546 1269 580
rect 1303 546 1319 580
rect 1253 497 1319 546
rect 1253 463 1269 497
rect 1303 463 1319 497
rect 1253 424 1319 463
rect 954 350 1017 354
rect 954 286 970 350
rect 1004 286 1017 350
rect 954 270 1017 286
rect 1053 257 1116 380
rect 1253 380 1269 424
rect 1303 380 1319 424
rect 1353 580 1419 649
rect 1353 546 1369 580
rect 1403 546 1419 580
rect 1353 506 1419 546
rect 1353 472 1369 506
rect 1403 472 1419 506
rect 1353 438 1419 472
rect 1353 404 1369 438
rect 1403 404 1419 438
rect 1353 388 1419 404
rect 1453 580 1509 596
rect 1453 546 1469 580
rect 1503 546 1509 580
rect 1453 497 1509 546
rect 1453 463 1469 497
rect 1503 463 1509 497
rect 1453 424 1509 463
rect 1151 350 1218 354
rect 1151 286 1169 350
rect 1203 286 1218 350
rect 1151 270 1218 286
rect 1253 257 1319 380
rect 1453 380 1469 424
rect 1503 380 1509 424
rect 1354 350 1418 354
rect 1354 286 1368 350
rect 1402 286 1418 350
rect 1354 270 1418 286
rect 1053 236 1105 257
rect 1253 236 1305 257
rect 868 176 869 210
rect 903 176 919 210
rect 868 120 919 176
rect 868 86 869 120
rect 903 86 919 120
rect 868 70 919 86
rect 953 210 1005 226
rect 953 176 962 210
rect 996 176 1005 210
rect 953 123 1005 176
rect 953 89 962 123
rect 996 89 1005 123
rect 953 17 1005 89
rect 1043 210 1105 236
rect 1043 176 1055 210
rect 1089 176 1105 210
rect 1043 120 1105 176
rect 1043 86 1055 120
rect 1089 86 1105 120
rect 1043 70 1105 86
rect 1141 210 1205 226
rect 1141 176 1155 210
rect 1189 176 1205 210
rect 1141 123 1205 176
rect 1141 89 1155 123
rect 1189 89 1205 123
rect 1141 17 1205 89
rect 1239 210 1305 236
rect 1453 226 1509 380
rect 1547 580 1609 649
rect 1547 546 1559 580
rect 1593 546 1609 580
rect 1547 497 1609 546
rect 1547 463 1559 497
rect 1593 463 1609 497
rect 1547 414 1609 463
rect 1547 380 1559 414
rect 1593 380 1609 414
rect 1547 364 1609 380
rect 1239 176 1255 210
rect 1289 176 1305 210
rect 1239 120 1305 176
rect 1239 86 1255 120
rect 1289 86 1305 120
rect 1239 70 1305 86
rect 1341 210 1409 226
rect 1341 176 1357 210
rect 1391 176 1409 210
rect 1341 123 1409 176
rect 1341 89 1357 123
rect 1391 89 1409 123
rect 1341 17 1409 89
rect 1443 210 1509 226
rect 1443 176 1459 210
rect 1493 176 1509 210
rect 1443 120 1509 176
rect 1443 86 1459 120
rect 1493 86 1509 120
rect 1443 70 1509 86
rect 1543 210 1609 226
rect 1543 176 1545 210
rect 1579 176 1609 210
rect 1543 120 1609 176
rect 1543 86 1545 120
rect 1579 86 1609 120
rect 1543 17 1609 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 129 414 163 424
rect 129 390 163 414
rect 319 422 353 424
rect 319 390 353 422
rect 509 414 543 424
rect 509 390 543 414
rect 229 320 263 350
rect 229 316 263 320
rect 417 320 451 350
rect 417 316 451 320
rect 699 414 733 424
rect 699 390 733 414
rect 605 320 639 350
rect 605 316 639 320
rect 879 414 913 424
rect 879 390 913 414
rect 788 320 822 350
rect 788 316 822 320
rect 1069 414 1103 424
rect 1069 390 1103 414
rect 970 320 1004 350
rect 970 316 1004 320
rect 1269 414 1303 424
rect 1269 390 1303 414
rect 1169 320 1203 350
rect 1169 316 1203 320
rect 1469 414 1503 424
rect 1469 390 1503 414
rect 1368 320 1402 350
rect 1368 316 1402 320
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 117 424 1515 430
rect 117 390 129 424
rect 163 390 319 424
rect 353 390 509 424
rect 543 390 699 424
rect 733 390 879 424
rect 913 390 1069 424
rect 1103 390 1269 424
rect 1303 390 1469 424
rect 1503 390 1515 424
rect 117 384 1515 390
rect 217 350 1414 356
rect 217 316 229 350
rect 263 316 417 350
rect 451 316 605 350
rect 639 316 788 350
rect 822 316 970 350
rect 1004 316 1169 350
rect 1203 316 1368 350
rect 1402 316 1414 350
rect 217 310 1414 316
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew
flabel nwell s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew
rlabel comment s 0 0 0 0 4 inv_16
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew
flabel metal1 s 117 384 1515 430 0 FreeSans 400 0 0 0 Y
port 6 nsew
flabel metal1 s 217 310 1414 356 0 FreeSans 400 0 0 0 A
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 1632 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1803336
string GDS_START 1789728
<< end >>
