magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 1921 325 1971 425
rect 2109 325 2159 425
rect 2289 325 2367 425
rect 1921 291 2367 325
rect 101 215 575 257
rect 665 215 1139 257
rect 1333 215 1807 257
rect 1879 215 2217 257
rect 2289 181 2367 291
rect 117 145 2367 181
rect 117 51 183 145
rect 305 51 371 145
rect 493 51 559 145
rect 681 51 747 145
rect 869 51 935 145
rect 1057 51 1123 145
rect 1349 51 1415 145
rect 1537 51 1603 145
rect 1725 51 1791 145
rect 1913 51 1979 145
rect 2101 51 2167 145
rect 2289 51 2367 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2484 561
rect 23 325 81 493
rect 125 359 175 527
rect 219 325 269 493
rect 313 359 363 527
rect 407 325 457 493
rect 501 359 551 527
rect 595 459 1217 493
rect 595 325 645 459
rect 23 291 645 325
rect 689 325 739 425
rect 783 359 833 459
rect 877 325 927 425
rect 971 359 1021 459
rect 1065 325 1115 425
rect 1159 359 1217 459
rect 1255 459 2451 493
rect 1255 359 1313 459
rect 1357 325 1407 425
rect 1451 359 1501 459
rect 1545 325 1595 425
rect 1639 359 1689 459
rect 1733 325 1783 425
rect 689 291 1783 325
rect 1827 291 1877 459
rect 2015 359 2065 459
rect 2203 359 2253 459
rect 2401 291 2451 459
rect 23 17 83 181
rect 217 17 271 111
rect 405 17 459 111
rect 593 17 647 111
rect 781 17 835 111
rect 969 17 1023 111
rect 1157 17 1315 111
rect 1449 17 1503 111
rect 1637 17 1691 111
rect 1825 17 1879 111
rect 2013 17 2067 111
rect 2201 17 2255 111
rect 2401 17 2451 181
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2484 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
<< metal1 >>
rect 0 561 2484 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2484 561
rect 0 496 2484 527
rect 0 17 2484 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2484 17
rect 0 -48 2484 -17
<< labels >>
rlabel locali s 101 215 575 257 6 A
port 1 nsew signal input
rlabel locali s 665 215 1139 257 6 B
port 2 nsew signal input
rlabel locali s 1333 215 1807 257 6 C
port 3 nsew signal input
rlabel locali s 1879 215 2217 257 6 D
port 4 nsew signal input
rlabel locali s 2289 325 2367 425 6 Y
port 5 nsew signal output
rlabel locali s 2289 181 2367 291 6 Y
port 5 nsew signal output
rlabel locali s 2289 51 2367 145 6 Y
port 5 nsew signal output
rlabel locali s 2109 325 2159 425 6 Y
port 5 nsew signal output
rlabel locali s 2101 51 2167 145 6 Y
port 5 nsew signal output
rlabel locali s 1921 325 1971 425 6 Y
port 5 nsew signal output
rlabel locali s 1921 291 2367 325 6 Y
port 5 nsew signal output
rlabel locali s 1913 51 1979 145 6 Y
port 5 nsew signal output
rlabel locali s 1725 51 1791 145 6 Y
port 5 nsew signal output
rlabel locali s 1537 51 1603 145 6 Y
port 5 nsew signal output
rlabel locali s 1349 51 1415 145 6 Y
port 5 nsew signal output
rlabel locali s 1057 51 1123 145 6 Y
port 5 nsew signal output
rlabel locali s 869 51 935 145 6 Y
port 5 nsew signal output
rlabel locali s 681 51 747 145 6 Y
port 5 nsew signal output
rlabel locali s 493 51 559 145 6 Y
port 5 nsew signal output
rlabel locali s 305 51 371 145 6 Y
port 5 nsew signal output
rlabel locali s 117 145 2367 181 6 Y
port 5 nsew signal output
rlabel locali s 117 51 183 145 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -48 2484 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 2484 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2484 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3497046
string GDS_START 3479092
<< end >>
