magic
tech sky130A
magscale 1 2
timestamp 1601050047
<< nwell >>
rect -38 332 2918 704
<< pwell >>
rect 0 0 2880 49
<< scpmos >>
rect 84 368 114 592
rect 281 392 311 592
rect 383 392 413 592
rect 484 424 514 592
rect 697 424 727 592
rect 819 424 849 592
rect 1118 424 1148 592
rect 1316 368 1346 592
rect 1421 424 1451 592
rect 1659 424 1689 592
rect 1865 424 1895 592
rect 2022 424 2052 592
rect 2159 392 2189 592
rect 2293 392 2323 592
rect 2491 368 2521 592
rect 2581 368 2611 592
rect 2671 368 2701 592
rect 2763 368 2793 592
<< nmoslvt >>
rect 102 74 132 222
rect 350 105 380 233
rect 436 105 466 233
rect 522 105 552 233
rect 674 105 704 233
rect 874 105 904 233
rect 1043 105 1073 233
rect 1410 74 1440 222
rect 1505 79 1535 207
rect 1710 79 1740 207
rect 1876 79 1906 207
rect 2042 79 2072 207
rect 2156 79 2186 207
rect 2282 79 2312 207
rect 2492 74 2522 222
rect 2578 74 2608 222
rect 2678 74 2708 222
rect 2766 74 2796 222
<< ndiff >>
rect 42 149 102 222
rect 42 115 57 149
rect 91 115 102 149
rect 42 74 102 115
rect 132 207 185 222
rect 132 173 143 207
rect 177 173 185 207
rect 132 120 185 173
rect 132 86 143 120
rect 177 86 185 120
rect 279 220 350 233
rect 279 186 291 220
rect 325 186 350 220
rect 279 152 350 186
rect 279 118 291 152
rect 325 118 350 152
rect 279 105 350 118
rect 380 152 436 233
rect 380 118 391 152
rect 425 118 436 152
rect 380 105 436 118
rect 466 221 522 233
rect 466 187 477 221
rect 511 187 522 221
rect 466 151 522 187
rect 466 117 477 151
rect 511 117 522 151
rect 466 105 522 117
rect 552 221 674 233
rect 552 187 629 221
rect 663 187 674 221
rect 552 105 674 187
rect 704 221 874 233
rect 704 187 797 221
rect 831 187 874 221
rect 704 105 874 187
rect 904 221 1043 233
rect 904 187 969 221
rect 1003 187 1043 221
rect 904 105 1043 187
rect 1073 162 1123 233
rect 1073 150 1183 162
rect 1073 116 1137 150
rect 1171 116 1183 150
rect 1360 132 1410 222
rect 1073 105 1183 116
rect 1271 120 1410 132
rect 132 74 185 86
rect 1271 86 1283 120
rect 1317 86 1410 120
rect 1271 74 1410 86
rect 1440 207 1490 222
rect 1921 221 1979 233
rect 1921 207 1933 221
rect 1440 176 1505 207
rect 1440 142 1451 176
rect 1485 142 1505 176
rect 1440 79 1505 142
rect 1535 199 1710 207
rect 1535 165 1661 199
rect 1695 165 1710 199
rect 1535 121 1710 165
rect 1535 87 1619 121
rect 1653 87 1710 121
rect 1535 79 1710 87
rect 1740 195 1876 207
rect 1740 161 1765 195
rect 1799 161 1876 195
rect 1740 125 1876 161
rect 1740 91 1765 125
rect 1799 91 1876 125
rect 1740 79 1876 91
rect 1906 187 1933 207
rect 1967 207 1979 221
rect 1967 187 2042 207
rect 1906 79 2042 187
rect 2072 182 2156 207
rect 2072 148 2085 182
rect 2119 148 2156 182
rect 2072 79 2156 148
rect 2186 85 2282 207
rect 2186 79 2221 85
rect 1440 74 1490 79
rect 2209 51 2221 79
rect 2255 79 2282 85
rect 2312 195 2367 207
rect 2312 161 2323 195
rect 2357 161 2367 195
rect 2312 125 2367 161
rect 2312 91 2323 125
rect 2357 91 2367 125
rect 2312 79 2367 91
rect 2421 112 2492 222
rect 2255 51 2267 79
rect 2421 78 2431 112
rect 2465 78 2492 112
rect 2421 74 2492 78
rect 2522 210 2578 222
rect 2522 176 2533 210
rect 2567 176 2578 210
rect 2522 120 2578 176
rect 2522 86 2533 120
rect 2567 86 2578 120
rect 2522 74 2578 86
rect 2608 210 2678 222
rect 2608 176 2619 210
rect 2653 176 2678 210
rect 2608 120 2678 176
rect 2608 86 2619 120
rect 2653 86 2678 120
rect 2608 74 2678 86
rect 2708 210 2766 222
rect 2708 176 2720 210
rect 2754 176 2766 210
rect 2708 121 2766 176
rect 2708 87 2720 121
rect 2754 87 2766 121
rect 2708 74 2766 87
rect 2796 123 2853 222
rect 2796 89 2807 123
rect 2841 89 2853 123
rect 2796 74 2853 89
rect 2421 66 2477 74
rect 2209 39 2267 51
<< pdiff >>
rect 2207 622 2275 634
rect 2207 592 2224 622
rect 27 580 84 592
rect 27 546 37 580
rect 71 546 84 580
rect 27 482 84 546
rect 27 448 37 482
rect 71 448 84 482
rect 27 368 84 448
rect 114 580 170 592
rect 114 546 127 580
rect 161 546 170 580
rect 114 501 170 546
rect 114 467 127 501
rect 161 467 170 501
rect 114 414 170 467
rect 114 380 127 414
rect 161 380 170 414
rect 224 580 281 592
rect 224 546 234 580
rect 268 546 281 580
rect 224 509 281 546
rect 224 475 234 509
rect 268 475 281 509
rect 224 438 281 475
rect 224 404 234 438
rect 268 404 281 438
rect 224 392 281 404
rect 311 580 383 592
rect 311 546 324 580
rect 358 546 383 580
rect 311 510 383 546
rect 311 476 324 510
rect 358 476 383 510
rect 311 440 383 476
rect 311 406 324 440
rect 358 406 383 440
rect 311 392 383 406
rect 413 580 484 592
rect 413 546 427 580
rect 461 546 484 580
rect 413 466 484 546
rect 413 432 427 466
rect 461 432 484 466
rect 413 424 484 432
rect 514 528 697 592
rect 514 494 527 528
rect 561 494 640 528
rect 674 494 697 528
rect 514 424 697 494
rect 727 476 819 592
rect 727 442 756 476
rect 790 442 819 476
rect 727 424 819 442
rect 849 470 1118 592
rect 849 436 872 470
rect 906 436 993 470
rect 1027 436 1118 470
rect 849 424 1118 436
rect 1148 538 1205 592
rect 1148 504 1161 538
rect 1195 504 1205 538
rect 1148 424 1205 504
rect 1259 566 1316 592
rect 1259 532 1269 566
rect 1303 532 1316 566
rect 413 392 466 424
rect 114 368 170 380
rect 1259 368 1316 532
rect 1346 424 1421 592
rect 1451 544 1659 592
rect 1451 510 1527 544
rect 1561 510 1612 544
rect 1646 510 1659 544
rect 1451 466 1659 510
rect 1451 432 1527 466
rect 1561 432 1612 466
rect 1646 432 1659 466
rect 1451 424 1659 432
rect 1689 547 1865 592
rect 1689 513 1797 547
rect 1831 513 1865 547
rect 1689 466 1865 513
rect 1689 432 1797 466
rect 1831 432 1865 466
rect 1689 424 1865 432
rect 1895 580 2022 592
rect 1895 546 1965 580
rect 1999 546 2022 580
rect 1895 470 2022 546
rect 1895 436 1965 470
rect 1999 436 2022 470
rect 1895 424 2022 436
rect 2052 476 2159 592
rect 2052 442 2082 476
rect 2116 442 2159 476
rect 2052 424 2159 442
rect 1346 414 1403 424
rect 1346 380 1359 414
rect 1393 380 1403 414
rect 1346 368 1403 380
rect 2106 392 2159 424
rect 2189 588 2224 592
rect 2258 592 2275 622
rect 2258 588 2293 592
rect 2189 392 2293 588
rect 2323 440 2380 592
rect 2434 578 2491 592
rect 2434 544 2444 578
rect 2478 544 2491 578
rect 2434 530 2491 544
rect 2323 406 2336 440
rect 2370 406 2380 440
rect 2323 392 2380 406
rect 2438 368 2491 530
rect 2521 419 2581 592
rect 2521 385 2534 419
rect 2568 385 2581 419
rect 2521 368 2581 385
rect 2611 578 2671 592
rect 2611 544 2624 578
rect 2658 544 2671 578
rect 2611 368 2671 544
rect 2701 580 2763 592
rect 2701 546 2715 580
rect 2749 546 2763 580
rect 2701 497 2763 546
rect 2701 463 2715 497
rect 2749 463 2763 497
rect 2701 414 2763 463
rect 2701 380 2715 414
rect 2749 380 2763 414
rect 2701 368 2763 380
rect 2793 580 2853 592
rect 2793 546 2809 580
rect 2843 546 2853 580
rect 2793 497 2853 546
rect 2793 463 2809 497
rect 2843 463 2853 497
rect 2793 414 2853 463
rect 2793 380 2809 414
rect 2843 380 2853 414
rect 2793 368 2853 380
<< ndiffc >>
rect 57 115 91 149
rect 143 173 177 207
rect 143 86 177 120
rect 291 186 325 220
rect 291 118 325 152
rect 391 118 425 152
rect 477 187 511 221
rect 477 117 511 151
rect 629 187 663 221
rect 797 187 831 221
rect 969 187 1003 221
rect 1137 116 1171 150
rect 1283 86 1317 120
rect 1451 142 1485 176
rect 1661 165 1695 199
rect 1619 87 1653 121
rect 1765 161 1799 195
rect 1765 91 1799 125
rect 1933 187 1967 221
rect 2085 148 2119 182
rect 2221 51 2255 85
rect 2323 161 2357 195
rect 2323 91 2357 125
rect 2431 78 2465 112
rect 2533 176 2567 210
rect 2533 86 2567 120
rect 2619 176 2653 210
rect 2619 86 2653 120
rect 2720 176 2754 210
rect 2720 87 2754 121
rect 2807 89 2841 123
<< pdiffc >>
rect 37 546 71 580
rect 37 448 71 482
rect 127 546 161 580
rect 127 467 161 501
rect 127 380 161 414
rect 234 546 268 580
rect 234 475 268 509
rect 234 404 268 438
rect 324 546 358 580
rect 324 476 358 510
rect 324 406 358 440
rect 427 546 461 580
rect 427 432 461 466
rect 527 494 561 528
rect 640 494 674 528
rect 756 442 790 476
rect 872 436 906 470
rect 993 436 1027 470
rect 1161 504 1195 538
rect 1269 532 1303 566
rect 1527 510 1561 544
rect 1612 510 1646 544
rect 1527 432 1561 466
rect 1612 432 1646 466
rect 1797 513 1831 547
rect 1797 432 1831 466
rect 1965 546 1999 580
rect 1965 436 1999 470
rect 2082 442 2116 476
rect 1359 380 1393 414
rect 2224 588 2258 622
rect 2444 544 2478 578
rect 2336 406 2370 440
rect 2534 385 2568 419
rect 2624 544 2658 578
rect 2715 546 2749 580
rect 2715 463 2749 497
rect 2715 380 2749 414
rect 2809 546 2843 580
rect 2809 463 2843 497
rect 2809 380 2843 414
<< poly >>
rect 84 592 114 618
rect 281 592 311 618
rect 383 592 413 618
rect 484 592 514 618
rect 697 592 727 618
rect 819 592 849 618
rect 1118 592 1148 618
rect 1316 592 1346 618
rect 1421 592 1451 618
rect 1659 592 1689 618
rect 1865 592 1895 618
rect 2022 592 2052 618
rect 2159 592 2189 618
rect 484 409 514 424
rect 697 409 727 424
rect 819 409 849 424
rect 1118 409 1148 424
rect 281 377 311 392
rect 383 377 413 392
rect 481 379 646 409
rect 694 392 730 409
rect 816 399 852 409
rect 84 353 114 368
rect 81 326 117 353
rect 81 310 230 326
rect 81 276 180 310
rect 214 276 230 310
rect 81 260 230 276
rect 278 324 314 377
rect 380 324 416 377
rect 278 308 466 324
rect 278 274 366 308
rect 400 274 466 308
rect 102 222 132 260
rect 278 258 466 274
rect 508 321 574 337
rect 508 287 524 321
rect 558 287 574 321
rect 508 271 574 287
rect 616 278 646 379
rect 688 376 754 392
rect 688 342 704 376
rect 738 342 754 376
rect 688 326 754 342
rect 796 370 1073 399
rect 796 369 1023 370
rect 796 278 826 369
rect 1007 336 1023 369
rect 1057 336 1073 370
rect 1115 353 1151 409
rect 1421 409 1451 424
rect 1659 409 1689 424
rect 1865 409 1895 424
rect 2022 409 2052 424
rect 1418 392 1454 409
rect 1418 376 1501 392
rect 1656 389 1692 409
rect 1862 392 1898 409
rect 1316 353 1346 368
rect 350 233 380 258
rect 436 233 466 258
rect 522 233 552 271
rect 616 248 826 278
rect 868 305 934 321
rect 868 271 884 305
rect 918 271 934 305
rect 868 255 934 271
rect 674 233 704 248
rect 874 233 904 255
rect 1007 251 1073 336
rect 1121 323 1349 353
rect 1418 342 1451 376
rect 1485 342 1501 376
rect 1418 326 1501 342
rect 1543 373 1820 389
rect 1543 339 1559 373
rect 1593 359 1820 373
rect 1593 339 1609 359
rect 1043 233 1073 251
rect 1175 278 1349 323
rect 1543 305 1609 339
rect 1175 248 1440 278
rect 1543 271 1559 305
rect 1593 271 1609 305
rect 1543 255 1609 271
rect 1682 295 1748 311
rect 1682 261 1698 295
rect 1732 261 1748 295
rect 1543 252 1573 255
rect 1175 234 1241 248
rect 1175 200 1191 234
rect 1225 200 1241 234
rect 1410 222 1440 248
rect 1505 222 1573 252
rect 1682 245 1748 261
rect 1790 278 1820 359
rect 1862 376 1928 392
rect 1862 342 1878 376
rect 1912 342 1928 376
rect 1862 326 1928 342
rect 1970 379 2055 409
rect 2293 592 2323 618
rect 2491 592 2521 618
rect 2581 592 2611 618
rect 2671 592 2701 618
rect 2763 592 2793 618
rect 1970 278 2000 379
rect 2159 377 2189 392
rect 2293 377 2323 392
rect 2156 360 2192 377
rect 2156 344 2248 360
rect 1790 248 2000 278
rect 2042 321 2108 337
rect 2042 287 2058 321
rect 2092 287 2108 321
rect 2042 271 2108 287
rect 2156 310 2198 344
rect 2232 310 2248 344
rect 2156 294 2248 310
rect 2290 356 2326 377
rect 2290 340 2356 356
rect 2491 353 2521 368
rect 2581 353 2611 368
rect 2671 353 2701 368
rect 2763 353 2793 368
rect 2290 306 2306 340
rect 2340 306 2356 340
rect 2488 310 2524 353
rect 2578 310 2614 353
rect 2668 326 2704 353
rect 2760 326 2796 353
rect 1175 184 1241 200
rect 350 79 380 105
rect 436 79 466 105
rect 522 79 552 105
rect 674 79 704 105
rect 874 79 904 105
rect 1043 79 1073 105
rect 1505 207 1535 222
rect 1710 207 1740 245
rect 1876 207 1906 248
rect 2042 207 2072 271
rect 2156 207 2186 294
rect 2290 290 2356 306
rect 2417 294 2614 310
rect 2290 252 2320 290
rect 2282 222 2320 252
rect 2417 260 2433 294
rect 2467 260 2614 294
rect 2656 310 2796 326
rect 2656 276 2672 310
rect 2706 276 2796 310
rect 2656 260 2796 276
rect 2417 244 2614 260
rect 2492 222 2522 244
rect 2578 222 2608 244
rect 2678 222 2708 260
rect 2766 222 2796 260
rect 2282 207 2312 222
rect 102 48 132 74
rect 1410 48 1440 74
rect 1505 53 1535 79
rect 1710 53 1740 79
rect 1876 53 1906 79
rect 2042 53 2072 79
rect 2156 53 2186 79
rect 2282 53 2312 79
rect 2492 48 2522 74
rect 2578 48 2608 74
rect 2678 48 2708 74
rect 2766 48 2796 74
<< polycont >>
rect 180 276 214 310
rect 366 274 400 308
rect 524 287 558 321
rect 704 342 738 376
rect 1023 336 1057 370
rect 884 271 918 305
rect 1451 342 1485 376
rect 1559 339 1593 373
rect 1559 271 1593 305
rect 1698 261 1732 295
rect 1191 200 1225 234
rect 1878 342 1912 376
rect 2058 287 2092 321
rect 2198 310 2232 344
rect 2306 306 2340 340
rect 2433 260 2467 294
rect 2672 276 2706 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2880 683
rect 21 580 72 649
rect 21 546 37 580
rect 71 546 72 580
rect 21 482 72 546
rect 21 448 37 482
rect 71 448 72 482
rect 21 432 72 448
rect 111 580 177 596
rect 111 546 127 580
rect 161 546 177 580
rect 111 501 177 546
rect 111 467 127 501
rect 161 467 177 501
rect 111 414 177 467
rect 111 398 127 414
rect 67 380 127 398
rect 161 380 177 414
rect 67 364 177 380
rect 218 580 268 596
rect 218 546 234 580
rect 218 509 268 546
rect 218 475 234 509
rect 218 438 268 475
rect 218 404 234 438
rect 67 294 130 364
rect 218 326 268 404
rect 308 580 374 649
rect 308 546 324 580
rect 358 546 374 580
rect 308 510 374 546
rect 308 476 324 510
rect 358 476 374 510
rect 308 440 374 476
rect 308 406 324 440
rect 358 406 374 440
rect 308 390 374 406
rect 411 580 1211 612
rect 411 546 427 580
rect 461 578 1211 580
rect 461 546 477 578
rect 411 466 477 546
rect 511 528 1111 544
rect 511 494 527 528
rect 561 494 640 528
rect 674 510 1111 528
rect 674 494 690 510
rect 511 478 690 494
rect 411 432 427 466
rect 461 432 477 466
rect 411 403 477 432
rect 25 276 130 294
rect 25 242 31 276
rect 65 242 130 276
rect 164 310 279 326
rect 164 276 180 310
rect 214 276 279 310
rect 164 260 279 276
rect 25 236 130 242
rect 96 226 130 236
rect 96 207 193 226
rect 96 192 143 207
rect 141 173 143 192
rect 177 173 193 207
rect 34 149 107 158
rect 34 115 57 149
rect 91 115 107 149
rect 34 17 107 115
rect 141 120 193 173
rect 141 86 143 120
rect 177 86 193 120
rect 245 224 279 260
rect 313 308 409 356
rect 313 274 366 308
rect 400 274 409 308
rect 313 258 409 274
rect 443 237 477 403
rect 511 321 579 430
rect 511 287 524 321
rect 558 287 579 321
rect 511 271 579 287
rect 245 220 341 224
rect 245 186 291 220
rect 325 186 341 220
rect 443 221 511 237
rect 443 203 477 221
rect 245 152 341 186
rect 461 187 477 203
rect 245 118 291 152
rect 325 118 341 152
rect 245 101 341 118
rect 375 152 425 169
rect 375 118 391 152
rect 141 70 193 86
rect 375 17 425 118
rect 461 151 511 187
rect 461 117 477 151
rect 545 153 579 271
rect 613 237 647 478
rect 724 442 756 476
rect 790 442 822 476
rect 724 426 822 442
rect 688 376 754 392
rect 688 342 704 376
rect 738 342 754 376
rect 688 326 754 342
rect 613 221 679 237
rect 613 187 629 221
rect 663 187 679 221
rect 713 153 747 326
rect 788 282 822 426
rect 856 436 872 470
rect 906 436 993 470
rect 1027 436 1043 470
rect 856 420 1043 436
rect 1077 454 1111 510
rect 1145 538 1211 578
rect 1145 504 1161 538
rect 1195 504 1211 538
rect 1253 566 1319 649
rect 2203 622 2279 649
rect 1253 532 1269 566
rect 1303 532 1319 566
rect 1253 516 1319 532
rect 1443 581 1915 615
rect 1145 488 1211 504
rect 1443 482 1477 581
rect 1245 454 1477 482
rect 1077 448 1477 454
rect 1077 420 1279 448
rect 881 305 919 321
rect 788 276 847 282
rect 788 242 799 276
rect 833 242 847 276
rect 788 237 847 242
rect 781 221 847 237
rect 781 187 797 221
rect 831 187 847 221
rect 881 271 884 305
rect 918 271 919 305
rect 881 153 919 271
rect 953 286 987 420
rect 1343 386 1359 414
rect 1021 380 1359 386
rect 1393 380 1409 414
rect 1021 370 1409 380
rect 1021 336 1023 370
rect 1057 352 1409 370
rect 1057 336 1073 352
rect 1021 320 1073 336
rect 1107 286 1309 305
rect 953 271 1309 286
rect 953 252 1141 271
rect 953 221 1019 252
rect 953 187 969 221
rect 1003 187 1019 221
rect 1175 234 1241 237
rect 1175 218 1191 234
rect 1053 200 1191 218
rect 1225 200 1241 234
rect 1053 184 1241 200
rect 1275 204 1309 271
rect 1343 272 1409 352
rect 1443 392 1477 448
rect 1511 544 1662 547
rect 1511 510 1527 544
rect 1561 510 1612 544
rect 1646 510 1662 544
rect 1511 466 1662 510
rect 1511 432 1527 466
rect 1561 432 1612 466
rect 1646 432 1662 466
rect 1511 426 1662 432
rect 1443 376 1501 392
rect 1443 342 1451 376
rect 1485 342 1501 376
rect 1443 326 1501 342
rect 1535 373 1594 389
rect 1535 339 1559 373
rect 1593 339 1594 373
rect 1535 305 1594 339
rect 1343 238 1501 272
rect 1053 153 1087 184
rect 1275 170 1401 204
rect 545 119 1087 153
rect 461 85 511 117
rect 1121 116 1137 150
rect 1171 116 1187 150
rect 1121 85 1187 116
rect 461 51 1187 85
rect 1267 120 1333 136
rect 1267 86 1283 120
rect 1317 86 1333 120
rect 1267 17 1333 86
rect 1367 85 1401 170
rect 1435 176 1501 238
rect 1435 142 1451 176
rect 1485 142 1501 176
rect 1435 126 1501 142
rect 1535 271 1559 305
rect 1593 271 1594 305
rect 1535 255 1594 271
rect 1535 85 1569 255
rect 1628 208 1662 426
rect 1696 295 1747 581
rect 1696 261 1698 295
rect 1732 261 1747 295
rect 1696 245 1747 261
rect 1781 513 1797 547
rect 1831 513 1847 547
rect 1781 466 1847 513
rect 1781 432 1797 466
rect 1831 432 1847 466
rect 1781 426 1847 432
rect 1781 211 1815 426
rect 1881 392 1915 581
rect 1628 202 1711 208
rect 1628 199 1663 202
rect 1628 165 1661 199
rect 1697 168 1711 202
rect 1695 165 1711 168
rect 1628 128 1711 165
rect 1367 51 1569 85
rect 1603 121 1711 128
rect 1603 87 1619 121
rect 1653 87 1711 121
rect 1603 78 1711 87
rect 1749 195 1815 211
rect 1749 161 1765 195
rect 1799 161 1815 195
rect 1749 125 1815 161
rect 1749 91 1765 125
rect 1799 91 1815 125
rect 1849 376 1915 392
rect 1849 342 1878 376
rect 1912 342 1915 376
rect 1849 326 1915 342
rect 1949 580 2015 596
rect 2203 588 2224 622
rect 2258 588 2279 622
rect 1949 546 1965 580
rect 1999 554 2015 580
rect 2428 578 2494 649
rect 1999 546 2394 554
rect 1949 520 2394 546
rect 2428 544 2444 578
rect 2478 544 2494 578
rect 2428 542 2494 544
rect 2608 578 2674 649
rect 2608 544 2624 578
rect 2658 544 2674 578
rect 2608 542 2674 544
rect 2714 580 2775 596
rect 2714 546 2715 580
rect 2749 546 2775 580
rect 1949 470 2015 520
rect 2360 508 2394 520
rect 1949 436 1965 470
rect 1999 436 2015 470
rect 1949 420 2015 436
rect 2062 476 2162 486
rect 2062 442 2082 476
rect 2116 442 2162 476
rect 2360 474 2680 508
rect 2062 426 2162 442
rect 1849 153 1883 326
rect 1949 237 1983 420
rect 1917 221 1983 237
rect 1917 187 1933 221
rect 1967 187 1983 221
rect 2017 321 2094 337
rect 2017 287 2058 321
rect 2092 287 2094 321
rect 2017 271 2094 287
rect 2017 153 2051 271
rect 2128 237 2162 426
rect 1849 119 2051 153
rect 2085 203 2162 237
rect 2196 406 2336 440
rect 2370 406 2386 440
rect 2196 390 2386 406
rect 2517 419 2584 440
rect 2196 344 2248 390
rect 2517 385 2534 419
rect 2568 385 2584 419
rect 2196 310 2198 344
rect 2232 310 2248 344
rect 2196 211 2248 310
rect 2290 340 2375 356
rect 2290 306 2306 340
rect 2340 306 2375 340
rect 2517 310 2584 385
rect 2646 326 2680 474
rect 2714 497 2775 546
rect 2714 463 2715 497
rect 2749 463 2775 497
rect 2714 414 2775 463
rect 2714 380 2715 414
rect 2749 380 2775 414
rect 2714 364 2775 380
rect 2809 580 2859 649
rect 2843 546 2859 580
rect 2809 497 2859 546
rect 2843 463 2859 497
rect 2809 414 2859 463
rect 2843 380 2859 414
rect 2809 364 2859 380
rect 2646 310 2707 326
rect 2290 290 2375 306
rect 2417 294 2483 310
rect 2417 260 2433 294
rect 2467 260 2483 294
rect 2085 182 2119 203
rect 2196 195 2373 211
rect 2196 169 2323 195
rect 2085 119 2119 148
rect 2153 161 2323 169
rect 2357 161 2373 195
rect 2417 202 2483 260
rect 2417 168 2431 202
rect 2465 168 2483 202
rect 2417 162 2483 168
rect 2517 210 2567 310
rect 2646 276 2672 310
rect 2706 276 2707 310
rect 2646 260 2707 276
rect 2741 301 2775 364
rect 2741 226 2855 301
rect 2517 176 2533 210
rect 2153 135 2373 161
rect 1749 85 1815 91
rect 2153 85 2187 135
rect 2307 125 2373 135
rect 1749 51 2187 85
rect 2221 85 2271 101
rect 2255 51 2271 85
rect 2307 91 2323 125
rect 2357 91 2373 125
rect 2307 75 2373 91
rect 2415 112 2481 128
rect 2415 78 2431 112
rect 2465 78 2481 112
rect 2221 17 2271 51
rect 2415 17 2481 78
rect 2517 120 2567 176
rect 2517 86 2533 120
rect 2517 70 2567 86
rect 2603 210 2669 226
rect 2603 176 2619 210
rect 2653 176 2669 210
rect 2603 120 2669 176
rect 2603 86 2619 120
rect 2653 86 2669 120
rect 2603 17 2669 86
rect 2703 210 2855 226
rect 2703 176 2720 210
rect 2754 176 2855 210
rect 2703 160 2855 176
rect 2703 121 2757 160
rect 2703 87 2720 121
rect 2754 87 2757 121
rect 2703 71 2757 87
rect 2791 123 2857 126
rect 2791 89 2807 123
rect 2841 89 2857 123
rect 2791 17 2857 89
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2880 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 31 242 65 276
rect 799 242 833 276
rect 1663 199 1697 202
rect 1663 168 1695 199
rect 1695 168 1697 199
rect 2431 168 2465 202
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
<< metal1 >>
rect 0 683 2880 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2880 683
rect 0 617 2880 649
rect 19 276 77 282
rect 19 242 31 276
rect 65 273 77 276
rect 787 276 845 282
rect 787 273 799 276
rect 65 245 799 273
rect 65 242 77 245
rect 19 236 77 242
rect 787 242 799 245
rect 833 242 845 276
rect 787 236 845 242
rect 1651 202 1709 208
rect 1651 168 1663 202
rect 1697 199 1709 202
rect 2419 202 2477 208
rect 2419 199 2431 202
rect 1697 171 2431 199
rect 1697 168 1709 171
rect 1651 162 1709 168
rect 2419 168 2431 171
rect 2465 168 2477 202
rect 2419 162 2477 168
rect 0 17 2880 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2880 17
rect 0 -49 2880 -17
<< labels >>
rlabel comment s 0 0 0 0 4 fah_2
flabel pwell s 0 0 2880 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 2880 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 2880 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 2880 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 2335 316 2369 350 0 FreeSans 340 0 0 0 CI
port 3 nsew
flabel corelocali s 2815 168 2849 202 0 FreeSans 340 0 0 0 SUM
port 9 nsew
flabel corelocali s 2815 242 2849 276 0 FreeSans 340 0 0 0 SUM
port 9 nsew
flabel corelocali s 2527 316 2561 350 0 FreeSans 340 0 0 0 COUT
port 8 nsew
flabel corelocali s 2527 390 2561 424 0 FreeSans 340 0 0 0 COUT
port 8 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 511 390 545 424 0 FreeSans 340 0 0 0 B
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 2880 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 2552342
string GDS_START 2532674
<< end >>
