magic
tech sky130A
magscale 1 2
timestamp 1599588244
<< locali >>
rect 25 224 110 358
rect 871 364 942 596
rect 212 224 278 352
rect 313 236 386 352
rect 444 224 551 358
rect 585 224 651 304
rect 697 224 765 309
rect 908 226 942 364
rect 871 70 942 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 23 581 518 615
rect 23 392 89 581
rect 144 386 210 547
rect 244 386 310 581
rect 344 426 410 547
rect 452 460 518 581
rect 564 460 630 649
rect 664 426 730 587
rect 344 392 730 426
rect 344 386 410 392
rect 144 190 178 386
rect 664 379 730 392
rect 771 379 837 649
rect 803 260 874 326
rect 803 190 837 260
rect 28 156 837 190
rect 28 70 94 156
rect 192 17 361 120
rect 459 66 626 156
rect 724 17 837 122
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
rlabel locali s 585 224 651 304 6 A1
port 1 nsew signal input
rlabel locali s 697 224 765 309 6 A2
port 2 nsew signal input
rlabel locali s 444 224 551 358 6 B1
port 3 nsew signal input
rlabel locali s 313 236 386 352 6 B2
port 4 nsew signal input
rlabel locali s 25 224 110 358 6 C1
port 5 nsew signal input
rlabel locali s 212 224 278 352 6 C2
port 6 nsew signal input
rlabel locali s 908 226 942 364 6 X
port 7 nsew signal output
rlabel locali s 871 364 942 596 6 X
port 7 nsew signal output
rlabel locali s 871 70 942 226 6 X
port 7 nsew signal output
rlabel metal1 s 0 -49 960 49 8 VGND
port 8 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 9 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 10 nsew power bidirectional
rlabel metal1 s 0 617 960 715 6 VPWR
port 11 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3479230
string GDS_START 3470454
<< end >>
