magic
tech sky130A
magscale 1 2
timestamp 1604502693
<< nwell >>
rect -38 261 1602 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 351 47 381 131
rect 458 47 488 119
rect 545 47 575 119
rect 640 47 670 131
rect 828 47 858 177
rect 1016 47 1046 177
rect 1100 47 1130 177
rect 1184 47 1214 177
rect 1286 47 1316 177
rect 1370 47 1400 177
rect 1454 47 1484 177
<< pmoshvt >>
rect 79 363 109 491
rect 163 363 193 491
rect 351 369 381 497
rect 447 413 477 497
rect 555 413 585 497
rect 627 413 657 497
rect 823 297 853 497
rect 923 297 953 497
rect 1088 297 1118 497
rect 1184 297 1214 497
rect 1286 297 1316 497
rect 1370 297 1400 497
rect 1454 297 1484 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 299 93 351 131
rect 299 59 307 93
rect 341 59 351 93
rect 299 47 351 59
rect 381 119 431 131
rect 776 133 828 177
rect 590 119 640 131
rect 381 47 458 119
rect 488 107 545 119
rect 488 73 499 107
rect 533 73 545 107
rect 488 47 545 73
rect 575 47 640 119
rect 670 106 722 131
rect 670 72 680 106
rect 714 72 722 106
rect 670 47 722 72
rect 776 99 784 133
rect 818 99 828 133
rect 776 47 828 99
rect 858 107 910 177
rect 858 73 868 107
rect 902 73 910 107
rect 858 47 910 73
rect 964 108 1016 177
rect 964 74 972 108
rect 1006 74 1016 108
rect 964 47 1016 74
rect 1046 47 1100 177
rect 1130 93 1184 177
rect 1130 59 1140 93
rect 1174 59 1184 93
rect 1130 47 1184 59
rect 1214 101 1286 177
rect 1214 67 1224 101
rect 1258 67 1286 101
rect 1214 47 1286 67
rect 1316 93 1370 177
rect 1316 59 1326 93
rect 1360 59 1370 93
rect 1316 47 1370 59
rect 1400 161 1454 177
rect 1400 127 1410 161
rect 1444 127 1454 161
rect 1400 93 1454 127
rect 1400 59 1410 93
rect 1444 59 1454 93
rect 1400 47 1454 59
rect 1484 161 1536 177
rect 1484 127 1494 161
rect 1528 127 1536 161
rect 1484 93 1536 127
rect 1484 59 1494 93
rect 1528 59 1536 93
rect 1484 47 1536 59
<< pdiff >>
rect 27 477 79 491
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 363 79 375
rect 109 461 163 491
rect 109 427 119 461
rect 153 427 163 461
rect 109 363 163 427
rect 193 477 245 491
rect 193 443 203 477
rect 237 443 245 477
rect 193 409 245 443
rect 193 375 203 409
rect 237 375 245 409
rect 193 363 245 375
rect 299 485 351 497
rect 299 451 307 485
rect 341 451 351 485
rect 299 369 351 451
rect 381 413 447 497
rect 477 473 555 497
rect 477 439 511 473
rect 545 439 555 473
rect 477 413 555 439
rect 585 413 627 497
rect 657 485 709 497
rect 657 451 667 485
rect 701 451 709 485
rect 657 413 709 451
rect 771 471 823 497
rect 771 437 779 471
rect 813 437 823 471
rect 381 369 431 413
rect 771 368 823 437
rect 771 334 779 368
rect 813 334 823 368
rect 771 297 823 334
rect 853 471 923 497
rect 853 437 866 471
rect 900 437 923 471
rect 853 297 923 437
rect 953 477 1088 497
rect 953 443 973 477
rect 1007 443 1088 477
rect 953 409 1088 443
rect 953 375 973 409
rect 1007 375 1088 409
rect 953 341 1088 375
rect 953 307 973 341
rect 1007 307 1088 341
rect 953 297 1088 307
rect 1118 485 1184 497
rect 1118 451 1134 485
rect 1168 451 1184 485
rect 1118 417 1184 451
rect 1118 383 1134 417
rect 1168 383 1184 417
rect 1118 297 1184 383
rect 1214 475 1286 497
rect 1214 441 1224 475
rect 1258 441 1286 475
rect 1214 297 1286 441
rect 1316 485 1370 497
rect 1316 451 1326 485
rect 1360 451 1370 485
rect 1316 297 1370 451
rect 1400 485 1454 497
rect 1400 451 1410 485
rect 1444 451 1454 485
rect 1400 417 1454 451
rect 1400 383 1410 417
rect 1444 383 1454 417
rect 1400 349 1454 383
rect 1400 315 1410 349
rect 1444 315 1454 349
rect 1400 297 1454 315
rect 1484 485 1536 497
rect 1484 451 1494 485
rect 1528 451 1536 485
rect 1484 417 1536 451
rect 1484 383 1494 417
rect 1528 383 1536 417
rect 1484 349 1536 383
rect 1484 315 1494 349
rect 1528 315 1536 349
rect 1484 297 1536 315
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 307 59 341 93
rect 499 73 533 107
rect 680 72 714 106
rect 784 99 818 133
rect 868 73 902 107
rect 972 74 1006 108
rect 1140 59 1174 93
rect 1224 67 1258 101
rect 1326 59 1360 93
rect 1410 127 1444 161
rect 1410 59 1444 93
rect 1494 127 1528 161
rect 1494 59 1528 93
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 427 153 461
rect 203 443 237 477
rect 203 375 237 409
rect 307 451 341 485
rect 511 439 545 473
rect 667 451 701 485
rect 779 437 813 471
rect 779 334 813 368
rect 866 437 900 471
rect 973 443 1007 477
rect 973 375 1007 409
rect 973 307 1007 341
rect 1134 451 1168 485
rect 1134 383 1168 417
rect 1224 441 1258 475
rect 1326 451 1360 485
rect 1410 451 1444 485
rect 1410 383 1444 417
rect 1410 315 1444 349
rect 1494 451 1528 485
rect 1494 383 1528 417
rect 1494 315 1528 349
<< poly >>
rect 79 491 109 517
rect 163 491 193 517
rect 351 497 381 523
rect 447 497 477 523
rect 555 497 585 523
rect 627 497 657 523
rect 823 497 853 523
rect 923 497 953 523
rect 1088 497 1118 523
rect 1184 497 1214 523
rect 1286 497 1316 523
rect 1370 497 1400 523
rect 1454 497 1484 523
rect 79 348 109 363
rect 46 318 109 348
rect 46 280 76 318
rect 21 264 76 280
rect 163 274 193 363
rect 21 230 32 264
rect 66 230 76 264
rect 21 214 76 230
rect 118 264 193 274
rect 118 230 134 264
rect 168 230 193 264
rect 118 220 193 230
rect 46 176 76 214
rect 46 146 109 176
rect 79 131 109 146
rect 163 131 193 220
rect 351 219 381 369
rect 447 337 477 413
rect 555 375 585 413
rect 423 321 477 337
rect 519 365 585 375
rect 519 331 535 365
rect 569 331 585 365
rect 519 321 585 331
rect 627 373 657 413
rect 627 357 715 373
rect 627 323 671 357
rect 705 323 715 357
rect 423 287 433 321
rect 467 287 477 321
rect 423 279 477 287
rect 627 307 715 323
rect 423 249 575 279
rect 324 203 390 219
rect 324 169 340 203
rect 374 169 390 203
rect 324 153 390 169
rect 448 191 503 207
rect 448 157 459 191
rect 493 157 503 191
rect 324 152 381 153
rect 351 131 381 152
rect 448 141 503 157
rect 458 119 488 141
rect 545 119 575 249
rect 627 183 657 307
rect 823 265 853 297
rect 923 265 953 297
rect 1088 265 1118 297
rect 1184 265 1214 297
rect 1286 265 1316 297
rect 1370 265 1400 297
rect 1454 265 1484 297
rect 711 249 858 265
rect 711 215 721 249
rect 755 215 858 249
rect 711 199 858 215
rect 900 249 954 265
rect 900 215 910 249
rect 944 222 954 249
rect 1088 249 1142 265
rect 944 215 1046 222
rect 900 199 1046 215
rect 1088 215 1098 249
rect 1132 215 1142 249
rect 1088 199 1142 215
rect 1184 249 1484 265
rect 1184 215 1198 249
rect 1232 215 1266 249
rect 1300 215 1484 249
rect 1184 199 1484 215
rect 627 153 670 183
rect 828 177 858 199
rect 923 192 1046 199
rect 1016 177 1046 192
rect 1100 177 1130 199
rect 1184 177 1214 199
rect 1286 177 1316 199
rect 1370 177 1400 199
rect 1454 177 1484 199
rect 640 131 670 153
rect 79 21 109 47
rect 163 21 193 47
rect 351 21 381 47
rect 458 21 488 47
rect 545 21 575 47
rect 640 21 670 47
rect 828 21 858 47
rect 1016 21 1046 47
rect 1100 21 1130 47
rect 1184 21 1214 47
rect 1286 21 1316 47
rect 1370 21 1400 47
rect 1454 21 1484 47
<< polycont >>
rect 32 230 66 264
rect 134 230 168 264
rect 535 331 569 365
rect 671 323 705 357
rect 433 287 467 321
rect 340 169 374 203
rect 459 157 493 191
rect 721 215 755 249
rect 910 215 944 249
rect 1098 215 1132 249
rect 1198 215 1232 249
rect 1266 215 1300 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 17 477 69 493
rect 17 443 35 477
rect 17 409 69 443
rect 103 461 169 527
rect 103 427 119 461
rect 153 427 169 461
rect 203 477 248 493
rect 237 443 248 477
rect 17 375 35 409
rect 203 409 248 443
rect 290 485 363 527
rect 667 485 739 527
rect 290 451 307 485
rect 341 451 363 485
rect 290 439 363 451
rect 495 473 633 485
rect 495 439 511 473
rect 545 439 633 473
rect 583 421 633 439
rect 701 451 739 485
rect 667 435 739 451
rect 779 471 823 487
rect 813 437 823 471
rect 583 418 636 421
rect 583 412 637 418
rect 69 391 156 393
rect 69 375 122 391
rect 17 359 122 375
rect 18 264 66 325
rect 18 255 32 264
rect 18 221 30 255
rect 64 221 66 230
rect 18 197 66 221
rect 122 280 156 357
rect 237 375 248 409
rect 203 317 248 375
rect 305 391 547 405
rect 596 403 637 412
rect 339 381 547 391
rect 339 371 569 381
rect 501 365 569 371
rect 409 321 467 337
rect 409 317 433 321
rect 203 287 433 317
rect 501 331 535 365
rect 501 315 569 331
rect 122 264 168 280
rect 122 230 134 264
rect 122 214 168 230
rect 203 271 467 287
rect 122 161 156 214
rect 17 127 156 161
rect 17 119 69 127
rect 17 85 35 119
rect 203 119 256 271
rect 513 207 547 315
rect 603 265 637 403
rect 779 373 823 437
rect 859 471 916 527
rect 859 437 866 471
rect 900 437 916 471
rect 859 402 916 437
rect 950 477 1007 493
rect 950 443 973 477
rect 950 409 1007 443
rect 671 368 823 373
rect 671 357 779 368
rect 705 334 779 357
rect 813 334 823 368
rect 705 323 823 334
rect 671 307 823 323
rect 789 265 823 307
rect 950 375 973 409
rect 950 341 1007 375
rect 1115 485 1168 527
rect 1115 451 1134 485
rect 1115 417 1168 451
rect 1115 383 1134 417
rect 1115 367 1168 383
rect 1208 475 1274 491
rect 1208 441 1224 475
rect 1258 441 1274 475
rect 1208 401 1274 441
rect 1308 485 1360 527
rect 1308 451 1326 485
rect 1308 435 1360 451
rect 1394 485 1460 493
rect 1394 451 1410 485
rect 1444 451 1460 485
rect 1394 417 1460 451
rect 1394 401 1410 417
rect 1208 383 1410 401
rect 1444 383 1460 417
rect 1208 367 1460 383
rect 1317 357 1460 367
rect 950 307 973 341
rect 1350 349 1460 357
rect 1007 307 1228 333
rect 950 299 1228 307
rect 603 249 755 265
rect 603 233 721 249
rect 306 169 340 203
rect 374 169 390 203
rect 306 153 390 169
rect 458 191 547 207
rect 458 157 459 191
rect 493 157 547 191
rect 458 141 547 157
rect 581 215 721 233
rect 581 199 755 215
rect 789 249 944 265
rect 789 215 910 249
rect 789 199 944 215
rect 17 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 237 85 256 119
rect 581 107 615 199
rect 789 149 823 199
rect 978 177 1012 299
rect 1046 255 1148 265
rect 1080 249 1148 255
rect 1080 221 1098 249
rect 1046 215 1098 221
rect 1132 215 1148 249
rect 1046 211 1148 215
rect 1182 258 1228 299
rect 1350 315 1410 349
rect 1444 315 1460 349
rect 1182 249 1316 258
rect 1182 215 1198 249
rect 1232 215 1266 249
rect 1300 215 1316 249
rect 1182 211 1316 215
rect 1182 177 1224 211
rect 1350 177 1460 315
rect 1494 485 1547 527
rect 1528 451 1547 485
rect 1494 417 1547 451
rect 1528 383 1547 417
rect 1494 349 1547 383
rect 1528 315 1547 349
rect 1494 297 1547 315
rect 978 165 1224 177
rect 203 69 256 85
rect 103 17 169 59
rect 290 59 307 93
rect 341 59 357 93
rect 483 73 499 107
rect 533 73 615 107
rect 779 133 823 149
rect 950 143 1224 165
rect 1258 161 1460 177
rect 1258 143 1410 161
rect 290 17 357 59
rect 663 72 680 106
rect 714 72 730 106
rect 779 99 784 133
rect 818 99 823 133
rect 779 83 823 99
rect 859 107 916 143
rect 663 17 730 72
rect 859 73 868 107
rect 902 73 916 107
rect 859 17 916 73
rect 950 108 1012 143
rect 1258 109 1292 143
rect 1394 127 1410 143
rect 1444 127 1460 161
rect 950 74 972 108
rect 1006 74 1012 108
rect 950 58 1012 74
rect 1118 93 1174 109
rect 1118 59 1140 93
rect 1118 17 1174 59
rect 1208 101 1292 109
rect 1208 67 1224 101
rect 1258 67 1292 101
rect 1208 51 1292 67
rect 1326 93 1360 109
rect 1326 17 1360 59
rect 1394 93 1460 127
rect 1394 59 1410 93
rect 1444 59 1460 93
rect 1394 51 1460 59
rect 1494 161 1547 177
rect 1528 127 1547 161
rect 1494 93 1547 127
rect 1528 59 1547 93
rect 1494 17 1547 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 122 357 156 391
rect 30 230 32 255
rect 32 230 64 255
rect 30 221 64 230
rect 305 357 339 391
rect 1046 221 1080 255
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
<< metal1 >>
rect 0 561 1564 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 0 496 1564 527
rect 110 391 168 397
rect 110 357 122 391
rect 156 388 168 391
rect 293 391 351 397
rect 293 388 305 391
rect 156 360 305 388
rect 156 357 168 360
rect 110 351 168 357
rect 293 357 305 360
rect 339 357 351 391
rect 293 351 351 357
rect 18 255 76 261
rect 18 221 30 255
rect 64 252 76 255
rect 1034 255 1092 261
rect 1034 252 1046 255
rect 64 224 1046 252
rect 64 221 76 224
rect 18 215 76 221
rect 1034 221 1046 224
rect 1080 221 1092 255
rect 1034 215 1092 221
rect 0 17 1564 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
rect 0 -48 1564 -17
<< labels >>
flabel corelocali s 30 289 64 323 0 FreeSans 200 0 0 0 CLK
port 1 nsew
flabel corelocali s 1317 357 1351 391 0 FreeSans 200 0 0 0 GCLK
port 7 nsew
flabel corelocali s 1409 153 1443 187 0 FreeSans 200 0 0 0 GCLK
port 7 nsew
flabel corelocali s 1409 425 1443 459 0 FreeSans 200 0 0 0 GCLK
port 7 nsew
flabel corelocali s 1409 357 1443 391 0 FreeSans 200 0 0 0 GCLK
port 7 nsew
flabel corelocali s 1409 221 1443 255 0 FreeSans 200 0 0 0 GCLK
port 7 nsew
flabel corelocali s 1231 425 1265 459 0 FreeSans 200 0 0 0 GCLK
port 7 nsew
flabel corelocali s 1409 289 1443 323 0 FreeSans 200 0 0 0 GCLK
port 7 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 200 0 0 0 CLK
port 1 nsew
flabel corelocali s 306 153 340 187 0 FreeSans 200 0 0 0 GATE
port 2 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel metal1 s 47 0 47 0 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel metal1 s 47 544 47 544 0 FreeSans 200 0 0 0 VPWR
port 6 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew
rlabel comment s 0 0 0 0 4 dlclkp_4
<< properties >>
string FIXED_BBOX 0 0 1564 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2598802
string GDS_START 2586004
<< end >>
