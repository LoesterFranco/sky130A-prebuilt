magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 644 561
rect 26 299 85 527
rect 137 333 203 493
rect 237 367 271 527
rect 305 333 371 493
rect 405 367 439 527
rect 473 337 539 493
rect 573 435 607 527
rect 473 333 627 337
rect 137 299 627 333
rect 21 215 523 265
rect 557 181 627 299
rect 153 145 627 181
rect 26 17 79 109
rect 153 51 187 145
rect 237 17 271 109
rect 321 51 355 145
rect 405 17 439 109
rect 489 51 523 145
rect 557 17 607 110
rect 0 -17 644 17
<< metal1 >>
rect 0 496 644 592
rect 0 -48 644 48
<< labels >>
rlabel locali s 21 215 523 265 6 A
port 1 nsew signal input
rlabel locali s 557 181 627 299 6 Y
port 2 nsew signal output
rlabel locali s 489 51 523 145 6 Y
port 2 nsew signal output
rlabel locali s 473 337 539 493 6 Y
port 2 nsew signal output
rlabel locali s 473 333 627 337 6 Y
port 2 nsew signal output
rlabel locali s 321 51 355 145 6 Y
port 2 nsew signal output
rlabel locali s 305 333 371 493 6 Y
port 2 nsew signal output
rlabel locali s 153 145 627 181 6 Y
port 2 nsew signal output
rlabel locali s 153 51 187 145 6 Y
port 2 nsew signal output
rlabel locali s 137 333 203 493 6 Y
port 2 nsew signal output
rlabel locali s 137 299 627 333 6 Y
port 2 nsew signal output
rlabel locali s 557 17 607 110 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 405 17 439 109 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 237 17 271 109 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 26 17 79 109 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 0 -17 644 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 644 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 573 435 607 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 405 367 439 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 237 367 271 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 26 299 85 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 0 527 644 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 496 644 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2230196
string GDS_START 2224246
<< end >>
