magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 113 333 179 493
rect 301 333 367 493
rect 489 333 555 493
rect 677 333 743 493
rect 865 333 931 493
rect 1053 333 1119 493
rect 1241 333 1307 493
rect 1429 333 1495 493
rect 1617 333 1683 493
rect 1805 333 1871 493
rect 1993 333 2059 493
rect 2181 333 2247 493
rect 113 299 2247 333
rect 67 211 1153 265
rect 1209 211 1291 299
rect 2193 265 2247 299
rect 1325 211 2139 265
rect 2193 211 2287 265
rect 1231 177 1291 211
rect 2193 177 2247 211
rect 1231 127 2247 177
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2392 561
rect 25 299 79 527
rect 213 367 267 527
rect 401 367 455 527
rect 589 367 643 527
rect 777 367 831 527
rect 965 367 1019 527
rect 1153 367 1207 527
rect 1341 367 1395 527
rect 1529 367 1583 527
rect 1717 367 1771 527
rect 1905 367 1959 527
rect 2093 367 2147 527
rect 2281 299 2335 527
rect 18 143 1197 177
rect 18 51 85 143
rect 119 17 173 109
rect 207 51 273 143
rect 307 17 361 109
rect 395 51 461 143
rect 495 17 549 109
rect 583 51 649 143
rect 683 17 737 109
rect 771 51 837 143
rect 871 17 925 109
rect 959 51 1025 143
rect 1059 17 1113 109
rect 1147 93 1197 143
rect 2291 93 2341 177
rect 1147 51 2341 93
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2392 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
<< metal1 >>
rect 0 561 2392 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2392 561
rect 0 496 2392 527
rect 0 17 2392 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2392 17
rect 0 -48 2392 -17
<< labels >>
rlabel locali s 1325 211 2139 265 6 A
port 1 nsew signal input
rlabel locali s 67 211 1153 265 6 B
port 2 nsew signal input
rlabel locali s 2193 265 2247 299 6 Y
port 3 nsew signal output
rlabel locali s 2193 211 2287 265 6 Y
port 3 nsew signal output
rlabel locali s 2193 177 2247 211 6 Y
port 3 nsew signal output
rlabel locali s 2181 333 2247 493 6 Y
port 3 nsew signal output
rlabel locali s 1993 333 2059 493 6 Y
port 3 nsew signal output
rlabel locali s 1805 333 1871 493 6 Y
port 3 nsew signal output
rlabel locali s 1617 333 1683 493 6 Y
port 3 nsew signal output
rlabel locali s 1429 333 1495 493 6 Y
port 3 nsew signal output
rlabel locali s 1241 333 1307 493 6 Y
port 3 nsew signal output
rlabel locali s 1231 177 1291 211 6 Y
port 3 nsew signal output
rlabel locali s 1231 127 2247 177 6 Y
port 3 nsew signal output
rlabel locali s 1209 211 1291 299 6 Y
port 3 nsew signal output
rlabel locali s 1053 333 1119 493 6 Y
port 3 nsew signal output
rlabel locali s 865 333 931 493 6 Y
port 3 nsew signal output
rlabel locali s 677 333 743 493 6 Y
port 3 nsew signal output
rlabel locali s 489 333 555 493 6 Y
port 3 nsew signal output
rlabel locali s 301 333 367 493 6 Y
port 3 nsew signal output
rlabel locali s 113 333 179 493 6 Y
port 3 nsew signal output
rlabel locali s 113 299 2247 333 6 Y
port 3 nsew signal output
rlabel metal1 s 0 -48 2392 48 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 496 2392 592 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2392 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3457254
string GDS_START 3440238
<< end >>
