magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 29 153 89 323
rect 326 329 455 391
rect 489 316 616 473
rect 554 155 616 316
rect 541 51 616 155
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 35 403 69 489
rect 103 437 179 527
rect 35 357 180 403
rect 133 227 180 357
rect 214 295 281 484
rect 327 433 455 527
rect 214 265 416 295
rect 214 261 501 265
rect 133 161 250 227
rect 284 189 501 261
rect 133 131 177 161
rect 18 17 85 118
rect 129 56 177 131
rect 284 122 328 189
rect 243 83 328 122
rect 243 54 277 83
rect 400 17 489 116
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 29 153 89 323 6 A_N
port 1 nsew signal input
rlabel locali s 326 329 455 391 6 B
port 2 nsew signal input
rlabel locali s 554 155 616 316 6 X
port 3 nsew signal output
rlabel locali s 541 51 616 155 6 X
port 3 nsew signal output
rlabel locali s 489 316 616 473 6 X
port 3 nsew signal output
rlabel metal1 s 0 -48 644 48 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1500784
string GDS_START 1495146
<< end >>
