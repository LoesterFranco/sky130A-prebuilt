magic
tech sky130A
magscale 1 2
timestamp 1601050056
<< nwell >>
rect -38 332 806 704
<< pwell >>
rect 0 0 768 49
<< scpmos >>
rect 97 368 133 592
rect 187 368 223 592
rect 350 384 386 584
rect 440 384 476 584
rect 542 384 578 584
rect 650 384 686 584
<< nmoslvt >>
rect 82 74 112 222
rect 168 74 198 222
rect 362 74 392 222
rect 454 74 484 222
rect 554 74 584 222
rect 654 74 684 222
<< ndiff >>
rect 27 210 82 222
rect 27 176 37 210
rect 71 176 82 210
rect 27 124 82 176
rect 27 90 37 124
rect 71 90 82 124
rect 27 74 82 90
rect 112 203 168 222
rect 112 169 123 203
rect 157 169 168 203
rect 112 120 168 169
rect 112 86 123 120
rect 157 86 168 120
rect 112 74 168 86
rect 198 140 248 222
rect 312 154 362 222
rect 198 124 253 140
rect 198 90 209 124
rect 243 90 253 124
rect 198 74 253 90
rect 307 131 362 154
rect 307 97 317 131
rect 351 97 362 131
rect 307 74 362 97
rect 392 210 454 222
rect 392 176 406 210
rect 440 176 454 210
rect 392 74 454 176
rect 484 210 554 222
rect 484 176 509 210
rect 543 176 554 210
rect 484 120 554 176
rect 484 86 509 120
rect 543 86 554 120
rect 484 74 554 86
rect 584 142 654 222
rect 584 108 609 142
rect 643 108 654 142
rect 584 74 654 108
rect 684 210 741 222
rect 684 176 695 210
rect 729 176 741 210
rect 684 120 741 176
rect 684 86 695 120
rect 729 86 741 120
rect 684 74 741 86
<< pdiff >>
rect 31 580 97 592
rect 31 546 43 580
rect 77 546 97 580
rect 31 497 97 546
rect 31 463 43 497
rect 77 463 97 497
rect 31 414 97 463
rect 31 380 43 414
rect 77 380 97 414
rect 31 368 97 380
rect 133 580 187 592
rect 133 546 143 580
rect 177 546 187 580
rect 133 497 187 546
rect 133 463 143 497
rect 177 463 187 497
rect 133 414 187 463
rect 133 380 143 414
rect 177 380 187 414
rect 133 368 187 380
rect 223 584 289 592
rect 223 580 350 584
rect 223 546 233 580
rect 267 571 350 580
rect 267 546 306 571
rect 223 537 306 546
rect 340 537 350 571
rect 223 508 350 537
rect 223 474 233 508
rect 267 499 350 508
rect 267 474 306 499
rect 223 465 306 474
rect 340 465 350 499
rect 223 384 350 465
rect 386 384 440 584
rect 476 572 542 584
rect 476 538 486 572
rect 520 538 542 572
rect 476 504 542 538
rect 476 470 486 504
rect 520 470 542 504
rect 476 436 542 470
rect 476 402 486 436
rect 520 402 542 436
rect 476 384 542 402
rect 578 384 650 584
rect 686 572 741 584
rect 686 538 696 572
rect 730 538 741 572
rect 686 504 741 538
rect 686 470 696 504
rect 730 470 741 504
rect 686 436 741 470
rect 686 402 696 436
rect 730 402 741 436
rect 686 384 741 402
rect 223 368 273 384
<< ndiffc >>
rect 37 176 71 210
rect 37 90 71 124
rect 123 169 157 203
rect 123 86 157 120
rect 209 90 243 124
rect 317 97 351 131
rect 406 176 440 210
rect 509 176 543 210
rect 509 86 543 120
rect 609 108 643 142
rect 695 176 729 210
rect 695 86 729 120
<< pdiffc >>
rect 43 546 77 580
rect 43 463 77 497
rect 43 380 77 414
rect 143 546 177 580
rect 143 463 177 497
rect 143 380 177 414
rect 233 546 267 580
rect 306 537 340 571
rect 233 474 267 508
rect 306 465 340 499
rect 486 538 520 572
rect 486 470 520 504
rect 486 402 520 436
rect 696 538 730 572
rect 696 470 730 504
rect 696 402 730 436
<< poly >>
rect 97 592 133 618
rect 187 592 223 618
rect 350 584 386 610
rect 440 584 476 610
rect 542 584 578 610
rect 650 584 686 610
rect 97 326 133 368
rect 187 326 223 368
rect 350 352 386 384
rect 440 352 476 384
rect 542 352 578 384
rect 309 336 392 352
rect 82 310 261 326
rect 82 278 211 310
rect 82 222 112 278
rect 168 276 211 278
rect 245 276 261 310
rect 309 302 325 336
rect 359 302 392 336
rect 309 286 392 302
rect 434 336 500 352
rect 434 302 450 336
rect 484 302 500 336
rect 434 286 500 302
rect 542 336 608 352
rect 542 302 558 336
rect 592 302 608 336
rect 542 286 608 302
rect 650 326 686 384
rect 650 310 747 326
rect 168 260 261 276
rect 168 222 198 260
rect 362 222 392 286
rect 454 222 484 286
rect 554 222 584 286
rect 650 276 697 310
rect 731 276 747 310
rect 650 260 747 276
rect 654 222 684 260
rect 82 48 112 74
rect 168 48 198 74
rect 362 48 392 74
rect 454 48 484 74
rect 554 48 584 74
rect 654 48 684 74
<< polycont >>
rect 211 276 245 310
rect 325 302 359 336
rect 450 302 484 336
rect 558 302 592 336
rect 697 276 731 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 27 580 93 649
rect 27 546 43 580
rect 77 546 93 580
rect 27 497 93 546
rect 27 463 43 497
rect 77 463 93 497
rect 27 414 93 463
rect 27 380 43 414
rect 77 380 93 414
rect 27 364 93 380
rect 127 580 193 596
rect 127 546 143 580
rect 177 546 193 580
rect 127 497 193 546
rect 127 463 143 497
rect 177 463 193 497
rect 127 414 193 463
rect 227 580 358 649
rect 227 546 233 580
rect 267 571 358 580
rect 267 546 306 571
rect 227 537 306 546
rect 340 537 358 571
rect 227 508 358 537
rect 227 474 233 508
rect 267 499 358 508
rect 267 474 306 499
rect 227 465 306 474
rect 340 465 358 499
rect 227 458 358 465
rect 470 572 536 588
rect 470 538 486 572
rect 520 538 536 572
rect 470 504 536 538
rect 470 470 486 504
rect 520 470 536 504
rect 470 436 536 470
rect 470 424 486 436
rect 127 380 143 414
rect 177 380 193 414
rect 127 364 193 380
rect 227 402 486 424
rect 520 402 536 436
rect 227 390 536 402
rect 680 572 746 649
rect 680 538 696 572
rect 730 538 746 572
rect 680 504 746 538
rect 680 470 696 504
rect 730 470 746 504
rect 680 436 746 470
rect 680 402 696 436
rect 730 402 746 436
rect 680 390 746 402
rect 127 226 161 364
rect 227 326 261 390
rect 195 310 261 326
rect 195 276 211 310
rect 245 276 261 310
rect 309 336 375 356
rect 309 302 325 336
rect 359 302 375 336
rect 309 286 375 302
rect 409 336 500 356
rect 409 302 450 336
rect 484 302 500 336
rect 409 286 500 302
rect 542 336 647 356
rect 542 302 558 336
rect 592 302 647 336
rect 542 286 647 302
rect 681 310 747 356
rect 195 260 261 276
rect 681 276 697 310
rect 731 276 747 310
rect 681 260 747 276
rect 227 226 261 260
rect 21 210 73 226
rect 21 176 37 210
rect 71 176 73 210
rect 21 124 73 176
rect 21 90 37 124
rect 71 90 73 124
rect 21 17 73 90
rect 107 203 173 226
rect 107 169 123 203
rect 157 169 173 203
rect 227 210 459 226
rect 227 176 406 210
rect 440 176 459 210
rect 107 164 173 169
rect 107 120 158 164
rect 401 160 459 176
rect 493 210 745 226
rect 493 176 509 210
rect 543 192 695 210
rect 543 176 559 192
rect 301 131 367 142
rect 107 86 123 120
rect 157 86 158 120
rect 107 70 158 86
rect 193 124 259 128
rect 193 90 209 124
rect 243 90 259 124
rect 193 17 259 90
rect 301 97 317 131
rect 351 104 367 131
rect 493 120 559 176
rect 729 176 745 210
rect 493 104 509 120
rect 351 97 509 104
rect 301 86 509 97
rect 543 86 559 120
rect 301 70 559 86
rect 593 142 659 158
rect 593 108 609 142
rect 643 108 659 142
rect 593 17 659 108
rect 695 120 745 176
rect 729 86 745 120
rect 695 70 745 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
rlabel comment s 0 0 0 0 4 o22a_2
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 127 168 161 202 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 768 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1282800
string GDS_START 1275870
<< end >>
