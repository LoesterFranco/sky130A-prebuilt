magic
tech sky130A
magscale 1 2
timestamp 1604502697
<< nwell >>
rect -38 261 406 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 120 67 150 177
rect 222 67 252 177
<< pmoshvt >>
rect 96 297 146 497
rect 202 297 252 497
<< ndiff >>
rect 63 133 120 177
rect 63 99 75 133
rect 109 99 120 133
rect 63 67 120 99
rect 150 67 222 177
rect 252 133 309 177
rect 252 99 263 133
rect 297 99 309 133
rect 252 67 309 99
<< pdiff >>
rect 39 485 96 497
rect 39 451 47 485
rect 81 451 96 485
rect 39 417 96 451
rect 39 383 47 417
rect 81 383 96 417
rect 39 297 96 383
rect 146 471 202 497
rect 146 437 157 471
rect 191 437 202 471
rect 146 351 202 437
rect 146 317 157 351
rect 191 317 202 351
rect 146 297 202 317
rect 252 485 325 497
rect 252 451 283 485
rect 317 451 325 485
rect 252 414 325 451
rect 252 380 283 414
rect 317 380 325 414
rect 252 343 325 380
rect 252 309 283 343
rect 317 309 325 343
rect 252 297 325 309
<< ndiffc >>
rect 75 99 109 133
rect 263 99 297 133
<< pdiffc >>
rect 47 451 81 485
rect 47 383 81 417
rect 157 437 191 471
rect 157 317 191 351
rect 283 451 317 485
rect 283 380 317 414
rect 283 309 317 343
<< poly >>
rect 96 497 146 523
rect 202 497 252 523
rect 96 263 146 297
rect 29 249 146 263
rect 29 215 86 249
rect 120 234 146 249
rect 202 234 252 297
rect 120 215 252 234
rect 29 199 252 215
rect 120 177 150 199
rect 222 177 252 199
rect 120 41 150 67
rect 222 41 252 67
<< polycont >>
rect 86 215 120 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 45 525 333 527
rect 45 485 111 525
rect 45 451 47 485
rect 81 451 111 485
rect 45 417 111 451
rect 45 383 47 417
rect 81 383 111 417
rect 45 367 111 383
rect 157 471 247 491
rect 191 437 247 471
rect 157 351 247 437
rect 29 249 120 333
rect 29 215 86 249
rect 29 199 120 215
rect 191 317 247 351
rect 157 150 247 317
rect 281 485 333 525
rect 281 451 283 485
rect 317 451 333 485
rect 281 414 333 451
rect 281 380 283 414
rect 317 380 333 414
rect 281 343 333 380
rect 281 309 283 343
rect 317 309 333 343
rect 281 291 333 309
rect 59 133 123 149
rect 59 99 75 133
rect 109 99 123 133
rect 59 17 123 99
rect 157 133 309 150
rect 157 99 263 133
rect 297 99 309 133
rect 157 63 309 99
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
<< metal1 >>
rect 0 561 368 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 0 496 368 527
rect 0 17 368 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
rect 0 -48 368 -17
<< labels >>
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew
flabel corelocali s 211 153 245 187 0 FreeSans 200 0 0 0 Y
port 6 nsew
flabel corelocali s 211 221 245 255 0 FreeSans 200 0 0 0 Y
port 6 nsew
flabel corelocali s 29 289 63 323 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 211 85 245 119 0 FreeSans 200 0 0 0 Y
port 6 nsew
flabel corelocali s 29 221 63 255 0 FreeSans 200 0 0 0 A
port 1 nsew
rlabel comment s 0 0 0 0 4 clkinvlp_2
<< properties >>
string FIXED_BBOX 0 0 368 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1821594
string GDS_START 1817988
<< end >>
