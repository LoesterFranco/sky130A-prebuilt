magic
tech sky130A
magscale 1 2
timestamp 1601050047
<< nwell >>
rect -38 332 1670 704
<< pwell >>
rect 0 0 1632 49
<< scpmos >>
rect 89 392 119 592
rect 189 392 219 592
rect 279 392 309 592
rect 369 392 399 592
rect 471 392 501 592
rect 561 392 591 592
rect 661 392 691 592
rect 761 392 791 592
rect 875 392 905 592
rect 965 392 995 592
rect 1055 392 1085 592
rect 1145 392 1175 592
rect 1246 368 1276 592
rect 1336 368 1366 592
rect 1426 368 1456 592
rect 1516 368 1546 592
<< nmoslvt >>
rect 84 125 114 253
rect 202 125 232 253
rect 288 125 318 253
rect 388 125 418 253
rect 474 125 504 253
rect 572 125 602 253
rect 658 125 688 253
rect 776 78 806 206
rect 876 78 906 206
rect 978 119 1008 247
rect 1064 119 1094 247
rect 1150 119 1180 247
rect 1252 99 1282 247
rect 1346 99 1376 247
rect 1432 99 1462 247
rect 1518 99 1548 247
<< ndiff >>
rect 27 241 84 253
rect 27 207 39 241
rect 73 207 84 241
rect 27 171 84 207
rect 27 137 39 171
rect 73 137 84 171
rect 27 125 84 137
rect 114 125 202 253
rect 232 173 288 253
rect 232 139 243 173
rect 277 139 288 173
rect 232 125 288 139
rect 318 173 388 253
rect 318 139 343 173
rect 377 139 388 173
rect 318 125 388 139
rect 418 173 474 253
rect 418 139 429 173
rect 463 139 474 173
rect 418 125 474 139
rect 504 171 572 253
rect 504 137 521 171
rect 555 137 572 171
rect 504 125 572 137
rect 602 173 658 253
rect 602 139 613 173
rect 647 139 658 173
rect 602 125 658 139
rect 688 206 738 253
rect 928 206 978 247
rect 688 125 776 206
rect 129 124 187 125
rect 129 90 141 124
rect 175 90 187 124
rect 129 78 187 90
rect 703 123 776 125
rect 703 89 715 123
rect 749 89 776 123
rect 703 78 776 89
rect 806 124 876 206
rect 806 90 817 124
rect 851 90 876 124
rect 806 78 876 90
rect 906 124 978 206
rect 906 90 917 124
rect 951 119 978 124
rect 1008 237 1064 247
rect 1008 203 1019 237
rect 1053 203 1064 237
rect 1008 169 1064 203
rect 1008 135 1019 169
rect 1053 135 1064 169
rect 1008 119 1064 135
rect 1094 176 1150 247
rect 1094 142 1105 176
rect 1139 142 1150 176
rect 1094 119 1150 142
rect 1180 219 1252 247
rect 1180 185 1207 219
rect 1241 185 1252 219
rect 1180 145 1252 185
rect 1180 119 1207 145
rect 951 90 963 119
rect 906 78 963 90
rect 703 77 761 78
rect 1195 111 1207 119
rect 1241 111 1252 145
rect 1195 99 1252 111
rect 1282 219 1346 247
rect 1282 185 1301 219
rect 1335 185 1346 219
rect 1282 145 1346 185
rect 1282 111 1301 145
rect 1335 111 1346 145
rect 1282 99 1346 111
rect 1376 151 1432 247
rect 1376 117 1387 151
rect 1421 117 1432 151
rect 1376 99 1432 117
rect 1462 235 1518 247
rect 1462 201 1473 235
rect 1507 201 1518 235
rect 1462 99 1518 201
rect 1548 163 1598 247
rect 1548 151 1605 163
rect 1548 117 1559 151
rect 1593 117 1605 151
rect 1548 99 1605 117
<< pdiff >>
rect 30 580 89 592
rect 30 546 42 580
rect 76 546 89 580
rect 30 509 89 546
rect 30 475 42 509
rect 76 475 89 509
rect 30 438 89 475
rect 30 404 42 438
rect 76 404 89 438
rect 30 392 89 404
rect 119 580 189 592
rect 119 546 132 580
rect 166 546 189 580
rect 119 493 189 546
rect 119 459 132 493
rect 166 459 189 493
rect 119 392 189 459
rect 219 531 279 592
rect 219 497 232 531
rect 266 497 279 531
rect 219 449 279 497
rect 219 415 232 449
rect 266 415 279 449
rect 219 392 279 415
rect 309 570 369 592
rect 309 536 322 570
rect 356 536 369 570
rect 309 392 369 536
rect 399 561 471 592
rect 399 527 413 561
rect 447 527 471 561
rect 399 392 471 527
rect 501 561 561 592
rect 501 527 514 561
rect 548 527 561 561
rect 501 392 561 527
rect 591 547 661 592
rect 591 513 614 547
rect 648 513 661 547
rect 591 477 661 513
rect 591 443 614 477
rect 648 443 661 477
rect 591 392 661 443
rect 691 561 761 592
rect 691 527 714 561
rect 748 527 761 561
rect 691 392 761 527
rect 791 561 875 592
rect 791 527 814 561
rect 848 527 875 561
rect 791 392 875 527
rect 905 561 965 592
rect 905 527 918 561
rect 952 527 965 561
rect 905 392 965 527
rect 995 460 1055 592
rect 995 426 1008 460
rect 1042 426 1055 460
rect 995 392 1055 426
rect 1085 561 1145 592
rect 1085 527 1098 561
rect 1132 527 1145 561
rect 1085 392 1145 527
rect 1175 580 1246 592
rect 1175 546 1188 580
rect 1222 546 1246 580
rect 1175 509 1246 546
rect 1175 475 1188 509
rect 1222 475 1246 509
rect 1175 438 1246 475
rect 1175 404 1188 438
rect 1222 404 1246 438
rect 1175 392 1246 404
rect 1193 368 1246 392
rect 1276 580 1336 592
rect 1276 546 1289 580
rect 1323 546 1336 580
rect 1276 499 1336 546
rect 1276 465 1289 499
rect 1323 465 1336 499
rect 1276 419 1336 465
rect 1276 385 1289 419
rect 1323 385 1336 419
rect 1276 368 1336 385
rect 1366 580 1426 592
rect 1366 546 1379 580
rect 1413 546 1426 580
rect 1366 487 1426 546
rect 1366 453 1379 487
rect 1413 453 1426 487
rect 1366 368 1426 453
rect 1456 580 1516 592
rect 1456 546 1469 580
rect 1503 546 1516 580
rect 1456 497 1516 546
rect 1456 463 1469 497
rect 1503 463 1516 497
rect 1456 414 1516 463
rect 1456 380 1469 414
rect 1503 380 1516 414
rect 1456 368 1516 380
rect 1546 580 1605 592
rect 1546 546 1559 580
rect 1593 546 1605 580
rect 1546 497 1605 546
rect 1546 463 1559 497
rect 1593 463 1605 497
rect 1546 414 1605 463
rect 1546 380 1559 414
rect 1593 380 1605 414
rect 1546 368 1605 380
<< ndiffc >>
rect 39 207 73 241
rect 39 137 73 171
rect 243 139 277 173
rect 343 139 377 173
rect 429 139 463 173
rect 521 137 555 171
rect 613 139 647 173
rect 141 90 175 124
rect 715 89 749 123
rect 817 90 851 124
rect 917 90 951 124
rect 1019 203 1053 237
rect 1019 135 1053 169
rect 1105 142 1139 176
rect 1207 185 1241 219
rect 1207 111 1241 145
rect 1301 185 1335 219
rect 1301 111 1335 145
rect 1387 117 1421 151
rect 1473 201 1507 235
rect 1559 117 1593 151
<< pdiffc >>
rect 42 546 76 580
rect 42 475 76 509
rect 42 404 76 438
rect 132 546 166 580
rect 132 459 166 493
rect 232 497 266 531
rect 232 415 266 449
rect 322 536 356 570
rect 413 527 447 561
rect 514 527 548 561
rect 614 513 648 547
rect 614 443 648 477
rect 714 527 748 561
rect 814 527 848 561
rect 918 527 952 561
rect 1008 426 1042 460
rect 1098 527 1132 561
rect 1188 546 1222 580
rect 1188 475 1222 509
rect 1188 404 1222 438
rect 1289 546 1323 580
rect 1289 465 1323 499
rect 1289 385 1323 419
rect 1379 546 1413 580
rect 1379 453 1413 487
rect 1469 546 1503 580
rect 1469 463 1503 497
rect 1469 380 1503 414
rect 1559 546 1593 580
rect 1559 463 1593 497
rect 1559 380 1593 414
<< poly >>
rect 89 592 119 618
rect 189 592 219 618
rect 279 592 309 618
rect 369 592 399 618
rect 471 592 501 618
rect 561 592 591 618
rect 661 592 691 618
rect 761 592 791 618
rect 875 592 905 618
rect 965 592 995 618
rect 1055 592 1085 618
rect 1145 592 1175 618
rect 1246 592 1276 618
rect 1336 592 1366 618
rect 1426 592 1456 618
rect 1516 592 1546 618
rect 89 377 119 392
rect 189 377 219 392
rect 279 377 309 392
rect 369 377 399 392
rect 471 377 501 392
rect 561 377 591 392
rect 661 377 691 392
rect 761 377 791 392
rect 875 377 905 392
rect 965 377 995 392
rect 1055 377 1085 392
rect 1145 377 1175 392
rect 86 298 122 377
rect 186 341 222 377
rect 276 341 312 377
rect 366 360 402 377
rect 360 344 426 360
rect 84 268 122 298
rect 192 325 318 341
rect 192 291 243 325
rect 277 291 318 325
rect 360 310 376 344
rect 410 310 426 344
rect 360 294 426 310
rect 192 275 318 291
rect 84 253 114 268
rect 202 253 232 275
rect 288 253 318 275
rect 388 253 418 294
rect 468 268 504 377
rect 558 341 594 377
rect 658 341 694 377
rect 758 341 794 377
rect 872 360 908 377
rect 962 360 998 377
rect 1052 360 1088 377
rect 848 344 914 360
rect 558 325 694 341
rect 558 291 574 325
rect 608 305 694 325
rect 736 325 806 341
rect 608 291 688 305
rect 558 275 688 291
rect 736 291 752 325
rect 786 291 806 325
rect 848 310 864 344
rect 898 310 914 344
rect 848 294 914 310
rect 962 344 1088 360
rect 962 310 994 344
rect 1028 324 1088 344
rect 1028 310 1094 324
rect 962 294 1094 310
rect 736 275 806 291
rect 474 253 504 268
rect 572 253 602 275
rect 658 253 688 275
rect 776 206 806 275
rect 876 206 906 294
rect 978 247 1008 294
rect 1064 247 1094 294
rect 1142 292 1178 377
rect 1246 353 1276 368
rect 1336 353 1366 368
rect 1426 353 1456 368
rect 1516 353 1546 368
rect 1243 335 1279 353
rect 1333 335 1369 353
rect 1423 335 1459 353
rect 1513 335 1549 353
rect 1228 319 1549 335
rect 1142 262 1180 292
rect 1228 285 1244 319
rect 1278 285 1312 319
rect 1346 285 1380 319
rect 1414 299 1549 319
rect 1414 285 1548 299
rect 1228 269 1548 285
rect 1150 247 1180 262
rect 1252 247 1282 269
rect 1346 247 1376 269
rect 1432 247 1462 269
rect 1518 247 1548 269
rect 84 51 114 125
rect 202 99 232 125
rect 288 99 318 125
rect 388 51 418 125
rect 84 21 418 51
rect 474 51 504 125
rect 572 99 602 125
rect 658 99 688 125
rect 978 93 1008 119
rect 1064 93 1094 119
rect 776 51 806 78
rect 474 21 806 51
rect 876 51 906 78
rect 1150 51 1180 119
rect 1252 73 1282 99
rect 1346 73 1376 99
rect 1432 73 1462 99
rect 1518 73 1548 99
rect 876 21 1180 51
<< polycont >>
rect 243 291 277 325
rect 376 310 410 344
rect 574 291 608 325
rect 752 291 786 325
rect 864 310 898 344
rect 994 310 1028 344
rect 1244 285 1278 319
rect 1312 285 1346 319
rect 1380 285 1414 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 26 580 76 649
rect 26 546 42 580
rect 26 509 76 546
rect 26 475 42 509
rect 26 438 76 475
rect 116 581 372 615
rect 116 580 182 581
rect 116 546 132 580
rect 166 546 182 580
rect 306 570 372 581
rect 116 493 182 546
rect 116 459 132 493
rect 166 459 182 493
rect 116 443 182 459
rect 219 531 270 547
rect 219 497 232 531
rect 266 497 270 531
rect 306 536 322 570
rect 356 536 372 570
rect 306 511 372 536
rect 412 561 464 649
rect 412 527 413 561
rect 447 527 464 561
rect 412 511 464 527
rect 498 581 764 615
rect 498 561 564 581
rect 498 527 514 561
rect 548 527 564 561
rect 698 561 764 581
rect 498 511 564 527
rect 598 513 614 547
rect 648 513 664 547
rect 219 477 270 497
rect 598 477 664 513
rect 698 527 714 561
rect 748 527 764 561
rect 698 511 764 527
rect 798 561 864 649
rect 798 527 814 561
rect 848 527 864 561
rect 798 511 864 527
rect 902 561 968 596
rect 902 527 918 561
rect 952 545 968 561
rect 1082 561 1148 596
rect 1082 545 1098 561
rect 952 527 1098 545
rect 1132 527 1148 561
rect 902 511 1148 527
rect 1188 580 1238 649
rect 1222 546 1238 580
rect 1188 509 1238 546
rect 219 449 614 477
rect 26 404 42 438
rect 219 415 232 449
rect 266 443 614 449
rect 648 460 1058 477
rect 648 443 1008 460
rect 266 415 282 443
rect 219 409 282 415
rect 992 426 1008 443
rect 1042 428 1058 460
rect 1222 475 1238 509
rect 1188 438 1238 475
rect 1042 426 1112 428
rect 26 388 76 404
rect 159 375 282 409
rect 421 375 914 409
rect 992 394 1112 426
rect 23 241 89 257
rect 23 207 39 241
rect 73 207 89 241
rect 23 171 89 207
rect 23 137 39 171
rect 73 137 89 171
rect 159 192 193 375
rect 421 360 455 375
rect 360 344 455 360
rect 227 325 293 341
rect 227 291 243 325
rect 277 291 293 325
rect 360 310 376 344
rect 410 310 455 344
rect 848 344 914 375
rect 360 294 455 310
rect 505 325 647 341
rect 227 260 293 291
rect 505 291 574 325
rect 608 291 647 325
rect 505 260 647 291
rect 227 226 647 260
rect 697 325 802 341
rect 697 291 752 325
rect 786 291 802 325
rect 848 310 864 344
rect 898 310 914 344
rect 848 294 914 310
rect 951 344 1044 360
rect 951 310 994 344
rect 1028 310 1044 344
rect 951 294 1044 310
rect 1078 335 1112 394
rect 1222 404 1238 438
rect 1188 388 1238 404
rect 1273 580 1339 596
rect 1273 546 1289 580
rect 1323 546 1339 580
rect 1273 499 1339 546
rect 1273 465 1289 499
rect 1323 465 1339 499
rect 1273 419 1339 465
rect 1379 580 1429 649
rect 1413 546 1429 580
rect 1379 487 1429 546
rect 1413 453 1429 487
rect 1379 437 1429 453
rect 1469 580 1503 596
rect 1469 497 1503 546
rect 1273 385 1289 419
rect 1323 403 1339 419
rect 1469 414 1503 463
rect 1323 385 1469 403
rect 1273 380 1469 385
rect 1273 369 1503 380
rect 1078 319 1430 335
rect 697 260 802 291
rect 951 260 985 294
rect 1078 285 1244 319
rect 1278 285 1312 319
rect 1346 285 1380 319
rect 1414 285 1430 319
rect 1469 330 1503 369
rect 1543 580 1609 649
rect 1543 546 1559 580
rect 1593 546 1609 580
rect 1543 497 1609 546
rect 1543 463 1559 497
rect 1593 463 1609 497
rect 1543 414 1609 463
rect 1543 380 1559 414
rect 1593 380 1609 414
rect 1543 364 1609 380
rect 1469 296 1607 330
rect 1078 269 1430 285
rect 1078 260 1112 269
rect 697 226 985 260
rect 1019 237 1112 260
rect 1053 226 1112 237
rect 1561 235 1607 296
rect 1019 192 1053 203
rect 1191 219 1241 235
rect 159 173 293 192
rect 159 158 243 173
rect 23 17 89 137
rect 227 139 243 158
rect 277 139 293 173
rect 125 90 141 124
rect 175 90 191 124
rect 227 121 293 139
rect 327 173 393 192
rect 327 139 343 173
rect 377 139 393 173
rect 125 87 191 90
rect 327 87 393 139
rect 125 53 393 87
rect 429 173 463 192
rect 429 17 463 139
rect 499 171 577 187
rect 499 137 521 171
rect 555 137 577 171
rect 499 87 577 137
rect 613 173 1053 192
rect 647 169 1053 173
rect 647 158 1019 169
rect 647 139 663 158
rect 613 121 663 139
rect 699 123 765 124
rect 699 89 715 123
rect 749 89 765 123
rect 699 87 765 89
rect 499 53 765 87
rect 801 90 817 124
rect 851 90 867 124
rect 801 17 867 90
rect 901 90 917 124
rect 951 90 967 124
rect 1019 119 1053 135
rect 1089 176 1155 192
rect 1089 142 1105 176
rect 1139 142 1155 176
rect 901 85 967 90
rect 1089 85 1155 142
rect 901 51 1155 85
rect 1191 185 1207 219
rect 1191 145 1241 185
rect 1191 111 1207 145
rect 1191 17 1241 111
rect 1285 219 1473 235
rect 1285 185 1301 219
rect 1335 201 1473 219
rect 1507 201 1607 235
rect 1285 145 1335 185
rect 1285 111 1301 145
rect 1285 95 1335 111
rect 1371 151 1437 167
rect 1371 117 1387 151
rect 1421 117 1437 151
rect 1371 17 1437 117
rect 1543 151 1609 167
rect 1543 117 1559 151
rect 1593 117 1609 151
rect 1543 17 1609 117
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
rlabel comment s 0 0 0 0 4 maj3_4
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 703 242 737 276 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 511 242 545 276 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 607 242 641 276 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 1567 242 1601 276 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 1632 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1896102
string GDS_START 1883796
<< end >>
