magic
tech sky130A
magscale 1 2
timestamp 1604502741
<< locali >>
rect 175 430 241 596
rect 387 430 453 596
rect 175 378 453 430
rect 47 364 453 378
rect 47 344 241 364
rect 47 202 81 344
rect 115 236 181 310
rect 217 236 295 310
rect 343 236 455 310
rect 489 236 555 310
rect 47 168 548 202
rect 482 70 548 168
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 75 412 141 649
rect 280 464 346 649
rect 487 364 553 649
rect 22 17 157 120
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
rlabel locali s 489 236 555 310 6 A
port 1 nsew signal input
rlabel locali s 343 236 455 310 6 B
port 2 nsew signal input
rlabel locali s 217 236 295 310 6 C
port 3 nsew signal input
rlabel locali s 115 236 181 310 6 D
port 4 nsew signal input
rlabel locali s 482 70 548 168 6 Y
port 5 nsew signal output
rlabel locali s 387 430 453 596 6 Y
port 5 nsew signal output
rlabel locali s 175 430 241 596 6 Y
port 5 nsew signal output
rlabel locali s 175 378 453 430 6 Y
port 5 nsew signal output
rlabel locali s 47 364 453 378 6 Y
port 5 nsew signal output
rlabel locali s 47 344 241 364 6 Y
port 5 nsew signal output
rlabel locali s 47 202 81 344 6 Y
port 5 nsew signal output
rlabel locali s 47 168 548 202 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -49 576 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 576 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 576 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 2071340
string GDS_START 2066088
<< end >>
