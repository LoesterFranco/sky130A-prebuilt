magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 295 398 368 596
rect 25 290 113 356
rect 261 364 368 398
rect 261 226 295 364
rect 409 326 455 578
rect 350 260 455 326
rect 489 260 555 356
rect 217 70 295 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 27 424 93 596
rect 127 458 261 649
rect 27 390 183 424
rect 149 326 183 390
rect 149 260 227 326
rect 149 256 183 260
rect 22 222 183 256
rect 504 390 554 649
rect 22 70 72 222
rect 108 17 174 188
rect 329 192 553 226
rect 329 70 363 192
rect 399 17 467 136
rect 503 70 553 192
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
rlabel locali s 489 260 555 356 6 A1
port 1 nsew signal input
rlabel locali s 409 326 455 578 6 A2
port 2 nsew signal input
rlabel locali s 350 260 455 326 6 A2
port 2 nsew signal input
rlabel locali s 25 290 113 356 6 B1_N
port 3 nsew signal input
rlabel locali s 295 398 368 596 6 Y
port 4 nsew signal output
rlabel locali s 261 364 368 398 6 Y
port 4 nsew signal output
rlabel locali s 261 226 295 364 6 Y
port 4 nsew signal output
rlabel locali s 217 70 295 226 6 Y
port 4 nsew signal output
rlabel metal1 s 0 -49 576 49 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 617 576 715 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 576 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1381908
string GDS_START 1375542
<< end >>
