magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 28 215 248 255
<< obsli1 >>
rect 0 527 1196 561
rect 19 323 85 493
rect 119 367 173 527
rect 207 323 273 493
rect 307 367 361 527
rect 395 323 461 493
rect 495 367 549 527
rect 583 323 649 493
rect 683 367 737 527
rect 771 323 837 493
rect 871 367 925 527
rect 959 323 1025 493
rect 19 289 319 323
rect 395 289 1025 323
rect 1059 297 1119 527
rect 284 249 319 289
rect 284 215 809 249
rect 284 181 319 215
rect 858 181 1025 289
rect 29 147 319 181
rect 395 147 1025 181
rect 29 51 89 147
rect 123 17 179 113
rect 213 51 267 147
rect 301 17 361 113
rect 395 51 461 147
rect 495 17 549 113
rect 583 51 649 147
rect 683 17 737 113
rect 771 51 837 147
rect 871 17 925 113
rect 959 51 1025 147
rect 1059 17 1109 177
rect 0 -17 1196 17
<< via1 >>
rect 1046 518 1098 570
rect 1110 518 1162 570
rect 410 212 462 264
rect 474 212 526 264
rect 1046 -26 1098 26
rect 1110 -26 1162 26
<< obsm1 >>
rect 0 570 1196 592
rect 0 518 1046 570
rect 1098 518 1110 570
rect 1162 518 1196 570
rect 0 496 1196 518
rect 404 212 410 264
rect 462 212 474 264
rect 526 252 532 264
rect 849 252 979 261
rect 526 224 979 252
rect 526 212 532 224
rect 849 215 979 224
rect 0 26 1196 48
rect 0 -26 1046 26
rect 1098 -26 1110 26
rect 1162 -26 1196 26
rect 0 -48 1196 -26
<< via2 >>
rect 1036 570 1092 572
rect 1116 570 1172 572
rect 1036 518 1046 570
rect 1046 518 1092 570
rect 1116 518 1162 570
rect 1162 518 1172 570
rect 1036 516 1092 518
rect 1116 516 1172 518
rect 387 264 443 266
rect 467 264 523 266
rect 387 212 410 264
rect 410 212 443 264
rect 467 212 474 264
rect 474 212 523 264
rect 387 210 443 212
rect 467 210 523 212
rect 1036 26 1092 28
rect 1116 26 1172 28
rect 1036 -26 1046 26
rect 1046 -26 1092 26
rect 1116 -26 1162 26
rect 1162 -26 1172 26
rect 1036 -28 1092 -26
rect 1116 -28 1172 -26
<< obsm2 >>
rect 1027 516 1036 572
rect 1092 570 1116 572
rect 1098 518 1110 570
rect 1092 516 1116 518
rect 1172 516 1181 572
rect 378 210 387 266
rect 443 264 467 266
rect 523 264 532 266
rect 462 212 467 264
rect 526 212 532 264
rect 443 210 467 212
rect 523 210 532 212
rect 1027 -28 1036 28
rect 1092 26 1116 28
rect 1098 -26 1110 26
rect 1092 -28 1116 -26
rect 1172 -28 1181 28
<< obsm3 >>
rect 1026 576 1182 577
rect 1026 512 1032 576
rect 1096 512 1112 576
rect 1176 512 1182 576
rect 1026 511 1182 512
rect 377 270 533 271
rect -143 206 -137 270
rect -73 206 -57 270
rect 7 206 13 270
rect 377 206 383 270
rect 447 206 463 270
rect 527 206 533 270
rect 377 205 533 206
rect 1026 32 1182 33
rect 1026 -32 1032 32
rect 1096 -32 1112 32
rect 1176 -32 1182 32
rect 1026 -33 1182 -32
<< via3 >>
rect 1032 572 1096 576
rect 1032 516 1036 572
rect 1036 516 1092 572
rect 1092 516 1096 572
rect 1032 512 1096 516
rect 1112 572 1176 576
rect 1112 516 1116 572
rect 1116 516 1172 572
rect 1172 516 1176 572
rect 1112 512 1176 516
rect -137 206 -73 270
rect -57 206 7 270
rect 383 266 447 270
rect 383 210 387 266
rect 387 210 443 266
rect 443 210 447 266
rect 383 206 447 210
rect 463 266 527 270
rect 463 210 467 266
rect 467 210 523 266
rect 523 210 527 266
rect 463 206 527 210
rect 1032 28 1096 32
rect 1032 -28 1036 28
rect 1036 -28 1092 28
rect 1092 -28 1096 28
rect 1032 -32 1096 -28
rect 1112 28 1176 32
rect 1112 -28 1116 28
rect 1116 -28 1172 28
rect 1172 -28 1176 28
rect 1112 -32 1176 -28
<< metal4 >>
rect 986 576 1222 723
rect 986 512 1032 576
rect 1096 512 1112 576
rect 1176 512 1222 576
rect 986 487 1222 512
rect 986 32 1222 57
rect 986 -32 1032 32
rect 1096 -32 1112 32
rect 1176 -32 1222 32
rect 986 -179 1222 -32
<< obsm4 >>
rect -228 270 8 390
rect -228 206 -137 270
rect -73 206 -57 270
rect 7 206 8 270
rect -228 154 8 206
rect 292 270 528 390
rect 292 206 383 270
rect 447 206 463 270
rect 527 206 528 270
rect 292 154 528 206
<< metal5 >>
rect -252 112 212 432
rect 872 635 1335 778
rect 912 575 1335 635
rect 872 432 1335 575
rect 872 -31 1335 112
rect 912 -91 1335 -31
rect 872 -234 1335 -91
<< obsm5 >>
rect 232 -221 552 765
rect 872 595 892 615
rect 872 -71 892 -51
<< labels >>
rlabel locali s 28 215 248 255 6 A
port 1 nsew signal input
rlabel metal5 s -252 112 212 432 4 X
port 2 nsew signal output
rlabel metal4 s 986 -179 1222 57 8 VGND
port 3 nsew ground input
rlabel metal5 s 912 -91 1335 -31 8 VGND
port 3 nsew ground input
rlabel metal5 s 872 -31 1335 112 6 VGND
port 3 nsew ground input
rlabel metal5 s 872 -234 1335 -91 8 VGND
port 3 nsew ground input
rlabel metal4 s 986 487 1222 723 6 VPWR
port 4 nsew power input
rlabel metal5 s 912 575 1335 635 6 VPWR
port 4 nsew power input
rlabel metal5 s 872 635 1335 778 6 VPWR
port 4 nsew power input
rlabel metal5 s 872 432 1335 575 6 VPWR
port 4 nsew power input
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 178158
string GDS_START 165970
<< end >>
