magic
tech sky130A
magscale 1 2
timestamp 1599588238
<< locali >>
rect 114 378 170 596
rect 114 310 180 378
rect 145 210 180 310
rect 145 70 211 210
rect 313 236 398 307
rect 440 236 551 310
rect 585 236 651 310
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 24 364 74 649
rect 204 409 270 649
rect 308 375 358 596
rect 59 17 109 226
rect 214 341 358 375
rect 398 378 448 596
rect 488 412 554 649
rect 594 378 644 596
rect 398 344 644 378
rect 214 244 279 341
rect 245 202 279 244
rect 245 168 459 202
rect 245 17 359 134
rect 393 70 459 168
rect 573 17 639 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel locali s 440 236 551 310 6 A1
port 1 nsew signal input
rlabel locali s 585 236 651 310 6 A2
port 2 nsew signal input
rlabel locali s 313 236 398 307 6 B1
port 3 nsew signal input
rlabel locali s 145 210 180 310 6 X
port 4 nsew signal output
rlabel locali s 145 70 211 210 6 X
port 4 nsew signal output
rlabel locali s 114 378 170 596 6 X
port 4 nsew signal output
rlabel locali s 114 310 180 378 6 X
port 4 nsew signal output
rlabel metal1 s 0 -49 672 49 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 617 672 715 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 4005364
string GDS_START 3998422
<< end >>
