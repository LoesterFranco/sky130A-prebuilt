magic
tech sky130A
magscale 1 2
timestamp 1601050082
<< locali >>
rect 111 424 177 547
rect 25 390 177 424
rect 25 236 76 390
rect 285 390 647 424
rect 117 270 183 356
rect 285 336 319 390
rect 249 286 319 336
rect 389 286 455 356
rect 505 310 647 390
rect 681 390 1013 424
rect 537 286 603 310
rect 681 286 747 390
rect 979 356 1013 390
rect 793 286 935 356
rect 979 286 1127 356
rect 218 236 1086 252
rect 25 218 1086 236
rect 25 202 252 218
rect 25 70 76 202
rect 218 70 252 202
rect 590 70 636 218
rect 1036 70 1086 218
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 21 596 453 615
rect 21 581 633 596
rect 21 458 71 581
rect 217 370 251 581
rect 291 492 363 547
rect 403 526 633 581
rect 671 526 721 649
rect 761 492 827 596
rect 867 526 901 649
rect 941 492 1007 596
rect 291 458 1007 492
rect 1047 390 1097 649
rect 112 17 182 168
rect 288 150 556 184
rect 288 70 354 150
rect 388 17 456 116
rect 490 66 556 150
rect 670 150 1000 184
rect 670 66 806 150
rect 840 17 906 116
rect 940 66 1000 150
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
rlabel locali s 979 356 1013 390 6 A1
port 1 nsew signal input
rlabel locali s 979 286 1127 356 6 A1
port 1 nsew signal input
rlabel locali s 681 390 1013 424 6 A1
port 1 nsew signal input
rlabel locali s 681 286 747 390 6 A1
port 1 nsew signal input
rlabel locali s 793 286 935 356 6 A2
port 2 nsew signal input
rlabel locali s 537 286 603 310 6 B1
port 3 nsew signal input
rlabel locali s 505 310 647 390 6 B1
port 3 nsew signal input
rlabel locali s 285 390 647 424 6 B1
port 3 nsew signal input
rlabel locali s 285 336 319 390 6 B1
port 3 nsew signal input
rlabel locali s 249 286 319 336 6 B1
port 3 nsew signal input
rlabel locali s 389 286 455 356 6 B2
port 4 nsew signal input
rlabel locali s 117 270 183 356 6 C1
port 5 nsew signal input
rlabel locali s 1036 70 1086 218 6 Y
port 6 nsew signal output
rlabel locali s 590 70 636 218 6 Y
port 6 nsew signal output
rlabel locali s 218 236 1086 252 6 Y
port 6 nsew signal output
rlabel locali s 218 70 252 202 6 Y
port 6 nsew signal output
rlabel locali s 111 424 177 547 6 Y
port 6 nsew signal output
rlabel locali s 25 390 177 424 6 Y
port 6 nsew signal output
rlabel locali s 25 236 76 390 6 Y
port 6 nsew signal output
rlabel locali s 25 218 1086 236 6 Y
port 6 nsew signal output
rlabel locali s 25 202 252 218 6 Y
port 6 nsew signal output
rlabel locali s 25 70 76 202 6 Y
port 6 nsew signal output
rlabel metal1 s 0 -49 1152 49 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1152 715 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 4128748
string GDS_START 4118786
<< end >>
