magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 17 288 122 493
rect 17 185 80 288
rect 17 70 118 185
rect 392 199 529 265
rect 1417 289 1543 345
rect 1417 199 1461 289
rect 1601 215 1739 265
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 166 443 233 527
rect 270 447 609 481
rect 662 447 743 481
rect 777 447 843 527
rect 930 455 1589 489
rect 1671 455 1810 527
rect 270 409 314 447
rect 709 413 743 447
rect 930 413 964 455
rect 160 375 314 409
rect 394 379 675 413
rect 709 379 964 413
rect 160 173 200 375
rect 247 307 597 341
rect 160 139 290 173
rect 162 17 212 105
rect 246 85 290 139
rect 324 119 358 307
rect 563 265 597 307
rect 641 339 675 379
rect 641 305 747 339
rect 690 275 747 305
rect 563 199 628 265
rect 414 131 656 165
rect 498 85 578 91
rect 246 51 578 85
rect 612 85 656 131
rect 690 119 724 275
rect 781 241 815 379
rect 861 289 964 343
rect 758 207 815 241
rect 758 85 792 207
rect 612 51 792 85
rect 826 17 860 173
rect 906 83 964 289
rect 999 119 1033 421
rect 1067 178 1101 455
rect 1854 421 1913 493
rect 1149 323 1232 409
rect 1349 387 1913 421
rect 1149 289 1315 323
rect 1152 199 1237 254
rect 1067 165 1121 178
rect 1067 144 1160 165
rect 1077 131 1160 144
rect 999 97 1043 119
rect 999 53 1082 97
rect 1126 64 1160 131
rect 1194 126 1237 199
rect 1281 85 1315 289
rect 1349 119 1383 387
rect 1806 375 1913 387
rect 1587 299 1823 341
rect 1789 265 1823 299
rect 1495 189 1557 255
rect 1789 199 1845 265
rect 1495 146 1536 189
rect 1789 181 1823 199
rect 1603 150 1823 181
rect 1595 147 1823 150
rect 1417 85 1520 93
rect 1281 51 1520 85
rect 1595 59 1653 147
rect 1879 117 1913 375
rect 1697 17 1787 113
rect 1853 51 1913 117
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< obsm1 >>
rect 701 320 759 329
rect 1191 320 1249 329
rect 701 292 1249 320
rect 701 283 759 292
rect 1191 283 1249 292
rect 895 184 953 193
rect 1191 184 1249 193
rect 1487 184 1545 193
rect 895 156 1545 184
rect 895 147 953 156
rect 1191 147 1249 156
rect 1487 147 1545 156
rect 997 116 1055 125
rect 1589 116 1647 125
rect 997 88 1647 116
rect 997 79 1055 88
rect 1589 79 1647 88
<< labels >>
rlabel locali s 1601 215 1739 265 6 A
port 1 nsew signal input
rlabel locali s 1417 289 1543 345 6 B
port 2 nsew signal input
rlabel locali s 1417 199 1461 289 6 B
port 2 nsew signal input
rlabel locali s 392 199 529 265 6 C
port 3 nsew signal input
rlabel locali s 17 288 122 493 6 X
port 4 nsew signal output
rlabel locali s 17 185 80 288 6 X
port 4 nsew signal output
rlabel locali s 17 70 118 185 6 X
port 4 nsew signal output
rlabel metal1 s 0 -48 1932 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 1932 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1932 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 793102
string GDS_START 780618
<< end >>
