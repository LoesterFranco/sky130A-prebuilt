magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 1326 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 79 47 109 177
rect 183 47 213 177
rect 267 47 297 177
rect 371 47 401 177
rect 455 47 485 177
rect 673 47 703 177
rect 757 47 787 177
rect 861 47 891 177
rect 1049 47 1079 177
rect 1143 47 1173 177
<< pmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 583 297 619 497
rect 677 297 713 497
rect 771 297 807 497
rect 865 297 901 497
rect 1067 297 1103 497
rect 1161 297 1197 497
<< ndiff >>
rect 27 165 79 177
rect 27 131 35 165
rect 69 131 79 165
rect 27 93 79 131
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 165 183 177
rect 109 131 129 165
rect 163 131 183 165
rect 109 47 183 131
rect 213 93 267 177
rect 213 59 223 93
rect 257 59 267 93
rect 213 47 267 59
rect 297 165 371 177
rect 297 131 317 165
rect 351 131 371 165
rect 297 47 371 131
rect 401 93 455 177
rect 401 59 411 93
rect 445 59 455 93
rect 401 47 455 59
rect 485 93 673 177
rect 485 59 590 93
rect 624 59 673 93
rect 485 47 673 59
rect 703 165 757 177
rect 703 131 713 165
rect 747 131 757 165
rect 703 93 757 131
rect 703 59 713 93
rect 747 59 757 93
rect 703 47 757 59
rect 787 93 861 177
rect 787 59 807 93
rect 841 59 861 93
rect 787 47 861 59
rect 891 165 1049 177
rect 891 131 917 165
rect 951 131 985 165
rect 1019 131 1049 165
rect 891 93 1049 131
rect 891 59 917 93
rect 951 59 985 93
rect 1019 59 1049 93
rect 891 47 1049 59
rect 1079 93 1143 177
rect 1079 59 1099 93
rect 1133 59 1143 93
rect 1079 47 1143 59
rect 1173 165 1253 177
rect 1173 131 1211 165
rect 1245 131 1253 165
rect 1173 93 1253 131
rect 1173 59 1211 93
rect 1245 59 1253 93
rect 1173 47 1253 59
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 417 175 497
rect 117 383 129 417
rect 163 383 175 417
rect 117 349 175 383
rect 117 315 129 349
rect 163 315 175 349
rect 117 297 175 315
rect 211 485 269 497
rect 211 451 223 485
rect 257 451 269 485
rect 211 417 269 451
rect 211 383 223 417
rect 257 383 269 417
rect 211 297 269 383
rect 305 485 363 497
rect 305 451 317 485
rect 351 451 363 485
rect 305 297 363 451
rect 399 485 453 497
rect 399 451 411 485
rect 445 451 453 485
rect 399 417 453 451
rect 399 383 411 417
rect 445 383 453 417
rect 399 297 453 383
rect 525 485 583 497
rect 525 451 533 485
rect 567 451 583 485
rect 525 417 583 451
rect 525 383 533 417
rect 567 383 583 417
rect 525 297 583 383
rect 619 417 677 497
rect 619 383 631 417
rect 665 383 677 417
rect 619 349 677 383
rect 619 315 631 349
rect 665 315 677 349
rect 619 297 677 315
rect 713 485 771 497
rect 713 451 725 485
rect 759 451 771 485
rect 713 417 771 451
rect 713 383 725 417
rect 759 383 771 417
rect 713 349 771 383
rect 713 315 725 349
rect 759 315 771 349
rect 713 297 771 315
rect 807 417 865 497
rect 807 383 819 417
rect 853 383 865 417
rect 807 349 865 383
rect 807 315 819 349
rect 853 315 865 349
rect 807 297 865 315
rect 901 485 959 497
rect 901 451 917 485
rect 951 451 959 485
rect 901 417 959 451
rect 901 383 917 417
rect 951 383 959 417
rect 901 297 959 383
rect 1013 485 1067 497
rect 1013 451 1021 485
rect 1055 451 1067 485
rect 1013 417 1067 451
rect 1013 383 1021 417
rect 1055 383 1067 417
rect 1013 297 1067 383
rect 1103 485 1161 497
rect 1103 451 1115 485
rect 1149 451 1161 485
rect 1103 417 1161 451
rect 1103 383 1115 417
rect 1149 383 1161 417
rect 1103 349 1161 383
rect 1103 315 1115 349
rect 1149 315 1161 349
rect 1103 297 1161 315
rect 1197 485 1255 497
rect 1197 451 1213 485
rect 1247 451 1255 485
rect 1197 417 1255 451
rect 1197 383 1213 417
rect 1247 383 1255 417
rect 1197 349 1255 383
rect 1197 315 1213 349
rect 1247 315 1255 349
rect 1197 297 1255 315
<< ndiffc >>
rect 35 131 69 165
rect 35 59 69 93
rect 129 131 163 165
rect 223 59 257 93
rect 317 131 351 165
rect 411 59 445 93
rect 590 59 624 93
rect 713 131 747 165
rect 713 59 747 93
rect 807 59 841 93
rect 917 131 951 165
rect 985 131 1019 165
rect 917 59 951 93
rect 985 59 1019 93
rect 1099 59 1133 93
rect 1211 131 1245 165
rect 1211 59 1245 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 383 163 417
rect 129 315 163 349
rect 223 451 257 485
rect 223 383 257 417
rect 317 451 351 485
rect 411 451 445 485
rect 411 383 445 417
rect 533 451 567 485
rect 533 383 567 417
rect 631 383 665 417
rect 631 315 665 349
rect 725 451 759 485
rect 725 383 759 417
rect 725 315 759 349
rect 819 383 853 417
rect 819 315 853 349
rect 917 451 951 485
rect 917 383 951 417
rect 1021 451 1055 485
rect 1021 383 1055 417
rect 1115 451 1149 485
rect 1115 383 1149 417
rect 1115 315 1149 349
rect 1213 451 1247 485
rect 1213 383 1247 417
rect 1213 315 1247 349
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 583 497 619 523
rect 677 497 713 523
rect 771 497 807 523
rect 865 497 901 523
rect 1067 497 1103 523
rect 1161 497 1197 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 583 282 619 297
rect 677 282 713 297
rect 771 282 807 297
rect 865 282 901 297
rect 1067 282 1103 297
rect 1161 282 1197 297
rect 79 265 119 282
rect 173 265 213 282
rect 79 249 213 265
rect 79 215 129 249
rect 163 215 213 249
rect 79 199 213 215
rect 79 177 109 199
rect 183 177 213 199
rect 267 265 307 282
rect 361 265 401 282
rect 267 249 401 265
rect 581 265 621 282
rect 675 265 715 282
rect 769 265 809 282
rect 863 265 903 282
rect 1065 265 1105 282
rect 1159 265 1199 282
rect 581 253 715 265
rect 267 215 297 249
rect 331 215 401 249
rect 267 199 401 215
rect 267 177 297 199
rect 371 177 401 199
rect 455 249 715 253
rect 455 223 623 249
rect 455 177 485 223
rect 581 215 623 223
rect 657 215 715 249
rect 581 199 715 215
rect 757 249 903 265
rect 757 215 811 249
rect 845 215 903 249
rect 757 199 903 215
rect 1049 249 1199 265
rect 1049 215 1101 249
rect 1135 215 1199 249
rect 1049 199 1199 215
rect 673 177 703 199
rect 757 177 787 199
rect 861 177 891 199
rect 1049 177 1079 199
rect 1143 177 1173 199
rect 79 21 109 47
rect 183 21 213 47
rect 267 21 297 47
rect 371 21 401 47
rect 455 21 485 47
rect 673 21 703 47
rect 757 21 787 47
rect 861 21 891 47
rect 1049 21 1079 47
rect 1143 21 1173 47
<< polycont >>
rect 129 215 163 249
rect 297 215 331 249
rect 623 215 657 249
rect 811 215 845 249
rect 1101 215 1135 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 18 485 273 493
rect 18 451 35 485
rect 69 459 223 485
rect 18 417 69 451
rect 257 451 273 485
rect 18 383 35 417
rect 18 349 69 383
rect 18 315 35 349
rect 18 299 69 315
rect 103 417 179 419
rect 103 383 129 417
rect 163 383 179 417
rect 103 349 179 383
rect 223 417 273 451
rect 317 485 351 527
rect 317 435 351 451
rect 385 485 461 491
rect 385 451 411 485
rect 445 451 461 485
rect 257 401 273 417
rect 385 417 461 451
rect 385 401 411 417
rect 257 383 411 401
rect 445 383 461 417
rect 223 367 461 383
rect 517 485 967 489
rect 517 451 533 485
rect 567 451 725 485
rect 759 451 917 485
rect 951 451 967 485
rect 517 417 567 451
rect 725 417 759 451
rect 917 417 967 451
rect 517 383 533 417
rect 517 367 567 383
rect 605 383 631 417
rect 665 383 681 417
rect 103 315 129 349
rect 163 333 179 349
rect 605 349 681 383
rect 605 333 631 349
rect 163 315 631 333
rect 665 315 681 349
rect 103 299 681 315
rect 725 349 759 383
rect 725 299 759 315
rect 803 383 819 417
rect 853 383 869 417
rect 803 349 869 383
rect 951 383 967 417
rect 917 367 967 383
rect 1014 485 1055 527
rect 1014 451 1021 485
rect 1014 417 1055 451
rect 1014 383 1021 417
rect 1014 367 1055 383
rect 1099 485 1165 492
rect 1099 451 1115 485
rect 1149 451 1165 485
rect 1099 417 1165 451
rect 1099 383 1115 417
rect 1149 383 1165 417
rect 803 315 819 349
rect 853 333 869 349
rect 1099 349 1165 383
rect 1099 333 1115 349
rect 853 315 1115 333
rect 1149 315 1165 349
rect 803 299 1165 315
rect 1209 485 1253 527
rect 1209 451 1213 485
rect 1247 451 1253 485
rect 1209 417 1253 451
rect 1209 383 1213 417
rect 1247 383 1253 417
rect 1209 349 1253 383
rect 1209 315 1213 349
rect 1247 315 1253 349
rect 1209 299 1253 315
rect 18 249 179 265
rect 18 215 129 249
rect 163 215 179 249
rect 213 249 363 265
rect 213 215 297 249
rect 331 215 363 249
rect 397 221 474 299
rect 531 249 673 265
rect 397 181 449 221
rect 531 215 623 249
rect 657 215 673 249
rect 744 249 986 265
rect 744 215 811 249
rect 845 215 986 249
rect 1040 249 1259 265
rect 1040 215 1101 249
rect 1135 215 1259 249
rect 18 165 69 181
rect 18 131 35 165
rect 103 165 449 181
rect 103 131 129 165
rect 163 131 317 165
rect 351 131 449 165
rect 497 165 1261 181
rect 497 143 713 165
rect 18 97 69 131
rect 497 97 531 143
rect 687 131 713 143
rect 747 143 917 165
rect 747 131 763 143
rect 18 93 531 97
rect 18 59 35 93
rect 69 59 223 93
rect 257 59 411 93
rect 445 59 531 93
rect 18 51 531 59
rect 574 93 650 109
rect 574 59 590 93
rect 624 59 650 93
rect 574 17 650 59
rect 687 93 763 131
rect 901 131 917 143
rect 951 131 985 165
rect 1019 143 1211 165
rect 1019 131 1035 143
rect 687 59 713 93
rect 747 59 763 93
rect 687 51 763 59
rect 807 93 841 109
rect 807 17 841 59
rect 901 93 1035 131
rect 1195 131 1211 143
rect 1245 131 1261 165
rect 901 59 917 93
rect 951 59 985 93
rect 1019 59 1035 93
rect 901 51 1035 59
rect 1071 93 1147 109
rect 1071 59 1099 93
rect 1133 59 1147 93
rect 1071 17 1147 59
rect 1195 93 1261 131
rect 1195 59 1211 93
rect 1245 59 1261 93
rect 1195 51 1261 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
flabel corelocali s 1130 221 1164 255 0 FreeSans 250 0 0 0 A1
port 1 nsew
flabel corelocali s 217 221 251 255 0 FreeSans 250 0 0 0 B1
port 4 nsew
flabel corelocali s 857 221 891 255 0 FreeSans 250 0 0 0 A2
port 2 nsew
flabel corelocali s 1040 221 1074 255 0 FreeSans 250 0 0 0 A1
port 1 nsew
flabel corelocali s 766 221 800 255 0 FreeSans 250 0 0 0 A2
port 2 nsew
flabel corelocali s 584 221 618 255 0 FreeSans 250 0 0 0 A3
port 3 nsew
flabel corelocali s 400 221 434 255 0 FreeSans 250 0 0 0 Y
port 10 nsew
flabel corelocali s 401 289 435 323 0 FreeSans 250 0 0 0 Y
port 10 nsew
flabel corelocali s 306 221 340 255 0 FreeSans 250 0 0 0 B1
port 4 nsew
flabel corelocali s 121 221 155 255 0 FreeSans 250 0 0 0 B2
port 5 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 250 0 0 0 B2
port 5 nsew
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew
rlabel comment s 0 0 0 0 4 o32ai_2
<< properties >>
string FIXED_BBOX 0 0 1288 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 591166
string GDS_START 580822
<< end >>
