magic
tech sky130A
magscale 1 2
timestamp 1601050082
<< locali >>
rect 99 294 165 360
rect 307 294 373 360
rect 985 284 1059 356
rect 1177 290 1415 356
rect 1449 290 1515 356
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 241 596 487 615
rect 61 581 487 596
rect 61 540 307 581
rect 25 472 301 506
rect 25 208 59 472
rect 151 404 233 438
rect 199 260 233 404
rect 267 428 301 472
rect 347 498 381 547
rect 421 532 487 581
rect 525 532 591 649
rect 705 532 771 649
rect 885 532 951 649
rect 988 498 1054 596
rect 1094 526 1144 649
rect 347 492 1054 498
rect 1184 492 1218 596
rect 347 464 1218 492
rect 347 462 381 464
rect 988 458 1218 464
rect 1258 458 1330 649
rect 505 428 861 430
rect 267 394 861 428
rect 1184 424 1218 458
rect 1370 424 1404 596
rect 505 364 861 394
rect 895 390 1143 424
rect 1184 390 1404 424
rect 1444 390 1510 649
rect 895 330 929 390
rect 411 296 929 330
rect 411 264 781 296
rect 411 260 465 264
rect 181 226 465 260
rect 1109 253 1143 390
rect 835 230 1035 237
rect 25 202 71 208
rect 25 168 31 202
rect 65 168 71 202
rect 25 162 71 168
rect 79 17 145 128
rect 181 78 217 226
rect 251 17 317 192
rect 351 78 387 226
rect 507 202 749 230
rect 423 17 473 192
rect 507 168 511 202
rect 545 196 749 202
rect 545 168 584 196
rect 507 78 584 168
rect 620 17 663 162
rect 699 81 749 196
rect 785 187 1035 230
rect 1109 187 1221 253
rect 1257 197 1507 249
rect 785 17 835 187
rect 1355 153 1421 163
rect 883 119 1421 153
rect 883 101 949 119
rect 1457 85 1507 197
rect 1073 51 1507 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 31 168 65 202
rect 511 168 545 202
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 19 202 77 208
rect 19 168 31 202
rect 65 199 77 202
rect 499 202 557 208
rect 499 199 511 202
rect 65 171 511 199
rect 65 168 77 171
rect 19 162 77 168
rect 499 168 511 171
rect 545 168 557 202
rect 499 162 557 168
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
rlabel locali s 1177 290 1415 356 6 A1
port 1 nsew signal input
rlabel locali s 1449 290 1515 356 6 A2
port 2 nsew signal input
rlabel locali s 985 284 1059 356 6 A3
port 3 nsew signal input
rlabel locali s 307 294 373 360 6 B1
port 4 nsew signal input
rlabel locali s 99 294 165 360 6 C1
port 5 nsew signal input
rlabel metal1 s 499 199 557 208 6 X
port 6 nsew signal output
rlabel metal1 s 499 162 557 171 6 X
port 6 nsew signal output
rlabel metal1 s 19 199 77 208 6 X
port 6 nsew signal output
rlabel metal1 s 19 171 557 199 6 X
port 6 nsew signal output
rlabel metal1 s 19 162 77 171 6 X
port 6 nsew signal output
rlabel metal1 s 0 -49 1536 49 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1536 715 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1536 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3594508
string GDS_START 3582222
<< end >>
