magic
tech sky130A
magscale 1 2
timestamp 1599588232
<< locali >>
rect 25 290 114 356
rect 162 290 257 356
rect 399 295 465 361
rect 505 295 573 361
rect 685 364 754 596
rect 720 226 754 364
rect 686 70 754 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 24 390 90 649
rect 210 513 276 596
rect 317 547 388 649
rect 554 547 644 649
rect 210 479 651 513
rect 210 390 276 479
rect 323 395 513 445
rect 323 356 357 395
rect 291 290 357 356
rect 617 327 651 479
rect 791 364 841 649
rect 323 261 357 290
rect 617 261 686 327
rect 23 222 261 256
rect 323 227 475 261
rect 23 70 73 222
rect 109 17 175 188
rect 211 70 261 222
rect 295 85 361 193
rect 409 119 475 227
rect 509 227 651 261
rect 509 85 543 227
rect 295 51 543 85
rect 577 17 643 193
rect 788 17 838 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel locali s 505 295 573 361 6 A1_N
port 1 nsew signal input
rlabel locali s 399 295 465 361 6 A2_N
port 2 nsew signal input
rlabel locali s 25 290 114 356 6 B1
port 3 nsew signal input
rlabel locali s 162 290 257 356 6 B2
port 4 nsew signal input
rlabel locali s 720 226 754 364 6 X
port 5 nsew signal output
rlabel locali s 686 70 754 226 6 X
port 5 nsew signal output
rlabel locali s 685 364 754 596 6 X
port 5 nsew signal output
rlabel metal1 s 0 -49 864 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 7 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 617 864 715 6 VPWR
port 9 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1252868
string GDS_START 1244816
<< end >>
