magic
tech sky130A
magscale 1 2
timestamp 1604502710
<< nwell >>
rect -38 351 2342 704
rect -38 332 272 351
rect 607 332 2342 351
rect 607 324 1412 332
rect 1108 311 1412 324
<< pwell >>
rect 0 0 2304 49
<< scpmos >>
rect 83 508 119 592
rect 173 508 209 592
rect 375 387 411 611
rect 465 387 501 611
rect 673 463 709 547
rect 763 463 799 547
rect 841 463 877 547
rect 968 463 1004 547
rect 1200 347 1236 547
rect 1290 347 1326 547
rect 1432 471 1468 555
rect 1516 471 1552 555
rect 1618 471 1654 555
rect 1708 471 1744 555
rect 1811 368 1847 592
rect 2082 424 2118 592
rect 2185 368 2221 592
<< nmoslvt >>
rect 95 78 125 162
rect 173 78 203 162
rect 384 119 414 267
rect 488 119 518 267
rect 702 119 732 203
rect 802 119 832 203
rect 880 119 910 203
rect 958 119 988 203
rect 1076 74 1106 202
rect 1194 74 1224 202
rect 1404 74 1434 158
rect 1482 74 1512 158
rect 1594 74 1624 158
rect 1672 74 1702 158
rect 1873 74 1903 222
rect 2088 74 2118 184
rect 2188 74 2218 222
<< ndiff >>
rect 318 228 384 267
rect 318 194 330 228
rect 364 194 384 228
rect 38 137 95 162
rect 38 103 50 137
rect 84 103 95 137
rect 38 78 95 103
rect 125 78 173 162
rect 203 137 264 162
rect 203 103 222 137
rect 256 103 264 137
rect 318 160 384 194
rect 318 126 330 160
rect 364 126 384 160
rect 318 119 384 126
rect 414 160 488 267
rect 414 126 434 160
rect 468 126 488 160
rect 414 119 488 126
rect 518 222 568 267
rect 518 161 584 222
rect 518 127 534 161
rect 568 127 584 161
rect 518 119 584 127
rect 645 179 702 203
rect 645 145 657 179
rect 691 145 702 179
rect 645 119 702 145
rect 732 179 802 203
rect 732 145 757 179
rect 791 145 802 179
rect 732 119 802 145
rect 832 119 880 203
rect 910 119 958 203
rect 988 202 1045 203
rect 1121 218 1179 230
rect 1121 202 1133 218
rect 988 119 1076 202
rect 318 118 369 119
rect 203 78 264 103
rect 429 118 473 119
rect 1003 82 1076 119
rect 1003 48 1015 82
rect 1049 74 1076 82
rect 1106 184 1133 202
rect 1167 202 1179 218
rect 1167 184 1194 202
rect 1106 74 1194 184
rect 1224 158 1274 202
rect 1816 210 1873 222
rect 1816 176 1828 210
rect 1862 176 1873 210
rect 1224 130 1404 158
rect 1224 96 1322 130
rect 1356 96 1404 130
rect 1224 74 1404 96
rect 1434 74 1482 158
rect 1512 128 1594 158
rect 1512 94 1536 128
rect 1570 94 1594 128
rect 1512 74 1594 94
rect 1624 74 1672 158
rect 1702 133 1759 158
rect 1702 99 1713 133
rect 1747 99 1759 133
rect 1702 74 1759 99
rect 1816 120 1873 176
rect 1816 86 1828 120
rect 1862 86 1873 120
rect 1816 74 1873 86
rect 1903 210 1974 222
rect 1903 176 1928 210
rect 1962 176 1974 210
rect 2133 210 2188 222
rect 2133 184 2141 210
rect 1903 120 1974 176
rect 1903 86 1928 120
rect 1962 86 1974 120
rect 1903 74 1974 86
rect 2031 145 2088 184
rect 2031 111 2043 145
rect 2077 111 2088 145
rect 2031 74 2088 111
rect 2118 176 2141 184
rect 2175 176 2188 210
rect 2118 120 2188 176
rect 2118 86 2141 120
rect 2175 86 2188 120
rect 2118 74 2188 86
rect 2218 210 2275 222
rect 2218 176 2229 210
rect 2263 176 2275 210
rect 2218 120 2275 176
rect 2218 86 2229 120
rect 2263 86 2275 120
rect 2218 74 2275 86
rect 1049 48 1061 74
rect 1003 36 1061 48
<< pdiff >>
rect 27 567 83 592
rect 27 533 39 567
rect 73 533 83 567
rect 27 508 83 533
rect 119 567 173 592
rect 119 533 129 567
rect 163 533 173 567
rect 119 508 173 533
rect 209 584 265 592
rect 209 550 219 584
rect 253 550 265 584
rect 209 508 265 550
rect 319 462 375 611
rect 307 437 375 462
rect 307 403 315 437
rect 349 403 375 437
rect 307 387 375 403
rect 411 584 465 611
rect 411 550 421 584
rect 455 550 465 584
rect 411 387 465 550
rect 501 437 557 611
rect 501 403 511 437
rect 545 403 557 437
rect 501 387 557 403
rect 892 585 953 597
rect 892 551 905 585
rect 939 551 953 585
rect 892 547 953 551
rect 1759 567 1811 592
rect 1759 555 1767 567
rect 1382 547 1432 555
rect 617 522 673 547
rect 617 488 629 522
rect 663 488 673 522
rect 617 463 673 488
rect 709 539 763 547
rect 709 505 719 539
rect 753 505 763 539
rect 709 463 763 505
rect 799 463 841 547
rect 877 463 968 547
rect 1004 520 1057 547
rect 1004 486 1015 520
rect 1049 486 1057 520
rect 1004 463 1057 486
rect 1144 535 1200 547
rect 1144 501 1156 535
rect 1190 501 1200 535
rect 1144 466 1200 501
rect 1144 432 1156 466
rect 1190 432 1200 466
rect 1144 398 1200 432
rect 1144 364 1156 398
rect 1190 364 1200 398
rect 1144 347 1200 364
rect 1236 535 1290 547
rect 1236 501 1246 535
rect 1280 501 1290 535
rect 1236 464 1290 501
rect 1236 430 1246 464
rect 1280 430 1290 464
rect 1236 393 1290 430
rect 1236 359 1246 393
rect 1280 359 1290 393
rect 1236 347 1290 359
rect 1326 523 1432 547
rect 1326 489 1361 523
rect 1395 489 1432 523
rect 1326 471 1432 489
rect 1468 471 1516 555
rect 1552 530 1618 555
rect 1552 496 1567 530
rect 1601 496 1618 530
rect 1552 471 1618 496
rect 1654 530 1708 555
rect 1654 496 1664 530
rect 1698 496 1708 530
rect 1654 471 1708 496
rect 1744 533 1767 555
rect 1801 533 1811 567
rect 1744 471 1811 533
rect 1326 347 1376 471
rect 1759 437 1767 471
rect 1801 437 1811 471
rect 1759 368 1811 437
rect 1847 580 1967 592
rect 1847 546 1857 580
rect 1891 546 1925 580
rect 1959 546 1967 580
rect 1847 497 1967 546
rect 1847 463 1857 497
rect 1891 463 1925 497
rect 1959 463 1967 497
rect 1847 414 1967 463
rect 2026 579 2082 592
rect 2026 545 2038 579
rect 2072 545 2082 579
rect 2026 471 2082 545
rect 2026 437 2038 471
rect 2072 437 2082 471
rect 2026 424 2082 437
rect 2118 580 2185 592
rect 2118 546 2135 580
rect 2169 546 2185 580
rect 2118 497 2185 546
rect 2118 463 2135 497
rect 2169 463 2185 497
rect 2118 424 2185 463
rect 1847 380 1857 414
rect 1891 380 1925 414
rect 1959 380 1967 414
rect 1847 368 1967 380
rect 2133 414 2185 424
rect 2133 380 2141 414
rect 2175 380 2185 414
rect 2133 368 2185 380
rect 2221 580 2277 592
rect 2221 546 2231 580
rect 2265 546 2277 580
rect 2221 497 2277 546
rect 2221 463 2231 497
rect 2265 463 2277 497
rect 2221 414 2277 463
rect 2221 380 2231 414
rect 2265 380 2277 414
rect 2221 368 2277 380
<< ndiffc >>
rect 330 194 364 228
rect 50 103 84 137
rect 222 103 256 137
rect 330 126 364 160
rect 434 126 468 160
rect 534 127 568 161
rect 657 145 691 179
rect 757 145 791 179
rect 1015 48 1049 82
rect 1133 184 1167 218
rect 1828 176 1862 210
rect 1322 96 1356 130
rect 1536 94 1570 128
rect 1713 99 1747 133
rect 1828 86 1862 120
rect 1928 176 1962 210
rect 1928 86 1962 120
rect 2043 111 2077 145
rect 2141 176 2175 210
rect 2141 86 2175 120
rect 2229 176 2263 210
rect 2229 86 2263 120
<< pdiffc >>
rect 39 533 73 567
rect 129 533 163 567
rect 219 550 253 584
rect 315 403 349 437
rect 421 550 455 584
rect 511 403 545 437
rect 905 551 939 585
rect 629 488 663 522
rect 719 505 753 539
rect 1015 486 1049 520
rect 1156 501 1190 535
rect 1156 432 1190 466
rect 1156 364 1190 398
rect 1246 501 1280 535
rect 1246 430 1280 464
rect 1246 359 1280 393
rect 1361 489 1395 523
rect 1567 496 1601 530
rect 1664 496 1698 530
rect 1767 533 1801 567
rect 1767 437 1801 471
rect 1857 546 1891 580
rect 1925 546 1959 580
rect 1857 463 1891 497
rect 1925 463 1959 497
rect 2038 545 2072 579
rect 2038 437 2072 471
rect 2135 546 2169 580
rect 2135 463 2169 497
rect 1857 380 1891 414
rect 1925 380 1959 414
rect 2141 380 2175 414
rect 2231 546 2265 580
rect 2231 463 2265 497
rect 2231 380 2265 414
<< poly >>
rect 83 592 119 618
rect 173 592 209 618
rect 375 611 411 637
rect 465 611 501 637
rect 572 615 1326 645
rect 83 470 119 508
rect 44 386 125 470
rect 44 352 60 386
rect 94 352 125 386
rect 44 318 125 352
rect 44 284 60 318
rect 94 284 125 318
rect 44 250 125 284
rect 44 216 60 250
rect 94 216 125 250
rect 44 200 125 216
rect 95 162 125 200
rect 173 428 209 508
rect 173 412 266 428
rect 173 378 216 412
rect 250 378 266 412
rect 572 440 602 615
rect 673 547 709 573
rect 763 547 799 615
rect 841 547 877 573
rect 968 547 1004 573
rect 1200 547 1236 573
rect 1290 547 1326 615
rect 1811 592 1847 618
rect 2082 592 2118 618
rect 2185 592 2221 618
rect 1432 555 1468 581
rect 1516 555 1552 581
rect 1618 555 1654 581
rect 1708 555 1744 581
rect 173 344 266 378
rect 375 355 411 387
rect 465 355 501 387
rect 572 355 608 440
rect 673 403 709 463
rect 763 437 799 463
rect 841 431 877 463
rect 968 431 1004 463
rect 841 415 926 431
rect 173 310 216 344
rect 250 310 266 344
rect 173 276 266 310
rect 357 339 423 355
rect 357 305 373 339
rect 407 305 423 339
rect 357 289 423 305
rect 465 339 608 355
rect 465 305 495 339
rect 529 307 608 339
rect 650 387 716 403
rect 841 401 876 415
rect 650 353 666 387
rect 700 367 716 387
rect 860 381 876 401
rect 910 381 926 415
rect 700 353 810 367
rect 650 337 810 353
rect 529 305 620 307
rect 465 295 620 305
rect 173 242 216 276
rect 250 242 266 276
rect 384 267 414 289
rect 465 282 732 295
rect 488 267 518 282
rect 579 278 732 282
rect 173 226 266 242
rect 173 162 203 226
rect 583 265 732 278
rect 702 203 732 265
rect 780 249 810 337
rect 860 347 926 381
rect 860 313 876 347
rect 910 313 926 347
rect 860 297 926 313
rect 968 415 1112 431
rect 968 381 1062 415
rect 1096 381 1112 415
rect 968 365 1112 381
rect 780 219 832 249
rect 802 203 832 219
rect 880 203 910 297
rect 968 248 998 365
rect 1432 439 1468 471
rect 1408 423 1474 439
rect 1408 389 1424 423
rect 1458 389 1474 423
rect 1408 373 1474 389
rect 1200 323 1236 347
rect 1046 307 1236 323
rect 1046 273 1062 307
rect 1096 293 1236 307
rect 1290 325 1326 347
rect 1290 295 1434 325
rect 1096 273 1112 293
rect 1046 257 1112 273
rect 958 218 998 248
rect 958 203 988 218
rect 1076 202 1106 257
rect 1194 230 1362 247
rect 384 93 414 119
rect 488 93 518 119
rect 702 93 732 119
rect 802 93 832 119
rect 880 93 910 119
rect 95 52 125 78
rect 173 51 203 78
rect 958 51 988 119
rect 173 21 988 51
rect 1194 217 1312 230
rect 1194 202 1224 217
rect 1296 196 1312 217
rect 1346 196 1362 230
rect 1296 180 1362 196
rect 1404 158 1434 295
rect 1516 246 1552 471
rect 1618 433 1654 471
rect 1482 230 1552 246
rect 1482 196 1502 230
rect 1536 196 1552 230
rect 1482 180 1552 196
rect 1594 417 1660 433
rect 1594 383 1610 417
rect 1644 383 1660 417
rect 1594 367 1660 383
rect 1482 158 1512 180
rect 1594 158 1624 367
rect 1708 319 1744 471
rect 1811 319 1847 368
rect 2082 319 2118 424
rect 2185 326 2221 368
rect 1666 303 2118 319
rect 1666 269 1682 303
rect 1716 269 2118 303
rect 1666 253 2118 269
rect 2160 310 2226 326
rect 2160 276 2176 310
rect 2210 276 2226 310
rect 2160 260 2226 276
rect 1672 158 1702 253
rect 1873 222 1903 253
rect 2088 184 2118 253
rect 2188 222 2218 260
rect 1076 48 1106 74
rect 1194 48 1224 74
rect 1404 48 1434 74
rect 1482 48 1512 74
rect 1594 48 1624 74
rect 1672 48 1702 74
rect 1873 48 1903 74
rect 2088 48 2118 74
rect 2188 48 2218 74
<< polycont >>
rect 60 352 94 386
rect 60 284 94 318
rect 60 216 94 250
rect 216 378 250 412
rect 216 310 250 344
rect 373 305 407 339
rect 495 305 529 339
rect 666 353 700 387
rect 876 381 910 415
rect 216 242 250 276
rect 876 313 910 347
rect 1062 381 1096 415
rect 1424 389 1458 423
rect 1062 273 1096 307
rect 1312 196 1346 230
rect 1502 196 1536 230
rect 1610 383 1644 417
rect 1682 269 1716 303
rect 2176 276 2210 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2304 683
rect 23 567 73 649
rect 23 533 39 567
rect 23 504 73 533
rect 113 567 169 596
rect 113 533 129 567
rect 163 533 169 567
rect 203 584 269 649
rect 203 550 219 584
rect 253 550 269 584
rect 405 584 471 649
rect 405 550 421 584
rect 455 550 471 584
rect 888 585 957 649
rect 888 551 905 585
rect 939 551 957 585
rect 113 525 169 533
rect 113 516 178 525
rect 613 522 669 551
rect 613 516 629 522
rect 113 504 629 516
rect 138 488 629 504
rect 663 488 669 522
rect 703 539 854 551
rect 703 505 719 539
rect 753 517 854 539
rect 998 520 1065 536
rect 998 517 1015 520
rect 753 505 1015 517
rect 138 482 669 488
rect 25 386 104 439
rect 25 352 60 386
rect 94 352 104 386
rect 25 318 104 352
rect 25 284 60 318
rect 94 284 104 318
rect 25 250 104 284
rect 25 216 60 250
rect 94 216 104 250
rect 25 200 104 216
rect 138 166 172 482
rect 629 471 669 482
rect 802 486 1015 505
rect 1049 486 1065 520
rect 802 483 1065 486
rect 294 437 365 448
rect 206 424 260 428
rect 206 412 223 424
rect 206 378 216 412
rect 257 390 260 424
rect 250 378 260 390
rect 206 344 260 378
rect 206 310 216 344
rect 250 310 260 344
rect 206 276 260 310
rect 206 242 216 276
rect 250 242 260 276
rect 206 226 260 242
rect 294 403 315 437
rect 349 403 365 437
rect 294 389 365 403
rect 495 437 595 448
rect 629 437 768 471
rect 495 403 511 437
rect 545 412 595 437
rect 545 403 604 412
rect 495 389 700 403
rect 294 228 328 389
rect 558 387 700 389
rect 558 380 666 387
rect 409 355 455 356
rect 362 339 455 355
rect 362 305 373 339
rect 407 305 455 339
rect 495 339 533 355
rect 362 262 455 305
rect 489 305 495 310
rect 529 305 533 339
rect 489 228 533 305
rect 294 194 330 228
rect 364 195 533 228
rect 567 353 666 380
rect 567 315 700 353
rect 364 194 508 195
rect 34 137 172 166
rect 34 103 50 137
rect 84 132 172 137
rect 206 137 256 166
rect 84 103 100 132
rect 34 74 100 103
rect 206 103 222 137
rect 294 160 384 194
rect 567 161 623 315
rect 734 274 768 437
rect 294 126 330 160
rect 364 126 384 160
rect 294 110 384 126
rect 418 126 434 160
rect 468 126 484 160
rect 206 17 256 103
rect 418 17 484 126
rect 518 127 534 161
rect 568 127 623 161
rect 518 85 623 127
rect 657 240 768 274
rect 657 179 707 240
rect 802 206 836 483
rect 978 470 1065 483
rect 1156 535 1206 649
rect 1190 501 1206 535
rect 691 145 707 179
rect 657 119 707 145
rect 741 179 836 206
rect 870 415 926 431
rect 870 381 876 415
rect 910 381 926 415
rect 870 347 926 381
rect 870 313 876 347
rect 910 313 926 347
rect 870 218 926 313
rect 978 323 1012 470
rect 1156 466 1206 501
rect 1190 432 1206 466
rect 1046 424 1122 431
rect 1046 415 1087 424
rect 1046 381 1062 415
rect 1121 390 1122 424
rect 1096 381 1122 390
rect 1046 365 1122 381
rect 1156 398 1206 432
rect 1190 364 1206 398
rect 1156 348 1206 364
rect 1246 535 1296 551
rect 1280 501 1296 535
rect 1246 464 1296 501
rect 1340 523 1533 539
rect 1340 489 1361 523
rect 1395 489 1533 523
rect 1340 473 1533 489
rect 1280 430 1296 464
rect 1246 393 1296 430
rect 1280 359 1296 393
rect 978 307 1112 323
rect 1246 314 1296 359
rect 978 289 1062 307
rect 1046 273 1062 289
rect 1096 273 1112 307
rect 1046 257 1112 273
rect 1149 280 1296 314
rect 1330 423 1465 439
rect 1330 389 1424 423
rect 1458 389 1465 423
rect 1330 373 1465 389
rect 1149 218 1183 280
rect 1330 246 1364 373
rect 1499 319 1533 473
rect 1567 530 1612 649
rect 1762 567 1805 649
rect 1601 496 1612 530
rect 1567 467 1612 496
rect 1652 530 1728 546
rect 1652 496 1664 530
rect 1698 496 1728 530
rect 1652 467 1728 496
rect 1567 424 1660 433
rect 1601 417 1660 424
rect 1601 390 1610 417
rect 1567 383 1610 390
rect 1644 383 1660 417
rect 1567 367 1660 383
rect 1694 387 1728 467
rect 1762 533 1767 567
rect 1801 533 1805 567
rect 1762 471 1805 533
rect 1762 437 1767 471
rect 1801 437 1805 471
rect 1762 421 1805 437
rect 1852 580 1990 597
rect 1852 546 1857 580
rect 1891 546 1925 580
rect 1959 546 1990 580
rect 1852 497 1990 546
rect 1852 463 1857 497
rect 1891 463 1925 497
rect 1959 463 1990 497
rect 1852 414 1990 463
rect 1694 353 1794 387
rect 1852 380 1857 414
rect 1891 380 1925 414
rect 1959 380 1990 414
rect 1852 362 1990 380
rect 870 184 1133 218
rect 1167 184 1183 218
rect 1217 230 1364 246
rect 1217 196 1312 230
rect 1346 196 1364 230
rect 741 145 757 179
rect 791 145 836 179
rect 1217 180 1364 196
rect 1398 303 1726 319
rect 1398 285 1682 303
rect 1217 150 1251 180
rect 741 119 836 145
rect 870 116 1251 150
rect 1398 146 1432 285
rect 1666 269 1682 285
rect 1716 269 1726 303
rect 1666 253 1726 269
rect 1486 230 1552 246
rect 1486 196 1502 230
rect 1536 214 1552 230
rect 1760 214 1794 353
rect 1536 196 1794 214
rect 1486 180 1794 196
rect 1285 130 1432 146
rect 870 85 904 116
rect 518 51 904 85
rect 1285 96 1322 130
rect 1356 96 1432 130
rect 999 48 1015 82
rect 1049 48 1065 82
rect 1285 80 1432 96
rect 1507 128 1599 136
rect 1507 94 1536 128
rect 1570 94 1599 128
rect 999 17 1065 48
rect 1507 17 1599 94
rect 1697 133 1794 180
rect 1697 99 1713 133
rect 1747 99 1794 133
rect 1697 70 1794 99
rect 1828 210 1878 226
rect 1862 176 1878 210
rect 1828 120 1878 176
rect 1862 86 1878 120
rect 1828 17 1878 86
rect 1912 210 1990 362
rect 1912 176 1928 210
rect 1962 176 1990 210
rect 1912 120 1990 176
rect 1912 86 1928 120
rect 1962 86 1990 120
rect 1912 70 1990 86
rect 2038 579 2088 595
rect 2072 545 2088 579
rect 2038 471 2088 545
rect 2072 437 2088 471
rect 2038 326 2088 437
rect 2122 580 2181 649
rect 2122 546 2135 580
rect 2169 546 2181 580
rect 2122 497 2181 546
rect 2122 463 2135 497
rect 2169 463 2181 497
rect 2122 414 2181 463
rect 2122 380 2141 414
rect 2175 380 2181 414
rect 2122 364 2181 380
rect 2215 580 2287 596
rect 2215 546 2231 580
rect 2265 546 2287 580
rect 2215 497 2287 546
rect 2215 463 2231 497
rect 2265 463 2287 497
rect 2215 414 2287 463
rect 2215 380 2231 414
rect 2265 380 2287 414
rect 2215 364 2287 380
rect 2038 310 2219 326
rect 2038 276 2176 310
rect 2210 276 2219 310
rect 2038 260 2219 276
rect 2038 145 2088 260
rect 2253 226 2287 364
rect 2038 111 2043 145
rect 2077 111 2088 145
rect 2038 70 2088 111
rect 2129 210 2179 226
rect 2129 176 2141 210
rect 2175 176 2179 210
rect 2129 120 2179 176
rect 2129 86 2141 120
rect 2175 86 2179 120
rect 2129 17 2179 86
rect 2213 210 2287 226
rect 2213 176 2229 210
rect 2263 176 2287 210
rect 2213 120 2287 176
rect 2213 86 2229 120
rect 2263 86 2287 120
rect 2213 70 2287 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2304 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 223 412 257 424
rect 223 390 250 412
rect 250 390 257 412
rect 1087 415 1121 424
rect 1087 390 1096 415
rect 1096 390 1121 415
rect 1567 390 1601 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
<< metal1 >>
rect 0 683 2304 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2304 683
rect 0 617 2304 649
rect 211 424 269 430
rect 211 390 223 424
rect 257 421 269 424
rect 1075 424 1133 430
rect 1075 421 1087 424
rect 257 393 1087 421
rect 257 390 269 393
rect 211 384 269 390
rect 1075 390 1087 393
rect 1121 421 1133 424
rect 1555 424 1613 430
rect 1555 421 1567 424
rect 1121 393 1567 421
rect 1121 390 1133 393
rect 1075 384 1133 390
rect 1555 390 1567 393
rect 1601 390 1613 424
rect 1555 384 1613 390
rect 0 17 2304 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2304 17
rect 0 -49 2304 -17
<< labels >>
flabel pwell s 0 0 2304 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 2304 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel comment s 932 630 932 630 0 FreeSans 300 0 0 0 no_jumper_check
flabel comment s 591 36 591 36 0 FreeSans 300 0 0 0 no_jumper_check
rlabel comment s 0 0 0 0 4 dfrbp_1
flabel metal1 s 223 390 257 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew
flabel metal1 s 0 617 2304 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 2304 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 2239 94 2273 128 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 2239 168 2273 202 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 2239 390 2273 424 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 31 390 65 424 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 1951 390 1985 424 0 FreeSans 340 0 0 0 Q_N
port 9 nsew
flabel corelocali s 1951 464 1985 498 0 FreeSans 340 0 0 0 Q_N
port 9 nsew
flabel corelocali s 1951 538 1985 572 0 FreeSans 340 0 0 0 Q_N
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 2304 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 2641038
string GDS_START 2623504
<< end >>
