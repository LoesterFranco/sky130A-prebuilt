magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 17 153 73 335
rect 206 153 285 335
rect 571 344 667 394
rect 631 318 667 344
rect 631 211 763 318
rect 2511 51 2600 493
rect 2940 299 3016 490
rect 2961 165 3016 299
rect 2940 55 3016 165
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3128 561
rect 17 405 69 493
rect 103 439 163 527
rect 207 451 449 493
rect 207 405 241 451
rect 494 417 537 493
rect 588 428 656 527
rect 17 369 241 405
rect 279 374 369 415
rect 110 255 172 335
rect 110 221 126 255
rect 160 221 172 255
rect 110 153 172 221
rect 17 17 86 119
rect 331 112 369 374
rect 413 354 537 417
rect 413 181 480 354
rect 701 391 735 465
rect 769 455 845 527
rect 889 427 958 493
rect 701 355 859 391
rect 514 255 590 310
rect 514 221 529 255
rect 563 221 590 255
rect 514 215 590 221
rect 413 143 543 181
rect 807 177 859 355
rect 195 56 369 112
rect 405 17 441 109
rect 492 51 543 143
rect 704 143 859 177
rect 903 284 958 427
rect 992 318 1036 493
rect 1086 427 1241 493
rect 1289 455 1355 527
rect 903 218 968 284
rect 588 17 656 111
rect 704 51 741 143
rect 903 117 937 218
rect 1002 184 1036 318
rect 1121 315 1173 391
rect 1207 279 1241 427
rect 1420 421 1473 490
rect 1531 425 1742 527
rect 1776 425 1947 492
rect 2009 447 2085 527
rect 1285 387 1473 421
rect 1913 413 1947 425
rect 2129 413 2172 490
rect 2227 447 2293 527
rect 1285 315 1319 387
rect 1438 323 1545 353
rect 1438 289 1489 323
rect 1523 289 1545 323
rect 1582 299 1751 391
rect 1097 255 1387 279
rect 1590 255 1672 265
rect 786 17 848 109
rect 892 51 937 117
rect 971 51 1036 184
rect 1080 245 1672 255
rect 1080 51 1178 245
rect 1212 161 1295 203
rect 1350 195 1672 245
rect 1707 179 1751 299
rect 1823 215 1879 381
rect 1913 379 2293 413
rect 1937 323 2215 345
rect 1937 289 1947 323
rect 1981 305 2215 323
rect 2249 305 2293 379
rect 1981 289 1992 305
rect 1937 283 1992 289
rect 2337 271 2389 493
rect 2434 297 2476 527
rect 1922 179 1978 249
rect 1212 127 1417 161
rect 1707 139 1978 179
rect 2028 237 2389 271
rect 2028 171 2073 237
rect 2121 169 2309 203
rect 1212 17 1319 93
rect 1355 51 1417 127
rect 1508 17 1655 138
rect 2121 89 2155 169
rect 1832 55 2155 89
rect 2244 17 2278 109
rect 2353 108 2389 237
rect 2312 51 2389 108
rect 2434 17 2476 177
rect 2643 297 2701 527
rect 2744 265 2781 493
rect 2815 327 2896 527
rect 2744 199 2917 265
rect 2643 17 2701 177
rect 2744 51 2781 199
rect 3050 297 3103 527
rect 2815 17 2896 165
rect 3050 17 3103 177
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3128 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 2881 527 2915 561
rect 2973 527 3007 561
rect 3065 527 3099 561
rect 126 221 160 255
rect 529 221 563 255
rect 1489 289 1523 323
rect 1947 289 1981 323
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
rect 2881 -17 2915 17
rect 2973 -17 3007 17
rect 3065 -17 3099 17
<< metal1 >>
rect 0 561 3128 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3128 561
rect 0 496 3128 527
rect 1477 323 1545 329
rect 1477 289 1489 323
rect 1523 320 1545 323
rect 1935 323 1993 329
rect 1935 320 1947 323
rect 1523 292 1947 320
rect 1523 289 1545 292
rect 1477 283 1545 289
rect 1935 289 1947 292
rect 1981 289 1993 323
rect 1935 283 1993 289
rect 114 255 172 261
rect 114 221 126 255
rect 160 252 172 255
rect 517 255 575 261
rect 517 252 529 255
rect 160 224 529 252
rect 160 221 172 224
rect 114 215 172 221
rect 517 221 529 224
rect 563 221 575 255
rect 517 215 575 221
rect 0 17 3128 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3128 17
rect 0 -48 3128 -17
<< obsm1 >>
rect 813 388 881 397
rect 1109 388 1177 397
rect 1629 388 1687 397
rect 813 360 1687 388
rect 813 351 881 360
rect 1109 351 1177 360
rect 1629 351 1687 360
rect 323 320 391 329
rect 990 320 1048 329
rect 323 292 1048 320
rect 323 283 391 292
rect 990 283 1048 292
rect 905 252 963 261
rect 1823 252 1891 261
rect 905 224 1891 252
rect 905 215 963 224
rect 1823 215 1891 224
<< labels >>
rlabel locali s 631 318 667 344 6 CLK
port 1 nsew signal input
rlabel locali s 631 211 763 318 6 CLK
port 1 nsew signal input
rlabel locali s 571 344 667 394 6 CLK
port 1 nsew signal input
rlabel locali s 206 153 285 335 6 D
port 2 nsew signal input
rlabel locali s 2961 165 3016 299 6 Q
port 3 nsew signal output
rlabel locali s 2940 299 3016 490 6 Q
port 3 nsew signal output
rlabel locali s 2940 55 3016 165 6 Q
port 3 nsew signal output
rlabel locali s 2511 51 2600 493 6 Q_N
port 4 nsew signal output
rlabel locali s 17 153 73 335 6 SCD
port 5 nsew signal input
rlabel metal1 s 517 252 575 261 6 SCE
port 6 nsew signal input
rlabel metal1 s 517 215 575 224 6 SCE
port 6 nsew signal input
rlabel metal1 s 114 252 172 261 6 SCE
port 6 nsew signal input
rlabel metal1 s 114 224 575 252 6 SCE
port 6 nsew signal input
rlabel metal1 s 114 215 172 224 6 SCE
port 6 nsew signal input
rlabel metal1 s 1935 320 1993 329 6 SET_B
port 7 nsew signal input
rlabel metal1 s 1935 283 1993 292 6 SET_B
port 7 nsew signal input
rlabel metal1 s 1477 320 1545 329 6 SET_B
port 7 nsew signal input
rlabel metal1 s 1477 292 1993 320 6 SET_B
port 7 nsew signal input
rlabel metal1 s 1477 283 1545 292 6 SET_B
port 7 nsew signal input
rlabel metal1 s 0 -48 3128 48 8 VGND
port 8 nsew ground bidirectional
rlabel metal1 s 0 496 3128 592 6 VPWR
port 9 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 3128 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 223638
string GDS_START 200350
<< end >>
