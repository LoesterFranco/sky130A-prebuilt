magic
tech sky130A
magscale 1 2
timestamp 1599588244
<< locali >>
rect 21 236 87 310
rect 121 236 263 310
rect 477 236 551 302
rect 585 236 651 430
rect 697 70 784 430
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 53 378 103 596
rect 143 412 209 649
rect 249 378 283 596
rect 53 344 283 378
rect 317 562 584 596
rect 317 404 389 562
rect 317 310 351 404
rect 453 370 516 528
rect 550 498 584 562
rect 621 532 699 649
rect 813 532 879 649
rect 550 464 894 498
rect 297 276 351 310
rect 385 336 516 370
rect 297 202 331 276
rect 58 17 124 202
rect 216 168 331 202
rect 385 202 435 336
rect 385 168 574 202
rect 216 70 296 168
rect 330 17 504 134
rect 538 70 574 168
rect 610 17 663 188
rect 818 270 894 464
rect 820 17 870 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
rlabel locali s 585 236 651 430 6 A1_N
port 1 nsew signal input
rlabel locali s 477 236 551 302 6 A2_N
port 2 nsew signal input
rlabel locali s 21 236 87 310 6 B1
port 3 nsew signal input
rlabel locali s 121 236 263 310 6 B2
port 4 nsew signal input
rlabel locali s 697 70 784 430 6 X
port 5 nsew signal output
rlabel metal1 s 0 -49 960 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 7 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 617 960 715 6 VPWR
port 9 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3540562
string GDS_START 3532212
<< end >>
