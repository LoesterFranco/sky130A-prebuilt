magic
tech sky130A
magscale 1 2
timestamp 1604502729
<< locali >>
rect 123 378 189 547
rect 23 344 189 378
rect 23 202 71 344
rect 121 236 195 310
rect 261 276 651 310
rect 261 244 327 276
rect 585 236 651 276
rect 330 202 396 210
rect 23 168 396 202
rect 23 70 89 168
rect 330 70 396 168
rect 530 62 647 196
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 23 581 263 615
rect 23 412 89 581
rect 229 378 263 581
rect 303 446 369 598
rect 403 480 469 649
rect 503 446 559 598
rect 303 412 559 446
rect 593 378 649 596
rect 229 344 649 378
rect 123 17 296 130
rect 430 17 496 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel locali s 530 62 647 196 6 A
port 1 nsew signal input
rlabel locali s 585 236 651 276 6 B
port 2 nsew signal input
rlabel locali s 261 276 651 310 6 B
port 2 nsew signal input
rlabel locali s 261 244 327 276 6 B
port 2 nsew signal input
rlabel locali s 121 236 195 310 6 C
port 3 nsew signal input
rlabel locali s 330 202 396 210 6 Y
port 4 nsew signal output
rlabel locali s 330 70 396 168 6 Y
port 4 nsew signal output
rlabel locali s 123 378 189 547 6 Y
port 4 nsew signal output
rlabel locali s 23 344 189 378 6 Y
port 4 nsew signal output
rlabel locali s 23 202 71 344 6 Y
port 4 nsew signal output
rlabel locali s 23 168 396 202 6 Y
port 4 nsew signal output
rlabel locali s 23 70 89 168 6 Y
port 4 nsew signal output
rlabel metal1 s 0 -49 672 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 617 672 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1574424
string GDS_START 1567546
<< end >>
