magic
tech sky130A
magscale 1 2
timestamp 1599588244
<< locali >>
rect 85 270 161 356
rect 1158 451 1224 593
rect 1158 417 1235 451
rect 889 236 1012 310
rect 1201 276 1235 417
rect 1201 242 1330 276
rect 1264 70 1330 242
rect 1535 236 1601 310
rect 2215 364 2287 596
rect 2253 226 2287 364
rect 2231 70 2287 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2304 683
rect 17 390 97 596
rect 131 390 197 649
rect 238 581 762 615
rect 17 236 51 390
rect 238 370 304 581
rect 195 236 236 336
rect 270 298 304 370
rect 338 513 652 547
rect 338 366 372 513
rect 406 445 655 479
rect 406 400 440 445
rect 338 332 419 366
rect 480 361 555 411
rect 270 264 349 298
rect 17 230 236 236
rect 17 196 249 230
rect 17 96 73 196
rect 109 96 181 162
rect 109 17 143 96
rect 215 85 249 196
rect 283 119 349 264
rect 385 265 419 332
rect 385 202 455 265
rect 385 168 415 202
rect 449 168 455 202
rect 385 119 455 168
rect 489 145 555 361
rect 589 350 655 445
rect 589 316 607 350
rect 641 316 655 350
rect 589 145 655 316
rect 489 85 523 145
rect 692 129 762 581
rect 808 361 875 593
rect 909 361 975 649
rect 1020 395 1086 593
rect 1269 417 1495 594
rect 808 202 842 361
rect 1046 261 1080 395
rect 1114 295 1167 361
rect 1046 227 1099 261
rect 215 51 523 85
rect 557 85 623 111
rect 808 85 947 202
rect 557 51 947 85
rect 981 17 1031 193
rect 1065 128 1099 227
rect 1133 208 1167 295
rect 1269 350 1322 376
rect 1269 316 1279 350
rect 1313 316 1322 350
rect 1269 310 1322 316
rect 1133 202 1223 208
rect 1133 168 1183 202
rect 1217 168 1223 202
rect 1133 162 1223 168
rect 1065 78 1230 128
rect 1364 226 1427 360
rect 1364 202 1415 226
rect 1364 168 1375 202
rect 1409 168 1415 202
rect 1461 192 1495 417
rect 1529 388 1563 649
rect 1603 498 1669 596
rect 1715 574 2091 608
rect 1715 532 1781 574
rect 1912 498 2006 540
rect 1603 464 2006 498
rect 1603 364 1669 464
rect 1635 226 1669 364
rect 1827 364 1872 430
rect 1912 364 2006 464
rect 1703 350 1793 356
rect 1703 316 1759 350
rect 1703 310 1793 316
rect 1703 260 1753 310
rect 1827 276 1861 364
rect 1972 318 2006 364
rect 2040 386 2091 574
rect 2130 420 2180 649
rect 2040 352 2125 386
rect 1787 242 1861 276
rect 1895 252 1938 318
rect 1972 252 2057 318
rect 1787 226 1821 242
rect 1364 162 1415 168
rect 1449 70 1515 192
rect 1549 17 1599 202
rect 1635 70 1703 226
rect 1755 85 1821 226
rect 1895 208 1929 252
rect 2091 218 2125 352
rect 1855 202 1929 208
rect 1889 168 1929 202
rect 1855 162 1929 168
rect 1963 184 2125 218
rect 2162 260 2219 326
rect 1963 119 1997 184
rect 2162 150 2196 260
rect 2031 116 2196 150
rect 2031 85 2065 116
rect 1755 51 2065 85
rect 2099 17 2179 82
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2304 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 415 168 449 202
rect 607 316 641 350
rect 1279 316 1313 350
rect 1183 168 1217 202
rect 1375 168 1409 202
rect 1759 316 1793 350
rect 1855 168 1889 202
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
<< metal1 >>
rect 0 683 2304 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2304 683
rect 0 617 2304 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 2304 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2304 17
rect 0 -49 2304 -17
<< obsm1 >>
rect 595 350 653 356
rect 595 316 607 350
rect 641 347 653 350
rect 1267 350 1325 356
rect 1267 347 1279 350
rect 641 319 1279 347
rect 641 316 653 319
rect 595 310 653 316
rect 1267 316 1279 319
rect 1313 347 1325 350
rect 1747 350 1805 356
rect 1747 347 1759 350
rect 1313 319 1759 347
rect 1313 316 1325 319
rect 1267 310 1325 316
rect 1747 316 1759 319
rect 1793 316 1805 350
rect 1747 310 1805 316
rect 403 202 461 208
rect 403 168 415 202
rect 449 199 461 202
rect 1171 202 1229 208
rect 1171 199 1183 202
rect 449 171 1183 199
rect 449 168 461 171
rect 403 162 461 168
rect 1171 168 1183 171
rect 1217 199 1229 202
rect 1363 202 1421 208
rect 1363 199 1375 202
rect 1217 171 1375 199
rect 1217 168 1229 171
rect 1171 162 1229 168
rect 1363 168 1375 171
rect 1409 199 1421 202
rect 1843 202 1901 208
rect 1843 199 1855 202
rect 1409 171 1855 199
rect 1409 168 1421 171
rect 1363 162 1421 168
rect 1843 168 1855 171
rect 1889 168 1901 202
rect 1843 162 1901 168
<< labels >>
rlabel locali s 85 270 161 356 6 A
port 1 nsew signal input
rlabel locali s 889 236 1012 310 6 B
port 2 nsew signal input
rlabel locali s 1535 236 1601 310 6 CI
port 3 nsew signal input
rlabel locali s 1264 70 1330 242 6 COUT_N
port 4 nsew signal output
rlabel locali s 1201 276 1235 417 6 COUT_N
port 4 nsew signal output
rlabel locali s 1201 242 1330 276 6 COUT_N
port 4 nsew signal output
rlabel locali s 1158 451 1224 593 6 COUT_N
port 4 nsew signal output
rlabel locali s 1158 417 1235 451 6 COUT_N
port 4 nsew signal output
rlabel locali s 2253 226 2287 364 6 SUM
port 5 nsew signal output
rlabel locali s 2231 70 2287 226 6 SUM
port 5 nsew signal output
rlabel locali s 2215 364 2287 596 6 SUM
port 5 nsew signal output
rlabel metal1 s 0 -49 2304 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 7 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 617 2304 715 6 VPWR
port 9 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2304 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 2542472
string GDS_START 2524718
<< end >>
