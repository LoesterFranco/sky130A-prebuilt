magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 3110 704
rect 1204 320 1416 332
<< pwell >>
rect 0 0 3072 49
<< scnmos >>
rect 113 74 143 158
rect 191 74 221 158
rect 389 111 419 195
rect 475 111 505 195
rect 553 111 583 195
rect 639 111 669 195
rect 910 125 940 209
rect 996 125 1026 209
rect 1068 125 1098 209
rect 1265 74 1295 222
rect 1462 74 1492 222
rect 1658 97 1688 181
rect 1794 97 1824 181
rect 1910 97 1940 181
rect 2061 74 2091 202
rect 2283 74 2313 202
rect 2355 74 2385 202
rect 2457 74 2487 158
rect 2535 74 2565 158
rect 2760 74 2790 158
rect 2958 74 2988 222
<< pmoshvt >>
rect 84 464 114 592
rect 162 464 192 592
rect 388 463 418 591
rect 524 463 554 591
rect 602 463 632 591
rect 692 463 722 591
rect 887 455 917 583
rect 1023 455 1053 583
rect 1101 455 1131 583
rect 1295 356 1325 580
rect 1565 368 1595 592
rect 1760 508 1790 592
rect 1860 508 1890 592
rect 1946 508 1976 592
rect 2050 398 2080 566
rect 2244 392 2274 592
rect 2431 392 2461 592
rect 2538 508 2568 592
rect 2622 508 2652 592
rect 2764 464 2794 592
rect 2958 368 2988 592
<< ndiff >>
rect 332 170 389 195
rect 27 146 113 158
rect 27 112 53 146
rect 87 112 113 146
rect 27 74 113 112
rect 143 74 191 158
rect 221 133 278 158
rect 221 99 232 133
rect 266 99 278 133
rect 332 136 344 170
rect 378 136 389 170
rect 332 111 389 136
rect 419 170 475 195
rect 419 136 430 170
rect 464 136 475 170
rect 419 111 475 136
rect 505 111 553 195
rect 583 170 639 195
rect 583 136 594 170
rect 628 136 639 170
rect 583 111 639 136
rect 669 170 740 195
rect 669 136 694 170
rect 728 136 740 170
rect 669 111 740 136
rect 221 74 278 99
rect 854 178 910 209
rect 854 144 865 178
rect 899 144 910 178
rect 854 125 910 144
rect 940 178 996 209
rect 940 144 951 178
rect 985 144 996 178
rect 940 125 996 144
rect 1026 125 1068 209
rect 1098 184 1154 209
rect 1098 150 1109 184
rect 1143 150 1154 184
rect 1098 125 1154 150
rect 1208 150 1265 222
rect 1208 116 1220 150
rect 1254 116 1265 150
rect 1208 74 1265 116
rect 1295 199 1351 222
rect 1295 165 1306 199
rect 1340 165 1351 199
rect 1295 120 1351 165
rect 1295 86 1306 120
rect 1340 86 1351 120
rect 1295 74 1351 86
rect 1405 127 1462 222
rect 1405 93 1417 127
rect 1451 93 1462 127
rect 1405 74 1462 93
rect 1492 210 1548 222
rect 1492 176 1503 210
rect 1537 176 1548 210
rect 2011 181 2061 202
rect 1492 120 1548 176
rect 1492 86 1503 120
rect 1537 86 1548 120
rect 1602 169 1658 181
rect 1602 135 1613 169
rect 1647 135 1658 169
rect 1602 97 1658 135
rect 1688 169 1794 181
rect 1688 135 1749 169
rect 1783 135 1794 169
rect 1688 97 1794 135
rect 1824 97 1910 181
rect 1940 120 2061 181
rect 1940 97 1966 120
rect 1492 74 1548 86
rect 1955 86 1966 97
rect 2000 86 2061 120
rect 1955 74 2061 86
rect 2091 179 2148 202
rect 2091 145 2102 179
rect 2136 145 2148 179
rect 2091 74 2148 145
rect 2226 120 2283 202
rect 2226 86 2238 120
rect 2272 86 2283 120
rect 2226 74 2283 86
rect 2313 74 2355 202
rect 2385 188 2442 202
rect 2385 154 2396 188
rect 2430 158 2442 188
rect 2901 210 2958 222
rect 2901 176 2913 210
rect 2947 176 2958 210
rect 2430 154 2457 158
rect 2385 120 2457 154
rect 2385 86 2396 120
rect 2430 86 2457 120
rect 2385 74 2457 86
rect 2487 74 2535 158
rect 2565 120 2760 158
rect 2565 86 2576 120
rect 2610 86 2701 120
rect 2735 86 2760 120
rect 2565 74 2760 86
rect 2790 133 2847 158
rect 2790 99 2801 133
rect 2835 99 2847 133
rect 2790 74 2847 99
rect 2901 120 2958 176
rect 2901 86 2913 120
rect 2947 86 2958 120
rect 2901 74 2958 86
rect 2988 210 3045 222
rect 2988 176 2999 210
rect 3033 176 3045 210
rect 2988 120 3045 176
rect 2988 86 2999 120
rect 3033 86 3045 120
rect 2988 74 3045 86
<< pdiff >>
rect 27 580 84 592
rect 27 546 37 580
rect 71 546 84 580
rect 27 510 84 546
rect 27 476 37 510
rect 71 476 84 510
rect 27 464 84 476
rect 114 464 162 592
rect 192 578 251 592
rect 192 544 205 578
rect 239 544 251 578
rect 192 464 251 544
rect 329 520 388 591
rect 329 486 341 520
rect 375 486 388 520
rect 329 463 388 486
rect 418 577 524 591
rect 418 543 477 577
rect 511 543 524 577
rect 418 463 524 543
rect 554 463 602 591
rect 632 579 692 591
rect 632 545 645 579
rect 679 545 692 579
rect 632 509 692 545
rect 632 475 645 509
rect 679 475 692 509
rect 632 463 692 475
rect 722 579 777 591
rect 722 545 735 579
rect 769 545 777 579
rect 722 509 777 545
rect 722 475 735 509
rect 769 475 777 509
rect 722 463 777 475
rect 831 516 887 583
rect 831 482 840 516
rect 874 482 887 516
rect 831 455 887 482
rect 917 570 1023 583
rect 917 536 976 570
rect 1010 536 1023 570
rect 917 455 1023 536
rect 1053 455 1101 583
rect 1131 571 1186 583
rect 1131 537 1144 571
rect 1178 537 1186 571
rect 1131 501 1186 537
rect 1131 467 1144 501
rect 1178 467 1186 501
rect 1131 455 1186 467
rect 1240 568 1295 580
rect 1240 534 1248 568
rect 1282 534 1295 568
rect 1240 356 1295 534
rect 1325 409 1380 580
rect 1510 574 1565 592
rect 1510 540 1518 574
rect 1552 540 1565 574
rect 1325 375 1338 409
rect 1372 375 1380 409
rect 1325 356 1380 375
rect 1510 368 1565 540
rect 1595 415 1650 592
rect 1704 580 1760 592
rect 1704 546 1713 580
rect 1747 546 1760 580
rect 1704 508 1760 546
rect 1790 567 1860 592
rect 1790 533 1813 567
rect 1847 533 1860 567
rect 1790 508 1860 533
rect 1890 508 1946 592
rect 1976 580 2032 592
rect 1976 546 1989 580
rect 2023 566 2032 580
rect 2189 580 2244 592
rect 2023 546 2050 566
rect 1976 508 2050 546
rect 1595 381 1608 415
rect 1642 381 1650 415
rect 1595 368 1650 381
rect 1997 398 2050 508
rect 2080 444 2135 566
rect 2080 410 2093 444
rect 2127 410 2135 444
rect 2080 398 2135 410
rect 2189 546 2197 580
rect 2231 546 2244 580
rect 2189 392 2244 546
rect 2274 392 2431 592
rect 2461 580 2538 592
rect 2461 546 2474 580
rect 2508 546 2538 580
rect 2461 512 2538 546
rect 2461 478 2474 512
rect 2508 508 2538 512
rect 2568 508 2622 592
rect 2652 580 2764 592
rect 2652 546 2694 580
rect 2728 546 2764 580
rect 2652 508 2764 546
rect 2508 478 2520 508
rect 2461 438 2520 478
rect 2461 404 2474 438
rect 2508 404 2520 438
rect 2461 392 2520 404
rect 2711 464 2764 508
rect 2794 580 2849 592
rect 2794 546 2807 580
rect 2841 546 2849 580
rect 2794 510 2849 546
rect 2794 476 2807 510
rect 2841 476 2849 510
rect 2794 464 2849 476
rect 2903 580 2958 592
rect 2903 546 2911 580
rect 2945 546 2958 580
rect 2903 497 2958 546
rect 2903 463 2911 497
rect 2945 463 2958 497
rect 2903 414 2958 463
rect 2903 380 2911 414
rect 2945 380 2958 414
rect 2903 368 2958 380
rect 2988 580 3045 592
rect 2988 546 3001 580
rect 3035 546 3045 580
rect 2988 497 3045 546
rect 2988 463 3001 497
rect 3035 463 3045 497
rect 2988 414 3045 463
rect 2988 380 3001 414
rect 3035 380 3045 414
rect 2988 368 3045 380
<< ndiffc >>
rect 53 112 87 146
rect 232 99 266 133
rect 344 136 378 170
rect 430 136 464 170
rect 594 136 628 170
rect 694 136 728 170
rect 865 144 899 178
rect 951 144 985 178
rect 1109 150 1143 184
rect 1220 116 1254 150
rect 1306 165 1340 199
rect 1306 86 1340 120
rect 1417 93 1451 127
rect 1503 176 1537 210
rect 1503 86 1537 120
rect 1613 135 1647 169
rect 1749 135 1783 169
rect 1966 86 2000 120
rect 2102 145 2136 179
rect 2238 86 2272 120
rect 2396 154 2430 188
rect 2913 176 2947 210
rect 2396 86 2430 120
rect 2576 86 2610 120
rect 2701 86 2735 120
rect 2801 99 2835 133
rect 2913 86 2947 120
rect 2999 176 3033 210
rect 2999 86 3033 120
<< pdiffc >>
rect 37 546 71 580
rect 37 476 71 510
rect 205 544 239 578
rect 341 486 375 520
rect 477 543 511 577
rect 645 545 679 579
rect 645 475 679 509
rect 735 545 769 579
rect 735 475 769 509
rect 840 482 874 516
rect 976 536 1010 570
rect 1144 537 1178 571
rect 1144 467 1178 501
rect 1248 534 1282 568
rect 1518 540 1552 574
rect 1338 375 1372 409
rect 1713 546 1747 580
rect 1813 533 1847 567
rect 1989 546 2023 580
rect 1608 381 1642 415
rect 2093 410 2127 444
rect 2197 546 2231 580
rect 2474 546 2508 580
rect 2474 478 2508 512
rect 2694 546 2728 580
rect 2474 404 2508 438
rect 2807 546 2841 580
rect 2807 476 2841 510
rect 2911 546 2945 580
rect 2911 463 2945 497
rect 2911 380 2945 414
rect 3001 546 3035 580
rect 3001 463 3035 497
rect 3001 380 3035 414
<< poly >>
rect 84 592 114 618
rect 162 592 192 618
rect 388 591 418 617
rect 524 591 554 617
rect 602 591 632 617
rect 689 606 920 636
rect 692 591 722 606
rect 884 598 920 606
rect 84 449 114 464
rect 162 449 192 464
rect 887 583 917 598
rect 1023 583 1053 609
rect 1101 583 1131 609
rect 81 356 117 449
rect 159 434 195 449
rect 388 448 418 463
rect 524 448 554 463
rect 602 448 632 463
rect 159 422 225 434
rect 159 406 261 422
rect 159 404 211 406
rect 195 372 211 404
rect 245 372 261 406
rect 81 340 149 356
rect 81 306 99 340
rect 133 306 149 340
rect 81 272 149 306
rect 195 338 261 372
rect 195 304 211 338
rect 245 304 261 338
rect 333 418 557 448
rect 333 330 363 418
rect 411 354 505 370
rect 599 367 635 448
rect 692 437 722 463
rect 1295 580 1325 606
rect 1565 592 1595 618
rect 1760 592 1790 618
rect 1860 592 1890 618
rect 1946 592 1976 618
rect 2244 592 2274 618
rect 2431 592 2461 618
rect 2538 592 2568 618
rect 2622 592 2652 618
rect 2764 592 2794 618
rect 2958 592 2988 618
rect 887 440 917 455
rect 1023 440 1053 455
rect 1101 440 1131 455
rect 195 288 261 304
rect 303 314 369 330
rect 81 238 99 272
rect 133 238 149 272
rect 303 280 319 314
rect 353 280 369 314
rect 411 320 427 354
rect 461 320 505 354
rect 411 304 505 320
rect 303 240 369 280
rect 81 222 149 238
rect 113 158 143 222
rect 191 210 419 240
rect 191 158 221 210
rect 389 195 419 210
rect 475 195 505 304
rect 547 351 635 367
rect 547 317 563 351
rect 597 317 635 351
rect 547 301 635 317
rect 766 373 832 389
rect 766 339 782 373
rect 816 339 832 373
rect 766 305 832 339
rect 553 195 583 301
rect 766 271 782 305
rect 816 271 832 305
rect 884 302 920 440
rect 1020 349 1056 440
rect 990 333 1056 349
rect 766 240 832 271
rect 639 237 832 240
rect 639 210 782 237
rect 639 195 669 210
rect 766 203 782 210
rect 816 203 832 237
rect 880 286 946 302
rect 880 252 896 286
rect 930 252 946 286
rect 990 299 1006 333
rect 1040 299 1056 333
rect 990 283 1056 299
rect 1098 417 1134 440
rect 1098 401 1164 417
rect 1098 367 1114 401
rect 1148 367 1164 401
rect 1098 333 1164 367
rect 1412 416 1478 432
rect 1412 382 1428 416
rect 1462 382 1478 416
rect 1295 341 1325 356
rect 1412 353 1478 382
rect 2050 566 2080 592
rect 1760 493 1790 508
rect 1860 493 1890 508
rect 1946 493 1976 508
rect 1757 467 1793 493
rect 1682 451 1793 467
rect 1857 451 1893 493
rect 1682 417 1698 451
rect 1732 437 1793 451
rect 1732 417 1748 437
rect 1682 401 1748 417
rect 1835 435 1901 451
rect 1835 401 1851 435
rect 1885 401 1901 435
rect 1835 385 1901 401
rect 1565 353 1595 368
rect 1835 353 1865 385
rect 1098 299 1114 333
rect 1148 299 1164 333
rect 1292 310 1328 341
rect 1412 323 1865 353
rect 1098 283 1164 299
rect 1265 294 1332 310
rect 880 236 946 252
rect 910 209 940 236
rect 996 209 1026 283
rect 1265 260 1282 294
rect 1316 260 1332 294
rect 1265 244 1332 260
rect 1068 209 1098 235
rect 1265 222 1295 244
rect 1462 222 1492 323
rect 766 169 832 203
rect 766 135 782 169
rect 816 135 832 169
rect 389 85 419 111
rect 475 85 505 111
rect 553 85 583 111
rect 639 85 669 111
rect 766 101 832 135
rect 113 48 143 74
rect 191 48 221 74
rect 766 67 782 101
rect 816 67 832 101
rect 766 51 832 67
rect 910 51 940 125
rect 996 99 1026 125
rect 1068 51 1098 125
rect 1658 181 1688 323
rect 1943 297 1979 493
rect 2050 383 2080 398
rect 2538 493 2568 508
rect 2622 493 2652 508
rect 2047 366 2083 383
rect 2244 377 2274 392
rect 2431 377 2461 392
rect 2027 350 2093 366
rect 2027 316 2043 350
rect 2077 316 2093 350
rect 2027 300 2093 316
rect 2241 305 2277 377
rect 1910 281 1979 297
rect 1794 253 1868 269
rect 1794 219 1818 253
rect 1852 219 1868 253
rect 1794 203 1868 219
rect 1910 247 1929 281
rect 1963 247 1979 281
rect 1910 231 1979 247
rect 1794 181 1824 203
rect 1910 181 1940 231
rect 2061 202 2091 300
rect 2143 289 2277 305
rect 2319 344 2385 360
rect 2428 351 2464 377
rect 2319 310 2335 344
rect 2369 310 2385 344
rect 2319 294 2385 310
rect 2143 255 2159 289
rect 2193 255 2227 289
rect 2261 255 2277 289
rect 2143 252 2277 255
rect 2143 222 2313 252
rect 2283 202 2313 222
rect 2355 202 2385 294
rect 2427 335 2493 351
rect 2427 301 2443 335
rect 2477 301 2493 335
rect 2427 285 2493 301
rect 2535 311 2571 493
rect 2619 476 2655 493
rect 2613 460 2679 476
rect 2613 426 2629 460
rect 2663 426 2679 460
rect 2764 449 2794 464
rect 2613 410 2679 426
rect 2535 295 2601 311
rect 910 21 1098 51
rect 1265 48 1295 74
rect 1462 48 1492 74
rect 1658 71 1688 97
rect 1794 71 1824 97
rect 1910 71 1940 97
rect 2457 158 2487 285
rect 2535 261 2551 295
rect 2585 261 2601 295
rect 2535 245 2601 261
rect 2643 203 2673 410
rect 2761 324 2797 449
rect 2958 353 2988 368
rect 2955 324 2991 353
rect 2761 276 2991 324
rect 2723 260 2991 276
rect 2723 226 2739 260
rect 2773 246 2991 260
rect 2773 226 2791 246
rect 2723 210 2791 226
rect 2958 222 2988 246
rect 2535 173 2673 203
rect 2535 158 2565 173
rect 2760 158 2790 210
rect 2061 48 2091 74
rect 2283 48 2313 74
rect 2355 48 2385 74
rect 2457 48 2487 74
rect 2535 48 2565 74
rect 2760 48 2790 74
rect 2958 48 2988 74
<< polycont >>
rect 211 372 245 406
rect 99 306 133 340
rect 211 304 245 338
rect 99 238 133 272
rect 319 280 353 314
rect 427 320 461 354
rect 563 317 597 351
rect 782 339 816 373
rect 782 271 816 305
rect 782 203 816 237
rect 896 252 930 286
rect 1006 299 1040 333
rect 1114 367 1148 401
rect 1428 382 1462 416
rect 1698 417 1732 451
rect 1851 401 1885 435
rect 1114 299 1148 333
rect 1282 260 1316 294
rect 782 135 816 169
rect 782 67 816 101
rect 2043 316 2077 350
rect 1818 219 1852 253
rect 1929 247 1963 281
rect 2335 310 2369 344
rect 2159 255 2193 289
rect 2227 255 2261 289
rect 2443 301 2477 335
rect 2629 426 2663 460
rect 2551 261 2585 295
rect 2739 226 2773 260
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3072 683
rect 17 580 87 596
rect 17 546 37 580
rect 71 546 87 580
rect 17 510 87 546
rect 189 578 239 649
rect 189 544 205 578
rect 189 526 239 544
rect 273 581 443 615
rect 17 476 37 510
rect 71 492 87 510
rect 273 492 307 581
rect 71 476 307 492
rect 17 458 307 476
rect 341 520 375 547
rect 17 162 51 458
rect 341 424 375 486
rect 409 492 443 581
rect 477 577 527 649
rect 511 543 527 577
rect 477 526 527 543
rect 629 579 679 595
rect 629 545 645 579
rect 629 509 679 545
rect 629 492 645 509
rect 409 475 645 492
rect 409 458 679 475
rect 195 406 477 424
rect 195 372 211 406
rect 245 390 477 406
rect 245 372 261 390
rect 85 340 161 356
rect 85 306 99 340
rect 133 306 161 340
rect 85 272 161 306
rect 85 238 99 272
rect 133 238 161 272
rect 85 222 161 238
rect 195 338 261 372
rect 195 304 211 338
rect 245 304 261 338
rect 195 230 261 304
rect 303 314 369 356
rect 303 280 319 314
rect 353 280 369 314
rect 411 354 477 390
rect 411 320 427 354
rect 461 320 477 354
rect 411 304 477 320
rect 511 351 611 367
rect 511 350 563 351
rect 545 317 563 350
rect 597 317 611 351
rect 545 316 611 317
rect 511 301 611 316
rect 303 264 369 280
rect 645 267 679 458
rect 578 233 679 267
rect 713 581 942 615
rect 713 579 769 581
rect 713 545 735 579
rect 713 509 769 545
rect 713 475 735 509
rect 713 459 769 475
rect 803 516 874 547
rect 803 482 840 516
rect 195 199 362 230
rect 195 196 378 199
rect 328 170 378 196
rect 17 146 118 162
rect 17 112 53 146
rect 87 112 118 146
rect 17 96 118 112
rect 216 133 282 162
rect 216 99 232 133
rect 266 99 282 133
rect 328 136 344 170
rect 328 107 378 136
rect 414 170 480 199
rect 414 136 430 170
rect 464 136 480 170
rect 216 17 282 99
rect 414 17 480 136
rect 578 170 644 233
rect 713 199 747 459
rect 803 451 874 482
rect 908 485 942 581
rect 976 570 1026 649
rect 1010 536 1026 570
rect 976 519 1026 536
rect 1128 571 1198 587
rect 1128 537 1144 571
rect 1178 537 1198 571
rect 1128 501 1198 537
rect 1232 568 1298 649
rect 1232 534 1248 568
rect 1282 534 1298 568
rect 1502 574 1568 649
rect 1502 540 1518 574
rect 1552 540 1568 574
rect 1502 534 1568 540
rect 1602 580 1763 596
rect 1602 546 1713 580
rect 1747 546 1763 580
rect 1797 567 1863 596
rect 1128 485 1144 501
rect 908 467 1144 485
rect 1178 500 1198 501
rect 1602 500 1636 546
rect 1797 533 1813 567
rect 1847 533 1863 567
rect 1973 580 2039 649
rect 1973 546 1989 580
rect 2023 546 2039 580
rect 2181 580 2247 649
rect 2181 546 2197 580
rect 2231 546 2247 580
rect 2474 580 2561 596
rect 2508 546 2561 580
rect 1797 512 1863 533
rect 2474 512 2561 546
rect 2666 580 2757 649
rect 2666 546 2694 580
rect 2728 546 2757 580
rect 2666 530 2757 546
rect 2791 580 2857 596
rect 2791 546 2807 580
rect 2841 546 2857 580
rect 1178 467 1636 500
rect 1767 478 1863 512
rect 1897 478 2440 512
rect 908 466 1636 467
rect 908 451 1232 466
rect 803 417 837 451
rect 578 136 594 170
rect 628 136 644 170
rect 578 107 644 136
rect 678 170 747 199
rect 678 136 694 170
rect 728 136 747 170
rect 678 107 747 136
rect 781 401 1164 417
rect 781 383 1114 401
rect 781 373 837 383
rect 781 339 782 373
rect 816 339 837 373
rect 1098 367 1114 383
rect 1148 367 1164 401
rect 781 305 837 339
rect 781 271 782 305
rect 816 271 837 305
rect 985 333 1056 349
rect 781 237 837 271
rect 781 203 782 237
rect 816 203 837 237
rect 880 286 946 302
rect 880 252 896 286
rect 930 252 946 286
rect 880 236 946 252
rect 985 299 1006 333
rect 1040 299 1056 333
rect 985 236 1056 299
rect 1098 333 1164 367
rect 1098 299 1114 333
rect 1148 299 1164 333
rect 1098 283 1164 299
rect 1198 249 1232 451
rect 1322 416 1478 432
rect 1322 409 1428 416
rect 1322 375 1338 409
rect 1372 382 1428 409
rect 1462 382 1478 416
rect 1372 375 1478 382
rect 1322 366 1478 375
rect 1322 352 1400 366
rect 781 202 837 203
rect 1093 215 1232 249
rect 1266 294 1332 310
rect 1266 260 1282 294
rect 1316 260 1332 294
rect 1266 236 1332 260
rect 781 178 915 202
rect 781 169 865 178
rect 781 135 782 169
rect 816 144 865 169
rect 899 144 915 178
rect 816 135 915 144
rect 781 121 915 135
rect 951 178 1001 202
rect 985 144 1001 178
rect 781 101 837 121
rect 781 67 782 101
rect 816 67 837 101
rect 781 51 837 67
rect 951 17 1001 144
rect 1093 184 1159 215
rect 1366 202 1400 352
rect 1524 330 1558 466
rect 1681 451 1733 467
rect 1681 432 1698 451
rect 1592 417 1698 432
rect 1732 417 1733 451
rect 1592 415 1733 417
rect 1592 381 1608 415
rect 1642 398 1733 415
rect 1642 381 1715 398
rect 1592 364 1715 381
rect 1524 296 1647 330
rect 1093 150 1109 184
rect 1143 150 1159 184
rect 1290 199 1400 202
rect 1093 121 1159 150
rect 1204 150 1256 181
rect 1204 116 1220 150
rect 1254 116 1256 150
rect 1204 17 1256 116
rect 1290 165 1306 199
rect 1340 168 1400 199
rect 1503 210 1553 226
rect 1537 176 1553 210
rect 1340 165 1356 168
rect 1290 120 1356 165
rect 1290 86 1306 120
rect 1340 86 1356 120
rect 1290 70 1356 86
rect 1401 127 1467 134
rect 1401 93 1417 127
rect 1451 93 1467 127
rect 1401 17 1467 93
rect 1503 120 1553 176
rect 1537 86 1553 120
rect 1597 169 1647 296
rect 1597 135 1613 169
rect 1597 119 1647 135
rect 1503 85 1553 86
rect 1681 85 1715 364
rect 1767 358 1801 478
rect 1897 444 1931 478
rect 1835 435 1931 444
rect 1835 401 1851 435
rect 1885 401 1931 435
rect 1835 392 1931 401
rect 2077 410 2093 444
rect 2127 410 2161 444
rect 2077 394 2161 410
rect 2027 358 2093 359
rect 1749 350 2093 358
rect 1749 324 2043 350
rect 1749 169 1783 324
rect 2027 316 2043 324
rect 2077 316 2093 350
rect 2027 307 2093 316
rect 2127 305 2161 394
rect 2312 344 2372 360
rect 2312 310 2335 344
rect 2369 310 2372 344
rect 1913 281 1979 290
rect 1749 119 1783 135
rect 1817 253 1868 269
rect 1817 219 1818 253
rect 1852 219 1868 253
rect 1913 247 1929 281
rect 1963 273 1979 281
rect 2127 289 2277 305
rect 2127 273 2159 289
rect 1963 255 2159 273
rect 2193 255 2227 289
rect 2261 255 2277 289
rect 1963 247 2277 255
rect 1913 239 2277 247
rect 2312 256 2372 310
rect 2406 347 2440 478
rect 2508 478 2561 512
rect 2474 438 2561 478
rect 2791 510 2857 546
rect 2791 476 2807 510
rect 2841 476 2857 510
rect 2508 404 2561 438
rect 2613 460 2857 476
rect 2613 426 2629 460
rect 2663 426 2857 460
rect 2613 415 2857 426
rect 2474 388 2561 404
rect 2527 381 2561 388
rect 2527 347 2757 381
rect 2406 335 2493 347
rect 2406 301 2443 335
rect 2477 301 2493 335
rect 2406 290 2493 301
rect 2535 295 2601 311
rect 2535 261 2551 295
rect 2585 261 2601 295
rect 2535 256 2601 261
rect 1913 238 1979 239
rect 1817 204 1868 219
rect 1817 170 2068 204
rect 1817 85 1851 170
rect 1503 51 1851 85
rect 1950 120 2000 136
rect 1950 86 1966 120
rect 1950 17 2000 86
rect 2034 85 2068 170
rect 2102 179 2136 239
rect 2312 222 2601 256
rect 2312 205 2346 222
rect 2102 119 2136 145
rect 2170 171 2346 205
rect 2635 188 2669 347
rect 2723 276 2757 347
rect 2809 350 2857 415
rect 2809 316 2815 350
rect 2849 316 2857 350
rect 2809 310 2857 316
rect 2723 260 2789 276
rect 2723 226 2739 260
rect 2773 226 2789 260
rect 2723 210 2789 226
rect 2170 85 2204 171
rect 2380 154 2396 188
rect 2430 154 2669 188
rect 2823 162 2857 310
rect 2034 51 2204 85
rect 2238 120 2288 137
rect 2272 86 2288 120
rect 2238 17 2288 86
rect 2380 120 2446 154
rect 2785 133 2857 162
rect 2380 86 2396 120
rect 2430 86 2446 120
rect 2380 70 2446 86
rect 2560 86 2576 120
rect 2610 86 2701 120
rect 2735 86 2751 120
rect 2560 17 2751 86
rect 2785 99 2801 133
rect 2835 99 2857 133
rect 2785 70 2857 99
rect 2895 580 2963 596
rect 2895 546 2911 580
rect 2945 546 2963 580
rect 2895 497 2963 546
rect 2895 463 2911 497
rect 2945 463 2963 497
rect 2895 414 2963 463
rect 2895 380 2911 414
rect 2945 380 2963 414
rect 2895 210 2963 380
rect 3001 580 3051 649
rect 3035 546 3051 580
rect 3001 497 3051 546
rect 3035 463 3051 497
rect 3001 414 3051 463
rect 3035 380 3051 414
rect 3001 364 3051 380
rect 2895 176 2913 210
rect 2947 176 2963 210
rect 2895 120 2963 176
rect 2895 86 2913 120
rect 2947 86 2963 120
rect 2895 70 2963 86
rect 2999 210 3049 226
rect 3033 176 3049 210
rect 2999 120 3049 176
rect 3033 86 3049 120
rect 2999 17 3049 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3072 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 511 316 545 350
rect 2815 316 2849 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
<< metal1 >>
rect 0 683 3072 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3072 683
rect 0 617 3072 649
rect 499 350 557 356
rect 499 316 511 350
rect 545 347 557 350
rect 2803 350 2861 356
rect 2803 347 2815 350
rect 545 319 2815 347
rect 545 316 557 319
rect 499 310 557 316
rect 2803 316 2815 319
rect 2849 316 2861 350
rect 2803 310 2861 316
rect 0 17 3072 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3072 17
rect 0 -49 3072 -17
<< labels >>
rlabel comment s 0 0 0 0 4 sedfxtp_1
flabel comment s 1725 342 1725 342 0 FreeSans 200 0 0 0 no_jumper_check
flabel pwell s 0 0 3072 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nwell s 0 617 3072 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 0 617 3072 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 3072 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 1279 242 1313 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 2911 94 2945 128 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2911 168 2945 202 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2911 242 2945 276 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2911 316 2945 350 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2911 390 2945 424 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2911 464 2945 498 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2911 538 2945 572 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 991 242 1025 276 0 FreeSans 340 0 0 0 SCD
port 4 nsew
flabel corelocali s 895 242 929 276 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 DE
port 3 nsew
flabel corelocali s 127 242 161 276 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 3072 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 522932
string GDS_START 500636
<< end >>
