magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 105 292 375 326
rect 105 258 139 292
rect 341 258 375 292
rect 19 211 139 258
rect 173 211 307 258
rect 341 211 409 258
rect 573 211 639 323
rect 787 323 841 493
rect 975 323 1029 493
rect 1163 323 1217 493
rect 1351 323 1405 493
rect 787 289 1405 323
rect 1309 173 1359 289
rect 781 139 1411 173
rect 781 51 847 139
rect 969 51 1035 139
rect 1157 51 1223 139
rect 1345 51 1411 139
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 19 394 85 493
rect 119 428 173 527
rect 207 394 273 493
rect 307 428 361 527
rect 395 459 649 493
rect 395 394 455 459
rect 19 360 455 394
rect 19 292 71 360
rect 409 292 455 360
rect 489 358 549 425
rect 489 177 539 358
rect 583 357 649 459
rect 697 299 747 527
rect 875 357 941 527
rect 1063 357 1129 527
rect 1251 357 1317 527
rect 1443 289 1505 527
rect 713 207 1227 255
rect 713 177 747 207
rect 41 17 107 177
rect 207 135 747 177
rect 207 55 273 135
rect 389 17 455 101
rect 489 51 549 135
rect 583 17 747 101
rect 881 17 935 105
rect 1069 17 1123 105
rect 1257 17 1311 105
rect 1445 17 1495 181
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
<< metal1 >>
rect 0 561 1564 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 0 496 1564 527
rect 0 17 1564 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
rect 0 -48 1564 -17
<< labels >>
rlabel locali s 173 211 307 258 6 A1
port 1 nsew signal input
rlabel locali s 341 258 375 292 6 A2
port 2 nsew signal input
rlabel locali s 341 211 409 258 6 A2
port 2 nsew signal input
rlabel locali s 105 292 375 326 6 A2
port 2 nsew signal input
rlabel locali s 105 258 139 292 6 A2
port 2 nsew signal input
rlabel locali s 19 211 139 258 6 A2
port 2 nsew signal input
rlabel locali s 573 211 639 323 6 B1
port 3 nsew signal input
rlabel locali s 1351 323 1405 493 6 X
port 4 nsew signal output
rlabel locali s 1345 51 1411 139 6 X
port 4 nsew signal output
rlabel locali s 1309 173 1359 289 6 X
port 4 nsew signal output
rlabel locali s 1163 323 1217 493 6 X
port 4 nsew signal output
rlabel locali s 1157 51 1223 139 6 X
port 4 nsew signal output
rlabel locali s 975 323 1029 493 6 X
port 4 nsew signal output
rlabel locali s 969 51 1035 139 6 X
port 4 nsew signal output
rlabel locali s 787 323 841 493 6 X
port 4 nsew signal output
rlabel locali s 787 289 1405 323 6 X
port 4 nsew signal output
rlabel locali s 781 139 1411 173 6 X
port 4 nsew signal output
rlabel locali s 781 51 847 139 6 X
port 4 nsew signal output
rlabel metal1 s 0 -48 1564 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 1564 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1564 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3328492
string GDS_START 3316088
<< end >>
