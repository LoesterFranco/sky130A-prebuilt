magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 20 238 146 372
rect 487 363 559 612
rect 506 151 559 363
rect 487 71 559 151
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 19 441 80 545
rect 115 476 181 649
rect 283 530 349 580
rect 19 406 261 441
rect 195 204 261 406
rect 19 164 261 204
rect 295 325 349 530
rect 387 380 453 649
rect 295 259 472 325
rect 19 61 82 164
rect 117 17 183 130
rect 295 61 344 259
rect 387 17 453 150
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
rlabel locali s 20 238 146 372 6 A
port 1 nsew signal input
rlabel locali s 506 151 559 363 6 Y
port 2 nsew signal output
rlabel locali s 487 363 559 612 6 Y
port 2 nsew signal output
rlabel locali s 487 71 559 151 6 Y
port 2 nsew signal output
rlabel metal1 s 0 -49 576 49 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 617 576 715 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 576 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3390492
string GDS_START 3384680
<< end >>
