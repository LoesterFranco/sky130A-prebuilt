magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 1574 704
<< pwell >>
rect 0 0 1536 49
<< scnmos >>
rect 93 74 123 222
rect 184 74 214 222
rect 298 74 328 222
rect 384 74 414 222
rect 484 74 514 222
rect 570 74 600 222
rect 670 74 700 222
rect 756 74 786 222
rect 870 74 900 222
rect 956 74 986 222
rect 1096 74 1126 222
rect 1196 74 1226 222
rect 1296 74 1326 222
<< pmoshvt >>
rect 96 368 126 592
rect 186 368 216 592
rect 276 368 306 592
rect 381 368 411 592
rect 471 368 501 592
rect 561 368 591 592
rect 651 368 681 592
rect 741 368 771 592
rect 943 368 973 592
rect 1033 368 1063 592
rect 1123 368 1153 592
rect 1213 368 1243 592
rect 1330 368 1360 536
rect 1420 368 1450 536
<< ndiff >>
rect 27 210 93 222
rect 27 176 39 210
rect 73 176 93 210
rect 27 120 93 176
rect 27 86 39 120
rect 73 86 93 120
rect 27 74 93 86
rect 123 210 184 222
rect 123 176 139 210
rect 173 176 184 210
rect 123 120 184 176
rect 123 86 139 120
rect 173 86 184 120
rect 123 74 184 86
rect 214 152 298 222
rect 214 118 239 152
rect 273 118 298 152
rect 214 74 298 118
rect 328 210 384 222
rect 328 176 339 210
rect 373 176 384 210
rect 328 120 384 176
rect 328 86 339 120
rect 373 86 384 120
rect 328 74 384 86
rect 414 146 484 222
rect 414 112 439 146
rect 473 112 484 146
rect 414 74 484 112
rect 514 210 570 222
rect 514 176 525 210
rect 559 176 570 210
rect 514 120 570 176
rect 514 86 525 120
rect 559 86 570 120
rect 514 74 570 86
rect 600 146 670 222
rect 600 112 611 146
rect 645 112 670 146
rect 600 74 670 112
rect 700 210 756 222
rect 700 176 711 210
rect 745 176 756 210
rect 700 120 756 176
rect 700 86 711 120
rect 745 86 756 120
rect 700 74 756 86
rect 786 123 870 222
rect 786 89 811 123
rect 845 89 870 123
rect 786 74 870 89
rect 900 210 956 222
rect 900 176 911 210
rect 945 176 956 210
rect 900 120 956 176
rect 900 86 911 120
rect 945 86 956 120
rect 900 74 956 86
rect 986 120 1096 222
rect 986 86 1024 120
rect 1058 86 1096 120
rect 986 74 1096 86
rect 1126 210 1196 222
rect 1126 176 1137 210
rect 1171 176 1196 210
rect 1126 120 1196 176
rect 1126 86 1137 120
rect 1171 86 1196 120
rect 1126 74 1196 86
rect 1226 202 1296 222
rect 1226 168 1237 202
rect 1271 168 1296 202
rect 1226 120 1296 168
rect 1226 86 1237 120
rect 1271 86 1296 120
rect 1226 74 1296 86
rect 1326 202 1509 222
rect 1326 168 1337 202
rect 1371 168 1463 202
rect 1497 168 1509 202
rect 1326 117 1509 168
rect 1326 83 1337 117
rect 1371 83 1463 117
rect 1497 83 1509 117
rect 1326 74 1509 83
<< pdiff >>
rect 27 580 96 592
rect 27 546 39 580
rect 73 546 96 580
rect 27 510 96 546
rect 27 476 39 510
rect 73 476 96 510
rect 27 440 96 476
rect 27 406 39 440
rect 73 406 96 440
rect 27 368 96 406
rect 126 542 186 592
rect 126 508 139 542
rect 173 508 186 542
rect 126 432 186 508
rect 126 398 139 432
rect 173 398 186 432
rect 126 368 186 398
rect 216 580 276 592
rect 216 546 229 580
rect 263 546 276 580
rect 216 508 276 546
rect 216 474 229 508
rect 263 474 276 508
rect 216 368 276 474
rect 306 542 381 592
rect 306 508 321 542
rect 355 508 381 542
rect 306 424 381 508
rect 306 390 321 424
rect 355 390 381 424
rect 306 368 381 390
rect 411 566 471 592
rect 411 532 424 566
rect 458 532 471 566
rect 411 368 471 532
rect 501 414 561 592
rect 501 380 514 414
rect 548 380 561 414
rect 501 368 561 380
rect 591 566 651 592
rect 591 532 604 566
rect 638 532 651 566
rect 591 368 651 532
rect 681 414 741 592
rect 681 380 694 414
rect 728 380 741 414
rect 681 368 741 380
rect 771 566 830 592
rect 771 532 784 566
rect 818 532 830 566
rect 771 368 830 532
rect 884 566 943 592
rect 884 532 896 566
rect 930 532 943 566
rect 884 368 943 532
rect 973 582 1033 592
rect 973 548 986 582
rect 1020 548 1033 582
rect 973 514 1033 548
rect 973 480 986 514
rect 1020 480 1033 514
rect 973 446 1033 480
rect 973 412 986 446
rect 1020 412 1033 446
rect 973 368 1033 412
rect 1063 582 1123 592
rect 1063 548 1076 582
rect 1110 548 1123 582
rect 1063 514 1123 548
rect 1063 480 1076 514
rect 1110 480 1123 514
rect 1063 368 1123 480
rect 1153 582 1213 592
rect 1153 548 1166 582
rect 1200 548 1213 582
rect 1153 514 1213 548
rect 1153 480 1166 514
rect 1200 480 1213 514
rect 1153 446 1213 480
rect 1153 412 1166 446
rect 1200 412 1213 446
rect 1153 368 1213 412
rect 1243 582 1312 592
rect 1243 548 1266 582
rect 1300 548 1312 582
rect 1243 536 1312 548
rect 1243 514 1330 536
rect 1243 480 1266 514
rect 1300 480 1330 514
rect 1243 446 1330 480
rect 1243 412 1266 446
rect 1300 412 1330 446
rect 1243 368 1330 412
rect 1360 524 1420 536
rect 1360 490 1373 524
rect 1407 490 1420 524
rect 1360 414 1420 490
rect 1360 380 1373 414
rect 1407 380 1420 414
rect 1360 368 1420 380
rect 1450 524 1509 536
rect 1450 490 1463 524
rect 1497 490 1509 524
rect 1450 449 1509 490
rect 1450 415 1463 449
rect 1497 415 1509 449
rect 1450 368 1509 415
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 139 176 173 210
rect 139 86 173 120
rect 239 118 273 152
rect 339 176 373 210
rect 339 86 373 120
rect 439 112 473 146
rect 525 176 559 210
rect 525 86 559 120
rect 611 112 645 146
rect 711 176 745 210
rect 711 86 745 120
rect 811 89 845 123
rect 911 176 945 210
rect 911 86 945 120
rect 1024 86 1058 120
rect 1137 176 1171 210
rect 1137 86 1171 120
rect 1237 168 1271 202
rect 1237 86 1271 120
rect 1337 168 1371 202
rect 1463 168 1497 202
rect 1337 83 1371 117
rect 1463 83 1497 117
<< pdiffc >>
rect 39 546 73 580
rect 39 476 73 510
rect 39 406 73 440
rect 139 508 173 542
rect 139 398 173 432
rect 229 546 263 580
rect 229 474 263 508
rect 321 508 355 542
rect 321 390 355 424
rect 424 532 458 566
rect 514 380 548 414
rect 604 532 638 566
rect 694 380 728 414
rect 784 532 818 566
rect 896 532 930 566
rect 986 548 1020 582
rect 986 480 1020 514
rect 986 412 1020 446
rect 1076 548 1110 582
rect 1076 480 1110 514
rect 1166 548 1200 582
rect 1166 480 1200 514
rect 1166 412 1200 446
rect 1266 548 1300 582
rect 1266 480 1300 514
rect 1266 412 1300 446
rect 1373 490 1407 524
rect 1373 380 1407 414
rect 1463 490 1497 524
rect 1463 415 1497 449
<< poly >>
rect 96 592 126 618
rect 186 592 216 618
rect 276 592 306 618
rect 381 592 411 618
rect 471 592 501 618
rect 561 592 591 618
rect 651 592 681 618
rect 741 592 771 618
rect 943 592 973 618
rect 1033 592 1063 618
rect 1123 592 1153 618
rect 1213 592 1243 618
rect 1330 536 1360 562
rect 1420 536 1450 562
rect 96 353 126 368
rect 186 353 216 368
rect 276 353 306 368
rect 381 353 411 368
rect 471 353 501 368
rect 561 353 591 368
rect 651 353 681 368
rect 741 353 771 368
rect 943 353 973 368
rect 1033 353 1063 368
rect 1123 353 1153 368
rect 1213 353 1243 368
rect 1330 353 1360 368
rect 1420 353 1450 368
rect 93 336 129 353
rect 183 336 219 353
rect 273 336 309 353
rect 378 336 414 353
rect 93 320 414 336
rect 93 286 109 320
rect 143 286 177 320
rect 211 286 245 320
rect 279 286 313 320
rect 347 286 414 320
rect 93 270 414 286
rect 93 222 123 270
rect 184 222 214 270
rect 298 222 328 270
rect 384 222 414 270
rect 468 330 504 353
rect 558 330 594 353
rect 648 330 684 353
rect 738 330 774 353
rect 468 314 786 330
rect 468 280 532 314
rect 566 280 600 314
rect 634 280 668 314
rect 702 280 736 314
rect 770 280 786 314
rect 940 310 976 353
rect 1030 310 1066 353
rect 1120 310 1156 353
rect 1210 310 1246 353
rect 468 264 786 280
rect 484 222 514 264
rect 570 222 600 264
rect 670 222 700 264
rect 756 222 786 264
rect 870 294 1246 310
rect 870 260 904 294
rect 938 260 972 294
rect 1006 260 1040 294
rect 1074 260 1108 294
rect 1142 260 1176 294
rect 1210 280 1246 294
rect 1327 352 1363 353
rect 1417 352 1453 353
rect 1327 322 1453 352
rect 1327 294 1447 322
rect 1210 260 1226 280
rect 1327 274 1369 294
rect 870 244 1226 260
rect 870 222 900 244
rect 956 222 986 244
rect 1096 222 1126 244
rect 1196 222 1226 244
rect 1296 260 1369 274
rect 1403 260 1447 294
rect 1296 244 1447 260
rect 1296 222 1326 244
rect 93 48 123 74
rect 184 48 214 74
rect 298 48 328 74
rect 384 48 414 74
rect 484 48 514 74
rect 570 48 600 74
rect 670 48 700 74
rect 756 48 786 74
rect 870 48 900 74
rect 956 48 986 74
rect 1096 48 1126 74
rect 1196 48 1226 74
rect 1296 48 1326 74
<< polycont >>
rect 109 286 143 320
rect 177 286 211 320
rect 245 286 279 320
rect 313 286 347 320
rect 532 280 566 314
rect 600 280 634 314
rect 668 280 702 314
rect 736 280 770 314
rect 904 260 938 294
rect 972 260 1006 294
rect 1040 260 1074 294
rect 1108 260 1142 294
rect 1176 260 1210 294
rect 1369 260 1403 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 23 581 474 615
rect 23 580 89 581
rect 23 546 39 580
rect 73 546 89 580
rect 229 580 263 581
rect 23 510 89 546
rect 23 476 39 510
rect 73 476 89 510
rect 23 440 89 476
rect 23 406 39 440
rect 73 406 89 440
rect 23 390 89 406
rect 123 542 189 547
rect 123 508 139 542
rect 173 508 189 542
rect 123 432 189 508
rect 408 566 474 581
rect 229 508 263 546
rect 229 458 263 474
rect 305 542 371 547
rect 305 508 321 542
rect 355 508 371 542
rect 408 532 424 566
rect 458 550 474 566
rect 588 566 654 582
rect 588 550 604 566
rect 458 532 604 550
rect 638 550 654 566
rect 768 566 834 582
rect 768 550 784 566
rect 638 532 784 550
rect 818 532 834 566
rect 408 516 834 532
rect 880 566 946 649
rect 880 532 896 566
rect 930 532 946 566
rect 880 516 946 532
rect 986 582 1020 598
rect 305 482 371 508
rect 986 514 1020 548
rect 305 480 986 482
rect 1060 582 1126 649
rect 1060 548 1076 582
rect 1110 548 1126 582
rect 1060 514 1126 548
rect 1060 480 1076 514
rect 1110 480 1126 514
rect 1162 582 1216 598
rect 1162 548 1166 582
rect 1200 548 1216 582
rect 1162 514 1216 548
rect 1162 480 1166 514
rect 1200 480 1216 514
rect 123 398 139 432
rect 173 424 189 432
rect 305 448 1020 480
rect 305 424 374 448
rect 173 398 321 424
rect 123 390 321 398
rect 355 390 374 424
rect 959 446 1020 448
rect 1162 446 1216 480
rect 409 380 514 414
rect 548 380 694 414
rect 728 380 744 414
rect 959 412 986 446
rect 1020 412 1166 446
rect 1200 412 1216 446
rect 1250 582 1316 649
rect 1250 548 1266 582
rect 1300 548 1316 582
rect 1250 514 1316 548
rect 1250 480 1266 514
rect 1300 480 1316 514
rect 1250 446 1316 480
rect 1250 412 1266 446
rect 1300 412 1316 446
rect 1357 524 1411 540
rect 1357 490 1373 524
rect 1407 490 1411 524
rect 1357 414 1411 490
rect 409 364 744 380
rect 1357 380 1373 414
rect 1407 380 1411 414
rect 1447 524 1513 649
rect 1447 490 1463 524
rect 1497 490 1513 524
rect 1447 449 1513 490
rect 1447 415 1463 449
rect 1497 415 1513 449
rect 1447 412 1513 415
rect 1357 378 1411 380
rect 25 320 363 356
rect 25 286 109 320
rect 143 286 177 320
rect 211 286 245 320
rect 279 286 313 320
rect 347 286 363 320
rect 25 270 363 286
rect 409 236 455 364
rect 778 344 1513 378
rect 778 330 839 344
rect 516 314 839 330
rect 516 280 532 314
rect 566 280 600 314
rect 634 280 668 314
rect 702 280 736 314
rect 770 280 839 314
rect 516 264 839 280
rect 888 294 1319 310
rect 888 260 904 294
rect 938 260 972 294
rect 1006 260 1040 294
rect 1074 260 1108 294
rect 1142 260 1176 294
rect 1210 260 1319 294
rect 888 244 1319 260
rect 1273 236 1319 244
rect 1353 294 1419 310
rect 1353 260 1369 294
rect 1403 260 1419 294
rect 1353 236 1419 260
rect 123 230 455 236
rect 23 210 89 226
rect 23 176 39 210
rect 73 176 89 210
rect 23 120 89 176
rect 23 86 39 120
rect 73 86 89 120
rect 23 17 89 86
rect 123 210 761 230
rect 123 176 139 210
rect 173 202 339 210
rect 173 176 189 202
rect 123 120 189 176
rect 323 176 339 202
rect 373 196 525 210
rect 373 176 389 196
rect 123 86 139 120
rect 173 86 189 120
rect 123 70 189 86
rect 223 152 289 168
rect 223 118 239 152
rect 273 118 289 152
rect 223 17 289 118
rect 323 120 389 176
rect 559 196 711 210
rect 323 86 339 120
rect 373 86 389 120
rect 323 70 389 86
rect 423 146 489 162
rect 423 112 439 146
rect 473 112 489 146
rect 423 17 489 112
rect 525 120 559 176
rect 695 176 711 196
rect 745 176 911 210
rect 945 176 1137 210
rect 1171 176 1187 210
rect 1479 202 1513 344
rect 525 70 559 86
rect 595 146 661 162
rect 595 112 611 146
rect 645 112 661 146
rect 595 17 661 112
rect 695 120 761 176
rect 695 86 711 120
rect 745 86 761 120
rect 695 70 761 86
rect 795 123 861 142
rect 795 89 811 123
rect 845 89 861 123
rect 795 17 861 89
rect 895 120 961 176
rect 895 86 911 120
rect 945 86 961 120
rect 895 70 961 86
rect 995 120 1087 136
rect 995 86 1024 120
rect 1058 86 1087 120
rect 995 17 1087 86
rect 1121 120 1187 176
rect 1121 86 1137 120
rect 1171 86 1187 120
rect 1121 70 1187 86
rect 1221 168 1237 202
rect 1271 168 1287 202
rect 1221 120 1287 168
rect 1221 86 1237 120
rect 1271 86 1287 120
rect 1221 17 1287 86
rect 1321 168 1337 202
rect 1371 168 1463 202
rect 1497 168 1513 202
rect 1321 117 1513 168
rect 1321 83 1337 117
rect 1371 83 1463 117
rect 1497 83 1513 117
rect 1321 70 1513 83
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
rlabel comment s 0 0 0 0 4 nor3b_4
flabel pwell s 0 0 1536 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 1536 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 1536 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 1536 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 1279 242 1313 276 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 1375 242 1409 276 0 FreeSans 340 0 0 0 C_N
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 1536 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1948140
string GDS_START 1936346
<< end >>
