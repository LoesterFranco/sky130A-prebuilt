magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1196 561
rect 24 364 81 527
rect 196 451 262 527
rect 726 439 782 527
rect 816 417 858 493
rect 892 451 958 527
rect 992 417 1030 493
rect 816 405 1030 417
rect 368 371 1030 405
rect 1064 376 1130 527
rect 787 340 1030 371
rect 115 303 739 337
rect 115 264 295 303
rect 25 203 295 264
rect 397 214 655 269
rect 689 198 739 303
rect 787 289 1167 340
rect 781 203 1051 255
rect 1085 169 1167 289
rect 806 123 1167 169
rect 110 17 176 89
rect 282 17 348 89
rect 454 17 520 89
rect 626 17 692 89
rect 0 -17 1196 17
<< obsli1 >>
rect 115 417 162 493
rect 296 455 692 493
rect 296 417 334 455
rect 115 383 334 417
rect 24 123 772 164
rect 726 89 772 123
rect 726 51 1130 89
<< metal1 >>
rect 0 496 1196 592
rect 0 -48 1196 48
<< labels >>
rlabel locali s 689 198 739 303 6 A1
port 1 nsew signal input
rlabel locali s 115 303 739 337 6 A1
port 1 nsew signal input
rlabel locali s 115 264 295 303 6 A1
port 1 nsew signal input
rlabel locali s 25 203 295 264 6 A1
port 1 nsew signal input
rlabel locali s 397 214 655 269 6 A2
port 2 nsew signal input
rlabel locali s 781 203 1051 255 6 B1
port 3 nsew signal input
rlabel locali s 1085 169 1167 289 6 Y
port 4 nsew signal output
rlabel locali s 992 417 1030 493 6 Y
port 4 nsew signal output
rlabel locali s 816 417 858 493 6 Y
port 4 nsew signal output
rlabel locali s 816 405 1030 417 6 Y
port 4 nsew signal output
rlabel locali s 806 123 1167 169 6 Y
port 4 nsew signal output
rlabel locali s 787 340 1030 371 6 Y
port 4 nsew signal output
rlabel locali s 787 289 1167 340 6 Y
port 4 nsew signal output
rlabel locali s 368 371 1030 405 6 Y
port 4 nsew signal output
rlabel locali s 626 17 692 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 454 17 520 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 282 17 348 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 110 17 176 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 1196 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1196 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 1064 376 1130 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 892 451 958 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 726 439 782 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 196 451 262 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 24 364 81 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 1196 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 1196 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1367280
string GDS_START 1359226
<< end >>
