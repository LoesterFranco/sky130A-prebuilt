magic
tech sky130A
magscale 1 2
timestamp 1604502697
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 90 47 120 177
rect 176 47 206 177
rect 378 47 408 177
rect 470 47 500 177
rect 568 47 598 177
rect 670 47 700 177
<< pmoshvt >>
rect 82 297 118 497
rect 178 297 214 497
rect 370 297 406 497
rect 452 297 488 497
rect 570 297 606 497
rect 666 297 702 497
<< ndiff >>
rect 27 161 90 177
rect 27 127 36 161
rect 70 127 90 161
rect 27 93 90 127
rect 27 59 36 93
rect 70 59 90 93
rect 27 47 90 59
rect 120 47 176 177
rect 206 165 259 177
rect 206 131 217 165
rect 251 131 259 165
rect 206 47 259 131
rect 315 93 378 177
rect 315 59 324 93
rect 358 59 378 93
rect 315 47 378 59
rect 408 163 470 177
rect 408 129 425 163
rect 459 129 470 163
rect 408 47 470 129
rect 500 89 568 177
rect 500 55 515 89
rect 549 55 568 89
rect 500 47 568 55
rect 598 157 670 177
rect 598 123 615 157
rect 649 123 670 157
rect 598 89 670 123
rect 598 55 615 89
rect 649 55 670 89
rect 598 47 670 55
rect 700 89 798 177
rect 700 55 725 89
rect 759 55 798 89
rect 700 47 798 55
<< pdiff >>
rect 27 477 82 497
rect 27 443 35 477
rect 69 443 82 477
rect 27 381 82 443
rect 27 347 35 381
rect 69 347 82 381
rect 27 297 82 347
rect 118 489 178 497
rect 118 455 131 489
rect 165 455 178 489
rect 118 421 178 455
rect 118 387 131 421
rect 165 387 178 421
rect 118 297 178 387
rect 214 464 370 497
rect 214 430 241 464
rect 275 430 314 464
rect 348 430 370 464
rect 214 395 370 430
rect 214 361 241 395
rect 275 361 314 395
rect 348 361 370 395
rect 214 297 370 361
rect 406 297 452 497
rect 488 489 570 497
rect 488 455 511 489
rect 545 455 570 489
rect 488 421 570 455
rect 488 387 511 421
rect 545 387 570 421
rect 488 297 570 387
rect 606 477 666 497
rect 606 443 619 477
rect 653 443 666 477
rect 606 297 666 443
rect 702 485 784 497
rect 702 451 715 485
rect 749 451 784 485
rect 702 297 784 451
<< ndiffc >>
rect 36 127 70 161
rect 36 59 70 93
rect 217 131 251 165
rect 324 59 358 93
rect 425 129 459 163
rect 515 55 549 89
rect 615 123 649 157
rect 615 55 649 89
rect 725 55 759 89
<< pdiffc >>
rect 35 443 69 477
rect 35 347 69 381
rect 131 455 165 489
rect 131 387 165 421
rect 241 430 275 464
rect 314 430 348 464
rect 241 361 275 395
rect 314 361 348 395
rect 511 455 545 489
rect 511 387 545 421
rect 619 443 653 477
rect 715 451 749 485
<< poly >>
rect 82 497 118 523
rect 178 497 214 523
rect 370 497 406 523
rect 452 497 488 523
rect 570 497 606 523
rect 666 497 702 523
rect 82 282 118 297
rect 178 282 214 297
rect 370 282 406 297
rect 452 282 488 297
rect 570 282 606 297
rect 666 282 702 297
rect 80 274 120 282
rect 21 249 120 274
rect 21 215 38 249
rect 72 215 120 249
rect 21 199 120 215
rect 90 177 120 199
rect 176 265 216 282
rect 368 277 408 282
rect 176 249 255 265
rect 176 215 196 249
rect 230 215 255 249
rect 176 199 255 215
rect 320 249 408 277
rect 320 215 345 249
rect 379 215 408 249
rect 320 199 408 215
rect 450 265 490 282
rect 450 249 522 265
rect 450 215 466 249
rect 500 215 522 249
rect 450 199 522 215
rect 568 264 608 282
rect 664 264 704 282
rect 568 249 717 264
rect 568 215 591 249
rect 625 215 659 249
rect 693 215 717 249
rect 568 199 717 215
rect 176 177 206 199
rect 378 177 408 199
rect 470 177 500 199
rect 568 177 598 199
rect 670 177 700 199
rect 90 21 120 47
rect 176 21 206 47
rect 378 21 408 47
rect 470 21 500 47
rect 568 21 598 47
rect 670 21 700 47
<< polycont >>
rect 38 215 72 249
rect 196 215 230 249
rect 345 215 379 249
rect 466 215 500 249
rect 591 215 625 249
rect 659 215 693 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 18 477 71 493
rect 18 443 35 477
rect 69 443 71 477
rect 18 381 71 443
rect 105 489 181 527
rect 105 455 131 489
rect 165 455 181 489
rect 105 421 181 455
rect 105 387 131 421
rect 165 387 181 421
rect 225 464 364 493
rect 225 430 241 464
rect 275 430 314 464
rect 348 430 364 464
rect 225 395 364 430
rect 18 347 35 381
rect 69 353 71 381
rect 225 361 241 395
rect 275 361 314 395
rect 348 361 364 395
rect 475 489 571 527
rect 475 455 511 489
rect 545 455 571 489
rect 475 421 571 455
rect 475 387 511 421
rect 545 387 571 421
rect 617 477 655 493
rect 617 443 619 477
rect 653 443 655 477
rect 689 485 765 527
rect 689 451 715 485
rect 749 451 765 485
rect 617 415 655 443
rect 617 381 807 415
rect 225 353 364 361
rect 69 347 364 353
rect 18 302 605 347
rect 17 249 72 265
rect 17 215 38 249
rect 17 199 72 215
rect 106 165 152 302
rect 571 265 605 302
rect 186 249 262 265
rect 186 215 196 249
rect 230 215 262 249
rect 186 199 262 215
rect 301 249 389 265
rect 301 215 345 249
rect 379 215 389 249
rect 301 199 389 215
rect 433 249 535 265
rect 433 215 466 249
rect 500 215 535 249
rect 433 199 535 215
rect 571 249 713 265
rect 571 215 591 249
rect 625 215 659 249
rect 693 215 713 249
rect 571 199 713 215
rect 19 161 152 165
rect 19 127 36 161
rect 70 127 152 161
rect 186 131 217 165
rect 251 163 475 165
rect 251 131 425 163
rect 186 129 425 131
rect 459 129 475 163
rect 753 157 807 381
rect 186 127 475 129
rect 19 93 152 127
rect 589 123 615 157
rect 649 123 807 157
rect 19 59 36 93
rect 70 85 152 93
rect 70 59 86 85
rect 19 51 86 59
rect 307 59 324 93
rect 358 59 374 93
rect 307 17 374 59
rect 508 89 555 105
rect 508 55 515 89
rect 549 55 555 89
rect 508 17 555 55
rect 589 89 665 123
rect 589 55 615 89
rect 649 55 665 89
rect 589 51 665 55
rect 709 55 725 89
rect 759 55 775 89
rect 709 17 775 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel corelocali s 30 221 64 255 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 210 221 244 255 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 310 221 344 255 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 488 221 522 255 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 766 153 800 187 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
rlabel comment s 0 0 0 0 4 o211a_2
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2574944
string GDS_START 2568348
<< end >>
