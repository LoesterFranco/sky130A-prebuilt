magic
tech sky130A
magscale 1 2
timestamp 1599588232
<< locali >>
rect 95 316 161 428
rect 217 364 317 430
rect 95 282 409 316
rect 359 250 409 282
rect 511 228 556 430
rect 660 236 743 310
rect 2799 430 2855 596
rect 2799 364 2951 430
rect 2865 298 2951 364
rect 2835 264 2951 298
rect 2835 230 2869 264
rect 2798 74 2869 230
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 2976 683
rect 23 498 73 596
rect 113 532 179 649
rect 287 532 477 582
rect 512 566 578 649
rect 443 498 624 532
rect 709 516 775 649
rect 815 579 1146 613
rect 815 516 865 579
rect 23 464 409 498
rect 23 462 73 464
rect 23 246 57 462
rect 359 366 409 464
rect 23 180 245 246
rect 443 216 477 498
rect 590 482 624 498
rect 917 482 983 545
rect 590 448 983 482
rect 1023 453 1073 545
rect 917 414 983 448
rect 592 364 843 414
rect 312 182 477 216
rect 592 202 626 364
rect 777 270 843 364
rect 884 380 983 414
rect 23 70 89 180
rect 123 17 214 136
rect 312 70 378 182
rect 492 17 558 148
rect 592 70 670 202
rect 704 17 770 202
rect 806 85 840 226
rect 884 169 918 380
rect 952 237 993 346
rect 1027 309 1061 453
rect 1112 451 1146 579
rect 1219 485 1269 649
rect 1303 581 1473 615
rect 1303 451 1337 581
rect 1112 417 1337 451
rect 1112 409 1146 417
rect 1095 343 1146 409
rect 1371 383 1405 547
rect 1188 349 1405 383
rect 1439 379 1473 581
rect 1507 413 1541 649
rect 1581 447 1647 551
rect 1687 481 1737 649
rect 1800 581 2087 615
rect 1800 463 1866 581
rect 1581 429 1753 447
rect 1900 429 1966 547
rect 2021 495 2087 581
rect 2216 529 2266 649
rect 2306 495 2372 596
rect 2021 461 2372 495
rect 2412 496 2462 596
rect 2502 530 2568 649
rect 2412 462 2561 496
rect 1581 413 1966 429
rect 2178 428 2372 461
rect 1719 395 1966 413
rect 1439 361 1685 379
rect 2000 361 2144 427
rect 2178 394 2493 428
rect 1188 343 1254 349
rect 1439 345 2034 361
rect 1310 309 1376 314
rect 1027 275 1376 309
rect 952 203 1034 237
rect 884 119 966 169
rect 1000 85 1034 203
rect 806 51 1034 85
rect 1068 77 1118 275
rect 1196 140 1262 241
rect 1310 208 1376 275
rect 1441 276 1511 311
rect 1441 242 1471 276
rect 1505 242 1511 276
rect 1551 245 1617 311
rect 1651 295 2034 345
rect 2178 314 2212 394
rect 2082 280 2212 314
rect 1551 208 1585 245
rect 1310 174 1585 208
rect 1636 177 2016 211
rect 1196 106 1404 140
rect 1226 17 1292 72
rect 1338 70 1404 106
rect 1502 17 1602 136
rect 1636 70 1702 177
rect 1738 17 1804 143
rect 1850 85 1916 143
rect 1950 119 2016 177
rect 2082 162 2116 280
rect 2289 276 2375 360
rect 2050 85 2116 162
rect 2189 192 2255 246
rect 2289 242 2335 276
rect 2369 242 2375 276
rect 2289 236 2375 242
rect 2427 226 2493 394
rect 2527 192 2561 462
rect 2189 158 2561 192
rect 1850 51 2116 85
rect 2328 17 2466 120
rect 2500 70 2561 158
rect 2607 330 2674 596
rect 2708 364 2765 649
rect 2889 464 2955 649
rect 2607 264 2801 330
rect 2607 94 2673 264
rect 2711 17 2761 230
rect 2903 17 2953 230
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 2976 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 1471 242 1505 276
rect 2335 242 2369 276
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
<< metal1 >>
rect 0 683 2976 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 2976 683
rect 0 617 2976 649
rect 0 616 50 617
rect 1459 276 1517 282
rect 1459 242 1471 276
rect 1505 273 1517 276
rect 2323 276 2381 282
rect 2323 273 2335 276
rect 1505 245 2335 273
rect 1505 242 1517 245
rect 1459 236 1517 242
rect 2323 242 2335 245
rect 2369 242 2381 276
rect 2323 236 2381 242
rect 0 49 50 50
rect 0 17 2976 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 2976 17
rect 0 -49 2976 -17
<< labels >>
rlabel locali s 217 364 317 430 6 D
port 1 nsew signal input
rlabel locali s 2865 298 2951 364 6 Q
port 2 nsew signal output
rlabel locali s 2835 264 2951 298 6 Q
port 2 nsew signal output
rlabel locali s 2835 230 2869 264 6 Q
port 2 nsew signal output
rlabel locali s 2799 430 2855 596 6 Q
port 2 nsew signal output
rlabel locali s 2799 364 2951 430 6 Q
port 2 nsew signal output
rlabel locali s 2798 74 2869 230 6 Q
port 2 nsew signal output
rlabel locali s 511 228 556 430 6 SCD
port 3 nsew signal input
rlabel locali s 359 250 409 282 6 SCE
port 4 nsew signal input
rlabel locali s 95 316 161 428 6 SCE
port 4 nsew signal input
rlabel locali s 95 282 409 316 6 SCE
port 4 nsew signal input
rlabel metal1 s 2323 273 2381 282 6 SET_B
port 5 nsew signal input
rlabel metal1 s 2323 236 2381 245 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1459 273 1517 282 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1459 245 2381 273 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1459 236 1517 245 6 SET_B
port 5 nsew signal input
rlabel locali s 660 236 743 310 6 CLK
port 6 nsew clock input
rlabel metal1 s 0 -49 2976 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 8 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 9 nsew power bidirectional
rlabel metal1 s 0 617 2976 715 6 VPWR
port 10 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2976 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 105368
string GDS_START 83718
<< end >>
