magic
tech sky130A
magscale 1 2
timestamp 1599588218
<< nwell >>
rect -38 335 2342 704
rect -38 332 258 335
rect 629 332 2342 335
rect 629 311 1386 332
<< pwell >>
rect 0 0 2304 49
<< scpmos >>
rect 81 527 117 611
rect 171 527 207 611
rect 367 387 403 611
rect 457 387 493 611
rect 663 463 699 547
rect 753 463 789 547
rect 837 463 873 547
rect 961 463 997 547
rect 1163 347 1199 547
rect 1264 362 1300 562
rect 1445 493 1481 577
rect 1529 493 1565 577
rect 1629 493 1665 577
rect 1771 493 1807 577
rect 1888 409 1924 577
rect 2095 368 2131 592
rect 2185 368 2221 592
<< nmoslvt >>
rect 87 78 117 162
rect 165 78 195 162
rect 363 119 393 267
rect 477 119 507 267
rect 687 138 717 222
rect 787 138 817 222
rect 865 138 895 222
rect 943 138 973 222
rect 1146 74 1176 222
rect 1241 74 1271 222
rect 1451 81 1481 165
rect 1529 81 1559 165
rect 1633 81 1663 165
rect 1711 81 1741 165
rect 1907 74 1937 222
rect 2105 74 2135 222
rect 2191 74 2221 222
<< ndiff >>
rect 306 230 363 267
rect 306 196 318 230
rect 352 196 363 230
rect 306 162 363 196
rect 30 137 87 162
rect 30 103 42 137
rect 76 103 87 137
rect 30 78 87 103
rect 117 78 165 162
rect 195 136 252 162
rect 195 102 206 136
rect 240 102 252 136
rect 306 128 318 162
rect 352 128 363 162
rect 306 119 363 128
rect 393 162 477 267
rect 393 128 418 162
rect 452 128 477 162
rect 393 119 477 128
rect 507 198 557 267
rect 507 162 564 198
rect 507 128 518 162
rect 552 128 564 162
rect 630 197 687 222
rect 630 163 642 197
rect 676 163 687 197
rect 630 138 687 163
rect 717 190 787 222
rect 717 156 742 190
rect 776 156 787 190
rect 717 138 787 156
rect 817 138 865 222
rect 895 138 943 222
rect 973 138 1146 222
rect 507 119 564 128
rect 195 78 252 102
rect 988 74 1146 138
rect 1176 189 1241 222
rect 1176 155 1187 189
rect 1221 155 1241 189
rect 1176 74 1241 155
rect 1271 165 1321 222
rect 1851 194 1907 222
rect 1271 153 1451 165
rect 1271 119 1287 153
rect 1321 119 1373 153
rect 1407 119 1451 153
rect 1271 81 1451 119
rect 1481 81 1529 165
rect 1559 127 1633 165
rect 1559 93 1579 127
rect 1613 93 1633 127
rect 1559 81 1633 93
rect 1663 81 1711 165
rect 1741 140 1797 165
rect 1741 106 1752 140
rect 1786 106 1797 140
rect 1741 81 1797 106
rect 1851 160 1862 194
rect 1896 160 1907 194
rect 1851 120 1907 160
rect 1851 86 1862 120
rect 1896 86 1907 120
rect 1271 74 1321 81
rect 988 73 1065 74
rect 988 39 1009 73
rect 1043 39 1065 73
rect 1851 74 1907 86
rect 1937 209 1994 222
rect 1937 175 1948 209
rect 1982 175 1994 209
rect 1937 120 1994 175
rect 1937 86 1948 120
rect 1982 86 1994 120
rect 1937 74 1994 86
rect 2048 210 2105 222
rect 2048 176 2060 210
rect 2094 176 2105 210
rect 2048 120 2105 176
rect 2048 86 2060 120
rect 2094 86 2105 120
rect 2048 74 2105 86
rect 2135 210 2191 222
rect 2135 176 2146 210
rect 2180 176 2191 210
rect 2135 120 2191 176
rect 2135 86 2146 120
rect 2180 86 2191 120
rect 2135 74 2191 86
rect 2221 210 2277 222
rect 2221 176 2232 210
rect 2266 176 2277 210
rect 2221 120 2277 176
rect 2221 86 2232 120
rect 2266 86 2277 120
rect 2221 74 2277 86
rect 988 27 1065 39
<< pdiff >>
rect 27 586 81 611
rect 27 552 37 586
rect 71 552 81 586
rect 27 527 81 552
rect 117 586 171 611
rect 117 552 127 586
rect 161 552 171 586
rect 117 527 171 552
rect 207 593 260 611
rect 207 559 217 593
rect 251 559 260 593
rect 207 527 260 559
rect 314 439 367 611
rect 314 405 323 439
rect 357 405 367 439
rect 314 387 367 405
rect 403 593 457 611
rect 403 559 413 593
rect 447 559 457 593
rect 403 387 457 559
rect 493 439 546 611
rect 493 405 503 439
rect 537 405 546 439
rect 493 387 546 405
rect 888 573 946 597
rect 888 547 900 573
rect 608 524 663 547
rect 608 490 618 524
rect 652 490 663 524
rect 608 463 663 490
rect 699 539 753 547
rect 699 505 709 539
rect 743 505 753 539
rect 699 463 753 505
rect 789 463 837 547
rect 873 539 900 547
rect 934 547 946 573
rect 2034 580 2095 592
rect 1395 562 1445 577
rect 1214 547 1264 562
rect 934 539 961 547
rect 873 463 961 539
rect 997 505 1053 547
rect 997 471 1007 505
rect 1041 471 1053 505
rect 997 463 1053 471
rect 1107 535 1163 547
rect 1107 501 1119 535
rect 1153 501 1163 535
rect 1107 467 1163 501
rect 1107 433 1119 467
rect 1153 433 1163 467
rect 1107 399 1163 433
rect 1107 365 1119 399
rect 1153 365 1163 399
rect 1107 347 1163 365
rect 1199 535 1264 547
rect 1199 501 1219 535
rect 1253 501 1264 535
rect 1199 421 1264 501
rect 1199 387 1219 421
rect 1253 387 1264 421
rect 1199 362 1264 387
rect 1300 545 1445 562
rect 1300 511 1319 545
rect 1353 511 1401 545
rect 1435 511 1445 545
rect 1300 493 1445 511
rect 1481 493 1529 577
rect 1565 552 1629 577
rect 1565 518 1575 552
rect 1609 518 1629 552
rect 1565 493 1629 518
rect 1665 539 1771 577
rect 1665 505 1701 539
rect 1735 505 1771 539
rect 1665 493 1771 505
rect 1807 552 1888 577
rect 1807 518 1834 552
rect 1868 518 1888 552
rect 1807 493 1888 518
rect 1300 362 1350 493
rect 1199 347 1249 362
rect 1822 409 1888 493
rect 1924 565 1980 577
rect 1924 531 1934 565
rect 1968 531 1980 565
rect 1924 456 1980 531
rect 1924 422 1934 456
rect 1968 422 1980 456
rect 1924 409 1980 422
rect 2034 546 2046 580
rect 2080 546 2095 580
rect 2034 497 2095 546
rect 2034 463 2046 497
rect 2080 463 2095 497
rect 2034 414 2095 463
rect 2034 380 2046 414
rect 2080 380 2095 414
rect 2034 368 2095 380
rect 2131 580 2185 592
rect 2131 546 2141 580
rect 2175 546 2185 580
rect 2131 497 2185 546
rect 2131 463 2141 497
rect 2175 463 2185 497
rect 2131 414 2185 463
rect 2131 380 2141 414
rect 2175 380 2185 414
rect 2131 368 2185 380
rect 2221 580 2277 592
rect 2221 546 2231 580
rect 2265 546 2277 580
rect 2221 497 2277 546
rect 2221 463 2231 497
rect 2265 463 2277 497
rect 2221 414 2277 463
rect 2221 380 2231 414
rect 2265 380 2277 414
rect 2221 368 2277 380
<< ndiffc >>
rect 318 196 352 230
rect 42 103 76 137
rect 206 102 240 136
rect 318 128 352 162
rect 418 128 452 162
rect 518 128 552 162
rect 642 163 676 197
rect 742 156 776 190
rect 1187 155 1221 189
rect 1287 119 1321 153
rect 1373 119 1407 153
rect 1579 93 1613 127
rect 1752 106 1786 140
rect 1862 160 1896 194
rect 1862 86 1896 120
rect 1009 39 1043 73
rect 1948 175 1982 209
rect 1948 86 1982 120
rect 2060 176 2094 210
rect 2060 86 2094 120
rect 2146 176 2180 210
rect 2146 86 2180 120
rect 2232 176 2266 210
rect 2232 86 2266 120
<< pdiffc >>
rect 37 552 71 586
rect 127 552 161 586
rect 217 559 251 593
rect 323 405 357 439
rect 413 559 447 593
rect 503 405 537 439
rect 618 490 652 524
rect 709 505 743 539
rect 900 539 934 573
rect 1007 471 1041 505
rect 1119 501 1153 535
rect 1119 433 1153 467
rect 1119 365 1153 399
rect 1219 501 1253 535
rect 1219 387 1253 421
rect 1319 511 1353 545
rect 1401 511 1435 545
rect 1575 518 1609 552
rect 1701 505 1735 539
rect 1834 518 1868 552
rect 1934 531 1968 565
rect 1934 422 1968 456
rect 2046 546 2080 580
rect 2046 463 2080 497
rect 2046 380 2080 414
rect 2141 546 2175 580
rect 2141 463 2175 497
rect 2141 380 2175 414
rect 2231 546 2265 580
rect 2231 463 2265 497
rect 2231 380 2265 414
<< poly >>
rect 81 611 117 637
rect 171 611 207 637
rect 367 611 403 637
rect 457 611 493 637
rect 561 615 1300 645
rect 81 402 117 527
rect 171 430 207 527
rect 44 386 117 402
rect 44 352 60 386
rect 94 352 117 386
rect 44 318 117 352
rect 44 284 60 318
rect 94 284 117 318
rect 44 250 117 284
rect 44 216 60 250
rect 94 216 117 250
rect 44 200 117 216
rect 87 162 117 200
rect 165 414 257 430
rect 165 380 207 414
rect 241 380 257 414
rect 165 346 257 380
rect 367 355 403 387
rect 457 355 493 387
rect 561 355 591 615
rect 663 547 699 573
rect 753 547 789 615
rect 837 547 873 573
rect 961 547 997 573
rect 1163 547 1199 573
rect 1264 562 1300 615
rect 1445 577 1481 603
rect 1529 577 1565 603
rect 1629 577 1665 603
rect 1771 577 1807 603
rect 1888 577 1924 603
rect 2095 592 2131 618
rect 2185 592 2221 618
rect 663 387 699 463
rect 753 431 789 463
rect 165 312 207 346
rect 241 312 257 346
rect 165 278 257 312
rect 349 339 415 355
rect 349 305 365 339
rect 399 305 415 339
rect 349 289 415 305
rect 457 339 591 355
rect 457 305 503 339
rect 537 306 591 339
rect 633 371 699 387
rect 633 337 649 371
rect 683 351 699 371
rect 837 425 873 463
rect 961 425 997 463
rect 837 409 905 425
rect 837 375 855 409
rect 889 375 905 409
rect 837 359 905 375
rect 961 409 1057 425
rect 961 375 1007 409
rect 1041 375 1057 409
rect 961 359 1057 375
rect 683 337 795 351
rect 633 326 795 337
rect 637 321 795 326
rect 765 311 795 321
rect 537 305 596 306
rect 457 301 596 305
rect 457 296 599 301
rect 457 290 603 296
rect 165 244 207 278
rect 241 244 257 278
rect 363 267 393 289
rect 457 282 608 290
rect 477 267 507 282
rect 568 278 608 282
rect 765 281 817 311
rect 570 275 608 278
rect 571 273 608 275
rect 165 228 257 244
rect 165 162 195 228
rect 572 237 717 273
rect 687 222 717 237
rect 787 222 817 281
rect 865 222 895 359
rect 961 267 991 359
rect 1445 461 1481 493
rect 1391 445 1481 461
rect 1391 411 1407 445
rect 1441 411 1481 445
rect 1391 395 1481 411
rect 1529 395 1565 493
rect 1629 455 1665 493
rect 1613 439 1679 455
rect 1613 405 1629 439
rect 1663 405 1679 439
rect 1264 347 1300 362
rect 1163 315 1199 347
rect 1264 317 1481 347
rect 943 237 991 267
rect 1071 299 1199 315
rect 1071 265 1087 299
rect 1121 285 1199 299
rect 1121 265 1176 285
rect 1071 249 1176 265
rect 943 222 973 237
rect 1146 222 1176 249
rect 1241 253 1409 269
rect 1241 239 1359 253
rect 1241 222 1271 239
rect 363 93 393 119
rect 477 93 507 119
rect 687 112 717 138
rect 787 112 817 138
rect 865 112 895 138
rect 87 52 117 78
rect 165 51 195 78
rect 943 51 973 138
rect 165 21 973 51
rect 1343 219 1359 239
rect 1393 219 1409 253
rect 1343 203 1409 219
rect 1451 165 1481 317
rect 1529 278 1559 395
rect 1613 389 1679 405
rect 1525 262 1591 278
rect 1525 228 1541 262
rect 1575 228 1591 262
rect 1525 212 1591 228
rect 1529 165 1559 212
rect 1633 165 1663 389
rect 1771 378 1807 493
rect 1741 362 1807 378
rect 1741 341 1757 362
rect 1711 328 1757 341
rect 1791 341 1807 362
rect 1888 341 1924 409
rect 1791 328 1937 341
rect 1711 311 1937 328
rect 1711 165 1741 311
rect 1907 222 1937 311
rect 1985 310 2051 326
rect 1985 276 2001 310
rect 2035 290 2051 310
rect 2095 290 2131 368
rect 2185 290 2221 368
rect 2035 276 2221 290
rect 1985 260 2221 276
rect 2105 222 2135 260
rect 2191 222 2221 260
rect 1146 48 1176 74
rect 1241 48 1271 74
rect 1451 55 1481 81
rect 1529 55 1559 81
rect 1633 55 1663 81
rect 1711 55 1741 81
rect 1907 48 1937 74
rect 2105 48 2135 74
rect 2191 48 2221 74
<< polycont >>
rect 60 352 94 386
rect 60 284 94 318
rect 60 216 94 250
rect 207 380 241 414
rect 207 312 241 346
rect 365 305 399 339
rect 503 305 537 339
rect 649 337 683 371
rect 855 375 889 409
rect 1007 375 1041 409
rect 207 244 241 278
rect 1407 411 1441 445
rect 1629 405 1663 439
rect 1087 265 1121 299
rect 1359 219 1393 253
rect 1541 228 1575 262
rect 1757 328 1791 362
rect 2001 276 2035 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2304 683
rect 21 586 87 649
rect 21 552 37 586
rect 71 552 87 586
rect 21 504 87 552
rect 127 586 167 611
rect 161 552 167 586
rect 201 593 267 649
rect 201 559 217 593
rect 251 559 267 593
rect 397 593 463 649
rect 397 559 413 593
rect 447 559 463 593
rect 884 573 950 649
rect 127 525 167 552
rect 603 525 675 545
rect 127 524 675 525
rect 127 504 618 524
rect 133 490 618 504
rect 652 490 675 524
rect 133 489 675 490
rect 709 539 850 572
rect 884 539 900 573
rect 934 539 950 573
rect 743 505 850 539
rect 1103 535 1169 649
rect 709 489 1007 505
rect 25 386 99 434
rect 25 352 60 386
rect 94 352 99 386
rect 25 318 99 352
rect 25 284 60 318
rect 94 284 99 318
rect 25 250 99 284
rect 25 216 60 250
rect 94 216 99 250
rect 25 200 99 216
rect 133 166 167 489
rect 641 455 675 489
rect 786 471 1007 489
rect 1041 471 1057 505
rect 786 464 1057 471
rect 1103 501 1119 535
rect 1153 501 1169 535
rect 1103 467 1169 501
rect 786 459 957 464
rect 291 439 373 455
rect 201 424 257 430
rect 201 414 223 424
rect 201 380 207 414
rect 241 380 257 390
rect 201 346 257 380
rect 201 312 207 346
rect 241 312 257 346
rect 201 278 257 312
rect 201 244 207 278
rect 241 244 257 278
rect 201 228 257 244
rect 291 405 323 439
rect 357 405 373 439
rect 291 389 373 405
rect 503 439 607 455
rect 537 405 607 439
rect 641 421 752 455
rect 503 397 611 405
rect 503 389 616 397
rect 291 230 325 389
rect 565 387 616 389
rect 565 379 684 387
rect 570 371 684 379
rect 409 355 455 356
rect 359 339 455 355
rect 359 305 365 339
rect 399 305 455 339
rect 503 339 540 355
rect 359 264 455 305
rect 489 305 503 310
rect 537 305 540 339
rect 489 230 540 305
rect 291 196 318 230
rect 352 196 540 230
rect 574 337 649 371
rect 683 337 684 371
rect 574 321 684 337
rect 26 137 167 166
rect 26 103 42 137
rect 76 132 167 137
rect 206 136 256 166
rect 76 103 92 132
rect 26 74 92 103
rect 240 102 256 136
rect 291 162 368 196
rect 574 162 608 321
rect 718 281 752 421
rect 291 128 318 162
rect 352 128 368 162
rect 291 112 368 128
rect 402 128 418 162
rect 452 128 468 162
rect 206 17 256 102
rect 402 17 468 128
rect 502 128 518 162
rect 552 128 608 162
rect 642 247 752 281
rect 642 197 692 247
rect 786 213 820 459
rect 676 163 692 197
rect 642 134 692 163
rect 726 190 820 213
rect 854 409 889 425
rect 854 375 855 409
rect 854 225 889 375
rect 923 315 957 459
rect 1103 433 1119 467
rect 1153 433 1169 467
rect 991 424 1057 430
rect 1025 409 1057 424
rect 991 375 1007 390
rect 1041 375 1057 409
rect 991 359 1057 375
rect 1103 399 1169 433
rect 1103 365 1119 399
rect 1153 365 1169 399
rect 1103 349 1169 365
rect 1203 535 1269 551
rect 1203 501 1219 535
rect 1253 501 1269 535
rect 1203 421 1269 501
rect 1203 387 1219 421
rect 1253 387 1269 421
rect 1203 371 1269 387
rect 1303 545 1525 561
rect 1303 511 1319 545
rect 1353 511 1401 545
rect 1435 511 1525 545
rect 1303 495 1525 511
rect 923 299 1137 315
rect 923 265 1087 299
rect 1121 265 1137 299
rect 923 259 1137 265
rect 1203 226 1237 371
rect 1303 337 1337 495
rect 1171 225 1237 226
rect 854 191 1237 225
rect 726 156 742 190
rect 776 156 820 190
rect 1171 189 1237 191
rect 726 134 820 156
rect 502 100 608 128
rect 854 123 1137 157
rect 854 100 888 123
rect 502 66 888 100
rect 984 73 1069 89
rect 984 39 1009 73
rect 1043 39 1069 73
rect 1103 85 1137 123
rect 1171 155 1187 189
rect 1221 155 1237 189
rect 1171 119 1237 155
rect 1271 303 1337 337
rect 1391 445 1457 461
rect 1391 411 1407 445
rect 1441 411 1457 445
rect 1271 169 1305 303
rect 1391 269 1457 411
rect 1491 346 1525 495
rect 1559 552 1625 649
rect 1559 518 1575 552
rect 1609 518 1625 552
rect 1559 489 1625 518
rect 1659 539 1777 555
rect 1659 505 1701 539
rect 1735 505 1777 539
rect 1659 489 1777 505
rect 1818 552 1884 649
rect 1818 518 1834 552
rect 1868 518 1884 552
rect 1818 489 1884 518
rect 1918 565 1984 581
rect 1918 531 1934 565
rect 1968 531 1984 565
rect 1743 455 1777 489
rect 1918 456 1984 531
rect 1561 439 1679 455
rect 1561 424 1629 439
rect 1561 390 1567 424
rect 1601 405 1629 424
rect 1663 405 1679 439
rect 1743 421 1875 455
rect 1601 390 1679 405
rect 1561 384 1679 390
rect 1741 362 1807 378
rect 1741 346 1757 362
rect 1491 328 1757 346
rect 1791 328 1807 362
rect 1491 312 1807 328
rect 1841 278 1875 421
rect 1918 422 1934 456
rect 1968 422 1984 456
rect 1918 406 1984 422
rect 1345 253 1491 269
rect 1345 219 1359 253
rect 1393 219 1491 253
rect 1345 203 1491 219
rect 1525 262 1875 278
rect 1525 228 1541 262
rect 1575 244 1875 262
rect 1932 326 1984 406
rect 2030 580 2096 649
rect 2030 546 2046 580
rect 2080 546 2096 580
rect 2030 497 2096 546
rect 2030 463 2046 497
rect 2080 463 2096 497
rect 2030 414 2096 463
rect 2030 380 2046 414
rect 2080 380 2096 414
rect 2030 364 2096 380
rect 2130 580 2196 596
rect 2130 546 2141 580
rect 2175 546 2196 580
rect 2130 497 2196 546
rect 2130 463 2141 497
rect 2175 463 2196 497
rect 2130 414 2196 463
rect 2130 380 2141 414
rect 2175 380 2196 414
rect 1932 310 2038 326
rect 1932 276 2001 310
rect 2035 276 2038 310
rect 1932 260 2038 276
rect 1575 228 1591 244
rect 1525 212 1591 228
rect 1271 153 1423 169
rect 1271 119 1287 153
rect 1321 119 1373 153
rect 1407 119 1423 153
rect 1457 85 1491 203
rect 1103 51 1491 85
rect 1554 127 1638 143
rect 1554 93 1579 127
rect 1613 93 1638 127
rect 984 17 1069 39
rect 1554 17 1638 93
rect 1736 140 1802 244
rect 1736 106 1752 140
rect 1786 106 1802 140
rect 1736 77 1802 106
rect 1846 194 1896 210
rect 1846 160 1862 194
rect 1846 120 1896 160
rect 1846 86 1862 120
rect 1846 17 1896 86
rect 1932 209 1998 260
rect 1932 175 1948 209
rect 1982 175 1998 209
rect 1932 120 1998 175
rect 1932 86 1948 120
rect 1982 86 1998 120
rect 1932 70 1998 86
rect 2044 210 2094 226
rect 2044 176 2060 210
rect 2044 120 2094 176
rect 2044 86 2060 120
rect 2044 17 2094 86
rect 2130 210 2196 380
rect 2231 580 2281 649
rect 2265 546 2281 580
rect 2231 497 2281 546
rect 2265 463 2281 497
rect 2231 414 2281 463
rect 2265 380 2281 414
rect 2231 364 2281 380
rect 2130 176 2146 210
rect 2180 176 2196 210
rect 2130 120 2196 176
rect 2130 86 2146 120
rect 2180 86 2196 120
rect 2130 70 2196 86
rect 2232 210 2282 226
rect 2266 176 2282 210
rect 2232 120 2282 176
rect 2266 86 2282 120
rect 2232 17 2282 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2304 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 223 414 257 424
rect 223 390 241 414
rect 241 390 257 414
rect 991 409 1025 424
rect 991 390 1007 409
rect 1007 390 1025 409
rect 1567 390 1601 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
<< metal1 >>
rect 0 683 2304 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2304 683
rect 0 617 2304 649
rect 211 424 269 430
rect 211 390 223 424
rect 257 421 269 424
rect 979 424 1037 430
rect 979 421 991 424
rect 257 393 991 421
rect 257 390 269 393
rect 211 384 269 390
rect 979 390 991 393
rect 1025 421 1037 424
rect 1555 424 1613 430
rect 1555 421 1567 424
rect 1025 393 1567 421
rect 1025 390 1037 393
rect 979 384 1037 390
rect 1555 390 1567 393
rect 1601 390 1613 424
rect 1555 384 1613 390
rect 0 17 2304 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2304 17
rect 0 -49 2304 -17
<< labels >>
flabel pwell s 0 0 2304 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 0 617 2304 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
rlabel comment s 0 0 0 0 4 dfrtp_2
flabel comment s 943 630 943 630 0 FreeSans 300 0 0 0 no_jumper_check
flabel comment s 552 36 552 36 0 FreeSans 300 0 0 0 no_jumper_check
flabel metal1 s 223 390 257 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew
flabel metal1 s 0 617 2304 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 2304 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 31 390 65 424 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 2143 94 2177 128 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 2143 168 2177 202 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 2143 242 2177 276 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 2143 316 2177 350 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 2143 390 2177 424 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 2143 464 2177 498 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 2143 538 2177 572 0 FreeSans 340 0 0 0 Q
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 2304 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 2867410
string GDS_START 2849740
<< end >>
