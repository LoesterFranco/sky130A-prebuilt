magic
tech sky130A
magscale 1 2
timestamp 1604502729
<< locali >>
rect 160 264 226 352
rect 268 310 615 360
rect 811 394 845 596
rect 975 394 1041 596
rect 811 360 1127 394
rect 268 298 334 310
rect 657 276 709 310
rect 601 264 709 276
rect 160 230 709 264
rect 1081 226 1127 360
rect 21 51 155 128
rect 811 192 1127 226
rect 811 70 845 192
rect 977 70 1027 192
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 22 268 72 596
rect 112 388 178 649
rect 214 506 280 596
rect 316 540 567 596
rect 601 506 667 596
rect 214 472 667 506
rect 214 394 280 472
rect 601 462 667 472
rect 701 462 767 649
rect 406 428 477 438
rect 406 394 777 428
rect 22 196 93 268
rect 743 326 777 394
rect 885 428 935 649
rect 1081 428 1131 649
rect 743 260 1035 326
rect 743 196 777 260
rect 22 162 382 196
rect 189 17 282 128
rect 316 62 382 162
rect 416 162 777 196
rect 416 70 482 162
rect 516 17 582 128
rect 618 70 668 162
rect 702 17 770 120
rect 881 17 931 158
rect 1063 17 1129 158
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
rlabel locali s 657 276 709 310 6 A
port 1 nsew signal input
rlabel locali s 601 264 709 276 6 A
port 1 nsew signal input
rlabel locali s 160 264 226 352 6 A
port 1 nsew signal input
rlabel locali s 160 230 709 264 6 A
port 1 nsew signal input
rlabel locali s 268 310 615 360 6 B
port 2 nsew signal input
rlabel locali s 268 298 334 310 6 B
port 2 nsew signal input
rlabel locali s 21 51 155 128 6 C_N
port 3 nsew signal input
rlabel locali s 1081 226 1127 360 6 X
port 4 nsew signal output
rlabel locali s 977 70 1027 192 6 X
port 4 nsew signal output
rlabel locali s 975 394 1041 596 6 X
port 4 nsew signal output
rlabel locali s 811 394 845 596 6 X
port 4 nsew signal output
rlabel locali s 811 360 1127 394 6 X
port 4 nsew signal output
rlabel locali s 811 192 1127 226 6 X
port 4 nsew signal output
rlabel locali s 811 70 845 192 6 X
port 4 nsew signal output
rlabel metal1 s 0 -49 1152 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 617 1152 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 844070
string GDS_START 833878
<< end >>
