magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1012 561
rect 103 425 175 527
rect 17 199 66 323
rect 291 379 357 527
rect 459 379 531 527
rect 638 323 704 425
rect 806 323 872 425
rect 638 289 872 323
rect 638 170 714 289
rect 748 204 995 255
rect 103 17 169 97
rect 275 17 341 97
rect 443 17 511 97
rect 638 127 995 170
rect 0 -17 1012 17
<< obsli1 >>
rect 17 391 69 493
rect 17 357 175 391
rect 100 265 175 357
rect 215 345 257 493
rect 391 345 425 493
rect 565 459 995 493
rect 565 345 599 459
rect 215 311 599 345
rect 738 357 772 459
rect 906 289 995 459
rect 100 199 604 265
rect 100 165 139 199
rect 17 131 139 165
rect 207 131 604 165
rect 17 51 69 131
rect 207 51 241 131
rect 375 51 409 131
rect 547 93 604 131
rect 547 51 995 93
<< metal1 >>
rect 0 496 1012 592
rect 0 -48 1012 48
<< labels >>
rlabel locali s 748 204 995 255 6 A
port 1 nsew signal input
rlabel locali s 17 199 66 323 6 TE
port 2 nsew signal input
rlabel locali s 806 323 872 425 6 Z
port 3 nsew signal output
rlabel locali s 638 323 704 425 6 Z
port 3 nsew signal output
rlabel locali s 638 289 872 323 6 Z
port 3 nsew signal output
rlabel locali s 638 170 714 289 6 Z
port 3 nsew signal output
rlabel locali s 638 127 995 170 6 Z
port 3 nsew signal output
rlabel locali s 443 17 511 97 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 275 17 341 97 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 103 17 169 97 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 1012 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1012 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 459 379 531 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 291 379 357 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 103 425 175 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 1012 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 1012 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1012 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2926804
string GDS_START 2918840
<< end >>
