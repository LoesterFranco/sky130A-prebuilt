magic
tech sky130A
magscale 1 2
timestamp 1604502710
<< nwell >>
rect -38 332 1190 704
<< pwell >>
rect 0 0 1152 49
<< scpmos >>
rect 91 368 127 592
rect 181 368 217 592
rect 343 368 379 592
rect 440 368 476 592
rect 533 368 569 592
rect 633 368 669 592
rect 743 368 779 592
rect 843 368 879 592
rect 933 368 969 592
rect 1023 368 1059 592
<< nmoslvt >>
rect 84 74 114 222
rect 170 74 200 222
rect 368 85 398 233
rect 454 85 484 233
rect 540 85 570 233
rect 651 85 681 233
rect 737 85 767 233
rect 843 85 873 233
rect 939 85 969 233
rect 1037 85 1067 233
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 189 170 222
rect 114 155 125 189
rect 159 155 170 189
rect 114 74 170 155
rect 200 210 257 222
rect 200 176 211 210
rect 245 176 257 210
rect 200 120 257 176
rect 200 86 211 120
rect 245 86 257 120
rect 200 74 257 86
rect 311 148 368 233
rect 311 114 323 148
rect 357 114 368 148
rect 311 85 368 114
rect 398 194 454 233
rect 398 160 409 194
rect 443 160 454 194
rect 398 85 454 160
rect 484 148 540 233
rect 484 114 495 148
rect 529 114 540 148
rect 484 85 540 114
rect 570 221 651 233
rect 570 187 601 221
rect 635 187 651 221
rect 570 153 651 187
rect 570 119 600 153
rect 634 119 651 153
rect 570 85 651 119
rect 681 220 737 233
rect 681 186 692 220
rect 726 186 737 220
rect 681 131 737 186
rect 681 97 692 131
rect 726 97 737 131
rect 681 85 737 97
rect 767 148 843 233
rect 767 114 792 148
rect 826 114 843 148
rect 767 85 843 114
rect 873 220 939 233
rect 873 186 892 220
rect 926 186 939 220
rect 873 131 939 186
rect 873 97 892 131
rect 926 97 939 131
rect 873 85 939 97
rect 969 148 1037 233
rect 969 114 992 148
rect 1026 114 1037 148
rect 969 85 1037 114
rect 1067 220 1125 233
rect 1067 186 1078 220
rect 1112 186 1125 220
rect 1067 131 1125 186
rect 1067 97 1078 131
rect 1112 97 1125 131
rect 1067 85 1125 97
<< pdiff >>
rect 35 580 91 592
rect 35 546 47 580
rect 81 546 91 580
rect 35 510 91 546
rect 35 476 47 510
rect 81 476 91 510
rect 35 440 91 476
rect 35 406 47 440
rect 81 406 91 440
rect 35 368 91 406
rect 127 580 181 592
rect 127 546 137 580
rect 171 546 181 580
rect 127 497 181 546
rect 127 463 137 497
rect 171 463 181 497
rect 127 414 181 463
rect 127 380 137 414
rect 171 380 181 414
rect 127 368 181 380
rect 217 576 343 592
rect 217 542 227 576
rect 261 542 299 576
rect 333 542 343 576
rect 217 368 343 542
rect 379 578 440 592
rect 379 544 389 578
rect 423 544 440 578
rect 379 368 440 544
rect 476 519 533 592
rect 476 485 489 519
rect 523 485 533 519
rect 476 368 533 485
rect 569 578 633 592
rect 569 544 589 578
rect 623 544 633 578
rect 569 368 633 544
rect 669 578 743 592
rect 669 544 689 578
rect 723 544 743 578
rect 669 368 743 544
rect 779 578 843 592
rect 779 544 789 578
rect 823 544 843 578
rect 779 368 843 544
rect 879 519 933 592
rect 879 485 889 519
rect 923 485 933 519
rect 879 368 933 485
rect 969 580 1023 592
rect 969 546 979 580
rect 1013 546 1023 580
rect 969 508 1023 546
rect 969 474 979 508
rect 1013 474 1023 508
rect 969 368 1023 474
rect 1059 580 1125 592
rect 1059 546 1079 580
rect 1113 546 1125 580
rect 1059 508 1125 546
rect 1059 474 1079 508
rect 1113 474 1125 508
rect 1059 368 1125 474
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 125 155 159 189
rect 211 176 245 210
rect 211 86 245 120
rect 323 114 357 148
rect 409 160 443 194
rect 495 114 529 148
rect 601 187 635 221
rect 600 119 634 153
rect 692 186 726 220
rect 692 97 726 131
rect 792 114 826 148
rect 892 186 926 220
rect 892 97 926 131
rect 992 114 1026 148
rect 1078 186 1112 220
rect 1078 97 1112 131
<< pdiffc >>
rect 47 546 81 580
rect 47 476 81 510
rect 47 406 81 440
rect 137 546 171 580
rect 137 463 171 497
rect 137 380 171 414
rect 227 542 261 576
rect 299 542 333 576
rect 389 544 423 578
rect 489 485 523 519
rect 589 544 623 578
rect 689 544 723 578
rect 789 544 823 578
rect 889 485 923 519
rect 979 546 1013 580
rect 979 474 1013 508
rect 1079 546 1113 580
rect 1079 474 1113 508
<< poly >>
rect 91 592 127 618
rect 181 592 217 618
rect 343 592 379 618
rect 440 592 476 618
rect 533 592 569 618
rect 633 592 669 618
rect 743 592 779 618
rect 843 592 879 618
rect 933 592 969 618
rect 1023 592 1059 618
rect 91 326 127 368
rect 21 318 127 326
rect 181 318 217 368
rect 343 336 379 368
rect 440 336 476 368
rect 533 336 569 368
rect 633 336 669 368
rect 743 336 779 368
rect 843 336 879 368
rect 933 336 969 368
rect 21 310 217 318
rect 21 276 37 310
rect 71 276 217 310
rect 21 260 217 276
rect 326 320 392 336
rect 326 286 342 320
rect 376 288 392 320
rect 446 320 570 336
rect 446 306 520 320
rect 376 286 398 288
rect 84 222 114 260
rect 170 222 200 260
rect 326 258 398 286
rect 368 233 398 258
rect 454 286 520 306
rect 554 286 570 320
rect 454 270 570 286
rect 615 320 681 336
rect 615 286 631 320
rect 665 286 681 320
rect 615 270 681 286
rect 729 320 795 336
rect 729 286 745 320
rect 779 286 795 320
rect 729 270 795 286
rect 843 320 969 336
rect 843 286 885 320
rect 919 286 969 320
rect 843 270 969 286
rect 1023 336 1059 368
rect 1023 320 1089 336
rect 1023 286 1039 320
rect 1073 286 1089 320
rect 1023 270 1089 286
rect 454 233 484 270
rect 540 233 570 270
rect 651 233 681 270
rect 737 233 767 270
rect 843 233 873 270
rect 939 233 969 270
rect 1037 233 1067 270
rect 84 48 114 74
rect 170 48 200 74
rect 368 59 398 85
rect 454 59 484 85
rect 540 59 570 85
rect 651 59 681 85
rect 737 59 767 85
rect 843 59 873 85
rect 939 59 969 85
rect 1037 59 1067 85
<< polycont >>
rect 37 276 71 310
rect 342 286 376 320
rect 520 286 554 320
rect 631 286 665 320
rect 745 286 779 320
rect 885 286 919 320
rect 1039 286 1073 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 31 580 81 649
rect 31 546 47 580
rect 31 510 81 546
rect 31 476 47 510
rect 31 440 81 476
rect 31 406 47 440
rect 31 390 81 406
rect 121 580 171 596
rect 121 546 137 580
rect 121 497 171 546
rect 211 576 339 649
rect 211 542 227 576
rect 261 542 299 576
rect 333 542 339 576
rect 211 526 339 542
rect 373 581 639 615
rect 373 578 439 581
rect 373 544 389 578
rect 423 544 439 578
rect 573 578 639 581
rect 373 526 439 544
rect 121 463 137 497
rect 473 519 539 547
rect 573 544 589 578
rect 623 544 639 578
rect 573 526 639 544
rect 673 578 739 649
rect 673 544 689 578
rect 723 544 739 578
rect 673 526 739 544
rect 773 581 1029 615
rect 773 578 839 581
rect 773 544 789 578
rect 823 544 839 578
rect 963 580 1029 581
rect 773 526 839 544
rect 473 492 489 519
rect 171 485 489 492
rect 523 492 539 519
rect 873 519 923 547
rect 873 492 889 519
rect 523 485 889 492
rect 171 463 923 485
rect 121 458 923 463
rect 963 546 979 580
rect 1013 546 1029 580
rect 963 508 1029 546
rect 963 474 979 508
rect 1013 474 1029 508
rect 963 458 1029 474
rect 1063 580 1129 649
rect 1063 546 1079 580
rect 1113 546 1129 580
rect 1063 508 1129 546
rect 1063 474 1079 508
rect 1113 474 1129 508
rect 1063 458 1129 474
rect 121 414 175 458
rect 121 380 137 414
rect 171 380 175 414
rect 21 310 87 356
rect 21 276 37 310
rect 71 276 87 310
rect 21 260 87 276
rect 23 210 73 226
rect 23 176 39 210
rect 23 120 73 176
rect 23 86 39 120
rect 121 189 175 380
rect 217 390 681 424
rect 217 320 455 390
rect 217 286 342 320
rect 376 286 455 320
rect 217 270 455 286
rect 504 320 570 356
rect 504 286 520 320
rect 554 286 570 320
rect 504 270 570 286
rect 615 320 681 390
rect 615 286 631 320
rect 665 286 681 320
rect 615 270 681 286
rect 729 390 1127 424
rect 729 320 795 390
rect 729 286 745 320
rect 779 286 795 320
rect 729 270 795 286
rect 869 320 935 356
rect 869 286 885 320
rect 919 286 935 320
rect 869 270 935 286
rect 985 320 1127 390
rect 985 286 1039 320
rect 1073 286 1127 320
rect 985 270 1127 286
rect 121 155 125 189
rect 159 155 175 189
rect 121 119 175 155
rect 211 221 656 236
rect 211 210 601 221
rect 245 202 601 210
rect 245 176 261 202
rect 211 120 261 176
rect 409 194 443 202
rect 23 85 73 86
rect 245 86 261 120
rect 211 85 261 86
rect 23 51 261 85
rect 307 148 373 164
rect 307 114 323 148
rect 357 114 373 148
rect 579 187 601 202
rect 635 187 656 221
rect 409 119 443 160
rect 479 148 545 164
rect 307 85 373 114
rect 479 114 495 148
rect 529 114 545 148
rect 579 153 656 187
rect 579 119 600 153
rect 634 119 656 153
rect 692 220 1129 236
rect 726 202 892 220
rect 726 186 742 202
rect 692 131 742 186
rect 876 186 892 202
rect 926 202 1078 220
rect 926 186 942 202
rect 479 85 545 114
rect 726 97 742 131
rect 692 85 742 97
rect 307 51 742 85
rect 776 148 842 164
rect 776 114 792 148
rect 826 114 842 148
rect 776 17 842 114
rect 876 131 942 186
rect 1112 186 1129 220
rect 876 97 892 131
rect 926 97 942 131
rect 876 81 942 97
rect 976 148 1042 164
rect 976 114 992 148
rect 1026 114 1042 148
rect 976 17 1042 114
rect 1078 131 1129 186
rect 1112 97 1129 131
rect 1078 81 1129 97
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
rlabel comment s 0 0 0 0 4 o221ai_2
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 127 168 161 202 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 127 242 161 276 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 127 390 161 424 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 127 464 161 498 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 127 538 161 572 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 C1
port 5 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 1152 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1172966
string GDS_START 1163076
<< end >>
