magic
tech sky130A
magscale 1 2
timestamp 1601050088
<< locali >>
rect 85 196 167 398
rect 313 290 381 356
rect 895 236 983 302
rect 1025 236 1127 302
rect 1341 236 1409 310
rect 3097 70 3165 430
rect 3287 395 3333 602
rect 3287 361 3433 395
rect 3340 226 3433 361
rect 3271 192 3433 226
rect 3271 70 3337 192
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3391 683
rect 3425 649 3456 683
rect 17 492 105 596
rect 213 526 263 649
rect 297 581 467 615
rect 297 492 331 581
rect 17 458 331 492
rect 17 146 51 458
rect 365 424 399 547
rect 433 492 467 581
rect 501 526 551 649
rect 653 492 709 594
rect 433 458 709 492
rect 201 390 527 424
rect 201 256 267 390
rect 461 303 527 390
rect 575 303 641 369
rect 675 269 709 458
rect 201 222 402 256
rect 17 84 116 146
rect 214 17 280 162
rect 336 109 402 222
rect 600 235 709 269
rect 743 581 973 615
rect 743 458 793 581
rect 436 17 502 201
rect 600 109 666 235
rect 743 201 777 458
rect 827 449 905 547
rect 939 485 973 581
rect 1007 519 1061 649
rect 1169 496 1261 585
rect 1297 530 1347 649
rect 1559 530 1625 649
rect 1761 530 1811 596
rect 1659 496 1811 530
rect 1845 506 1917 596
rect 2045 546 2111 649
rect 2264 546 2330 649
rect 1169 485 1693 496
rect 939 462 1693 485
rect 939 451 1295 462
rect 827 411 861 449
rect 700 109 777 201
rect 811 370 861 411
rect 1161 370 1227 417
rect 811 336 1227 370
rect 811 202 861 336
rect 1161 286 1227 336
rect 1261 252 1295 451
rect 1371 364 1531 428
rect 1164 218 1295 252
rect 1443 294 1531 364
rect 1581 330 1615 462
rect 1745 428 1811 461
rect 1649 364 1811 428
rect 1581 296 1743 330
rect 811 121 958 202
rect 811 73 861 121
rect 992 17 1058 202
rect 1164 121 1230 218
rect 1443 202 1477 294
rect 1283 17 1349 184
rect 1383 70 1477 202
rect 1511 17 1545 226
rect 1581 85 1647 226
rect 1693 119 1743 296
rect 1777 85 1811 364
rect 1845 372 1879 506
rect 1951 478 2544 512
rect 2578 504 2665 596
rect 2753 530 2861 649
rect 1951 472 1985 478
rect 1913 406 1985 472
rect 2152 410 2277 444
rect 1845 338 2188 372
rect 1845 119 1879 338
rect 2122 306 2188 338
rect 2243 304 2277 410
rect 2510 360 2544 478
rect 2631 377 2665 504
rect 2895 498 2967 596
rect 3007 532 3073 649
rect 3187 532 3253 649
rect 2895 476 3237 498
rect 2717 464 3237 476
rect 2717 411 3047 464
rect 2013 272 2079 304
rect 2243 272 2377 304
rect 1913 204 1971 269
rect 2013 238 2377 272
rect 2416 260 2476 360
rect 2510 294 2597 360
rect 2631 343 2773 377
rect 2895 360 3047 411
rect 2739 326 2773 343
rect 2639 260 2705 309
rect 1913 170 2172 204
rect 1913 85 1947 170
rect 1581 51 1947 85
rect 2054 17 2104 136
rect 2138 85 2172 170
rect 2206 119 2240 238
rect 2416 226 2705 260
rect 2739 260 2899 326
rect 2933 310 3047 360
rect 2416 204 2450 226
rect 2274 170 2450 204
rect 2739 188 2773 260
rect 2933 226 2967 310
rect 2274 85 2308 170
rect 2484 154 2773 188
rect 2138 51 2308 85
rect 2342 17 2392 136
rect 2484 70 2550 154
rect 2813 120 2867 224
rect 2664 17 2867 120
rect 2901 70 2967 226
rect 3013 17 3063 226
rect 3199 327 3237 464
rect 3367 429 3433 649
rect 3199 260 3302 327
rect 3201 17 3235 226
rect 3371 17 3423 158
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3456 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 3199 649 3233 683
rect 3295 649 3329 683
rect 3391 649 3425 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
<< metal1 >>
rect 0 683 3456 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3391 683
rect 3425 649 3456 683
rect 0 617 3456 649
rect 0 17 3456 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3456 17
rect 0 -49 3456 -17
<< obsm1 >>
rect 595 347 653 356
rect 2995 347 3053 356
rect 595 319 3053 347
rect 595 310 653 319
rect 2995 310 3053 319
<< labels >>
rlabel locali s 85 196 167 398 6 D
port 1 nsew signal input
rlabel locali s 313 290 381 356 6 DE
port 2 nsew signal input
rlabel locali s 3097 70 3165 430 6 Q
port 3 nsew signal output
rlabel locali s 3340 226 3433 361 6 Q_N
port 4 nsew signal output
rlabel locali s 3287 395 3333 602 6 Q_N
port 4 nsew signal output
rlabel locali s 3287 361 3433 395 6 Q_N
port 4 nsew signal output
rlabel locali s 3271 192 3433 226 6 Q_N
port 4 nsew signal output
rlabel locali s 3271 70 3337 192 6 Q_N
port 4 nsew signal output
rlabel locali s 1025 236 1127 302 6 SCD
port 5 nsew signal input
rlabel locali s 895 236 983 302 6 SCE
port 6 nsew signal input
rlabel locali s 1341 236 1409 310 6 CLK
port 7 nsew clock input
rlabel metal1 s 0 -49 3456 49 8 VGND
port 8 nsew ground bidirectional
rlabel metal1 s 0 617 3456 715 6 VPWR
port 9 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 3456 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 384728
string GDS_START 361276
<< end >>
