magic
tech sky130A
magscale 1 2
timestamp 1601050058
<< locali >>
rect 17 459 351 493
rect 17 425 29 459
rect 63 425 121 459
rect 155 425 213 459
rect 247 425 305 459
rect 339 425 351 459
rect 17 309 351 425
rect 201 205 351 309
<< viali >>
rect 29 425 63 459
rect 121 425 155 459
rect 213 425 247 459
rect 305 425 339 459
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 17 171 167 275
rect 17 17 351 171
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
<< metal1 >>
rect 0 561 368 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 0 496 368 527
rect 14 459 354 468
rect 14 428 29 459
rect 17 425 29 428
rect 63 425 121 459
rect 155 425 213 459
rect 247 425 305 459
rect 339 428 354 459
rect 339 425 351 428
rect 17 416 351 425
rect 0 17 368 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
rect 0 -48 368 -17
<< labels >>
rlabel viali s 305 425 339 459 6 KAPWR
port 1 nsew power bidirectional abutment
rlabel viali s 213 425 247 459 6 KAPWR
port 1 nsew power bidirectional abutment
rlabel viali s 121 425 155 459 6 KAPWR
port 1 nsew power bidirectional abutment
rlabel viali s 29 425 63 459 6 KAPWR
port 1 nsew power bidirectional abutment
rlabel locali s 201 205 351 309 6 KAPWR
port 1 nsew power bidirectional abutment
rlabel locali s 17 309 351 493 6 KAPWR
port 1 nsew power bidirectional abutment
rlabel metal1 s 17 416 351 428 6 KAPWR
port 1 nsew power bidirectional abutment
rlabel metal1 s 14 428 354 468 6 KAPWR
port 1 nsew power bidirectional abutment
rlabel metal1 s 0 -48 368 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 496 368 592 6 VPWR
port 3 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 368 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2284204
string GDS_START 2280944
<< end >>
