magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 276 561
rect 17 312 71 493
rect 105 375 171 527
rect 17 152 51 312
rect 189 197 255 271
rect 17 51 69 152
rect 105 17 171 93
rect 0 -17 276 17
<< obsli1 >>
rect 207 341 241 493
rect 108 307 241 341
rect 108 278 142 307
rect 85 212 142 278
rect 108 161 142 212
rect 108 127 241 161
rect 207 51 241 127
<< metal1 >>
rect 0 496 276 592
rect 0 -48 276 48
<< labels >>
rlabel locali s 189 197 255 271 6 A
port 1 nsew signal input
rlabel locali s 17 312 71 493 6 X
port 2 nsew signal output
rlabel locali s 17 152 51 312 6 X
port 2 nsew signal output
rlabel locali s 17 51 69 152 6 X
port 2 nsew signal output
rlabel locali s 105 17 171 93 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 0 -17 276 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 276 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 105 375 171 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 0 527 276 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 496 276 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 276 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3116952
string GDS_START 3113202
<< end >>
