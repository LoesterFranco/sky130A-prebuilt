magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 710 704
<< pwell >>
rect 0 0 672 49
<< scnmos >>
rect 152 74 182 222
rect 230 74 260 222
rect 338 74 368 222
rect 440 74 470 222
rect 558 74 588 222
<< pmoshvt >>
rect 149 368 179 592
rect 239 368 269 592
rect 365 368 395 592
rect 460 368 490 592
rect 551 368 581 592
<< ndiff >>
rect 27 202 152 222
rect 27 168 39 202
rect 73 168 107 202
rect 141 168 152 202
rect 27 120 152 168
rect 27 86 39 120
rect 73 86 107 120
rect 141 86 152 120
rect 27 74 152 86
rect 182 74 230 222
rect 260 74 338 222
rect 368 202 440 222
rect 368 168 381 202
rect 415 168 440 202
rect 368 120 440 168
rect 368 86 381 120
rect 415 86 440 120
rect 368 74 440 86
rect 470 120 558 222
rect 470 86 490 120
rect 524 86 558 120
rect 470 74 558 86
rect 588 202 645 222
rect 588 168 599 202
rect 633 168 645 202
rect 588 120 645 168
rect 588 86 599 120
rect 633 86 645 120
rect 588 74 645 86
<< pdiff >>
rect 80 582 149 592
rect 80 548 92 582
rect 126 548 149 582
rect 80 514 149 548
rect 80 480 92 514
rect 126 480 149 514
rect 80 446 149 480
rect 80 412 92 446
rect 126 412 149 446
rect 80 368 149 412
rect 179 580 239 592
rect 179 546 192 580
rect 226 546 239 580
rect 179 497 239 546
rect 179 463 192 497
rect 226 463 239 497
rect 179 414 239 463
rect 179 380 192 414
rect 226 380 239 414
rect 179 368 239 380
rect 269 582 365 592
rect 269 548 313 582
rect 347 548 365 582
rect 269 514 365 548
rect 269 480 313 514
rect 347 480 365 514
rect 269 446 365 480
rect 269 412 313 446
rect 347 412 365 446
rect 269 368 365 412
rect 395 580 460 592
rect 395 546 413 580
rect 447 546 460 580
rect 395 497 460 546
rect 395 463 413 497
rect 447 463 460 497
rect 395 414 460 463
rect 395 380 413 414
rect 447 380 460 414
rect 395 368 460 380
rect 490 368 551 592
rect 581 580 640 592
rect 581 546 594 580
rect 628 546 640 580
rect 581 497 640 546
rect 581 463 594 497
rect 628 463 640 497
rect 581 414 640 463
rect 581 380 594 414
rect 628 380 640 414
rect 581 368 640 380
<< ndiffc >>
rect 39 168 73 202
rect 107 168 141 202
rect 39 86 73 120
rect 107 86 141 120
rect 381 168 415 202
rect 381 86 415 120
rect 490 86 524 120
rect 599 168 633 202
rect 599 86 633 120
<< pdiffc >>
rect 92 548 126 582
rect 92 480 126 514
rect 92 412 126 446
rect 192 546 226 580
rect 192 463 226 497
rect 192 380 226 414
rect 313 548 347 582
rect 313 480 347 514
rect 313 412 347 446
rect 413 546 447 580
rect 413 463 447 497
rect 413 380 447 414
rect 594 546 628 580
rect 594 463 628 497
rect 594 380 628 414
<< poly >>
rect 149 592 179 618
rect 239 592 269 618
rect 365 592 395 618
rect 460 592 490 618
rect 551 592 581 618
rect 149 353 179 368
rect 239 353 269 368
rect 365 353 395 368
rect 460 353 490 368
rect 551 353 581 368
rect 146 310 182 353
rect 236 310 272 353
rect 362 310 398 353
rect 457 310 493 353
rect 548 310 584 353
rect 116 294 182 310
rect 116 260 132 294
rect 166 260 182 294
rect 116 244 182 260
rect 224 294 290 310
rect 224 260 240 294
rect 274 260 290 294
rect 224 244 290 260
rect 332 294 398 310
rect 332 260 348 294
rect 382 260 398 294
rect 332 244 398 260
rect 440 294 506 310
rect 440 260 456 294
rect 490 260 506 294
rect 440 244 506 260
rect 548 294 651 310
rect 548 260 601 294
rect 635 260 651 294
rect 548 244 651 260
rect 152 222 182 244
rect 230 222 260 244
rect 338 222 368 244
rect 440 222 470 244
rect 558 222 588 244
rect 152 48 182 74
rect 230 48 260 74
rect 338 48 368 74
rect 440 48 470 74
rect 558 48 588 74
<< polycont >>
rect 132 260 166 294
rect 240 260 274 294
rect 348 260 382 294
rect 456 260 490 294
rect 601 260 635 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 76 582 142 649
rect 76 548 92 582
rect 126 548 142 582
rect 76 514 142 548
rect 76 480 92 514
rect 126 480 142 514
rect 76 446 142 480
rect 76 412 92 446
rect 126 412 142 446
rect 176 580 263 596
rect 176 546 192 580
rect 226 546 263 580
rect 176 497 263 546
rect 176 463 192 497
rect 226 463 263 497
rect 176 414 263 463
rect 176 380 192 414
rect 226 380 263 414
rect 297 582 363 649
rect 297 548 313 582
rect 347 548 363 582
rect 297 514 363 548
rect 297 480 313 514
rect 347 480 363 514
rect 297 446 363 480
rect 297 412 313 446
rect 347 412 363 446
rect 397 580 463 596
rect 397 546 413 580
rect 447 546 463 580
rect 397 497 463 546
rect 397 463 413 497
rect 447 463 463 497
rect 397 414 463 463
rect 176 378 263 380
rect 397 380 413 414
rect 447 380 463 414
rect 397 378 463 380
rect 23 344 463 378
rect 578 580 644 649
rect 578 546 594 580
rect 628 546 644 580
rect 578 497 644 546
rect 578 463 594 497
rect 628 463 644 497
rect 578 414 644 463
rect 578 380 594 414
rect 628 380 644 414
rect 578 364 644 380
rect 23 202 57 344
rect 116 294 182 310
rect 116 260 132 294
rect 166 260 182 294
rect 116 236 182 260
rect 217 294 285 310
rect 217 260 240 294
rect 274 260 285 294
rect 23 168 39 202
rect 73 168 107 202
rect 141 168 157 202
rect 23 120 157 168
rect 23 86 39 120
rect 73 86 107 120
rect 141 86 157 120
rect 217 88 285 260
rect 319 294 398 310
rect 319 260 348 294
rect 382 260 398 294
rect 319 236 398 260
rect 440 294 551 310
rect 440 260 456 294
rect 490 260 551 294
rect 440 236 551 260
rect 585 294 651 310
rect 585 260 601 294
rect 635 260 651 294
rect 585 236 651 260
rect 365 168 381 202
rect 415 168 599 202
rect 633 168 649 202
rect 365 120 431 168
rect 583 120 649 168
rect 23 70 157 86
rect 365 86 381 120
rect 415 86 431 120
rect 365 70 431 86
rect 465 86 490 120
rect 524 86 549 120
rect 465 17 549 86
rect 583 86 599 120
rect 633 86 649 120
rect 583 70 649 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o2111ai_1
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 223 390 257 424 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 223 464 257 498 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 223 538 257 572 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 127 242 161 276 0 FreeSans 340 0 0 0 D1
port 5 nsew
flabel corelocali s 223 94 257 128 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 223 168 257 202 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 223 242 257 276 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 319 242 353 276 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 511 242 545 276 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 607 242 641 276 0 FreeSans 340 0 0 0 A1
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 672 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1336918
string GDS_START 1330058
<< end >>
