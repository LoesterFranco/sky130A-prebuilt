magic
tech sky130A
magscale 1 2
timestamp 1599588218
<< nwell >>
rect -38 332 1094 704
<< pwell >>
rect 0 0 1056 49
<< scpmos >>
rect 102 392 138 560
rect 216 392 252 592
rect 360 392 396 592
rect 492 392 528 592
rect 582 392 618 592
rect 737 368 773 592
rect 827 368 863 592
rect 934 368 970 536
<< nmoslvt >>
rect 84 74 114 184
rect 282 82 312 230
rect 360 82 390 230
rect 468 82 498 230
rect 570 82 600 230
rect 738 82 768 230
rect 824 82 854 230
rect 942 120 972 230
<< ndiff >>
rect 225 218 282 230
rect 225 184 237 218
rect 271 184 282 218
rect 27 146 84 184
rect 27 112 39 146
rect 73 112 84 146
rect 27 74 84 112
rect 114 146 171 184
rect 114 112 125 146
rect 159 112 171 146
rect 114 74 171 112
rect 225 128 282 184
rect 225 94 237 128
rect 271 94 282 128
rect 225 82 282 94
rect 312 82 360 230
rect 390 82 468 230
rect 498 82 570 230
rect 600 150 738 230
rect 600 116 611 150
rect 645 116 738 150
rect 600 82 738 116
rect 768 218 824 230
rect 768 184 779 218
rect 813 184 824 218
rect 768 82 824 184
rect 854 120 942 230
rect 972 176 1029 230
rect 972 142 983 176
rect 1017 142 1029 176
rect 972 120 1029 142
rect 854 82 927 120
rect 869 48 881 82
rect 915 48 927 82
rect 869 36 927 48
<< pdiff >>
rect 160 580 216 592
rect 160 560 172 580
rect 46 548 102 560
rect 46 514 58 548
rect 92 514 102 548
rect 46 440 102 514
rect 46 406 58 440
rect 92 406 102 440
rect 46 392 102 406
rect 138 546 172 560
rect 206 546 216 580
rect 138 492 216 546
rect 138 458 172 492
rect 206 458 216 492
rect 138 392 216 458
rect 252 580 360 592
rect 252 546 302 580
rect 336 546 360 580
rect 252 509 360 546
rect 252 475 302 509
rect 336 475 360 509
rect 252 438 360 475
rect 252 404 302 438
rect 336 404 360 438
rect 252 392 360 404
rect 396 580 492 592
rect 396 546 429 580
rect 463 546 492 580
rect 396 499 492 546
rect 396 465 429 499
rect 463 465 492 499
rect 396 392 492 465
rect 528 580 582 592
rect 528 546 538 580
rect 572 546 582 580
rect 528 510 582 546
rect 528 476 538 510
rect 572 476 582 510
rect 528 440 582 476
rect 528 406 538 440
rect 572 406 582 440
rect 528 392 582 406
rect 618 584 737 592
rect 618 550 656 584
rect 690 550 737 584
rect 618 498 737 550
rect 618 464 656 498
rect 690 464 737 498
rect 618 392 737 464
rect 687 368 737 392
rect 773 580 827 592
rect 773 546 783 580
rect 817 546 827 580
rect 773 499 827 546
rect 773 465 783 499
rect 817 465 827 499
rect 773 418 827 465
rect 773 384 783 418
rect 817 384 827 418
rect 773 368 827 384
rect 863 580 919 592
rect 863 546 873 580
rect 907 546 919 580
rect 863 536 919 546
rect 863 470 934 536
rect 863 436 873 470
rect 907 436 934 470
rect 863 368 934 436
rect 970 524 1029 536
rect 970 490 981 524
rect 1015 490 1029 524
rect 970 414 1029 490
rect 970 380 981 414
rect 1015 380 1029 414
rect 970 368 1029 380
<< ndiffc >>
rect 237 184 271 218
rect 39 112 73 146
rect 125 112 159 146
rect 237 94 271 128
rect 611 116 645 150
rect 779 184 813 218
rect 983 142 1017 176
rect 881 48 915 82
<< pdiffc >>
rect 58 514 92 548
rect 58 406 92 440
rect 172 546 206 580
rect 172 458 206 492
rect 302 546 336 580
rect 302 475 336 509
rect 302 404 336 438
rect 429 546 463 580
rect 429 465 463 499
rect 538 546 572 580
rect 538 476 572 510
rect 538 406 572 440
rect 656 550 690 584
rect 656 464 690 498
rect 783 546 817 580
rect 783 465 817 499
rect 783 384 817 418
rect 873 546 907 580
rect 873 436 907 470
rect 981 490 1015 524
rect 981 380 1015 414
<< poly >>
rect 216 592 252 618
rect 360 592 396 618
rect 492 592 528 618
rect 582 592 618 618
rect 737 592 773 618
rect 827 592 863 618
rect 102 560 138 586
rect 102 356 138 392
rect 44 340 132 356
rect 44 306 60 340
rect 94 306 132 340
rect 216 334 252 392
rect 44 290 132 306
rect 186 318 252 334
rect 360 318 396 392
rect 492 350 528 392
rect 582 350 618 392
rect 934 536 970 562
rect 462 334 528 350
rect 84 184 114 290
rect 186 284 202 318
rect 236 298 252 318
rect 354 302 420 318
rect 236 284 312 298
rect 186 268 312 284
rect 282 230 312 268
rect 354 268 370 302
rect 404 268 420 302
rect 462 300 478 334
rect 512 300 528 334
rect 462 284 528 300
rect 570 334 651 350
rect 737 334 773 368
rect 827 334 863 368
rect 570 300 601 334
rect 635 300 651 334
rect 570 284 651 300
rect 705 318 863 334
rect 705 284 721 318
rect 755 284 863 318
rect 354 252 420 268
rect 360 230 390 252
rect 468 230 498 284
rect 570 230 600 284
rect 705 268 863 284
rect 934 318 970 368
rect 934 302 1031 318
rect 934 268 981 302
rect 1015 268 1031 302
rect 738 230 768 268
rect 824 230 854 268
rect 934 252 1031 268
rect 942 230 972 252
rect 942 94 972 120
rect 84 48 114 74
rect 282 56 312 82
rect 360 56 390 82
rect 468 56 498 82
rect 570 56 600 82
rect 738 56 768 82
rect 824 56 854 82
<< polycont >>
rect 60 306 94 340
rect 202 284 236 318
rect 370 268 404 302
rect 478 300 512 334
rect 601 300 635 334
rect 721 284 755 318
rect 981 268 1015 302
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 156 580 222 649
rect 42 548 108 564
rect 42 514 58 548
rect 92 514 108 548
rect 42 440 108 514
rect 156 546 172 580
rect 206 546 222 580
rect 156 492 222 546
rect 156 458 172 492
rect 206 458 222 492
rect 286 580 352 596
rect 286 546 302 580
rect 336 546 352 580
rect 286 509 352 546
rect 286 475 302 509
rect 336 475 352 509
rect 42 406 58 440
rect 92 424 108 440
rect 286 438 352 475
rect 413 580 479 649
rect 413 546 429 580
rect 463 546 479 580
rect 413 499 479 546
rect 413 465 429 499
rect 463 465 479 499
rect 413 458 479 465
rect 522 580 588 596
rect 522 546 538 580
rect 572 546 588 580
rect 522 510 588 546
rect 522 476 538 510
rect 572 476 588 510
rect 92 406 187 424
rect 42 390 187 406
rect 25 340 110 356
rect 25 306 60 340
rect 94 306 110 340
rect 25 290 110 306
rect 153 334 187 390
rect 286 404 302 438
rect 336 424 352 438
rect 522 440 588 476
rect 640 584 706 649
rect 640 550 656 584
rect 690 550 706 584
rect 640 498 706 550
rect 640 464 656 498
rect 690 464 706 498
rect 640 458 706 464
rect 767 580 839 596
rect 767 546 783 580
rect 817 546 839 580
rect 767 499 839 546
rect 767 465 783 499
rect 817 465 839 499
rect 522 424 538 440
rect 336 406 538 424
rect 572 424 588 440
rect 572 406 733 424
rect 336 404 733 406
rect 286 390 733 404
rect 286 388 352 390
rect 153 318 252 334
rect 153 284 202 318
rect 236 284 252 318
rect 153 268 252 284
rect 153 256 187 268
rect 23 222 187 256
rect 286 234 320 388
rect 462 334 551 356
rect 23 146 73 222
rect 221 218 320 234
rect 23 112 39 146
rect 23 70 73 112
rect 109 146 175 188
rect 109 112 125 146
rect 159 112 175 146
rect 109 17 175 112
rect 221 184 237 218
rect 271 184 320 218
rect 354 302 420 318
rect 354 268 370 302
rect 404 268 420 302
rect 462 300 478 334
rect 512 300 551 334
rect 462 284 551 300
rect 585 334 651 356
rect 585 300 601 334
rect 635 300 651 334
rect 585 284 651 300
rect 699 334 733 390
rect 767 418 839 465
rect 873 580 923 649
rect 907 546 923 580
rect 873 470 923 546
rect 907 436 923 470
rect 873 420 923 436
rect 964 524 1033 540
rect 964 490 981 524
rect 1015 490 1033 524
rect 767 384 783 418
rect 817 384 839 418
rect 964 414 1033 490
rect 964 386 981 414
rect 767 368 839 384
rect 699 318 771 334
rect 699 284 721 318
rect 755 284 771 318
rect 699 268 771 284
rect 354 234 420 268
rect 805 234 839 368
rect 354 200 729 234
rect 221 128 320 184
rect 221 94 237 128
rect 271 94 320 128
rect 221 78 320 94
rect 595 150 661 166
rect 595 116 611 150
rect 645 116 661 150
rect 695 150 729 200
rect 763 218 839 234
rect 763 184 779 218
rect 813 184 839 218
rect 873 380 981 386
rect 1015 380 1033 414
rect 873 352 1033 380
rect 873 150 907 352
rect 965 302 1031 318
rect 965 268 981 302
rect 1015 268 1031 302
rect 965 236 1031 268
rect 967 176 1033 202
rect 967 150 983 176
rect 695 142 983 150
rect 1017 142 1033 176
rect 695 116 1033 142
rect 595 17 661 116
rect 865 48 881 82
rect 915 48 931 82
rect 865 17 931 48
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 683 1056 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 0 617 1056 649
rect 0 17 1056 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -49 1056 -17
<< labels >>
flabel pwell s 0 0 1056 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nwell s 0 617 1056 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
rlabel comment s 0 0 0 0 4 and4bb_2
flabel metal1 s 0 617 1056 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 1056 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 799 390 833 424 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 799 464 833 498 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 799 538 833 572 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 991 242 1025 276 0 FreeSans 340 0 0 0 B_N
port 2 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 D
port 4 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 C
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 1056 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3240880
string GDS_START 3232492
<< end >>
