magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 103 93 133 177
rect 221 47 251 177
rect 304 47 334 177
rect 401 47 431 177
rect 497 47 527 177
<< pmoshvt >>
rect 106 297 142 381
rect 213 297 249 497
rect 307 297 343 497
rect 403 297 439 497
rect 499 297 535 497
<< ndiff >>
rect 40 139 103 177
rect 40 105 48 139
rect 82 105 103 139
rect 40 93 103 105
rect 133 93 221 177
rect 148 59 156 93
rect 190 59 221 93
rect 148 47 221 59
rect 251 47 304 177
rect 334 47 401 177
rect 431 47 497 177
rect 527 166 617 177
rect 527 132 571 166
rect 605 132 617 166
rect 527 98 617 132
rect 527 64 571 98
rect 605 64 617 98
rect 527 47 617 64
<< pdiff >>
rect 159 485 213 497
rect 159 451 167 485
rect 201 451 213 485
rect 159 417 213 451
rect 159 383 167 417
rect 201 383 213 417
rect 159 381 213 383
rect 52 369 106 381
rect 52 335 60 369
rect 94 335 106 369
rect 52 297 106 335
rect 142 349 213 381
rect 142 315 167 349
rect 201 315 213 349
rect 142 297 213 315
rect 249 485 307 497
rect 249 451 261 485
rect 295 451 307 485
rect 249 417 307 451
rect 249 383 261 417
rect 295 383 307 417
rect 249 349 307 383
rect 249 315 261 349
rect 295 315 307 349
rect 249 297 307 315
rect 343 485 403 497
rect 343 451 355 485
rect 389 451 403 485
rect 343 417 403 451
rect 343 383 355 417
rect 389 383 403 417
rect 343 297 403 383
rect 439 484 499 497
rect 439 450 451 484
rect 485 450 499 484
rect 439 416 499 450
rect 439 382 451 416
rect 485 382 499 416
rect 439 348 499 382
rect 439 314 451 348
rect 485 314 499 348
rect 439 297 499 314
rect 535 485 617 497
rect 535 451 575 485
rect 609 451 617 485
rect 535 417 617 451
rect 535 383 575 417
rect 609 383 617 417
rect 535 297 617 383
<< ndiffc >>
rect 48 105 82 139
rect 156 59 190 93
rect 571 132 605 166
rect 571 64 605 98
<< pdiffc >>
rect 167 451 201 485
rect 167 383 201 417
rect 60 335 94 369
rect 167 315 201 349
rect 261 451 295 485
rect 261 383 295 417
rect 261 315 295 349
rect 355 451 389 485
rect 355 383 389 417
rect 451 450 485 484
rect 451 382 485 416
rect 451 314 485 348
rect 575 451 609 485
rect 575 383 609 417
<< poly >>
rect 213 497 249 523
rect 307 497 343 523
rect 403 497 439 523
rect 499 497 535 523
rect 106 381 142 407
rect 106 282 142 297
rect 213 282 249 297
rect 307 282 343 297
rect 403 282 439 297
rect 499 282 535 297
rect 104 265 144 282
rect 211 265 251 282
rect 305 265 345 282
rect 401 265 441 282
rect 497 265 537 282
rect 68 249 144 265
rect 68 215 85 249
rect 119 215 144 249
rect 68 199 144 215
rect 186 249 262 265
rect 186 215 202 249
rect 236 215 262 249
rect 186 199 262 215
rect 304 249 358 265
rect 304 215 314 249
rect 348 215 358 249
rect 304 199 358 215
rect 401 249 455 265
rect 401 215 411 249
rect 445 215 455 249
rect 401 199 455 215
rect 497 249 551 265
rect 497 215 507 249
rect 541 215 551 249
rect 497 199 551 215
rect 103 177 133 199
rect 221 177 251 199
rect 304 177 334 199
rect 401 177 431 199
rect 497 177 527 199
rect 103 67 133 93
rect 221 21 251 47
rect 304 21 334 47
rect 401 21 431 47
rect 497 21 527 47
<< polycont >>
rect 85 215 119 249
rect 202 215 236 249
rect 314 215 348 249
rect 411 215 445 249
rect 507 215 541 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 151 485 201 527
rect 151 451 167 485
rect 151 417 201 451
rect 17 369 101 385
rect 17 335 60 369
rect 94 335 101 369
rect 17 319 101 335
rect 151 383 167 417
rect 151 349 201 383
rect 17 165 51 319
rect 151 315 167 349
rect 151 299 201 315
rect 235 485 311 493
rect 235 451 261 485
rect 295 451 311 485
rect 235 417 311 451
rect 235 383 261 417
rect 295 383 311 417
rect 235 349 311 383
rect 345 485 400 527
rect 345 451 355 485
rect 389 451 400 485
rect 345 417 400 451
rect 345 383 355 417
rect 389 383 400 417
rect 345 367 400 383
rect 435 484 501 493
rect 435 450 451 484
rect 485 450 501 484
rect 435 416 501 450
rect 435 382 451 416
rect 485 382 501 416
rect 235 315 261 349
rect 295 333 311 349
rect 435 348 501 382
rect 575 485 618 527
rect 609 451 618 485
rect 575 417 618 451
rect 609 383 618 417
rect 575 367 618 383
rect 435 333 451 348
rect 295 315 451 333
rect 235 314 451 315
rect 485 333 501 348
rect 485 314 627 333
rect 235 299 627 314
rect 85 249 164 265
rect 119 215 164 249
rect 85 199 164 215
rect 202 249 266 265
rect 236 215 266 249
rect 202 199 266 215
rect 300 249 352 265
rect 300 215 314 249
rect 348 215 352 249
rect 300 192 352 215
rect 17 139 274 165
rect 308 153 352 192
rect 386 249 445 265
rect 386 215 411 249
rect 386 153 445 215
rect 479 249 541 265
rect 479 215 507 249
rect 479 199 541 215
rect 17 105 48 139
rect 82 131 274 139
rect 82 105 94 131
rect 17 89 94 105
rect 240 119 274 131
rect 479 119 520 199
rect 575 167 627 299
rect 133 93 206 97
rect 133 59 156 93
rect 190 59 206 93
rect 240 85 520 119
rect 555 166 627 167
rect 555 132 571 166
rect 605 132 627 166
rect 555 98 627 132
rect 133 17 206 59
rect 555 64 571 98
rect 605 64 627 98
rect 555 51 627 64
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel corelocali s 581 85 615 119 0 FreeSans 250 0 0 0 Y
port 9 nsew
flabel corelocali s 305 221 339 255 0 FreeSans 250 0 0 0 C
port 3 nsew
flabel corelocali s 213 221 247 255 0 FreeSans 250 0 0 0 D
port 4 nsew
flabel corelocali s 121 221 155 255 0 FreeSans 250 0 0 0 A_N
port 1 nsew
flabel corelocali s 397 221 431 255 0 FreeSans 250 0 0 0 B
port 2 nsew
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
rlabel comment s 0 0 0 0 4 nand4b_1
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2321804
string GDS_START 2315926
<< end >>
