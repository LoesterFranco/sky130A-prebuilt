magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 89 47 119 177
rect 173 47 203 177
rect 279 47 309 177
<< pmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 281 297 317 497
<< ndiff >>
rect 27 99 89 177
rect 27 65 35 99
rect 69 65 89 99
rect 27 47 89 65
rect 119 47 173 177
rect 203 47 279 177
rect 309 161 371 177
rect 309 127 329 161
rect 363 127 371 161
rect 309 93 371 127
rect 309 59 329 93
rect 363 59 371 93
rect 309 47 371 59
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 485 175 497
rect 117 451 129 485
rect 163 451 175 485
rect 117 417 175 451
rect 117 383 129 417
rect 163 383 175 417
rect 117 349 175 383
rect 117 315 129 349
rect 163 315 175 349
rect 117 297 175 315
rect 211 485 281 497
rect 211 451 223 485
rect 257 451 281 485
rect 211 417 281 451
rect 211 383 223 417
rect 257 383 281 417
rect 211 297 281 383
rect 317 485 371 497
rect 317 451 329 485
rect 363 451 371 485
rect 317 417 371 451
rect 317 383 329 417
rect 363 383 371 417
rect 317 349 371 383
rect 317 315 329 349
rect 363 315 371 349
rect 317 297 371 315
<< ndiffc >>
rect 35 65 69 99
rect 329 127 363 161
rect 329 59 363 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 451 163 485
rect 129 383 163 417
rect 129 315 163 349
rect 223 451 257 485
rect 223 383 257 417
rect 329 451 363 485
rect 329 383 363 417
rect 329 315 363 349
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 281 497 317 523
rect 81 282 117 297
rect 175 282 211 297
rect 281 282 317 297
rect 79 265 119 282
rect 22 249 119 265
rect 22 215 32 249
rect 66 215 119 249
rect 22 199 119 215
rect 89 177 119 199
rect 173 265 213 282
rect 279 265 319 282
rect 173 249 237 265
rect 173 215 183 249
rect 217 215 237 249
rect 173 199 237 215
rect 279 249 368 265
rect 279 215 324 249
rect 358 215 368 249
rect 279 199 368 215
rect 173 177 203 199
rect 279 177 309 199
rect 89 21 119 47
rect 173 21 203 47
rect 279 21 309 47
<< polycont >>
rect 32 215 66 249
rect 183 215 217 249
rect 324 215 358 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 18 485 69 527
rect 18 451 35 485
rect 18 417 69 451
rect 18 383 35 417
rect 18 349 69 383
rect 18 315 35 349
rect 18 299 69 315
rect 103 485 179 493
rect 103 451 129 485
rect 163 451 179 485
rect 103 417 179 451
rect 103 383 129 417
rect 163 383 179 417
rect 103 349 179 383
rect 223 485 269 527
rect 257 451 269 485
rect 223 417 269 451
rect 257 383 269 417
rect 223 367 269 383
rect 303 485 379 493
rect 303 451 329 485
rect 363 451 379 485
rect 303 417 379 451
rect 303 383 329 417
rect 363 383 379 417
rect 103 315 129 349
rect 163 333 179 349
rect 303 349 379 383
rect 303 333 329 349
rect 163 315 329 333
rect 363 315 379 349
rect 103 299 379 315
rect 22 249 66 265
rect 22 215 32 249
rect 22 149 66 215
rect 103 119 149 299
rect 183 249 257 265
rect 217 215 257 249
rect 183 153 257 215
rect 295 249 381 265
rect 295 215 324 249
rect 358 215 381 249
rect 295 199 381 215
rect 303 161 379 165
rect 303 127 329 161
rect 363 127 379 161
rect 303 119 379 127
rect 18 99 69 115
rect 18 65 35 99
rect 18 17 69 65
rect 103 93 379 119
rect 103 59 329 93
rect 363 59 379 93
rect 103 51 379 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
flabel corelocali s 118 85 152 119 0 FreeSans 250 0 0 0 Y
port 8 nsew
flabel corelocali s 308 221 342 255 0 FreeSans 250 0 0 0 A
port 1 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 250 0 0 0 C
port 3 nsew
flabel corelocali s 215 221 249 255 0 FreeSans 250 0 0 0 B
port 2 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
rlabel comment s 0 0 0 0 4 nand3_1
<< properties >>
string FIXED_BBOX 0 0 460 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2242692
string GDS_START 2238094
<< end >>
