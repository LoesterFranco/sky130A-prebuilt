magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 644 561
rect 142 299 192 527
rect 226 333 292 493
rect 326 367 383 527
rect 417 333 483 493
rect 541 367 584 527
rect 226 299 627 333
rect 85 199 155 265
rect 193 199 247 265
rect 301 153 351 265
rect 385 153 437 265
rect 585 165 627 299
rect 131 17 197 97
rect 539 51 627 165
rect 0 -17 644 17
<< obsli1 >>
rect 17 319 102 385
rect 17 165 51 319
rect 17 131 267 165
rect 471 199 551 265
rect 17 89 95 131
rect 231 119 267 131
rect 471 119 505 199
rect 231 85 505 119
<< metal1 >>
rect 0 496 644 592
rect 0 -48 644 48
<< labels >>
rlabel locali s 85 199 155 265 6 A_N
port 1 nsew signal input
rlabel locali s 385 153 437 265 6 B
port 2 nsew signal input
rlabel locali s 301 153 351 265 6 C
port 3 nsew signal input
rlabel locali s 193 199 247 265 6 D
port 4 nsew signal input
rlabel locali s 585 165 627 299 6 Y
port 5 nsew signal output
rlabel locali s 539 51 627 165 6 Y
port 5 nsew signal output
rlabel locali s 417 333 483 493 6 Y
port 5 nsew signal output
rlabel locali s 226 333 292 493 6 Y
port 5 nsew signal output
rlabel locali s 226 299 627 333 6 Y
port 5 nsew signal output
rlabel locali s 131 17 197 97 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 644 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 644 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 541 367 584 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 326 367 383 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 142 299 192 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 644 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 644 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1869494
string GDS_START 1863680
<< end >>
