magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 552 561
rect 17 425 256 483
rect 290 367 346 527
rect 121 265 166 323
rect 388 299 443 493
rect 17 199 87 265
rect 121 199 286 265
rect 409 152 443 299
rect 477 286 535 527
rect 106 17 172 97
rect 274 17 350 97
rect 388 83 443 152
rect 477 17 535 183
rect 0 -17 552 17
<< obsli1 >>
rect 21 357 254 391
rect 21 299 87 357
rect 220 333 254 357
rect 220 299 354 333
rect 320 265 354 299
rect 320 199 375 265
rect 320 165 354 199
rect 21 131 354 165
rect 21 61 72 131
rect 206 61 240 131
<< metal1 >>
rect 0 496 552 592
rect 0 -48 552 48
<< labels >>
rlabel locali s 121 265 166 323 6 A
port 1 nsew signal input
rlabel locali s 121 199 286 265 6 A
port 1 nsew signal input
rlabel locali s 17 425 256 483 6 B
port 2 nsew signal input
rlabel locali s 17 199 87 265 6 C
port 3 nsew signal input
rlabel locali s 409 152 443 299 6 X
port 4 nsew signal output
rlabel locali s 388 299 443 493 6 X
port 4 nsew signal output
rlabel locali s 388 83 443 152 6 X
port 4 nsew signal output
rlabel locali s 477 17 535 183 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 274 17 350 97 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 106 17 172 97 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 552 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 552 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 477 286 535 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 290 367 346 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 552 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 552 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 552 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1037274
string GDS_START 1031660
<< end >>
