magic
tech sky130A
magscale 1 2
timestamp 1604502705
<< nwell >>
rect -38 332 806 704
<< pwell >>
rect 0 0 768 49
<< scnmos >>
rect 79 47 689 202
<< scpmos >>
rect 79 368 689 619
<< ndiff >>
rect 27 190 79 202
rect 27 156 35 190
rect 69 156 79 190
rect 27 93 79 156
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 689 190 741 202
rect 689 156 699 190
rect 733 156 741 190
rect 689 93 741 156
rect 689 59 699 93
rect 733 59 741 93
rect 689 47 741 59
<< pdiff >>
rect 27 607 79 619
rect 27 573 35 607
rect 69 573 79 607
rect 27 510 79 573
rect 27 476 35 510
rect 69 476 79 510
rect 27 414 79 476
rect 27 380 35 414
rect 69 380 79 414
rect 27 368 79 380
rect 689 607 741 619
rect 689 573 699 607
rect 733 573 741 607
rect 689 510 741 573
rect 689 476 699 510
rect 733 476 741 510
rect 689 414 741 476
rect 689 380 699 414
rect 733 380 741 414
rect 689 368 741 380
<< ndiffc >>
rect 35 156 69 190
rect 35 59 69 93
rect 699 156 733 190
rect 699 59 733 93
<< pdiffc >>
rect 35 573 69 607
rect 35 476 69 510
rect 35 380 69 414
rect 699 573 733 607
rect 699 476 733 510
rect 699 380 733 414
<< poly >>
rect 79 619 689 645
rect 79 342 689 368
rect 52 320 186 342
rect 52 286 68 320
rect 102 286 136 320
rect 170 286 186 320
rect 404 320 538 342
rect 52 270 186 286
rect 228 284 362 300
rect 228 250 244 284
rect 278 250 312 284
rect 346 250 362 284
rect 404 286 420 320
rect 454 286 488 320
rect 522 286 538 320
rect 404 270 538 286
rect 580 284 714 300
rect 228 228 362 250
rect 580 250 596 284
rect 630 250 664 284
rect 698 250 714 284
rect 580 228 714 250
rect 79 202 689 228
rect 79 21 689 47
<< polycont >>
rect 68 286 102 320
rect 136 286 170 320
rect 244 250 278 284
rect 312 250 346 284
rect 420 286 454 320
rect 488 286 522 320
rect 596 250 630 284
rect 664 250 698 284
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 17 607 751 649
rect 17 573 35 607
rect 69 573 699 607
rect 733 573 751 607
rect 17 510 751 573
rect 17 476 35 510
rect 69 476 699 510
rect 733 476 751 510
rect 17 414 751 476
rect 17 380 35 414
rect 69 380 699 414
rect 733 380 751 414
rect 17 354 751 380
rect 17 286 68 320
rect 102 286 136 320
rect 170 286 190 320
rect 17 215 190 286
rect 224 284 366 354
rect 224 250 244 284
rect 278 250 312 284
rect 346 250 366 284
rect 400 286 420 320
rect 454 286 488 320
rect 522 286 542 320
rect 400 215 542 286
rect 576 284 751 354
rect 576 250 596 284
rect 630 250 664 284
rect 698 250 751 284
rect 17 214 542 215
rect 17 190 751 214
rect 17 156 35 190
rect 69 156 699 190
rect 733 156 751 190
rect 17 93 751 156
rect 17 59 35 93
rect 69 59 699 93
rect 733 59 751 93
rect 17 17 751 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 1 nsew
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 4 nsew
rlabel comment s 0 0 0 0 4 decaphe_8
flabel nbase s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 3 nsew
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 768 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2465784
string GDS_START 2461832
<< end >>
