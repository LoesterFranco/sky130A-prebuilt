magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 17 206 73 493
rect 17 51 85 206
rect 211 215 311 261
rect 397 255 431 478
rect 345 215 431 255
rect 465 215 535 323
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 107 372 253 527
rect 296 338 362 493
rect 120 295 362 338
rect 120 181 177 295
rect 476 383 620 527
rect 120 143 277 181
rect 123 17 157 109
rect 205 51 277 143
rect 311 143 542 181
rect 311 111 353 143
rect 396 17 430 109
rect 476 51 542 143
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 465 215 535 323 6 A1
port 1 nsew signal input
rlabel locali s 397 255 431 478 6 A2
port 2 nsew signal input
rlabel locali s 345 215 431 255 6 A2
port 2 nsew signal input
rlabel locali s 211 215 311 261 6 B1
port 3 nsew signal input
rlabel locali s 17 206 73 493 6 X
port 4 nsew signal output
rlabel locali s 17 51 85 206 6 X
port 4 nsew signal output
rlabel metal1 s 0 -48 644 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 969130
string GDS_START 963366
<< end >>
