magic
tech sky130A
magscale 1 2
timestamp 1604502729
<< locali >>
rect 17 364 89 596
rect 17 226 51 364
rect 217 342 263 356
rect 193 284 263 342
rect 301 286 367 356
rect 17 70 91 226
rect 601 236 743 302
rect 777 236 843 302
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 123 390 189 649
rect 331 490 564 649
rect 230 390 476 456
rect 598 414 664 556
rect 85 260 159 326
rect 125 250 159 260
rect 410 252 476 390
rect 125 216 292 250
rect 125 17 224 182
rect 258 85 292 216
rect 326 218 476 252
rect 529 380 664 414
rect 774 380 840 649
rect 326 119 376 218
rect 529 184 563 380
rect 497 85 563 184
rect 258 51 563 85
rect 599 168 841 202
rect 599 68 649 168
rect 683 17 749 134
rect 791 68 841 168
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel locali s 217 342 263 356 6 A1_N
port 1 nsew signal input
rlabel locali s 193 284 263 342 6 A1_N
port 1 nsew signal input
rlabel locali s 301 286 367 356 6 A2_N
port 2 nsew signal input
rlabel locali s 777 236 843 302 6 B1
port 3 nsew signal input
rlabel locali s 601 236 743 302 6 B2
port 4 nsew signal input
rlabel locali s 17 364 89 596 6 X
port 5 nsew signal output
rlabel locali s 17 226 51 364 6 X
port 5 nsew signal output
rlabel locali s 17 70 91 226 6 X
port 5 nsew signal output
rlabel metal1 s 0 -49 864 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 864 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1260800
string GDS_START 1252926
<< end >>
