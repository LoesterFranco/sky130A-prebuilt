magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 87 293 377 327
rect 87 265 123 293
rect 17 199 123 265
rect 341 265 377 293
rect 173 199 307 259
rect 341 199 393 265
rect 495 323 549 493
rect 683 323 737 493
rect 871 323 925 493
rect 495 289 995 323
rect 895 177 995 289
rect 495 143 995 177
rect 495 51 549 143
rect 683 51 737 143
rect 871 51 925 143
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 19 361 79 527
rect 113 395 173 493
rect 207 429 273 527
rect 307 395 361 493
rect 395 432 461 527
rect 113 361 461 395
rect 427 253 461 361
rect 583 357 649 527
rect 771 357 837 527
rect 959 357 1025 527
rect 427 211 861 253
rect 427 165 461 211
rect 19 17 85 165
rect 203 131 461 165
rect 203 51 269 131
rect 388 17 454 97
rect 583 17 649 109
rect 771 17 837 109
rect 959 17 1025 109
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
rlabel locali s 173 199 307 259 6 A
port 1 nsew signal input
rlabel locali s 341 265 377 293 6 B
port 2 nsew signal input
rlabel locali s 341 199 393 265 6 B
port 2 nsew signal input
rlabel locali s 87 293 377 327 6 B
port 2 nsew signal input
rlabel locali s 87 265 123 293 6 B
port 2 nsew signal input
rlabel locali s 17 199 123 265 6 B
port 2 nsew signal input
rlabel locali s 895 177 995 289 6 X
port 3 nsew signal output
rlabel locali s 871 323 925 493 6 X
port 3 nsew signal output
rlabel locali s 871 51 925 143 6 X
port 3 nsew signal output
rlabel locali s 683 323 737 493 6 X
port 3 nsew signal output
rlabel locali s 683 51 737 143 6 X
port 3 nsew signal output
rlabel locali s 495 323 549 493 6 X
port 3 nsew signal output
rlabel locali s 495 289 995 323 6 X
port 3 nsew signal output
rlabel locali s 495 143 995 177 6 X
port 3 nsew signal output
rlabel locali s 495 51 549 143 6 X
port 3 nsew signal output
rlabel metal1 s 0 -48 1104 48 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 496 1104 592 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1104 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3336940
string GDS_START 3328550
<< end >>
