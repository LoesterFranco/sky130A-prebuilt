magic
tech sky130A
magscale 1 2
timestamp 1601050088
<< locali >>
rect 137 394 171 596
rect 301 394 367 596
rect 25 360 367 394
rect 25 226 71 360
rect 485 287 551 356
rect 697 290 839 356
rect 25 192 338 226
rect 889 252 981 356
rect 132 70 166 192
rect 288 70 338 192
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 31 428 97 649
rect 211 428 261 649
rect 407 390 457 649
rect 495 581 725 615
rect 495 390 545 581
rect 127 260 441 326
rect 374 253 441 260
rect 585 256 651 547
rect 691 424 725 581
rect 765 458 815 649
rect 855 424 905 596
rect 945 458 1011 649
rect 1051 424 1101 596
rect 691 390 1101 424
rect 1051 388 1101 390
rect 585 253 844 256
rect 374 222 844 253
rect 374 219 651 222
rect 30 17 96 158
rect 202 17 252 158
rect 374 17 424 185
rect 472 90 522 219
rect 558 17 624 185
rect 692 85 758 188
rect 792 119 844 222
rect 880 184 1102 218
rect 880 85 914 184
rect 692 51 914 85
rect 950 17 1016 150
rect 1052 70 1102 184
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
rlabel locali s 697 290 839 356 6 A1
port 1 nsew signal input
rlabel locali s 889 252 981 356 6 A2
port 2 nsew signal input
rlabel locali s 485 287 551 356 6 B1
port 3 nsew signal input
rlabel locali s 301 394 367 596 6 X
port 4 nsew signal output
rlabel locali s 288 70 338 192 6 X
port 4 nsew signal output
rlabel locali s 137 394 171 596 6 X
port 4 nsew signal output
rlabel locali s 132 70 166 192 6 X
port 4 nsew signal output
rlabel locali s 25 360 367 394 6 X
port 4 nsew signal output
rlabel locali s 25 226 71 360 6 X
port 4 nsew signal output
rlabel locali s 25 192 338 226 6 X
port 4 nsew signal output
rlabel metal1 s 0 -49 1152 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 617 1152 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3962942
string GDS_START 3953422
<< end >>
