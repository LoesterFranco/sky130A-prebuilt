magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 644 561
rect 21 357 87 527
rect 382 435 448 527
rect 199 393 259 425
rect 482 393 529 493
rect 199 357 529 393
rect 24 289 419 323
rect 24 211 90 289
rect 124 215 284 255
rect 320 215 419 289
rect 123 17 157 109
rect 305 17 339 109
rect 487 119 529 357
rect 563 314 625 527
rect 563 153 626 280
rect 0 -17 644 17
<< obsli1 >>
rect 121 459 343 493
rect 121 357 165 459
rect 305 427 343 459
rect 21 143 453 177
rect 21 51 87 143
rect 193 51 259 143
rect 387 85 453 143
rect 563 85 625 119
rect 387 51 625 85
<< metal1 >>
rect 0 496 644 592
rect 0 -48 644 48
<< labels >>
rlabel locali s 320 215 419 289 6 A1
port 1 nsew signal input
rlabel locali s 24 289 419 323 6 A1
port 1 nsew signal input
rlabel locali s 24 211 90 289 6 A1
port 1 nsew signal input
rlabel locali s 124 215 284 255 6 A2
port 2 nsew signal input
rlabel locali s 563 153 626 280 6 B1
port 3 nsew signal input
rlabel locali s 487 119 529 357 6 Y
port 4 nsew signal output
rlabel locali s 482 393 529 493 6 Y
port 4 nsew signal output
rlabel locali s 199 393 259 425 6 Y
port 4 nsew signal output
rlabel locali s 199 357 529 393 6 Y
port 4 nsew signal output
rlabel locali s 305 17 339 109 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 123 17 157 109 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 644 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 644 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 563 314 625 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 382 435 448 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 21 357 87 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 644 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 644 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1359170
string GDS_START 1352726
<< end >>
