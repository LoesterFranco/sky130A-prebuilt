magic
tech sky130A
magscale 1 2
timestamp 1601050088
<< locali >>
rect 85 196 161 398
rect 303 264 369 356
rect 893 236 957 302
rect 991 236 1082 349
rect 1279 236 1345 310
rect 3092 430 3141 596
rect 3092 310 3239 430
rect 3092 226 3141 310
rect 3075 70 3141 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3264 683
rect 17 492 102 596
rect 210 526 260 649
rect 294 581 464 615
rect 294 492 328 581
rect 17 458 328 492
rect 17 162 51 458
rect 362 424 396 547
rect 430 492 464 581
rect 498 526 548 649
rect 650 492 700 595
rect 430 458 700 492
rect 195 390 477 424
rect 195 230 261 390
rect 411 304 477 390
rect 511 303 614 369
rect 666 269 700 458
rect 634 235 700 269
rect 734 581 968 615
rect 734 459 790 581
rect 195 196 373 230
rect 634 201 668 235
rect 734 201 768 459
rect 825 451 900 547
rect 934 485 968 581
rect 1002 519 1052 649
rect 1160 508 1226 587
rect 1272 542 1339 649
rect 1551 542 1617 649
rect 1753 538 1803 596
rect 1651 508 1803 538
rect 1160 504 1803 508
rect 1837 504 1909 596
rect 2043 546 2109 649
rect 2262 546 2330 649
rect 1160 485 1685 504
rect 934 474 1685 485
rect 934 451 1245 474
rect 825 417 859 451
rect 17 70 113 162
rect 211 17 277 162
rect 323 109 373 196
rect 409 17 475 201
rect 573 135 668 201
rect 702 109 768 201
rect 802 383 1177 417
rect 802 202 859 383
rect 1124 283 1177 383
rect 1211 213 1245 451
rect 1379 306 1523 440
rect 1573 330 1607 474
rect 1729 440 1801 470
rect 1641 404 1801 440
rect 1641 364 1763 404
rect 1837 366 1871 504
rect 1943 478 2546 512
rect 1943 470 1977 478
rect 1905 404 1977 470
rect 2150 410 2225 444
rect 802 121 943 202
rect 802 51 859 121
rect 977 17 1043 202
rect 1135 179 1245 213
rect 1379 202 1413 306
rect 1573 296 1695 330
rect 1135 121 1201 179
rect 1247 17 1299 136
rect 1335 70 1413 202
rect 1447 17 1497 226
rect 1533 85 1599 226
rect 1645 119 1695 296
rect 1729 85 1763 364
rect 1797 332 2157 366
rect 1797 119 1831 332
rect 2091 306 2157 332
rect 2191 304 2225 410
rect 1983 272 2049 298
rect 2191 272 2360 304
rect 1865 204 1931 269
rect 1983 238 2360 272
rect 2408 272 2474 360
rect 2512 351 2546 478
rect 2580 385 2650 596
rect 2738 530 2846 649
rect 2880 494 2950 596
rect 2702 460 2950 494
rect 2702 419 2768 460
rect 2816 385 2882 426
rect 2616 351 2882 385
rect 2512 306 2582 351
rect 2624 272 2690 317
rect 2408 238 2690 272
rect 1865 170 2141 204
rect 1865 85 1899 170
rect 1533 51 1899 85
rect 2020 17 2073 136
rect 2107 85 2141 170
rect 2175 119 2225 238
rect 2408 204 2442 238
rect 2724 204 2758 351
rect 2816 292 2882 351
rect 2916 356 2950 460
rect 2992 390 3058 649
rect 3175 464 3241 649
rect 2916 310 3047 356
rect 2916 258 2950 310
rect 2259 170 2442 204
rect 2478 170 2758 204
rect 2863 224 2950 258
rect 2259 85 2293 170
rect 2107 51 2293 85
rect 2327 17 2377 136
rect 2478 70 2544 170
rect 2642 17 2829 136
rect 2863 70 2929 224
rect 2975 17 3041 190
rect 3175 17 3241 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3264 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 3199 649 3233 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
<< metal1 >>
rect 0 683 3264 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3264 683
rect 0 617 3264 649
rect 0 17 3264 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3264 17
rect 0 -49 3264 -17
<< obsm1 >>
rect 499 347 557 356
rect 2995 347 3053 356
rect 499 319 3053 347
rect 499 310 557 319
rect 2995 310 3053 319
<< labels >>
rlabel locali s 85 196 161 398 6 D
port 1 nsew signal input
rlabel locali s 303 264 369 356 6 DE
port 2 nsew signal input
rlabel locali s 3092 430 3141 596 6 Q
port 3 nsew signal output
rlabel locali s 3092 310 3239 430 6 Q
port 3 nsew signal output
rlabel locali s 3092 226 3141 310 6 Q
port 3 nsew signal output
rlabel locali s 3075 70 3141 226 6 Q
port 3 nsew signal output
rlabel locali s 991 236 1082 349 6 SCD
port 4 nsew signal input
rlabel locali s 893 236 957 302 6 SCE
port 5 nsew signal input
rlabel locali s 1279 236 1345 310 6 CLK
port 6 nsew clock input
rlabel metal1 s 0 -49 3264 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 617 3264 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 3264 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 428070
string GDS_START 406500
<< end >>
