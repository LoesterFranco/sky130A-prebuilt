magic
tech sky130A
magscale 1 2
timestamp 1604502701
<< nwell >>
rect -38 332 998 704
<< pwell >>
rect 0 0 960 49
<< scpmos >>
rect 86 392 116 592
rect 170 392 200 592
rect 372 368 402 592
rect 472 368 502 592
rect 562 368 592 592
rect 652 368 682 592
rect 742 368 772 592
rect 842 368 872 592
<< nmoslvt >>
rect 153 74 183 202
rect 239 74 269 202
rect 369 74 399 222
rect 455 74 485 222
rect 641 74 671 222
rect 727 74 757 222
rect 846 74 876 222
<< ndiff >>
rect 319 202 369 222
rect 27 84 153 202
rect 27 50 65 84
rect 99 74 153 84
rect 183 136 239 202
rect 183 102 194 136
rect 228 102 239 136
rect 183 74 239 102
rect 269 136 369 202
rect 269 102 294 136
rect 328 102 369 136
rect 269 74 369 102
rect 399 136 455 222
rect 399 102 410 136
rect 444 102 455 136
rect 399 74 455 102
rect 485 84 641 222
rect 485 74 513 84
rect 99 50 138 74
rect 27 38 138 50
rect 500 50 513 74
rect 547 74 641 84
rect 671 160 727 222
rect 671 126 682 160
rect 716 126 727 160
rect 671 74 727 126
rect 757 100 846 222
rect 757 74 784 100
rect 547 50 560 74
rect 500 38 560 50
rect 772 66 784 74
rect 818 74 846 100
rect 876 210 933 222
rect 876 176 887 210
rect 921 176 933 210
rect 876 120 933 176
rect 876 86 887 120
rect 921 86 933 120
rect 876 74 933 86
rect 818 66 831 74
rect 772 54 831 66
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 510 86 546
rect 27 476 39 510
rect 73 476 86 510
rect 27 392 86 476
rect 116 392 170 592
rect 200 580 259 592
rect 200 546 213 580
rect 247 546 259 580
rect 200 511 259 546
rect 200 477 213 511
rect 247 477 259 511
rect 200 442 259 477
rect 200 408 213 442
rect 247 408 259 442
rect 200 392 259 408
rect 313 580 372 592
rect 313 546 325 580
rect 359 546 372 580
rect 313 510 372 546
rect 313 476 325 510
rect 359 476 372 510
rect 313 368 372 476
rect 402 579 472 592
rect 402 545 415 579
rect 449 545 472 579
rect 402 368 472 545
rect 502 580 562 592
rect 502 546 515 580
rect 549 546 562 580
rect 502 510 562 546
rect 502 476 515 510
rect 549 476 562 510
rect 502 368 562 476
rect 592 531 652 592
rect 592 497 605 531
rect 639 497 652 531
rect 592 420 652 497
rect 592 386 605 420
rect 639 386 652 420
rect 592 368 652 386
rect 682 580 742 592
rect 682 546 695 580
rect 729 546 742 580
rect 682 472 742 546
rect 682 438 695 472
rect 729 438 742 472
rect 682 368 742 438
rect 772 546 842 592
rect 772 512 785 546
rect 819 512 842 546
rect 772 368 842 512
rect 872 580 933 592
rect 872 546 886 580
rect 920 546 933 580
rect 872 472 933 546
rect 872 438 886 472
rect 920 438 933 472
rect 872 368 933 438
<< ndiffc >>
rect 65 50 99 84
rect 194 102 228 136
rect 294 102 328 136
rect 410 102 444 136
rect 513 50 547 84
rect 682 126 716 160
rect 784 66 818 100
rect 887 176 921 210
rect 887 86 921 120
<< pdiffc >>
rect 39 546 73 580
rect 39 476 73 510
rect 213 546 247 580
rect 213 477 247 511
rect 213 408 247 442
rect 325 546 359 580
rect 325 476 359 510
rect 415 545 449 579
rect 515 546 549 580
rect 515 476 549 510
rect 605 497 639 531
rect 605 386 639 420
rect 695 546 729 580
rect 695 438 729 472
rect 785 512 819 546
rect 886 546 920 580
rect 886 438 920 472
<< poly >>
rect 86 592 116 618
rect 170 592 200 618
rect 372 592 402 618
rect 472 592 502 618
rect 562 592 592 618
rect 652 592 682 618
rect 742 592 772 618
rect 842 592 872 618
rect 86 377 116 392
rect 170 377 200 392
rect 83 299 119 377
rect 167 347 261 377
rect 372 353 402 368
rect 472 353 502 368
rect 562 353 592 368
rect 652 353 682 368
rect 742 353 772 368
rect 842 353 872 368
rect 83 283 183 299
rect 83 249 133 283
rect 167 249 183 283
rect 83 233 183 249
rect 153 202 183 233
rect 231 290 261 347
rect 369 336 405 353
rect 469 336 505 353
rect 369 320 505 336
rect 231 274 297 290
rect 231 240 247 274
rect 281 240 297 274
rect 231 224 297 240
rect 369 286 385 320
rect 419 286 453 320
rect 487 286 505 320
rect 369 270 505 286
rect 559 336 595 353
rect 649 336 685 353
rect 559 320 685 336
rect 559 286 575 320
rect 609 286 685 320
rect 739 310 775 353
rect 839 310 875 353
rect 559 270 685 286
rect 727 294 875 310
rect 239 202 269 224
rect 369 222 399 270
rect 455 222 485 270
rect 641 222 671 270
rect 727 260 779 294
rect 813 274 875 294
rect 813 260 876 274
rect 727 244 876 260
rect 727 222 757 244
rect 846 222 876 244
rect 153 48 183 74
rect 239 48 269 74
rect 369 48 399 74
rect 455 48 485 74
rect 641 48 671 74
rect 727 48 757 74
rect 846 48 876 74
<< polycont >>
rect 133 249 167 283
rect 247 240 281 274
rect 385 286 419 320
rect 453 286 487 320
rect 575 286 609 320
rect 779 260 813 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 23 580 89 649
rect 23 546 39 580
rect 73 546 89 580
rect 23 510 89 546
rect 23 476 39 510
rect 73 476 89 510
rect 23 460 89 476
rect 213 580 263 596
rect 247 546 263 580
rect 213 511 263 546
rect 247 477 263 511
rect 213 442 263 477
rect 309 580 359 596
rect 309 546 325 580
rect 309 510 359 546
rect 399 579 465 649
rect 399 545 415 579
rect 449 545 465 579
rect 399 528 465 545
rect 499 581 735 615
rect 499 580 565 581
rect 499 546 515 580
rect 549 546 565 580
rect 679 580 735 581
rect 309 476 325 510
rect 499 510 565 546
rect 499 494 515 510
rect 359 476 515 494
rect 549 476 565 510
rect 309 460 565 476
rect 605 531 639 547
rect 49 408 213 426
rect 247 426 263 442
rect 247 408 571 426
rect 49 392 571 408
rect 49 168 83 392
rect 117 324 503 358
rect 117 283 183 324
rect 369 320 503 324
rect 117 249 133 283
rect 167 249 183 283
rect 117 233 183 249
rect 231 274 297 290
rect 231 240 247 274
rect 281 240 297 274
rect 369 286 385 320
rect 419 286 453 320
rect 487 286 503 320
rect 369 270 503 286
rect 537 336 571 392
rect 605 420 639 497
rect 679 546 695 580
rect 729 546 735 580
rect 679 472 735 546
rect 769 546 835 649
rect 769 512 785 546
rect 819 512 835 546
rect 769 506 835 512
rect 869 580 937 596
rect 869 546 886 580
rect 920 546 937 580
rect 869 472 937 546
rect 679 438 695 472
rect 729 438 886 472
rect 920 438 937 472
rect 639 386 937 404
rect 605 370 937 386
rect 537 320 625 336
rect 537 286 575 320
rect 609 286 625 320
rect 537 270 625 286
rect 697 294 829 310
rect 231 236 297 240
rect 697 260 779 294
rect 813 260 829 294
rect 697 236 829 260
rect 231 202 829 236
rect 871 210 937 370
rect 871 176 887 210
rect 921 176 937 210
rect 871 168 937 176
rect 49 136 244 168
rect 49 134 194 136
rect 178 102 194 134
rect 228 102 244 136
rect 23 84 142 100
rect 23 50 65 84
rect 99 50 142 84
rect 178 70 244 102
rect 278 136 344 168
rect 278 102 294 136
rect 328 102 344 136
rect 23 17 142 50
rect 278 17 344 102
rect 394 136 632 168
rect 394 102 410 136
rect 444 134 632 136
rect 444 102 460 134
rect 394 70 460 102
rect 496 84 564 100
rect 496 50 513 84
rect 547 50 564 84
rect 598 85 632 134
rect 666 160 937 168
rect 666 126 682 160
rect 716 134 937 160
rect 716 126 732 134
rect 666 119 732 126
rect 871 120 937 134
rect 768 85 784 100
rect 598 66 784 85
rect 818 66 835 100
rect 871 86 887 120
rect 921 86 937 120
rect 871 70 937 86
rect 598 51 835 66
rect 496 17 564 50
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
rlabel comment s 0 0 0 0 4 xor2_2
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 703 242 737 276 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 895 94 929 128 0 FreeSans 340 0 0 0 X
port 7 nsew
flabel corelocali s 895 168 929 202 0 FreeSans 340 0 0 0 X
port 7 nsew
flabel corelocali s 895 242 929 276 0 FreeSans 340 0 0 0 X
port 7 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 X
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 960 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 558652
string GDS_START 550956
<< end >>
