magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 1510 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 93 47 123 177
rect 177 47 207 177
rect 271 47 301 177
rect 365 47 395 177
rect 469 47 499 177
rect 657 47 687 177
rect 751 47 781 177
rect 845 47 875 177
rect 949 47 979 177
rect 1033 47 1063 177
rect 1127 47 1157 177
rect 1221 47 1251 177
rect 1325 47 1355 177
<< pmoshvt >>
rect 85 297 121 497
rect 179 297 215 497
rect 273 297 309 497
rect 367 297 403 497
rect 461 297 497 497
rect 659 297 695 497
rect 753 297 789 497
rect 847 297 883 497
rect 941 297 977 497
rect 1035 297 1071 497
rect 1129 297 1165 497
rect 1223 297 1259 497
rect 1317 297 1353 497
<< ndiff >>
rect 27 163 93 177
rect 27 129 39 163
rect 73 129 93 163
rect 27 95 93 129
rect 27 61 39 95
rect 73 61 93 95
rect 27 47 93 61
rect 123 95 177 177
rect 123 61 133 95
rect 167 61 177 95
rect 123 47 177 61
rect 207 163 271 177
rect 207 129 227 163
rect 261 129 271 163
rect 207 95 271 129
rect 207 61 227 95
rect 261 61 271 95
rect 207 47 271 61
rect 301 95 365 177
rect 301 61 321 95
rect 355 61 365 95
rect 301 47 365 61
rect 395 163 469 177
rect 395 129 415 163
rect 449 129 469 163
rect 395 95 469 129
rect 395 61 415 95
rect 449 61 469 95
rect 395 47 469 61
rect 499 95 657 177
rect 499 61 509 95
rect 543 61 613 95
rect 647 61 657 95
rect 499 47 657 61
rect 687 163 751 177
rect 687 129 707 163
rect 741 129 751 163
rect 687 95 751 129
rect 687 61 707 95
rect 741 61 751 95
rect 687 47 751 61
rect 781 95 845 177
rect 781 61 801 95
rect 835 61 845 95
rect 781 47 845 61
rect 875 163 949 177
rect 875 129 895 163
rect 929 129 949 163
rect 875 95 949 129
rect 875 61 895 95
rect 929 61 949 95
rect 875 47 949 61
rect 979 95 1033 177
rect 979 61 989 95
rect 1023 61 1033 95
rect 979 47 1033 61
rect 1063 163 1127 177
rect 1063 129 1083 163
rect 1117 129 1127 163
rect 1063 95 1127 129
rect 1063 61 1083 95
rect 1117 61 1127 95
rect 1063 47 1127 61
rect 1157 95 1221 177
rect 1157 61 1177 95
rect 1211 61 1221 95
rect 1157 47 1221 61
rect 1251 163 1325 177
rect 1251 129 1271 163
rect 1305 129 1325 163
rect 1251 95 1325 129
rect 1251 61 1271 95
rect 1305 61 1325 95
rect 1251 47 1325 61
rect 1355 95 1407 177
rect 1355 61 1365 95
rect 1399 61 1407 95
rect 1355 47 1407 61
<< pdiff >>
rect 27 477 85 497
rect 27 443 39 477
rect 73 443 85 477
rect 27 409 85 443
rect 27 375 39 409
rect 73 375 85 409
rect 27 341 85 375
rect 27 307 39 341
rect 73 307 85 341
rect 27 297 85 307
rect 121 477 179 497
rect 121 443 133 477
rect 167 443 179 477
rect 121 409 179 443
rect 121 375 133 409
rect 167 375 179 409
rect 121 297 179 375
rect 215 477 273 497
rect 215 443 227 477
rect 261 443 273 477
rect 215 409 273 443
rect 215 375 227 409
rect 261 375 273 409
rect 215 297 273 375
rect 309 477 367 497
rect 309 443 321 477
rect 355 443 367 477
rect 309 297 367 443
rect 403 477 461 497
rect 403 443 415 477
rect 449 443 461 477
rect 403 409 461 443
rect 403 375 415 409
rect 449 375 461 409
rect 403 297 461 375
rect 497 477 551 497
rect 497 443 509 477
rect 543 443 551 477
rect 497 297 551 443
rect 605 477 659 497
rect 605 443 613 477
rect 647 443 659 477
rect 605 297 659 443
rect 695 409 753 497
rect 695 375 707 409
rect 741 375 753 409
rect 695 297 753 375
rect 789 477 847 497
rect 789 443 801 477
rect 835 443 847 477
rect 789 297 847 443
rect 883 409 941 497
rect 883 375 895 409
rect 929 375 941 409
rect 883 297 941 375
rect 977 477 1035 497
rect 977 443 989 477
rect 1023 443 1035 477
rect 977 409 1035 443
rect 977 375 989 409
rect 1023 375 1035 409
rect 977 297 1035 375
rect 1071 409 1129 497
rect 1071 375 1083 409
rect 1117 375 1129 409
rect 1071 341 1129 375
rect 1071 307 1083 341
rect 1117 307 1129 341
rect 1071 297 1129 307
rect 1165 477 1223 497
rect 1165 443 1177 477
rect 1211 443 1223 477
rect 1165 409 1223 443
rect 1165 375 1177 409
rect 1211 375 1223 409
rect 1165 297 1223 375
rect 1259 409 1317 497
rect 1259 375 1271 409
rect 1305 375 1317 409
rect 1259 341 1317 375
rect 1259 307 1271 341
rect 1305 307 1317 341
rect 1259 297 1317 307
rect 1353 477 1407 497
rect 1353 443 1365 477
rect 1399 443 1407 477
rect 1353 409 1407 443
rect 1353 375 1365 409
rect 1399 375 1407 409
rect 1353 297 1407 375
<< ndiffc >>
rect 39 129 73 163
rect 39 61 73 95
rect 133 61 167 95
rect 227 129 261 163
rect 227 61 261 95
rect 321 61 355 95
rect 415 129 449 163
rect 415 61 449 95
rect 509 61 543 95
rect 613 61 647 95
rect 707 129 741 163
rect 707 61 741 95
rect 801 61 835 95
rect 895 129 929 163
rect 895 61 929 95
rect 989 61 1023 95
rect 1083 129 1117 163
rect 1083 61 1117 95
rect 1177 61 1211 95
rect 1271 129 1305 163
rect 1271 61 1305 95
rect 1365 61 1399 95
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 133 443 167 477
rect 133 375 167 409
rect 227 443 261 477
rect 227 375 261 409
rect 321 443 355 477
rect 415 443 449 477
rect 415 375 449 409
rect 509 443 543 477
rect 613 443 647 477
rect 707 375 741 409
rect 801 443 835 477
rect 895 375 929 409
rect 989 443 1023 477
rect 989 375 1023 409
rect 1083 375 1117 409
rect 1083 307 1117 341
rect 1177 443 1211 477
rect 1177 375 1211 409
rect 1271 375 1305 409
rect 1271 307 1305 341
rect 1365 443 1399 477
rect 1365 375 1399 409
<< poly >>
rect 85 497 121 523
rect 179 497 215 523
rect 273 497 309 523
rect 367 497 403 523
rect 461 497 497 523
rect 659 497 695 523
rect 753 497 789 523
rect 847 497 883 523
rect 941 497 977 523
rect 1035 497 1071 523
rect 1129 497 1165 523
rect 1223 497 1259 523
rect 1317 497 1353 523
rect 85 282 121 297
rect 179 282 215 297
rect 273 282 309 297
rect 367 282 403 297
rect 461 282 497 297
rect 659 282 695 297
rect 753 282 789 297
rect 847 282 883 297
rect 941 282 977 297
rect 1035 282 1071 297
rect 1129 282 1165 297
rect 1223 282 1259 297
rect 1317 282 1353 297
rect 83 265 123 282
rect 22 249 123 265
rect 22 215 38 249
rect 72 215 123 249
rect 22 199 123 215
rect 93 177 123 199
rect 177 265 217 282
rect 271 265 311 282
rect 365 265 405 282
rect 459 265 499 282
rect 177 249 499 265
rect 177 215 271 249
rect 305 215 349 249
rect 383 215 427 249
rect 461 215 499 249
rect 177 199 499 215
rect 177 177 207 199
rect 271 177 301 199
rect 365 177 395 199
rect 469 177 499 199
rect 657 265 697 282
rect 751 265 791 282
rect 845 265 885 282
rect 939 265 979 282
rect 657 249 979 265
rect 657 215 673 249
rect 707 215 751 249
rect 785 215 829 249
rect 863 215 979 249
rect 657 199 979 215
rect 657 177 687 199
rect 751 177 781 199
rect 845 177 875 199
rect 949 177 979 199
rect 1033 265 1073 282
rect 1127 265 1167 282
rect 1221 265 1261 282
rect 1315 265 1355 282
rect 1033 249 1355 265
rect 1033 215 1049 249
rect 1083 215 1127 249
rect 1161 215 1205 249
rect 1239 215 1283 249
rect 1317 215 1355 249
rect 1033 199 1355 215
rect 1033 177 1063 199
rect 1127 177 1157 199
rect 1221 177 1251 199
rect 1325 177 1355 199
rect 93 21 123 47
rect 177 21 207 47
rect 271 21 301 47
rect 365 21 395 47
rect 469 21 499 47
rect 657 21 687 47
rect 751 21 781 47
rect 845 21 875 47
rect 949 21 979 47
rect 1033 21 1063 47
rect 1127 21 1157 47
rect 1221 21 1251 47
rect 1325 21 1355 47
<< polycont >>
rect 38 215 72 249
rect 271 215 305 249
rect 349 215 383 249
rect 427 215 461 249
rect 673 215 707 249
rect 751 215 785 249
rect 829 215 863 249
rect 1049 215 1083 249
rect 1127 215 1161 249
rect 1205 215 1239 249
rect 1283 215 1317 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 22 477 81 493
rect 22 443 39 477
rect 73 443 81 477
rect 22 409 81 443
rect 22 375 39 409
rect 73 375 81 409
rect 22 341 81 375
rect 125 477 175 527
rect 125 443 133 477
rect 167 443 175 477
rect 125 409 175 443
rect 125 375 133 409
rect 167 375 175 409
rect 125 359 175 375
rect 219 477 269 493
rect 219 443 227 477
rect 261 443 269 477
rect 219 409 269 443
rect 313 477 363 527
rect 313 443 321 477
rect 355 443 363 477
rect 313 427 363 443
rect 407 477 457 493
rect 407 443 415 477
rect 449 443 457 477
rect 219 375 227 409
rect 261 393 269 409
rect 407 409 457 443
rect 501 477 551 527
rect 501 443 509 477
rect 543 443 551 477
rect 501 427 551 443
rect 605 477 1407 493
rect 605 443 613 477
rect 647 459 801 477
rect 647 443 655 459
rect 605 427 655 443
rect 793 443 801 459
rect 835 459 989 477
rect 835 443 843 459
rect 793 427 843 443
rect 981 443 989 459
rect 1023 459 1177 477
rect 1023 443 1031 459
rect 407 393 415 409
rect 261 375 415 393
rect 449 393 457 409
rect 699 409 749 425
rect 699 393 707 409
rect 449 375 707 393
rect 741 393 749 409
rect 887 409 937 425
rect 887 393 895 409
rect 741 375 895 393
rect 929 375 937 409
rect 219 359 937 375
rect 981 409 1031 443
rect 1169 443 1177 459
rect 1211 459 1365 477
rect 1211 443 1219 459
rect 981 375 989 409
rect 1023 375 1031 409
rect 981 359 1031 375
rect 1075 409 1125 425
rect 1075 375 1083 409
rect 1117 375 1125 409
rect 22 307 39 341
rect 73 325 81 341
rect 1075 341 1125 375
rect 1169 409 1219 443
rect 1357 443 1365 459
rect 1399 443 1407 477
rect 1169 375 1177 409
rect 1211 375 1219 409
rect 1169 359 1219 375
rect 1263 409 1313 425
rect 1263 375 1271 409
rect 1305 375 1313 409
rect 73 307 1031 325
rect 22 291 1031 307
rect 1075 307 1083 341
rect 1117 325 1125 341
rect 1263 341 1313 375
rect 1357 409 1407 443
rect 1357 375 1365 409
rect 1399 375 1407 409
rect 1357 359 1407 375
rect 1263 325 1271 341
rect 1117 307 1271 325
rect 1305 325 1313 341
rect 1305 307 1449 325
rect 1075 291 1449 307
rect 22 249 89 257
rect 22 215 38 249
rect 72 215 89 249
rect 133 181 167 291
rect 997 257 1031 291
rect 242 249 554 257
rect 242 215 271 249
rect 305 215 349 249
rect 383 215 427 249
rect 461 215 554 249
rect 657 249 940 257
rect 657 215 673 249
rect 707 215 751 249
rect 785 215 829 249
rect 863 215 940 249
rect 997 249 1344 257
rect 997 215 1049 249
rect 1083 215 1127 249
rect 1161 215 1205 249
rect 1239 215 1283 249
rect 1317 215 1344 249
rect 1381 181 1449 291
rect 22 163 167 181
rect 22 129 39 163
rect 73 147 167 163
rect 201 163 1449 181
rect 73 129 89 147
rect 22 95 89 129
rect 201 129 227 163
rect 261 145 415 163
rect 261 129 277 145
rect 22 61 39 95
rect 73 61 89 95
rect 22 51 89 61
rect 133 95 167 111
rect 133 17 167 61
rect 201 95 277 129
rect 389 129 415 145
rect 449 145 707 163
rect 449 129 465 145
rect 201 61 227 95
rect 261 61 277 95
rect 201 51 277 61
rect 321 95 355 111
rect 321 17 355 61
rect 389 95 465 129
rect 681 129 707 145
rect 741 145 895 163
rect 741 129 757 145
rect 389 61 415 95
rect 449 61 465 95
rect 389 51 465 61
rect 509 95 647 111
rect 543 61 613 95
rect 509 17 647 61
rect 681 95 757 129
rect 869 129 895 145
rect 929 145 1083 163
rect 929 129 945 145
rect 681 61 707 95
rect 741 61 757 95
rect 681 51 757 61
rect 801 95 835 111
rect 801 17 835 61
rect 869 95 945 129
rect 1057 129 1083 145
rect 1117 145 1271 163
rect 1117 129 1133 145
rect 869 61 895 95
rect 929 61 945 95
rect 869 51 945 61
rect 989 95 1023 111
rect 989 17 1023 61
rect 1057 95 1133 129
rect 1245 129 1271 145
rect 1305 145 1449 163
rect 1305 129 1321 145
rect 1057 61 1083 95
rect 1117 61 1133 95
rect 1057 51 1133 61
rect 1177 95 1211 111
rect 1177 17 1211 61
rect 1245 95 1321 129
rect 1245 61 1271 95
rect 1305 61 1321 95
rect 1245 51 1321 61
rect 1365 95 1399 111
rect 1365 17 1399 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< labels >>
flabel corelocali s 395 221 429 255 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 488 221 522 255 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 303 221 337 255 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 400 0 0 0 C_N
port 3 nsew
flabel corelocali s 763 221 797 255 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel corelocali s 1408 221 1442 255 0 FreeSans 400 0 0 0 Y
port 8 nsew
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
rlabel comment s 0 0 0 0 4 nor3b_4
<< properties >>
string FIXED_BBOX 0 0 1472 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2474650
string GDS_START 2464006
<< end >>
