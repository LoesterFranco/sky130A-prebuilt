magic
tech sky130A
magscale 1 2
timestamp 1601050056
<< nwell >>
rect -38 332 902 704
<< pwell >>
rect 0 0 864 49
<< scpmos >>
rect 84 424 120 592
rect 323 368 359 568
rect 407 368 443 568
rect 491 368 527 568
rect 599 368 635 568
rect 737 368 773 592
<< nmoslvt >>
rect 84 74 114 184
rect 198 74 228 184
rect 413 74 443 184
rect 527 74 557 184
rect 613 74 643 184
rect 742 74 772 222
<< ndiff >>
rect 692 184 742 222
rect 27 146 84 184
rect 27 112 39 146
rect 73 112 84 146
rect 27 74 84 112
rect 114 146 198 184
rect 114 112 139 146
rect 173 112 198 146
rect 114 74 198 112
rect 228 159 413 184
rect 228 125 239 159
rect 273 125 368 159
rect 402 125 413 159
rect 228 74 413 125
rect 443 139 527 184
rect 443 105 468 139
rect 502 105 527 139
rect 443 74 527 105
rect 557 146 613 184
rect 557 112 568 146
rect 602 112 613 146
rect 557 74 613 112
rect 643 136 742 184
rect 643 102 675 136
rect 709 102 742 136
rect 643 74 742 102
rect 772 210 829 222
rect 772 176 783 210
rect 817 176 829 210
rect 772 120 829 176
rect 772 86 783 120
rect 817 86 829 120
rect 772 74 829 86
<< pdiff >>
rect 28 580 84 592
rect 28 546 40 580
rect 74 546 84 580
rect 28 470 84 546
rect 28 436 40 470
rect 74 436 84 470
rect 28 424 84 436
rect 120 580 186 592
rect 120 546 140 580
rect 174 546 186 580
rect 671 580 737 592
rect 671 568 683 580
rect 120 508 186 546
rect 120 474 140 508
rect 174 474 186 508
rect 120 424 186 474
rect 267 556 323 568
rect 267 522 279 556
rect 313 522 323 556
rect 267 485 323 522
rect 267 451 279 485
rect 313 451 323 485
rect 267 414 323 451
rect 267 380 279 414
rect 313 380 323 414
rect 267 368 323 380
rect 359 368 407 568
rect 443 368 491 568
rect 527 368 599 568
rect 635 546 683 568
rect 717 546 737 580
rect 635 508 737 546
rect 635 474 683 508
rect 717 474 737 508
rect 635 368 737 474
rect 773 580 829 592
rect 773 546 783 580
rect 817 546 829 580
rect 773 497 829 546
rect 773 463 783 497
rect 817 463 829 497
rect 773 414 829 463
rect 773 380 783 414
rect 817 380 829 414
rect 773 368 829 380
<< ndiffc >>
rect 39 112 73 146
rect 139 112 173 146
rect 239 125 273 159
rect 368 125 402 159
rect 468 105 502 139
rect 568 112 602 146
rect 675 102 709 136
rect 783 176 817 210
rect 783 86 817 120
<< pdiffc >>
rect 40 546 74 580
rect 40 436 74 470
rect 140 546 174 580
rect 140 474 174 508
rect 279 522 313 556
rect 279 451 313 485
rect 279 380 313 414
rect 683 546 717 580
rect 683 474 717 508
rect 783 546 817 580
rect 783 463 817 497
rect 783 380 817 414
<< poly >>
rect 84 592 120 618
rect 323 568 359 594
rect 407 568 443 594
rect 491 568 527 594
rect 599 568 635 594
rect 737 592 773 618
rect 84 356 120 424
rect 48 340 120 356
rect 48 306 64 340
rect 98 326 120 340
rect 162 366 228 382
rect 162 332 178 366
rect 212 353 228 366
rect 323 353 359 368
rect 212 332 359 353
rect 98 306 114 326
rect 162 323 359 332
rect 162 316 228 323
rect 48 290 114 306
rect 84 184 114 290
rect 198 184 228 316
rect 407 275 443 368
rect 377 259 443 275
rect 377 225 393 259
rect 427 225 443 259
rect 491 302 527 368
rect 599 336 635 368
rect 599 320 665 336
rect 737 326 773 368
rect 491 286 557 302
rect 491 252 507 286
rect 541 252 557 286
rect 599 286 615 320
rect 649 286 665 320
rect 599 270 665 286
rect 713 310 779 326
rect 713 276 729 310
rect 763 276 779 310
rect 491 236 557 252
rect 377 209 443 225
rect 413 184 443 209
rect 527 184 557 236
rect 613 184 643 270
rect 713 260 779 276
rect 742 222 772 260
rect 84 48 114 74
rect 198 48 228 74
rect 413 48 443 74
rect 527 48 557 74
rect 613 48 643 74
rect 742 48 772 74
<< polycont >>
rect 64 306 98 340
rect 178 332 212 366
rect 393 225 427 259
rect 507 252 541 286
rect 615 286 649 320
rect 729 276 763 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 24 580 90 596
rect 24 546 40 580
rect 74 546 90 580
rect 24 470 90 546
rect 24 436 40 470
rect 74 436 90 470
rect 124 580 190 649
rect 124 546 140 580
rect 174 546 190 580
rect 667 580 733 649
rect 124 508 190 546
rect 124 474 140 508
rect 174 474 190 508
rect 124 458 190 474
rect 263 556 329 572
rect 263 522 279 556
rect 313 522 329 556
rect 263 485 329 522
rect 24 424 90 436
rect 263 451 279 485
rect 313 451 329 485
rect 667 546 683 580
rect 717 546 733 580
rect 667 508 733 546
rect 667 474 683 508
rect 717 474 733 508
rect 667 458 733 474
rect 767 580 847 596
rect 767 546 783 580
rect 817 546 847 580
rect 767 497 847 546
rect 767 463 783 497
rect 817 463 847 497
rect 263 424 329 451
rect 24 390 196 424
rect 162 382 196 390
rect 263 414 733 424
rect 162 366 228 382
rect 25 340 114 356
rect 25 306 64 340
rect 98 306 114 340
rect 25 290 114 306
rect 162 332 178 366
rect 212 332 228 366
rect 162 316 228 332
rect 263 380 279 414
rect 313 390 733 414
rect 313 380 329 390
rect 162 256 196 316
rect 23 222 196 256
rect 23 146 89 222
rect 23 112 39 146
rect 73 112 89 146
rect 23 70 89 112
rect 123 146 189 188
rect 263 175 329 380
rect 377 259 455 356
rect 377 225 393 259
rect 427 225 455 259
rect 491 286 557 356
rect 491 252 507 286
rect 541 252 557 286
rect 599 320 665 356
rect 599 286 615 320
rect 649 286 665 320
rect 599 270 665 286
rect 699 326 733 390
rect 767 414 847 463
rect 767 380 783 414
rect 817 380 847 414
rect 767 364 847 380
rect 699 310 779 326
rect 699 276 729 310
rect 763 276 779 310
rect 491 236 557 252
rect 699 260 779 276
rect 699 236 733 260
rect 377 209 455 225
rect 591 202 733 236
rect 813 226 847 364
rect 767 210 847 226
rect 591 188 625 202
rect 123 112 139 146
rect 173 112 189 146
rect 123 17 189 112
rect 223 159 418 175
rect 223 125 239 159
rect 273 125 368 159
rect 402 125 418 159
rect 223 109 418 125
rect 452 139 518 175
rect 452 105 468 139
rect 502 105 518 139
rect 452 17 518 105
rect 552 146 625 188
rect 767 176 783 210
rect 817 176 847 210
rect 552 112 568 146
rect 602 112 625 146
rect 552 70 625 112
rect 659 136 725 168
rect 659 102 675 136
rect 709 102 725 136
rect 659 17 725 102
rect 767 120 847 176
rect 767 86 783 120
rect 817 86 847 120
rect 767 70 847 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
rlabel comment s 0 0 0 0 4 or4b_1
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 D_N
port 4 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 511 242 545 276 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 415 242 449 276 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 799 390 833 424 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 799 464 833 498 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 799 538 833 572 0 FreeSans 340 0 0 0 X
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 864 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 837484
string GDS_START 830176
<< end >>
