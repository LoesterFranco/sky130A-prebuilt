magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 2668 561
rect 103 439 153 527
rect 538 428 606 527
rect 17 153 69 335
rect 109 153 165 335
rect 211 153 267 335
rect 474 215 540 320
rect 581 318 617 392
rect 719 455 785 527
rect 581 211 713 318
rect 581 145 620 211
rect 17 17 96 119
rect 365 17 401 109
rect 1189 455 1255 527
rect 538 17 606 111
rect 1401 425 1592 527
rect 1839 447 1905 527
rect 2027 447 2093 527
rect 1328 289 1403 353
rect 726 17 788 109
rect 1777 305 2015 345
rect 1777 283 1822 305
rect 2224 297 2266 527
rect 1122 17 1219 93
rect 1347 17 1526 161
rect 2044 17 2078 109
rect 2224 17 2266 177
rect 2300 51 2366 493
rect 2515 315 2549 527
rect 2583 299 2651 490
rect 2614 165 2651 299
rect 2508 17 2549 165
rect 2583 55 2651 165
rect 0 -17 2668 17
<< obsli1 >>
rect 17 405 69 493
rect 187 451 409 493
rect 187 405 221 451
rect 454 417 504 493
rect 17 369 221 405
rect 259 374 339 415
rect 301 323 339 374
rect 301 289 305 323
rect 301 141 339 289
rect 373 354 504 417
rect 373 181 440 354
rect 651 391 685 465
rect 819 427 888 493
rect 651 357 765 391
rect 651 355 799 357
rect 373 143 503 181
rect 747 177 799 355
rect 299 133 339 141
rect 295 131 339 133
rect 295 129 334 131
rect 292 127 334 129
rect 289 126 334 127
rect 288 124 334 126
rect 286 123 334 124
rect 284 122 332 123
rect 281 121 332 122
rect 279 120 332 121
rect 276 118 332 120
rect 276 112 331 118
rect 175 56 331 112
rect 452 51 503 143
rect 654 143 799 177
rect 833 284 888 427
rect 922 323 966 493
rect 1006 427 1151 493
rect 1075 357 1083 391
rect 922 318 949 323
rect 932 289 949 318
rect 1041 315 1083 357
rect 833 255 898 284
rect 833 221 857 255
rect 891 221 898 255
rect 833 218 898 221
rect 654 51 691 143
rect 833 117 867 218
rect 932 184 966 289
rect 1117 279 1151 427
rect 1310 421 1353 490
rect 1626 425 1787 492
rect 1185 387 1353 421
rect 1753 413 1787 425
rect 1939 413 1982 490
rect 1185 315 1219 387
rect 1438 357 1501 391
rect 1535 357 1601 391
rect 1438 299 1601 357
rect 1017 255 1287 279
rect 1460 255 1532 265
rect 822 51 867 117
rect 901 51 966 184
rect 1000 245 1532 255
rect 1000 51 1088 245
rect 1122 161 1195 203
rect 1250 195 1532 245
rect 1567 179 1601 299
rect 1673 255 1719 381
rect 1753 379 2093 413
rect 2049 305 2093 379
rect 2127 271 2179 493
rect 1673 221 1685 255
rect 1673 215 1719 221
rect 1762 179 1808 249
rect 1122 127 1307 161
rect 1255 51 1307 127
rect 1567 139 1808 179
rect 1858 237 2179 271
rect 1858 171 1893 237
rect 1931 169 2109 203
rect 1931 89 1965 169
rect 1682 55 1965 89
rect 2143 108 2179 237
rect 2112 51 2179 108
rect 2412 265 2454 493
rect 2412 199 2580 265
rect 2412 51 2454 199
<< obsli1c >>
rect 305 289 339 323
rect 765 357 799 391
rect 1041 357 1075 391
rect 949 289 983 323
rect 857 221 891 255
rect 1501 357 1535 391
rect 1685 221 1719 255
<< metal1 >>
rect 0 496 2668 592
rect 1316 320 1374 329
rect 1765 320 1823 329
rect 1316 292 1823 320
rect 1316 283 1374 292
rect 1765 283 1823 292
rect 110 252 168 261
rect 477 252 535 261
rect 110 224 535 252
rect 110 215 168 224
rect 477 215 535 224
rect 0 -48 2668 48
<< obsm1 >>
rect 753 391 811 397
rect 753 357 765 391
rect 799 388 811 391
rect 1029 391 1087 397
rect 1029 388 1041 391
rect 799 360 1041 388
rect 799 357 811 360
rect 753 351 811 357
rect 1029 357 1041 360
rect 1075 388 1087 391
rect 1489 391 1547 397
rect 1489 388 1501 391
rect 1075 360 1501 388
rect 1075 357 1087 360
rect 1029 351 1087 357
rect 1489 357 1501 360
rect 1535 357 1547 391
rect 1489 351 1547 357
rect 293 323 351 329
rect 293 289 305 323
rect 339 320 351 323
rect 937 323 995 329
rect 937 320 949 323
rect 339 292 949 320
rect 339 289 351 292
rect 293 283 351 289
rect 937 289 949 292
rect 983 289 995 323
rect 937 283 995 289
rect 845 255 903 261
rect 845 221 857 255
rect 891 252 903 255
rect 1673 255 1731 261
rect 1673 252 1685 255
rect 891 224 1685 252
rect 891 221 903 224
rect 845 215 903 221
rect 1673 221 1685 224
rect 1719 221 1731 255
rect 1673 215 1731 221
<< labels >>
rlabel locali s 211 153 267 335 6 D
port 1 nsew signal input
rlabel locali s 2614 165 2651 299 6 Q
port 2 nsew signal output
rlabel locali s 2583 299 2651 490 6 Q
port 2 nsew signal output
rlabel locali s 2583 55 2651 165 6 Q
port 2 nsew signal output
rlabel locali s 2300 51 2366 493 6 Q_N
port 3 nsew signal output
rlabel locali s 17 153 69 335 6 SCD
port 4 nsew signal input
rlabel locali s 109 153 165 335 6 SCE
port 5 nsew signal input
rlabel locali s 474 215 540 320 6 SCE
port 5 nsew signal input
rlabel metal1 s 477 252 535 261 6 SCE
port 5 nsew signal input
rlabel metal1 s 477 215 535 224 6 SCE
port 5 nsew signal input
rlabel metal1 s 110 252 168 261 6 SCE
port 5 nsew signal input
rlabel metal1 s 110 224 535 252 6 SCE
port 5 nsew signal input
rlabel metal1 s 110 215 168 224 6 SCE
port 5 nsew signal input
rlabel locali s 1328 289 1403 353 6 SET_B
port 6 nsew signal input
rlabel locali s 1777 305 2015 345 6 SET_B
port 6 nsew signal input
rlabel locali s 1777 283 1822 305 6 SET_B
port 6 nsew signal input
rlabel metal1 s 1765 320 1823 329 6 SET_B
port 6 nsew signal input
rlabel metal1 s 1765 283 1823 292 6 SET_B
port 6 nsew signal input
rlabel metal1 s 1316 320 1374 329 6 SET_B
port 6 nsew signal input
rlabel metal1 s 1316 292 1823 320 6 SET_B
port 6 nsew signal input
rlabel metal1 s 1316 283 1374 292 6 SET_B
port 6 nsew signal input
rlabel locali s 581 318 617 392 6 CLK
port 7 nsew clock input
rlabel locali s 581 211 713 318 6 CLK
port 7 nsew clock input
rlabel locali s 581 145 620 211 6 CLK
port 7 nsew clock input
rlabel locali s 2508 17 2549 165 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 2224 17 2266 177 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 2044 17 2078 109 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 1347 17 1526 161 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 1122 17 1219 93 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 726 17 788 109 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 538 17 606 111 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 365 17 401 109 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 17 17 96 119 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 0 -17 2668 17 8 VGND
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 2668 48 8 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 2515 315 2549 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 2224 297 2266 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 2027 447 2093 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 1839 447 1905 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 1401 425 1592 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 1189 455 1255 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 719 455 785 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 538 428 606 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 103 439 153 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 0 527 2668 561 6 VPWR
port 9 nsew power bidirectional abutment
rlabel metal1 s 0 496 2668 592 6 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2668 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 99194
string GDS_START 77522
<< end >>
