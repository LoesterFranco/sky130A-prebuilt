magic
tech sky130A
magscale 1 2
timestamp 1601050088
<< locali >>
rect 121 332 359 367
rect 121 298 541 332
rect 313 162 420 253
rect 475 252 541 298
rect 589 296 655 430
rect 879 330 929 355
rect 757 252 929 330
rect 757 203 844 252
rect 2705 282 2757 596
rect 2705 70 2771 282
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2880 683
rect 23 435 89 596
rect 123 469 313 649
rect 421 503 487 615
rect 619 537 685 649
rect 723 525 799 615
rect 941 559 1007 649
rect 1149 525 1199 545
rect 723 503 1199 525
rect 421 489 1199 503
rect 1239 498 1374 545
rect 1430 532 1497 649
rect 1538 498 1604 545
rect 1239 495 1604 498
rect 421 469 799 489
rect 689 466 799 469
rect 23 401 541 435
rect 23 253 57 401
rect 475 366 541 401
rect 23 187 228 253
rect 23 70 73 187
rect 689 262 723 466
rect 1149 461 1199 489
rect 1340 464 1604 495
rect 1650 464 1716 649
rect 757 424 833 432
rect 757 390 799 424
rect 757 366 833 390
rect 867 423 917 455
rect 867 389 997 423
rect 1031 393 1115 455
rect 1149 427 1306 461
rect 1031 389 1233 393
rect 963 355 997 389
rect 575 228 723 262
rect 963 289 1043 355
rect 1077 327 1233 389
rect 575 169 609 228
rect 963 218 997 289
rect 1077 244 1124 327
rect 1272 293 1306 427
rect 878 184 997 218
rect 1031 197 1124 244
rect 1158 259 1306 293
rect 1031 184 1084 197
rect 878 169 914 184
rect 109 17 175 153
rect 221 85 287 128
rect 454 119 609 169
rect 643 85 683 156
rect 221 51 683 85
rect 733 17 793 156
rect 829 119 914 169
rect 948 17 1000 150
rect 1034 93 1084 184
rect 1158 130 1223 259
rect 1340 225 1374 464
rect 1263 191 1374 225
rect 1408 218 1463 415
rect 1497 315 1531 464
rect 1565 424 1703 430
rect 1565 390 1663 424
rect 1697 390 1703 424
rect 1565 359 1703 390
rect 1750 343 1823 551
rect 1864 504 2078 570
rect 2112 546 2248 649
rect 2282 512 2348 596
rect 1864 368 1920 504
rect 1497 252 1684 315
rect 1750 226 1784 343
rect 1957 267 2010 466
rect 1718 218 1784 226
rect 1263 129 1329 191
rect 1408 184 1784 218
rect 1403 116 1684 150
rect 1718 119 1784 184
rect 1818 201 2010 267
rect 2044 240 2078 504
rect 2112 478 2348 512
rect 2112 350 2170 478
rect 2222 424 2288 444
rect 2222 390 2239 424
rect 2273 390 2288 424
rect 2222 384 2288 390
rect 2389 388 2455 649
rect 2489 388 2555 596
rect 2112 316 2446 350
rect 2112 274 2170 316
rect 2204 240 2378 282
rect 2044 222 2378 240
rect 2044 206 2238 222
rect 1403 93 1451 116
rect 1034 53 1451 93
rect 1650 85 1684 116
rect 1818 85 1852 201
rect 2044 162 2078 206
rect 2412 188 2446 316
rect 1886 96 2078 162
rect 1521 17 1616 82
rect 1650 51 1852 85
rect 2151 17 2217 162
rect 2309 154 2446 188
rect 2521 326 2555 388
rect 2601 364 2667 649
rect 2521 260 2671 326
rect 2791 364 2857 649
rect 2309 70 2375 154
rect 2421 17 2487 120
rect 2521 70 2573 260
rect 2619 17 2669 226
rect 2807 17 2857 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2880 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 799 390 833 424
rect 1663 390 1697 424
rect 2239 390 2273 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
<< metal1 >>
rect 0 683 2880 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2880 683
rect 0 617 2880 649
rect 787 424 845 430
rect 787 390 799 424
rect 833 421 845 424
rect 1651 424 1709 430
rect 1651 421 1663 424
rect 833 393 1663 421
rect 833 390 845 393
rect 787 384 845 390
rect 1651 390 1663 393
rect 1697 421 1709 424
rect 2227 424 2285 430
rect 2227 421 2239 424
rect 1697 393 2239 421
rect 1697 390 1709 393
rect 1651 384 1709 390
rect 2227 390 2239 393
rect 2273 390 2285 424
rect 2227 384 2285 390
rect 0 17 2880 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2880 17
rect 0 -49 2880 -17
<< labels >>
rlabel locali s 313 162 420 253 6 D
port 1 nsew signal input
rlabel locali s 2705 282 2757 596 6 Q
port 2 nsew signal output
rlabel locali s 2705 70 2771 282 6 Q
port 2 nsew signal output
rlabel metal1 s 2227 421 2285 430 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 2227 384 2285 393 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 1651 421 1709 430 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 1651 384 1709 393 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 787 421 845 430 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 787 393 2285 421 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 787 384 845 393 6 RESET_B
port 3 nsew signal input
rlabel locali s 589 296 655 430 6 SCD
port 4 nsew signal input
rlabel locali s 475 252 541 298 6 SCE
port 5 nsew signal input
rlabel locali s 121 332 359 367 6 SCE
port 5 nsew signal input
rlabel locali s 121 298 541 332 6 SCE
port 5 nsew signal input
rlabel locali s 879 330 929 355 6 CLK
port 6 nsew clock input
rlabel locali s 757 252 929 330 6 CLK
port 6 nsew clock input
rlabel locali s 757 203 844 252 6 CLK
port 6 nsew clock input
rlabel metal1 s 0 -49 2880 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 617 2880 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2880 666
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 210386
string GDS_START 189392
<< end >>
