magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 116 333 192 493
rect 304 333 380 493
rect 492 333 568 493
rect 680 333 756 493
rect 868 333 944 493
rect 1056 333 1132 493
rect 1244 333 1320 493
rect 1432 333 1508 493
rect 116 299 1508 333
rect 17 215 1225 263
rect 1403 181 1508 299
rect 116 143 1508 181
rect 116 51 192 143
rect 304 51 380 143
rect 492 51 568 143
rect 680 51 756 143
rect 868 51 944 143
rect 1056 51 1132 143
rect 1244 51 1320 143
rect 1432 51 1508 143
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 40 297 82 527
rect 236 367 270 527
rect 424 367 458 527
rect 612 367 646 527
rect 800 367 834 527
rect 988 367 1022 527
rect 1176 367 1210 527
rect 1364 367 1398 527
rect 1552 367 1594 527
rect 36 17 82 177
rect 236 17 270 109
rect 424 17 458 109
rect 612 17 646 109
rect 800 17 834 109
rect 988 17 1022 109
rect 1176 17 1210 109
rect 1364 17 1398 109
rect 1552 17 1594 177
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
<< metal1 >>
rect 0 561 1656 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 0 496 1656 527
rect 0 17 1656 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
rect 0 -48 1656 -17
<< labels >>
rlabel locali s 17 215 1225 263 6 A
port 1 nsew signal input
rlabel locali s 1432 333 1508 493 6 Y
port 2 nsew signal output
rlabel locali s 1432 51 1508 143 6 Y
port 2 nsew signal output
rlabel locali s 1403 181 1508 299 6 Y
port 2 nsew signal output
rlabel locali s 1244 333 1320 493 6 Y
port 2 nsew signal output
rlabel locali s 1244 51 1320 143 6 Y
port 2 nsew signal output
rlabel locali s 1056 333 1132 493 6 Y
port 2 nsew signal output
rlabel locali s 1056 51 1132 143 6 Y
port 2 nsew signal output
rlabel locali s 868 333 944 493 6 Y
port 2 nsew signal output
rlabel locali s 868 51 944 143 6 Y
port 2 nsew signal output
rlabel locali s 680 333 756 493 6 Y
port 2 nsew signal output
rlabel locali s 680 51 756 143 6 Y
port 2 nsew signal output
rlabel locali s 492 333 568 493 6 Y
port 2 nsew signal output
rlabel locali s 492 51 568 143 6 Y
port 2 nsew signal output
rlabel locali s 304 333 380 493 6 Y
port 2 nsew signal output
rlabel locali s 304 51 380 143 6 Y
port 2 nsew signal output
rlabel locali s 116 333 192 493 6 Y
port 2 nsew signal output
rlabel locali s 116 299 1508 333 6 Y
port 2 nsew signal output
rlabel locali s 116 143 1508 181 6 Y
port 2 nsew signal output
rlabel locali s 116 51 192 143 6 Y
port 2 nsew signal output
rlabel metal1 s 0 -48 1656 48 8 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 496 1656 592 6 VPWR
port 4 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1656 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2097992
string GDS_START 2085580
<< end >>
