magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 736 561
rect 120 366 185 527
rect 17 215 97 264
rect 447 367 569 527
rect 607 313 719 493
rect 116 17 182 113
rect 646 128 719 313
rect 448 17 569 113
rect 603 51 719 128
rect 0 -17 736 17
<< obsli1 >>
rect 17 332 86 493
rect 239 358 329 493
rect 17 298 201 332
rect 131 259 201 298
rect 131 205 221 259
rect 294 250 329 358
rect 363 333 413 493
rect 363 299 553 333
rect 519 265 553 299
rect 294 215 484 250
rect 131 181 201 205
rect 17 147 201 181
rect 294 171 329 215
rect 519 198 610 265
rect 519 181 553 198
rect 17 51 82 147
rect 235 51 329 171
rect 363 147 553 181
rect 363 51 413 147
<< metal1 >>
rect 0 496 736 592
rect 0 -48 736 48
<< labels >>
rlabel locali s 17 215 97 264 6 A
port 1 nsew signal input
rlabel locali s 646 128 719 313 6 X
port 2 nsew signal output
rlabel locali s 607 313 719 493 6 X
port 2 nsew signal output
rlabel locali s 603 51 719 128 6 X
port 2 nsew signal output
rlabel locali s 448 17 569 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 116 17 182 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 0 -17 736 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 736 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 447 367 569 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 120 366 185 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 0 527 736 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 496 736 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3129812
string GDS_START 3123692
<< end >>
