magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 489 333 549 493
rect 683 333 737 493
rect 871 333 925 493
rect 1059 333 1113 493
rect 1247 333 1301 493
rect 1435 333 1489 493
rect 489 295 1489 333
rect 105 215 264 261
rect 1392 181 1489 295
rect 495 143 1489 181
rect 495 56 549 143
rect 683 56 737 143
rect 871 56 925 143
rect 1059 56 1113 143
rect 1247 56 1301 143
rect 1435 56 1489 143
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 19 299 79 527
rect 113 333 179 493
rect 213 367 267 527
rect 307 333 361 493
rect 113 299 361 333
rect 114 295 361 299
rect 395 295 455 527
rect 583 367 649 527
rect 771 367 837 527
rect 959 367 1025 527
rect 1147 367 1213 527
rect 1335 367 1401 527
rect 307 261 361 295
rect 307 215 1337 261
rect 307 181 361 215
rect 1523 293 1589 527
rect 119 143 361 181
rect 19 17 85 122
rect 119 56 173 143
rect 207 17 273 109
rect 307 56 361 143
rect 395 17 461 109
rect 583 17 649 109
rect 771 17 837 109
rect 959 17 1025 109
rect 1147 17 1213 109
rect 1335 17 1401 109
rect 1523 17 1589 122
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
<< metal1 >>
rect 0 561 1656 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 0 496 1656 527
rect 0 17 1656 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
rect 0 -48 1656 -17
<< labels >>
rlabel locali s 105 215 264 261 6 A
port 1 nsew signal input
rlabel locali s 1435 333 1489 493 6 X
port 2 nsew signal output
rlabel locali s 1435 56 1489 143 6 X
port 2 nsew signal output
rlabel locali s 1392 181 1489 295 6 X
port 2 nsew signal output
rlabel locali s 1247 333 1301 493 6 X
port 2 nsew signal output
rlabel locali s 1247 56 1301 143 6 X
port 2 nsew signal output
rlabel locali s 1059 333 1113 493 6 X
port 2 nsew signal output
rlabel locali s 1059 56 1113 143 6 X
port 2 nsew signal output
rlabel locali s 871 333 925 493 6 X
port 2 nsew signal output
rlabel locali s 871 56 925 143 6 X
port 2 nsew signal output
rlabel locali s 683 333 737 493 6 X
port 2 nsew signal output
rlabel locali s 683 56 737 143 6 X
port 2 nsew signal output
rlabel locali s 495 143 1489 181 6 X
port 2 nsew signal output
rlabel locali s 495 56 549 143 6 X
port 2 nsew signal output
rlabel locali s 489 333 549 493 6 X
port 2 nsew signal output
rlabel locali s 489 295 1489 333 6 X
port 2 nsew signal output
rlabel metal1 s 0 -48 1656 48 8 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 496 1656 592 6 VPWR
port 4 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1656 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3365784
string GDS_START 3354012
<< end >>
