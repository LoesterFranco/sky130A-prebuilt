magic
tech sky130A
timestamp 1599587575
<< properties >>
string gencell xind4_02
string parameter m=1
string library sky130
<< end >>
