magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 2024 561
rect 31 359 81 527
rect 199 359 249 527
rect 367 359 417 527
rect 535 359 585 527
rect 703 359 851 527
rect 885 325 935 493
rect 969 359 1019 527
rect 1053 325 1103 493
rect 1137 359 1187 527
rect 1325 325 1375 425
rect 1493 325 1543 425
rect 885 291 1543 325
rect 1661 359 1711 527
rect 1829 359 1879 527
rect 85 215 365 257
rect 419 215 701 257
rect 1175 181 1231 291
rect 1293 215 1575 257
rect 1609 215 2001 257
rect 459 17 493 111
rect 627 17 661 111
rect 883 129 1231 181
rect 1333 17 1367 111
rect 1501 17 1535 111
rect 1669 17 1703 111
rect 1837 17 1871 111
rect 0 -17 2024 17
<< obsli1 >>
rect 115 325 165 493
rect 283 325 333 493
rect 451 325 501 493
rect 619 325 669 493
rect 1235 459 1627 493
rect 1235 359 1291 459
rect 1409 359 1459 459
rect 17 291 783 325
rect 1577 325 1627 459
rect 1745 325 1795 493
rect 1913 325 1975 493
rect 1577 291 1975 325
rect 17 181 51 291
rect 749 257 783 291
rect 749 215 1141 257
rect 17 129 341 181
rect 375 145 761 181
rect 375 95 425 145
rect 20 51 425 95
rect 527 51 593 145
rect 695 51 761 145
rect 812 95 849 167
rect 1265 147 1971 181
rect 1265 95 1299 147
rect 1401 145 1971 147
rect 812 51 1299 95
rect 1401 51 1467 145
rect 1569 51 1635 145
rect 1737 51 1803 145
rect 1905 51 1971 145
<< metal1 >>
rect 0 496 2024 592
rect 0 -48 2024 48
<< labels >>
rlabel locali s 419 215 701 257 6 A1_N
port 1 nsew signal input
rlabel locali s 85 215 365 257 6 A2_N
port 2 nsew signal input
rlabel locali s 1609 215 2001 257 6 B1
port 3 nsew signal input
rlabel locali s 1293 215 1575 257 6 B2
port 4 nsew signal input
rlabel locali s 1493 325 1543 425 6 Y
port 5 nsew signal output
rlabel locali s 1325 325 1375 425 6 Y
port 5 nsew signal output
rlabel locali s 1175 181 1231 291 6 Y
port 5 nsew signal output
rlabel locali s 1053 325 1103 493 6 Y
port 5 nsew signal output
rlabel locali s 885 325 935 493 6 Y
port 5 nsew signal output
rlabel locali s 885 291 1543 325 6 Y
port 5 nsew signal output
rlabel locali s 883 129 1231 181 6 Y
port 5 nsew signal output
rlabel locali s 1837 17 1871 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1669 17 1703 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1501 17 1535 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1333 17 1367 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 627 17 661 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 459 17 493 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 2024 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 2024 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1829 359 1879 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1661 359 1711 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1137 359 1187 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 969 359 1019 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 703 359 851 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 535 359 585 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 367 359 417 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 199 359 249 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 31 359 81 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 2024 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 2024 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2024 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 739742
string GDS_START 724980
<< end >>
