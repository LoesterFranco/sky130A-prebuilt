magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 1958 704
<< pwell >>
rect 0 0 1920 49
<< scnmos >>
rect 84 74 114 158
rect 170 74 200 158
rect 260 74 290 158
rect 346 74 376 158
rect 446 74 476 158
rect 532 74 562 158
rect 618 74 648 158
rect 704 74 734 158
rect 790 74 820 158
rect 876 74 906 158
rect 976 74 1006 158
rect 1062 74 1092 158
rect 1162 74 1192 158
rect 1248 74 1278 158
rect 1348 74 1378 158
rect 1434 74 1464 158
rect 1534 74 1564 158
rect 1620 74 1650 158
rect 1720 74 1750 158
rect 1806 74 1836 158
<< pmoshvt >>
rect 87 368 117 592
rect 177 368 207 592
rect 267 368 297 592
rect 357 368 387 592
rect 449 368 479 592
rect 539 368 569 592
rect 629 368 659 592
rect 719 368 749 592
rect 809 368 839 592
rect 899 368 929 592
rect 989 368 1019 592
rect 1079 368 1109 592
rect 1169 368 1199 592
rect 1259 368 1289 592
rect 1349 368 1379 592
rect 1439 368 1469 592
rect 1529 368 1559 592
rect 1619 368 1649 592
rect 1713 368 1743 592
rect 1803 368 1833 592
<< ndiff >>
rect 27 133 84 158
rect 27 99 39 133
rect 73 99 84 133
rect 27 74 84 99
rect 114 133 170 158
rect 114 99 125 133
rect 159 99 170 133
rect 114 74 170 99
rect 200 133 260 158
rect 200 99 211 133
rect 245 99 260 133
rect 200 74 260 99
rect 290 133 346 158
rect 290 99 301 133
rect 335 99 346 133
rect 290 74 346 99
rect 376 133 446 158
rect 376 99 387 133
rect 421 99 446 133
rect 376 74 446 99
rect 476 133 532 158
rect 476 99 487 133
rect 521 99 532 133
rect 476 74 532 99
rect 562 120 618 158
rect 562 86 573 120
rect 607 86 618 120
rect 562 74 618 86
rect 648 133 704 158
rect 648 99 659 133
rect 693 99 704 133
rect 648 74 704 99
rect 734 129 790 158
rect 734 95 745 129
rect 779 95 790 129
rect 734 74 790 95
rect 820 133 876 158
rect 820 99 831 133
rect 865 99 876 133
rect 820 74 876 99
rect 906 132 976 158
rect 906 98 917 132
rect 951 98 976 132
rect 906 74 976 98
rect 1006 133 1062 158
rect 1006 99 1017 133
rect 1051 99 1062 133
rect 1006 74 1062 99
rect 1092 120 1162 158
rect 1092 86 1103 120
rect 1137 86 1162 120
rect 1092 74 1162 86
rect 1192 133 1248 158
rect 1192 99 1203 133
rect 1237 99 1248 133
rect 1192 74 1248 99
rect 1278 120 1348 158
rect 1278 86 1289 120
rect 1323 86 1348 120
rect 1278 74 1348 86
rect 1378 133 1434 158
rect 1378 99 1389 133
rect 1423 99 1434 133
rect 1378 74 1434 99
rect 1464 120 1534 158
rect 1464 86 1475 120
rect 1509 86 1534 120
rect 1464 74 1534 86
rect 1564 133 1620 158
rect 1564 99 1575 133
rect 1609 99 1620 133
rect 1564 74 1620 99
rect 1650 120 1720 158
rect 1650 86 1661 120
rect 1695 86 1720 120
rect 1650 74 1720 86
rect 1750 133 1806 158
rect 1750 99 1761 133
rect 1795 99 1806 133
rect 1750 74 1806 99
rect 1836 133 1893 158
rect 1836 99 1847 133
rect 1881 99 1893 133
rect 1836 74 1893 99
<< pdiff >>
rect 28 580 87 592
rect 28 546 40 580
rect 74 546 87 580
rect 28 510 87 546
rect 28 476 40 510
rect 74 476 87 510
rect 28 440 87 476
rect 28 406 40 440
rect 74 406 87 440
rect 28 368 87 406
rect 117 580 177 592
rect 117 546 130 580
rect 164 546 177 580
rect 117 510 177 546
rect 117 476 130 510
rect 164 476 177 510
rect 117 440 177 476
rect 117 406 130 440
rect 164 406 177 440
rect 117 368 177 406
rect 207 580 267 592
rect 207 546 220 580
rect 254 546 267 580
rect 207 508 267 546
rect 207 474 220 508
rect 254 474 267 508
rect 207 368 267 474
rect 297 580 357 592
rect 297 546 310 580
rect 344 546 357 580
rect 297 510 357 546
rect 297 476 310 510
rect 344 476 357 510
rect 297 440 357 476
rect 297 406 310 440
rect 344 406 357 440
rect 297 368 357 406
rect 387 580 449 592
rect 387 546 400 580
rect 434 546 449 580
rect 387 508 449 546
rect 387 474 400 508
rect 434 474 449 508
rect 387 368 449 474
rect 479 580 539 592
rect 479 546 492 580
rect 526 546 539 580
rect 479 497 539 546
rect 479 463 492 497
rect 526 463 539 497
rect 479 414 539 463
rect 479 380 492 414
rect 526 380 539 414
rect 479 368 539 380
rect 569 580 629 592
rect 569 546 582 580
rect 616 546 629 580
rect 569 508 629 546
rect 569 474 582 508
rect 616 474 629 508
rect 569 440 629 474
rect 569 406 582 440
rect 616 406 629 440
rect 569 368 629 406
rect 659 580 719 592
rect 659 546 672 580
rect 706 546 719 580
rect 659 497 719 546
rect 659 463 672 497
rect 706 463 719 497
rect 659 414 719 463
rect 659 380 672 414
rect 706 380 719 414
rect 659 368 719 380
rect 749 580 809 592
rect 749 546 762 580
rect 796 546 809 580
rect 749 510 809 546
rect 749 476 762 510
rect 796 476 809 510
rect 749 440 809 476
rect 749 406 762 440
rect 796 406 809 440
rect 749 368 809 406
rect 839 580 899 592
rect 839 546 852 580
rect 886 546 899 580
rect 839 497 899 546
rect 839 463 852 497
rect 886 463 899 497
rect 839 414 899 463
rect 839 380 852 414
rect 886 380 899 414
rect 839 368 899 380
rect 929 580 989 592
rect 929 546 942 580
rect 976 546 989 580
rect 929 510 989 546
rect 929 476 942 510
rect 976 476 989 510
rect 929 440 989 476
rect 929 406 942 440
rect 976 406 989 440
rect 929 368 989 406
rect 1019 580 1079 592
rect 1019 546 1032 580
rect 1066 546 1079 580
rect 1019 497 1079 546
rect 1019 463 1032 497
rect 1066 463 1079 497
rect 1019 414 1079 463
rect 1019 380 1032 414
rect 1066 380 1079 414
rect 1019 368 1079 380
rect 1109 580 1169 592
rect 1109 546 1122 580
rect 1156 546 1169 580
rect 1109 510 1169 546
rect 1109 476 1122 510
rect 1156 476 1169 510
rect 1109 440 1169 476
rect 1109 406 1122 440
rect 1156 406 1169 440
rect 1109 368 1169 406
rect 1199 580 1259 592
rect 1199 546 1212 580
rect 1246 546 1259 580
rect 1199 497 1259 546
rect 1199 463 1212 497
rect 1246 463 1259 497
rect 1199 414 1259 463
rect 1199 380 1212 414
rect 1246 380 1259 414
rect 1199 368 1259 380
rect 1289 580 1349 592
rect 1289 546 1302 580
rect 1336 546 1349 580
rect 1289 510 1349 546
rect 1289 476 1302 510
rect 1336 476 1349 510
rect 1289 440 1349 476
rect 1289 406 1302 440
rect 1336 406 1349 440
rect 1289 368 1349 406
rect 1379 580 1439 592
rect 1379 546 1392 580
rect 1426 546 1439 580
rect 1379 497 1439 546
rect 1379 463 1392 497
rect 1426 463 1439 497
rect 1379 414 1439 463
rect 1379 380 1392 414
rect 1426 380 1439 414
rect 1379 368 1439 380
rect 1469 580 1529 592
rect 1469 546 1482 580
rect 1516 546 1529 580
rect 1469 510 1529 546
rect 1469 476 1482 510
rect 1516 476 1529 510
rect 1469 440 1529 476
rect 1469 406 1482 440
rect 1516 406 1529 440
rect 1469 368 1529 406
rect 1559 580 1619 592
rect 1559 546 1572 580
rect 1606 546 1619 580
rect 1559 497 1619 546
rect 1559 463 1572 497
rect 1606 463 1619 497
rect 1559 414 1619 463
rect 1559 380 1572 414
rect 1606 380 1619 414
rect 1559 368 1619 380
rect 1649 580 1713 592
rect 1649 546 1662 580
rect 1696 546 1713 580
rect 1649 510 1713 546
rect 1649 476 1662 510
rect 1696 476 1713 510
rect 1649 440 1713 476
rect 1649 406 1662 440
rect 1696 406 1713 440
rect 1649 368 1713 406
rect 1743 580 1803 592
rect 1743 546 1756 580
rect 1790 546 1803 580
rect 1743 497 1803 546
rect 1743 463 1756 497
rect 1790 463 1803 497
rect 1743 414 1803 463
rect 1743 380 1756 414
rect 1790 380 1803 414
rect 1743 368 1803 380
rect 1833 580 1892 592
rect 1833 546 1846 580
rect 1880 546 1892 580
rect 1833 510 1892 546
rect 1833 476 1846 510
rect 1880 476 1892 510
rect 1833 440 1892 476
rect 1833 406 1846 440
rect 1880 406 1892 440
rect 1833 368 1892 406
<< ndiffc >>
rect 39 99 73 133
rect 125 99 159 133
rect 211 99 245 133
rect 301 99 335 133
rect 387 99 421 133
rect 487 99 521 133
rect 573 86 607 120
rect 659 99 693 133
rect 745 95 779 129
rect 831 99 865 133
rect 917 98 951 132
rect 1017 99 1051 133
rect 1103 86 1137 120
rect 1203 99 1237 133
rect 1289 86 1323 120
rect 1389 99 1423 133
rect 1475 86 1509 120
rect 1575 99 1609 133
rect 1661 86 1695 120
rect 1761 99 1795 133
rect 1847 99 1881 133
<< pdiffc >>
rect 40 546 74 580
rect 40 476 74 510
rect 40 406 74 440
rect 130 546 164 580
rect 130 476 164 510
rect 130 406 164 440
rect 220 546 254 580
rect 220 474 254 508
rect 310 546 344 580
rect 310 476 344 510
rect 310 406 344 440
rect 400 546 434 580
rect 400 474 434 508
rect 492 546 526 580
rect 492 463 526 497
rect 492 380 526 414
rect 582 546 616 580
rect 582 474 616 508
rect 582 406 616 440
rect 672 546 706 580
rect 672 463 706 497
rect 672 380 706 414
rect 762 546 796 580
rect 762 476 796 510
rect 762 406 796 440
rect 852 546 886 580
rect 852 463 886 497
rect 852 380 886 414
rect 942 546 976 580
rect 942 476 976 510
rect 942 406 976 440
rect 1032 546 1066 580
rect 1032 463 1066 497
rect 1032 380 1066 414
rect 1122 546 1156 580
rect 1122 476 1156 510
rect 1122 406 1156 440
rect 1212 546 1246 580
rect 1212 463 1246 497
rect 1212 380 1246 414
rect 1302 546 1336 580
rect 1302 476 1336 510
rect 1302 406 1336 440
rect 1392 546 1426 580
rect 1392 463 1426 497
rect 1392 380 1426 414
rect 1482 546 1516 580
rect 1482 476 1516 510
rect 1482 406 1516 440
rect 1572 546 1606 580
rect 1572 463 1606 497
rect 1572 380 1606 414
rect 1662 546 1696 580
rect 1662 476 1696 510
rect 1662 406 1696 440
rect 1756 546 1790 580
rect 1756 463 1790 497
rect 1756 380 1790 414
rect 1846 546 1880 580
rect 1846 476 1880 510
rect 1846 406 1880 440
<< poly >>
rect 87 592 117 618
rect 177 592 207 618
rect 267 592 297 618
rect 357 592 387 618
rect 449 592 479 618
rect 539 592 569 618
rect 629 592 659 618
rect 719 592 749 618
rect 809 592 839 618
rect 899 592 929 618
rect 989 592 1019 618
rect 1079 592 1109 618
rect 1169 592 1199 618
rect 1259 592 1289 618
rect 1349 592 1379 618
rect 1439 592 1469 618
rect 1529 592 1559 618
rect 1619 592 1649 618
rect 1713 592 1743 618
rect 1803 592 1833 618
rect 87 353 117 368
rect 177 353 207 368
rect 267 353 297 368
rect 357 353 387 368
rect 449 353 479 368
rect 539 353 569 368
rect 629 353 659 368
rect 719 353 749 368
rect 809 353 839 368
rect 899 353 929 368
rect 989 353 1019 368
rect 1079 353 1109 368
rect 1169 353 1199 368
rect 1259 353 1289 368
rect 1349 353 1379 368
rect 1439 353 1469 368
rect 1529 353 1559 368
rect 1619 353 1649 368
rect 1713 353 1743 368
rect 1803 353 1833 368
rect 84 336 120 353
rect 174 336 210 353
rect 264 336 300 353
rect 354 336 390 353
rect 84 320 390 336
rect 84 286 100 320
rect 134 286 168 320
rect 202 286 236 320
rect 270 286 304 320
rect 338 286 390 320
rect 84 270 390 286
rect 446 304 482 353
rect 536 304 572 353
rect 626 304 662 353
rect 716 304 752 353
rect 806 304 842 353
rect 896 304 932 353
rect 986 304 1022 353
rect 1076 304 1112 353
rect 1166 304 1202 353
rect 1256 304 1292 353
rect 1346 304 1382 353
rect 1436 304 1472 353
rect 1526 304 1562 353
rect 1616 304 1652 353
rect 1710 304 1746 353
rect 1800 304 1836 353
rect 446 288 1836 304
rect 84 158 114 270
rect 170 158 200 270
rect 260 158 290 270
rect 346 158 376 270
rect 446 254 578 288
rect 612 254 750 288
rect 784 254 918 288
rect 952 254 1101 288
rect 1135 254 1289 288
rect 1323 254 1475 288
rect 1509 254 1661 288
rect 1695 254 1836 288
rect 446 238 1836 254
rect 446 158 476 238
rect 532 158 562 238
rect 618 158 648 238
rect 704 158 734 238
rect 790 158 820 238
rect 876 158 906 238
rect 976 158 1006 238
rect 1062 158 1092 238
rect 1162 158 1192 238
rect 1248 158 1278 238
rect 1348 158 1378 238
rect 1434 158 1464 238
rect 1534 158 1564 238
rect 1620 158 1650 238
rect 1720 158 1750 238
rect 1806 158 1836 238
rect 84 48 114 74
rect 170 48 200 74
rect 260 48 290 74
rect 346 48 376 74
rect 446 48 476 74
rect 532 48 562 74
rect 618 48 648 74
rect 704 48 734 74
rect 790 48 820 74
rect 876 48 906 74
rect 976 48 1006 74
rect 1062 48 1092 74
rect 1162 48 1192 74
rect 1248 48 1278 74
rect 1348 48 1378 74
rect 1434 48 1464 74
rect 1534 48 1564 74
rect 1620 48 1650 74
rect 1720 48 1750 74
rect 1806 48 1836 74
<< polycont >>
rect 100 286 134 320
rect 168 286 202 320
rect 236 286 270 320
rect 304 286 338 320
rect 578 254 612 288
rect 750 254 784 288
rect 918 254 952 288
rect 1101 254 1135 288
rect 1289 254 1323 288
rect 1475 254 1509 288
rect 1661 254 1695 288
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 24 580 74 649
rect 24 546 40 580
rect 24 510 74 546
rect 24 476 40 510
rect 24 440 74 476
rect 24 406 40 440
rect 24 390 74 406
rect 114 580 180 596
rect 114 546 130 580
rect 164 546 180 580
rect 114 510 180 546
rect 114 476 130 510
rect 164 476 180 510
rect 114 440 180 476
rect 220 580 254 649
rect 220 508 254 546
rect 220 458 254 474
rect 294 580 360 596
rect 294 546 310 580
rect 344 546 360 580
rect 294 510 360 546
rect 294 476 310 510
rect 344 476 360 510
rect 114 406 130 440
rect 164 424 180 440
rect 294 440 360 476
rect 400 580 450 649
rect 434 546 450 580
rect 400 508 450 546
rect 434 474 450 508
rect 400 458 450 474
rect 486 580 532 596
rect 486 546 492 580
rect 526 546 532 580
rect 486 497 532 546
rect 486 463 492 497
rect 526 463 532 497
rect 294 424 310 440
rect 164 406 310 424
rect 344 424 360 440
rect 486 424 532 463
rect 344 406 427 424
rect 114 390 427 406
rect 25 320 359 356
rect 25 286 100 320
rect 134 286 168 320
rect 202 286 236 320
rect 270 286 304 320
rect 338 286 359 320
rect 25 270 359 286
rect 393 282 427 390
rect 478 380 492 424
rect 526 380 532 424
rect 566 580 632 649
rect 566 546 582 580
rect 616 546 632 580
rect 566 508 632 546
rect 566 474 582 508
rect 616 474 632 508
rect 566 440 632 474
rect 566 406 582 440
rect 616 406 632 440
rect 668 580 709 596
rect 668 546 672 580
rect 706 546 709 580
rect 668 497 709 546
rect 668 463 672 497
rect 706 463 709 497
rect 668 424 709 463
rect 393 276 442 282
rect 393 242 402 276
rect 436 242 442 276
rect 393 236 442 242
rect 393 230 427 236
rect 109 196 427 230
rect 23 133 73 162
rect 23 99 39 133
rect 23 17 73 99
rect 109 133 159 196
rect 109 99 125 133
rect 109 70 159 99
rect 195 133 245 162
rect 195 99 211 133
rect 195 17 245 99
rect 285 133 335 196
rect 285 99 301 133
rect 285 70 335 99
rect 371 133 437 162
rect 371 99 387 133
rect 421 99 437 133
rect 371 17 437 99
rect 478 133 532 380
rect 668 380 672 424
rect 706 380 709 424
rect 746 580 812 649
rect 746 546 762 580
rect 796 546 812 580
rect 746 510 812 546
rect 746 476 762 510
rect 796 476 812 510
rect 746 440 812 476
rect 746 406 762 440
rect 796 406 812 440
rect 846 580 886 596
rect 846 546 852 580
rect 846 497 886 546
rect 846 463 852 497
rect 846 424 886 463
rect 668 372 709 380
rect 846 390 849 424
rect 883 414 886 424
rect 926 580 992 649
rect 926 546 942 580
rect 976 546 992 580
rect 926 510 992 546
rect 926 476 942 510
rect 976 476 992 510
rect 926 440 992 476
rect 926 406 942 440
rect 976 406 992 440
rect 1028 580 1070 596
rect 1028 546 1032 580
rect 1066 546 1070 580
rect 1028 497 1070 546
rect 1028 463 1032 497
rect 1066 463 1070 497
rect 1028 424 1070 463
rect 846 380 852 390
rect 846 372 886 380
rect 1028 380 1032 424
rect 1066 380 1070 424
rect 1106 580 1172 649
rect 1106 546 1122 580
rect 1156 546 1172 580
rect 1106 510 1172 546
rect 1106 476 1122 510
rect 1156 476 1172 510
rect 1106 440 1172 476
rect 1106 406 1122 440
rect 1156 406 1172 440
rect 1208 580 1249 596
rect 1208 546 1212 580
rect 1246 546 1249 580
rect 1208 497 1249 546
rect 1208 463 1212 497
rect 1246 463 1249 497
rect 1208 424 1249 463
rect 1028 372 1070 380
rect 1208 380 1212 424
rect 1246 380 1249 424
rect 1286 580 1352 649
rect 1286 546 1302 580
rect 1336 546 1352 580
rect 1286 510 1352 546
rect 1286 476 1302 510
rect 1336 476 1352 510
rect 1286 440 1352 476
rect 1286 406 1302 440
rect 1336 406 1352 440
rect 1389 580 1430 596
rect 1389 546 1392 580
rect 1426 546 1430 580
rect 1389 497 1430 546
rect 1389 463 1392 497
rect 1426 463 1430 497
rect 1389 424 1430 463
rect 1208 372 1249 380
rect 1389 380 1392 424
rect 1426 380 1430 424
rect 1466 580 1532 649
rect 1466 546 1482 580
rect 1516 546 1532 580
rect 1466 510 1532 546
rect 1466 476 1482 510
rect 1516 476 1532 510
rect 1466 440 1532 476
rect 1466 406 1482 440
rect 1516 406 1532 440
rect 1568 580 1610 596
rect 1568 546 1572 580
rect 1606 546 1610 580
rect 1568 497 1610 546
rect 1568 463 1572 497
rect 1606 463 1610 497
rect 1568 424 1610 463
rect 1389 372 1430 380
rect 1568 380 1572 424
rect 1606 380 1610 424
rect 1646 580 1712 649
rect 1646 546 1662 580
rect 1696 546 1712 580
rect 1646 510 1712 546
rect 1646 476 1662 510
rect 1696 476 1712 510
rect 1646 440 1712 476
rect 1646 406 1662 440
rect 1696 406 1712 440
rect 1750 580 1794 596
rect 1750 546 1756 580
rect 1790 546 1794 580
rect 1750 497 1794 546
rect 1750 463 1756 497
rect 1790 463 1794 497
rect 1750 424 1794 463
rect 1568 372 1610 380
rect 1750 380 1756 424
rect 1790 380 1794 424
rect 1830 580 1896 649
rect 1830 546 1846 580
rect 1880 546 1896 580
rect 1830 510 1896 546
rect 1830 476 1846 510
rect 1880 476 1896 510
rect 1830 440 1896 476
rect 1830 406 1846 440
rect 1880 406 1896 440
rect 1750 372 1794 380
rect 655 338 709 372
rect 834 338 886 372
rect 1005 338 1070 372
rect 1187 338 1249 372
rect 1373 338 1430 372
rect 1559 338 1610 372
rect 1745 366 1794 372
rect 567 288 621 304
rect 567 242 578 288
rect 612 242 621 288
rect 567 238 621 242
rect 478 99 487 133
rect 521 99 532 133
rect 478 70 532 99
rect 573 120 607 136
rect 573 17 607 86
rect 655 133 700 338
rect 734 288 800 304
rect 734 242 750 288
rect 784 242 800 288
rect 734 238 800 242
rect 834 149 868 338
rect 902 288 968 304
rect 902 242 918 288
rect 952 242 968 288
rect 902 238 968 242
rect 655 99 659 133
rect 693 99 700 133
rect 655 70 700 99
rect 734 129 779 145
rect 734 95 745 129
rect 734 17 779 95
rect 815 133 868 149
rect 815 99 831 133
rect 865 99 868 133
rect 815 70 868 99
rect 902 132 967 148
rect 902 98 917 132
rect 951 98 967 132
rect 902 17 967 98
rect 1005 133 1051 338
rect 1085 288 1151 304
rect 1085 242 1101 288
rect 1135 242 1151 288
rect 1085 238 1151 242
rect 1005 99 1017 133
rect 1005 70 1051 99
rect 1087 120 1153 136
rect 1087 86 1103 120
rect 1137 86 1153 120
rect 1087 17 1153 86
rect 1187 133 1237 338
rect 1273 288 1339 304
rect 1273 242 1289 288
rect 1323 242 1339 288
rect 1273 238 1339 242
rect 1187 99 1203 133
rect 1187 70 1237 99
rect 1273 120 1339 136
rect 1273 86 1289 120
rect 1323 86 1339 120
rect 1273 17 1339 86
rect 1373 133 1423 338
rect 1459 288 1525 304
rect 1459 242 1475 288
rect 1509 242 1525 288
rect 1459 238 1525 242
rect 1373 99 1389 133
rect 1373 70 1423 99
rect 1459 120 1525 136
rect 1459 86 1475 120
rect 1509 86 1525 120
rect 1459 17 1525 86
rect 1559 133 1609 338
rect 1645 288 1711 304
rect 1645 242 1661 288
rect 1695 242 1711 288
rect 1645 238 1711 242
rect 1559 99 1575 133
rect 1559 70 1609 99
rect 1645 120 1711 136
rect 1645 86 1661 120
rect 1695 86 1711 120
rect 1645 17 1711 86
rect 1745 133 1795 366
rect 1745 99 1761 133
rect 1745 70 1795 99
rect 1831 133 1897 149
rect 1831 99 1847 133
rect 1881 99 1897 133
rect 1831 17 1897 99
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 492 414 526 424
rect 492 390 526 414
rect 402 242 436 276
rect 672 414 706 424
rect 672 390 706 414
rect 849 414 883 424
rect 849 390 852 414
rect 852 390 883 414
rect 1032 414 1066 424
rect 1032 390 1066 414
rect 1212 414 1246 424
rect 1212 390 1246 414
rect 1392 414 1426 424
rect 1392 390 1426 414
rect 1572 414 1606 424
rect 1572 390 1606 414
rect 1756 414 1790 424
rect 1756 390 1790 414
rect 578 254 612 276
rect 578 242 612 254
rect 750 254 784 276
rect 750 242 784 254
rect 918 254 952 276
rect 918 242 952 254
rect 1101 254 1135 276
rect 1101 242 1135 254
rect 1289 254 1323 276
rect 1289 242 1323 254
rect 1475 254 1509 276
rect 1475 242 1509 254
rect 1661 254 1695 276
rect 1661 242 1695 254
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
<< metal1 >>
rect 0 683 1920 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 0 617 1920 649
rect 478 424 1818 430
rect 478 390 492 424
rect 526 390 672 424
rect 706 390 849 424
rect 883 390 1032 424
rect 1066 390 1212 424
rect 1246 390 1392 424
rect 1426 390 1572 424
rect 1606 390 1756 424
rect 1790 390 1818 424
rect 478 384 1818 390
rect 388 276 1728 282
rect 388 242 402 276
rect 436 242 578 276
rect 612 242 750 276
rect 784 242 918 276
rect 952 242 1101 276
rect 1135 242 1289 276
rect 1323 242 1475 276
rect 1509 242 1661 276
rect 1695 242 1728 276
rect 388 236 1728 242
rect 0 17 1920 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
rect 0 -49 1920 -17
<< labels >>
rlabel comment s 0 0 0 0 4 clkbuf_16
flabel pwell s 0 0 1920 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew
flabel nwell s 0 617 1920 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew
flabel metal1 s 0 617 1920 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew
flabel metal1 s 0 0 1920 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew
flabel metal1 s 478 384 1818 430 0 FreeSans 400 0 0 0 X
port 6 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 1920 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3328040
string GDS_START 3312114
<< end >>
