magic
tech sky130A
magscale 1 2
timestamp 1599588238
<< locali >>
rect 106 294 172 360
rect 329 236 364 547
rect 409 270 551 356
rect 601 236 647 282
rect 329 202 647 236
rect 329 192 549 202
rect 297 70 363 192
rect 499 70 549 192
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 22 260 72 596
rect 112 394 178 649
rect 224 581 470 615
rect 224 364 290 581
rect 229 260 295 310
rect 22 226 295 260
rect 404 424 470 581
rect 510 458 560 649
rect 600 424 650 596
rect 404 390 650 424
rect 600 364 650 390
rect 22 90 156 226
rect 197 17 263 192
rect 397 17 463 158
rect 583 17 649 168
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel locali s 409 270 551 356 6 A
port 1 nsew signal input
rlabel locali s 106 294 172 360 6 B_N
port 2 nsew signal input
rlabel locali s 601 236 647 282 6 Y
port 3 nsew signal output
rlabel locali s 499 70 549 192 6 Y
port 3 nsew signal output
rlabel locali s 329 236 364 547 6 Y
port 3 nsew signal output
rlabel locali s 329 202 647 236 6 Y
port 3 nsew signal output
rlabel locali s 329 192 549 202 6 Y
port 3 nsew signal output
rlabel locali s 297 70 363 192 6 Y
port 3 nsew signal output
rlabel metal1 s 0 -49 672 49 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 617 672 715 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1931412
string GDS_START 1925004
<< end >>
