magic
tech sky130A
magscale 1 2
timestamp 1599588218
<< nwell >>
rect -38 332 806 704
<< pwell >>
rect 0 0 768 49
<< scpmos >>
rect 86 392 122 592
rect 182 392 218 592
rect 272 392 308 592
rect 533 368 569 536
rect 640 368 676 592
<< nmoslvt >>
rect 92 136 122 264
rect 164 136 194 264
rect 272 136 302 264
rect 539 74 569 184
rect 634 74 664 222
<< ndiff >>
rect 39 235 92 264
rect 39 201 47 235
rect 81 201 92 235
rect 39 136 92 201
rect 122 136 164 264
rect 194 252 272 264
rect 194 218 209 252
rect 243 218 272 252
rect 194 178 272 218
rect 194 144 209 178
rect 243 144 272 178
rect 194 136 272 144
rect 302 184 355 264
rect 584 184 634 222
rect 302 150 313 184
rect 347 150 355 184
rect 302 136 355 150
rect 482 146 539 184
rect 482 112 494 146
rect 528 112 539 146
rect 482 74 539 112
rect 569 150 634 184
rect 569 116 584 150
rect 618 116 634 150
rect 569 74 634 116
rect 664 210 717 222
rect 664 176 675 210
rect 709 176 717 210
rect 664 120 717 176
rect 664 86 675 120
rect 709 86 717 120
rect 664 74 717 86
<< pdiff >>
rect 34 580 86 592
rect 34 546 42 580
rect 76 546 86 580
rect 34 509 86 546
rect 34 475 42 509
rect 76 475 86 509
rect 34 438 86 475
rect 34 404 42 438
rect 76 404 86 438
rect 34 392 86 404
rect 122 580 182 592
rect 122 546 135 580
rect 169 546 182 580
rect 122 508 182 546
rect 122 474 135 508
rect 169 474 182 508
rect 122 392 182 474
rect 218 580 272 592
rect 218 546 228 580
rect 262 546 272 580
rect 218 510 272 546
rect 218 476 228 510
rect 262 476 272 510
rect 218 440 272 476
rect 218 406 228 440
rect 262 406 272 440
rect 218 392 272 406
rect 308 580 360 592
rect 308 546 318 580
rect 352 546 360 580
rect 584 566 640 592
rect 308 509 360 546
rect 584 536 596 566
rect 308 475 318 509
rect 352 475 360 509
rect 308 438 360 475
rect 308 404 318 438
rect 352 404 360 438
rect 308 392 360 404
rect 481 414 533 536
rect 481 380 489 414
rect 523 380 533 414
rect 481 368 533 380
rect 569 532 596 536
rect 630 532 640 566
rect 569 368 640 532
rect 676 580 728 592
rect 676 546 686 580
rect 720 546 728 580
rect 676 497 728 546
rect 676 463 686 497
rect 720 463 728 497
rect 676 414 728 463
rect 676 380 686 414
rect 720 380 728 414
rect 676 368 728 380
<< ndiffc >>
rect 47 201 81 235
rect 209 218 243 252
rect 209 144 243 178
rect 313 150 347 184
rect 494 112 528 146
rect 584 116 618 150
rect 675 176 709 210
rect 675 86 709 120
<< pdiffc >>
rect 42 546 76 580
rect 42 475 76 509
rect 42 404 76 438
rect 135 546 169 580
rect 135 474 169 508
rect 228 546 262 580
rect 228 476 262 510
rect 228 406 262 440
rect 318 546 352 580
rect 318 475 352 509
rect 318 404 352 438
rect 489 380 523 414
rect 596 532 630 566
rect 686 546 720 580
rect 686 463 720 497
rect 686 380 720 414
<< poly >>
rect 86 592 122 618
rect 182 592 218 618
rect 272 592 308 618
rect 640 592 676 618
rect 533 536 569 562
rect 86 279 122 392
rect 182 356 218 392
rect 92 264 122 279
rect 164 340 230 356
rect 164 306 180 340
rect 214 306 230 340
rect 164 290 230 306
rect 272 309 308 392
rect 383 338 449 354
rect 383 309 399 338
rect 272 304 399 309
rect 433 304 449 338
rect 533 310 569 368
rect 640 330 676 368
rect 164 264 194 290
rect 272 279 449 304
rect 272 264 302 279
rect 383 270 449 279
rect 383 236 399 270
rect 433 236 449 270
rect 503 294 569 310
rect 503 260 519 294
rect 553 260 569 294
rect 617 314 683 330
rect 617 280 633 314
rect 667 280 683 314
rect 617 264 683 280
rect 503 244 569 260
rect 383 220 449 236
rect 539 184 569 244
rect 634 222 664 264
rect 92 114 122 136
rect 21 98 122 114
rect 164 110 194 136
rect 272 110 302 136
rect 21 64 37 98
rect 71 64 122 98
rect 21 48 122 64
rect 539 48 569 74
rect 634 48 664 74
<< polycont >>
rect 180 306 214 340
rect 399 304 433 338
rect 399 236 433 270
rect 519 260 553 294
rect 633 280 667 314
rect 37 64 71 98
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 26 580 92 596
rect 26 546 42 580
rect 76 546 92 580
rect 26 509 92 546
rect 26 475 42 509
rect 76 475 92 509
rect 26 438 92 475
rect 132 580 172 649
rect 132 546 135 580
rect 169 546 172 580
rect 132 508 172 546
rect 132 474 135 508
rect 169 474 172 508
rect 132 458 172 474
rect 212 580 278 596
rect 212 546 228 580
rect 262 546 278 580
rect 212 510 278 546
rect 212 476 228 510
rect 262 476 278 510
rect 26 404 42 438
rect 76 424 92 438
rect 212 440 278 476
rect 212 424 228 440
rect 76 406 228 424
rect 262 406 278 440
rect 76 404 278 406
rect 26 390 278 404
rect 315 580 352 596
rect 315 546 318 580
rect 315 509 352 546
rect 580 566 646 649
rect 580 532 596 566
rect 630 532 646 566
rect 580 516 646 532
rect 686 580 751 596
rect 720 546 751 580
rect 315 475 318 509
rect 686 497 751 546
rect 352 475 651 482
rect 315 448 651 475
rect 315 438 352 448
rect 315 404 318 438
rect 26 388 92 390
rect 315 388 352 404
rect 131 340 263 356
rect 131 306 180 340
rect 214 306 263 340
rect 131 290 263 306
rect 31 235 97 268
rect 315 256 349 388
rect 415 380 489 414
rect 523 380 539 414
rect 415 364 539 380
rect 415 354 449 364
rect 31 201 47 235
rect 81 219 97 235
rect 189 252 349 256
rect 81 201 155 219
rect 31 168 155 201
rect 21 98 87 134
rect 21 64 37 98
rect 71 64 87 98
rect 21 51 87 64
rect 121 17 155 168
rect 189 218 209 252
rect 243 222 349 252
rect 383 338 449 354
rect 383 304 399 338
rect 433 304 449 338
rect 617 330 651 448
rect 720 463 751 497
rect 686 414 751 463
rect 720 380 751 414
rect 686 364 751 380
rect 617 314 683 330
rect 383 270 449 304
rect 383 236 399 270
rect 433 236 449 270
rect 503 294 569 310
rect 503 260 519 294
rect 553 260 569 294
rect 617 280 633 314
rect 667 280 683 314
rect 617 264 683 280
rect 503 236 569 260
rect 243 218 263 222
rect 383 220 449 236
rect 717 226 751 364
rect 189 178 263 218
rect 415 188 449 220
rect 659 210 751 226
rect 189 144 209 178
rect 243 144 263 178
rect 189 132 263 144
rect 297 184 363 186
rect 297 150 313 184
rect 347 150 363 184
rect 297 17 363 150
rect 415 146 544 188
rect 415 112 494 146
rect 528 112 544 146
rect 415 70 544 112
rect 580 150 623 179
rect 580 116 584 150
rect 618 116 623 150
rect 580 17 623 116
rect 659 176 675 210
rect 709 176 751 210
rect 659 120 751 176
rect 659 86 675 120
rect 709 86 751 120
rect 659 70 751 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
rlabel comment s 0 0 0 0 4 a21bo_1
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 703 390 737 424 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 703 464 737 498 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 703 538 737 572 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 511 242 545 276 0 FreeSans 340 0 0 0 B1_N
port 3 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 31 94 65 128 0 FreeSans 340 0 0 0 A2
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 768 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3939132
string GDS_START 3932040
<< end >>
