magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 17 425 276 483
rect 111 265 176 323
rect 466 299 531 493
rect 17 199 77 265
rect 111 199 316 265
rect 494 152 531 299
rect 466 83 531 152
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 21 357 274 391
rect 320 367 414 527
rect 21 299 77 357
rect 240 333 274 357
rect 240 299 422 333
rect 378 265 422 299
rect 378 199 460 265
rect 378 165 422 199
rect 21 131 422 165
rect 565 286 623 527
rect 21 61 72 131
rect 106 17 182 97
rect 226 61 260 131
rect 294 17 418 97
rect 565 17 623 183
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 111 265 176 323 6 A
port 1 nsew signal input
rlabel locali s 111 199 316 265 6 A
port 1 nsew signal input
rlabel locali s 17 425 276 483 6 B
port 2 nsew signal input
rlabel locali s 17 199 77 265 6 C
port 3 nsew signal input
rlabel locali s 494 152 531 299 6 X
port 4 nsew signal output
rlabel locali s 466 299 531 493 6 X
port 4 nsew signal output
rlabel locali s 466 83 531 152 6 X
port 4 nsew signal output
rlabel metal1 s 0 -48 644 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 465000
string GDS_START 458956
<< end >>
