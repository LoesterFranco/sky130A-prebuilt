magic
tech sky130A
magscale 1 2
timestamp 1604502701
<< nwell >>
rect -38 332 1670 704
<< pwell >>
rect 0 0 1632 49
<< scpmos >>
rect 89 368 119 592
rect 179 368 209 592
rect 269 368 299 592
rect 359 368 389 592
rect 459 368 489 592
rect 549 368 579 592
rect 639 368 669 592
rect 739 368 769 592
rect 951 368 981 592
rect 1059 368 1089 592
rect 1161 368 1191 592
rect 1251 368 1281 592
<< nmoslvt >>
rect 84 74 114 222
rect 184 74 214 222
rect 270 74 300 222
rect 370 74 400 222
rect 456 74 486 222
rect 542 74 572 222
rect 628 74 658 222
rect 718 74 748 222
rect 804 74 834 222
rect 890 74 920 222
rect 976 74 1006 222
rect 1062 74 1092 222
rect 1260 84 1290 232
rect 1346 84 1376 232
rect 1432 84 1462 232
rect 1518 84 1548 232
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 136 184 222
rect 114 102 139 136
rect 173 102 184 136
rect 114 74 184 102
rect 214 210 270 222
rect 214 176 225 210
rect 259 176 270 210
rect 214 120 270 176
rect 214 86 225 120
rect 259 86 270 120
rect 214 74 270 86
rect 300 144 370 222
rect 300 110 325 144
rect 359 110 370 144
rect 300 74 370 110
rect 400 210 456 222
rect 400 176 411 210
rect 445 176 456 210
rect 400 120 456 176
rect 400 86 411 120
rect 445 86 456 120
rect 400 74 456 86
rect 486 144 542 222
rect 486 110 497 144
rect 531 110 542 144
rect 486 74 542 110
rect 572 210 628 222
rect 572 176 583 210
rect 617 176 628 210
rect 572 120 628 176
rect 572 86 583 120
rect 617 86 628 120
rect 572 74 628 86
rect 658 144 718 222
rect 658 110 669 144
rect 703 110 718 144
rect 658 74 718 110
rect 748 210 804 222
rect 748 176 759 210
rect 793 176 804 210
rect 748 120 804 176
rect 748 86 759 120
rect 793 86 804 120
rect 748 74 804 86
rect 834 120 890 222
rect 834 86 845 120
rect 879 86 890 120
rect 834 74 890 86
rect 920 207 976 222
rect 920 173 931 207
rect 965 173 976 207
rect 920 74 976 173
rect 1006 136 1062 222
rect 1006 102 1017 136
rect 1051 102 1062 136
rect 1006 74 1062 102
rect 1092 189 1149 222
rect 1092 155 1103 189
rect 1137 155 1149 189
rect 1092 74 1149 155
rect 1203 220 1260 232
rect 1203 186 1215 220
rect 1249 186 1260 220
rect 1203 130 1260 186
rect 1203 96 1215 130
rect 1249 96 1260 130
rect 1203 84 1260 96
rect 1290 194 1346 232
rect 1290 160 1301 194
rect 1335 160 1346 194
rect 1290 84 1346 160
rect 1376 149 1432 232
rect 1376 115 1387 149
rect 1421 115 1432 149
rect 1376 84 1432 115
rect 1462 194 1518 232
rect 1462 160 1473 194
rect 1507 160 1518 194
rect 1462 84 1518 160
rect 1548 220 1605 232
rect 1548 186 1559 220
rect 1593 186 1605 220
rect 1548 130 1605 186
rect 1548 96 1559 130
rect 1593 96 1605 130
rect 1548 84 1605 96
<< pdiff >>
rect 30 580 89 592
rect 30 546 42 580
rect 76 546 89 580
rect 30 510 89 546
rect 30 476 42 510
rect 76 476 89 510
rect 30 440 89 476
rect 30 406 42 440
rect 76 406 89 440
rect 30 368 89 406
rect 119 580 179 592
rect 119 546 132 580
rect 166 546 179 580
rect 119 508 179 546
rect 119 474 132 508
rect 166 474 179 508
rect 119 368 179 474
rect 209 580 269 592
rect 209 546 222 580
rect 256 546 269 580
rect 209 510 269 546
rect 209 476 222 510
rect 256 476 269 510
rect 209 440 269 476
rect 209 406 222 440
rect 256 406 269 440
rect 209 368 269 406
rect 299 580 359 592
rect 299 546 312 580
rect 346 546 359 580
rect 299 508 359 546
rect 299 474 312 508
rect 346 474 359 508
rect 299 368 359 474
rect 389 580 459 592
rect 389 546 402 580
rect 436 546 459 580
rect 389 510 459 546
rect 389 476 402 510
rect 436 476 459 510
rect 389 440 459 476
rect 389 406 402 440
rect 436 406 459 440
rect 389 368 459 406
rect 489 531 549 592
rect 489 497 502 531
rect 536 497 549 531
rect 489 440 549 497
rect 489 406 502 440
rect 536 406 549 440
rect 489 368 549 406
rect 579 580 639 592
rect 579 546 592 580
rect 626 546 639 580
rect 579 508 639 546
rect 579 474 592 508
rect 626 474 639 508
rect 579 368 639 474
rect 669 531 739 592
rect 669 497 692 531
rect 726 497 739 531
rect 669 440 739 497
rect 669 406 692 440
rect 726 406 739 440
rect 669 368 739 406
rect 769 580 838 592
rect 769 546 792 580
rect 826 546 838 580
rect 769 492 838 546
rect 769 458 792 492
rect 826 458 838 492
rect 769 368 838 458
rect 892 580 951 592
rect 892 546 904 580
rect 938 546 951 580
rect 892 492 951 546
rect 892 458 904 492
rect 938 458 951 492
rect 892 368 951 458
rect 981 580 1059 592
rect 981 546 1004 580
rect 1038 546 1059 580
rect 981 510 1059 546
rect 981 476 1004 510
rect 1038 476 1059 510
rect 981 440 1059 476
rect 981 406 1004 440
rect 1038 406 1059 440
rect 981 368 1059 406
rect 1089 580 1161 592
rect 1089 546 1104 580
rect 1138 546 1161 580
rect 1089 492 1161 546
rect 1089 458 1104 492
rect 1138 458 1161 492
rect 1089 368 1161 458
rect 1191 580 1251 592
rect 1191 546 1204 580
rect 1238 546 1251 580
rect 1191 510 1251 546
rect 1191 476 1204 510
rect 1238 476 1251 510
rect 1191 440 1251 476
rect 1191 406 1204 440
rect 1238 406 1251 440
rect 1191 368 1251 406
rect 1281 580 1454 592
rect 1281 546 1294 580
rect 1328 546 1408 580
rect 1442 546 1454 580
rect 1281 508 1454 546
rect 1281 474 1294 508
rect 1328 474 1408 508
rect 1442 474 1454 508
rect 1281 368 1454 474
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 139 102 173 136
rect 225 176 259 210
rect 225 86 259 120
rect 325 110 359 144
rect 411 176 445 210
rect 411 86 445 120
rect 497 110 531 144
rect 583 176 617 210
rect 583 86 617 120
rect 669 110 703 144
rect 759 176 793 210
rect 759 86 793 120
rect 845 86 879 120
rect 931 173 965 207
rect 1017 102 1051 136
rect 1103 155 1137 189
rect 1215 186 1249 220
rect 1215 96 1249 130
rect 1301 160 1335 194
rect 1387 115 1421 149
rect 1473 160 1507 194
rect 1559 186 1593 220
rect 1559 96 1593 130
<< pdiffc >>
rect 42 546 76 580
rect 42 476 76 510
rect 42 406 76 440
rect 132 546 166 580
rect 132 474 166 508
rect 222 546 256 580
rect 222 476 256 510
rect 222 406 256 440
rect 312 546 346 580
rect 312 474 346 508
rect 402 546 436 580
rect 402 476 436 510
rect 402 406 436 440
rect 502 497 536 531
rect 502 406 536 440
rect 592 546 626 580
rect 592 474 626 508
rect 692 497 726 531
rect 692 406 726 440
rect 792 546 826 580
rect 792 458 826 492
rect 904 546 938 580
rect 904 458 938 492
rect 1004 546 1038 580
rect 1004 476 1038 510
rect 1004 406 1038 440
rect 1104 546 1138 580
rect 1104 458 1138 492
rect 1204 546 1238 580
rect 1204 476 1238 510
rect 1204 406 1238 440
rect 1294 546 1328 580
rect 1408 546 1442 580
rect 1294 474 1328 508
rect 1408 474 1442 508
<< poly >>
rect 89 592 119 618
rect 179 592 209 618
rect 269 592 299 618
rect 359 592 389 618
rect 459 592 489 618
rect 549 592 579 618
rect 639 592 669 618
rect 739 592 769 618
rect 951 592 981 618
rect 1059 592 1089 618
rect 1161 592 1191 618
rect 1251 592 1281 618
rect 89 353 119 368
rect 179 353 209 368
rect 269 353 299 368
rect 359 353 389 368
rect 459 353 489 368
rect 549 353 579 368
rect 639 353 669 368
rect 739 353 769 368
rect 951 353 981 368
rect 1059 353 1089 368
rect 1161 353 1191 368
rect 1251 353 1281 368
rect 86 336 122 353
rect 176 336 212 353
rect 266 336 302 353
rect 356 336 392 353
rect 456 345 492 353
rect 546 345 582 353
rect 636 345 672 353
rect 736 345 772 353
rect 84 320 400 336
rect 84 286 100 320
rect 134 286 168 320
rect 202 286 236 320
rect 270 286 304 320
rect 338 286 400 320
rect 84 270 400 286
rect 84 222 114 270
rect 184 222 214 270
rect 270 222 300 270
rect 370 222 400 270
rect 456 320 772 345
rect 948 336 984 353
rect 1056 336 1092 353
rect 456 286 472 320
rect 506 286 540 320
rect 574 286 608 320
rect 642 286 676 320
rect 710 315 772 320
rect 890 320 1092 336
rect 710 286 750 315
rect 456 270 750 286
rect 890 286 906 320
rect 940 286 974 320
rect 1008 286 1042 320
rect 1076 286 1092 320
rect 890 270 1092 286
rect 1158 336 1194 353
rect 1248 336 1284 353
rect 1158 320 1376 336
rect 1158 286 1190 320
rect 1224 286 1258 320
rect 1292 286 1326 320
rect 1360 300 1376 320
rect 1360 286 1548 300
rect 1158 270 1548 286
rect 456 222 486 270
rect 542 222 572 270
rect 628 222 658 270
rect 718 222 748 270
rect 890 267 920 270
rect 804 237 920 267
rect 804 222 834 237
rect 890 222 920 237
rect 976 222 1006 270
rect 1062 222 1092 270
rect 1260 232 1290 270
rect 1346 232 1376 270
rect 1432 232 1462 270
rect 1518 232 1548 270
rect 84 48 114 74
rect 184 48 214 74
rect 270 48 300 74
rect 370 48 400 74
rect 456 48 486 74
rect 542 48 572 74
rect 628 48 658 74
rect 718 48 748 74
rect 804 48 834 74
rect 890 48 920 74
rect 976 48 1006 74
rect 1062 48 1092 74
rect 1260 58 1290 84
rect 1346 58 1376 84
rect 1432 58 1462 84
rect 1518 58 1548 84
<< polycont >>
rect 100 286 134 320
rect 168 286 202 320
rect 236 286 270 320
rect 304 286 338 320
rect 472 286 506 320
rect 540 286 574 320
rect 608 286 642 320
rect 676 286 710 320
rect 906 286 940 320
rect 974 286 1008 320
rect 1042 286 1076 320
rect 1190 286 1224 320
rect 1258 286 1292 320
rect 1326 286 1360 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 26 580 92 596
rect 26 546 42 580
rect 76 546 92 580
rect 26 510 92 546
rect 26 476 42 510
rect 76 476 92 510
rect 26 440 92 476
rect 132 580 166 649
rect 132 508 166 546
rect 132 458 166 474
rect 206 580 272 596
rect 206 546 222 580
rect 256 546 272 580
rect 206 510 272 546
rect 206 476 222 510
rect 256 476 272 510
rect 26 406 42 440
rect 76 424 92 440
rect 206 440 272 476
rect 312 580 346 649
rect 312 508 346 546
rect 312 458 346 474
rect 386 581 842 615
rect 386 580 452 581
rect 386 546 402 580
rect 436 546 452 580
rect 592 580 642 581
rect 386 510 452 546
rect 386 476 402 510
rect 436 476 452 510
rect 206 424 222 440
rect 76 406 222 424
rect 256 424 272 440
rect 386 440 452 476
rect 386 424 402 440
rect 256 406 402 424
rect 436 406 452 440
rect 26 390 452 406
rect 486 531 552 547
rect 486 497 502 531
rect 536 497 552 531
rect 486 440 552 497
rect 626 546 642 580
rect 776 580 842 581
rect 592 508 642 546
rect 626 474 642 508
rect 592 458 642 474
rect 676 531 742 547
rect 676 497 692 531
rect 726 497 742 531
rect 486 406 502 440
rect 536 424 552 440
rect 676 440 742 497
rect 776 546 792 580
rect 826 546 842 580
rect 776 492 842 546
rect 776 458 792 492
rect 826 458 842 492
rect 888 580 954 649
rect 888 546 904 580
rect 938 546 954 580
rect 888 492 954 546
rect 888 458 904 492
rect 938 458 954 492
rect 988 580 1054 596
rect 988 546 1004 580
rect 1038 546 1054 580
rect 988 510 1054 546
rect 988 476 1004 510
rect 1038 476 1054 510
rect 676 424 692 440
rect 536 406 692 424
rect 726 424 742 440
rect 988 440 1054 476
rect 1088 580 1154 649
rect 1088 546 1104 580
rect 1138 546 1154 580
rect 1088 492 1154 546
rect 1088 458 1104 492
rect 1138 458 1154 492
rect 1188 580 1254 596
rect 1188 546 1204 580
rect 1238 546 1254 580
rect 1188 510 1254 546
rect 1188 476 1204 510
rect 1238 476 1254 510
rect 988 424 1004 440
rect 726 406 1004 424
rect 1038 424 1054 440
rect 1188 440 1254 476
rect 1288 580 1458 649
rect 1288 546 1294 580
rect 1328 546 1408 580
rect 1442 546 1458 580
rect 1288 508 1458 546
rect 1288 474 1294 508
rect 1328 474 1408 508
rect 1442 474 1458 508
rect 1288 458 1458 474
rect 1188 424 1204 440
rect 1038 406 1204 424
rect 1238 424 1254 440
rect 1509 424 1607 578
rect 1238 406 1607 424
rect 486 390 1607 406
rect 25 320 359 356
rect 25 286 100 320
rect 134 286 168 320
rect 202 286 236 320
rect 270 286 304 320
rect 338 286 359 320
rect 25 270 359 286
rect 409 320 839 356
rect 409 286 472 320
rect 506 286 540 320
rect 574 286 608 320
rect 642 286 676 320
rect 710 286 839 320
rect 409 270 839 286
rect 889 320 1127 356
rect 889 286 906 320
rect 940 286 974 320
rect 1008 286 1042 320
rect 1076 286 1127 320
rect 889 270 1127 286
rect 1174 320 1415 356
rect 1174 286 1190 320
rect 1224 286 1258 320
rect 1292 286 1326 320
rect 1360 286 1415 320
rect 1174 270 1415 286
rect 1473 310 1607 390
rect 1473 236 1509 310
rect 23 210 1153 236
rect 23 176 39 210
rect 73 202 225 210
rect 73 176 89 202
rect 23 120 89 176
rect 259 202 411 210
rect 259 176 275 202
rect 23 86 39 120
rect 73 86 89 120
rect 23 70 89 86
rect 123 136 189 168
rect 123 102 139 136
rect 173 102 189 136
rect 123 17 189 102
rect 225 120 275 176
rect 445 202 583 210
rect 259 86 275 120
rect 225 70 275 86
rect 309 144 375 168
rect 309 110 325 144
rect 359 110 375 144
rect 309 17 375 110
rect 411 120 445 176
rect 617 202 759 210
rect 411 70 445 86
rect 481 144 547 168
rect 481 110 497 144
rect 531 110 547 144
rect 481 17 547 110
rect 583 120 617 176
rect 793 207 1153 210
rect 793 176 931 207
rect 759 173 931 176
rect 965 202 1153 207
rect 965 173 981 202
rect 583 70 617 86
rect 653 144 719 168
rect 653 110 669 144
rect 703 110 719 144
rect 653 17 719 110
rect 759 164 981 173
rect 1087 189 1153 202
rect 759 120 793 164
rect 1017 136 1051 168
rect 759 70 793 86
rect 829 120 1017 130
rect 829 86 845 120
rect 879 102 1017 120
rect 1087 155 1103 189
rect 1137 155 1153 189
rect 1087 119 1153 155
rect 1199 220 1265 236
rect 1199 186 1215 220
rect 1249 186 1265 220
rect 1199 130 1265 186
rect 879 86 1051 102
rect 829 85 1051 86
rect 1199 96 1215 130
rect 1249 96 1265 130
rect 1301 202 1509 236
rect 1301 194 1335 202
rect 1473 194 1509 202
rect 1301 119 1335 160
rect 1371 149 1437 168
rect 1199 85 1265 96
rect 1371 115 1387 149
rect 1421 115 1437 149
rect 1507 160 1509 194
rect 1473 119 1509 160
rect 1543 220 1609 236
rect 1543 186 1559 220
rect 1593 186 1609 220
rect 1543 130 1609 186
rect 1371 85 1437 115
rect 1543 96 1559 130
rect 1593 96 1609 130
rect 1543 85 1609 96
rect 829 51 1609 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o211ai_4
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 1087 316 1121 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 1183 316 1217 350 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 1279 316 1313 350 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 1375 316 1409 350 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 1567 316 1601 350 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 1567 390 1601 424 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 1567 464 1601 498 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 1567 538 1601 572 0 FreeSans 340 0 0 0 Y
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 1632 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1080700
string GDS_START 1066836
<< end >>
