magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1288 561
rect 96 374 162 527
rect 196 340 232 493
rect 268 374 334 527
rect 368 340 406 493
rect 440 440 506 527
rect 657 439 723 527
rect 858 439 911 527
rect 17 287 406 340
rect 1203 383 1269 527
rect 17 161 73 287
rect 508 289 856 337
rect 508 199 566 289
rect 611 207 748 255
rect 790 207 856 289
rect 898 299 1258 337
rect 898 207 969 299
rect 1006 207 1141 265
rect 1178 207 1258 299
rect 17 127 321 161
rect 119 123 321 127
rect 19 17 85 93
rect 119 51 153 123
rect 187 17 253 89
rect 287 51 321 123
rect 355 17 428 93
rect 934 17 997 105
rect 1131 17 1169 105
rect 0 -17 1288 17
<< obsli1 >>
rect 540 405 612 493
rect 757 405 824 493
rect 1031 405 1097 493
rect 440 371 1097 405
rect 440 253 474 371
rect 107 213 474 253
rect 440 163 474 213
rect 440 127 704 163
rect 834 139 1269 173
rect 834 93 900 139
rect 466 51 900 93
rect 1031 51 1097 139
rect 1203 51 1269 139
<< metal1 >>
rect 0 496 1288 592
rect 0 -48 1288 48
<< labels >>
rlabel locali s 1178 207 1258 299 6 A1
port 1 nsew signal input
rlabel locali s 898 299 1258 337 6 A1
port 1 nsew signal input
rlabel locali s 898 207 969 299 6 A1
port 1 nsew signal input
rlabel locali s 1006 207 1141 265 6 A2
port 2 nsew signal input
rlabel locali s 790 207 856 289 6 B1
port 3 nsew signal input
rlabel locali s 508 289 856 337 6 B1
port 3 nsew signal input
rlabel locali s 508 199 566 289 6 B1
port 3 nsew signal input
rlabel locali s 611 207 748 255 6 C1
port 4 nsew signal input
rlabel locali s 368 340 406 493 6 X
port 5 nsew signal output
rlabel locali s 287 51 321 123 6 X
port 5 nsew signal output
rlabel locali s 196 340 232 493 6 X
port 5 nsew signal output
rlabel locali s 119 123 321 127 6 X
port 5 nsew signal output
rlabel locali s 119 51 153 123 6 X
port 5 nsew signal output
rlabel locali s 17 287 406 340 6 X
port 5 nsew signal output
rlabel locali s 17 161 73 287 6 X
port 5 nsew signal output
rlabel locali s 17 127 321 161 6 X
port 5 nsew signal output
rlabel locali s 1131 17 1169 105 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 934 17 997 105 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 355 17 428 93 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 187 17 253 89 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 19 17 85 93 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 1288 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1288 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1203 383 1269 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 858 439 911 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 657 439 723 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 440 440 506 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 268 374 334 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 96 374 162 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 1288 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 1288 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1288 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1330034
string GDS_START 1321038
<< end >>
