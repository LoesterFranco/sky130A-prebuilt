magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 90 47 120 177
rect 162 47 192 177
rect 287 47 317 177
rect 383 47 413 177
rect 479 47 509 177
rect 585 47 615 177
<< pmoshvt >>
rect 82 297 118 497
rect 178 297 214 497
rect 289 297 325 497
rect 385 297 421 497
rect 481 297 517 497
rect 577 297 613 497
<< ndiff >>
rect 27 161 90 177
rect 27 127 35 161
rect 69 127 90 161
rect 27 93 90 127
rect 27 59 35 93
rect 69 59 90 93
rect 27 47 90 59
rect 120 47 162 177
rect 192 89 287 177
rect 192 55 227 89
rect 261 55 287 89
rect 192 47 287 55
rect 317 153 383 177
rect 317 119 338 153
rect 372 119 383 153
rect 317 47 383 119
rect 413 89 479 177
rect 413 55 434 89
rect 468 55 479 89
rect 413 47 479 55
rect 509 169 585 177
rect 509 135 530 169
rect 564 135 585 169
rect 509 101 585 135
rect 509 67 530 101
rect 564 67 585 101
rect 509 47 585 67
rect 615 89 672 177
rect 615 55 626 89
rect 660 55 672 89
rect 615 47 672 55
<< pdiff >>
rect 27 485 82 497
rect 27 451 35 485
rect 69 451 82 485
rect 27 417 82 451
rect 27 383 35 417
rect 69 383 82 417
rect 27 297 82 383
rect 118 477 178 497
rect 118 443 131 477
rect 165 443 178 477
rect 118 409 178 443
rect 118 375 131 409
rect 165 375 178 409
rect 118 297 178 375
rect 214 489 289 497
rect 214 455 234 489
rect 268 455 289 489
rect 214 421 289 455
rect 214 387 234 421
rect 268 387 289 421
rect 214 297 289 387
rect 325 477 385 497
rect 325 443 338 477
rect 372 443 385 477
rect 325 409 385 443
rect 325 375 338 409
rect 372 375 385 409
rect 325 297 385 375
rect 421 489 481 497
rect 421 455 434 489
rect 468 455 481 489
rect 421 421 481 455
rect 421 387 434 421
rect 468 387 481 421
rect 421 297 481 387
rect 517 477 577 497
rect 517 443 530 477
rect 564 443 577 477
rect 517 409 577 443
rect 517 375 530 409
rect 564 375 577 409
rect 517 341 577 375
rect 517 307 530 341
rect 564 307 577 341
rect 517 297 577 307
rect 613 489 672 497
rect 613 455 626 489
rect 660 455 672 489
rect 613 421 672 455
rect 613 387 626 421
rect 660 387 672 421
rect 613 297 672 387
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 227 55 261 89
rect 338 119 372 153
rect 434 55 468 89
rect 530 135 564 169
rect 530 67 564 101
rect 626 55 660 89
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 131 443 165 477
rect 131 375 165 409
rect 234 455 268 489
rect 234 387 268 421
rect 338 443 372 477
rect 338 375 372 409
rect 434 455 468 489
rect 434 387 468 421
rect 530 443 564 477
rect 530 375 564 409
rect 530 307 564 341
rect 626 455 660 489
rect 626 387 660 421
<< poly >>
rect 82 497 118 523
rect 178 497 214 523
rect 289 497 325 523
rect 385 497 421 523
rect 481 497 517 523
rect 577 497 613 523
rect 82 282 118 297
rect 178 282 214 297
rect 289 282 325 297
rect 385 282 421 297
rect 481 282 517 297
rect 577 282 613 297
rect 80 265 120 282
rect 176 265 216 282
rect 287 265 327 282
rect 383 265 423 282
rect 479 265 519 282
rect 575 265 615 282
rect 43 249 120 265
rect 43 215 53 249
rect 87 215 120 249
rect 43 199 120 215
rect 90 177 120 199
rect 162 249 226 265
rect 162 215 172 249
rect 206 215 226 249
rect 162 199 226 215
rect 287 249 615 265
rect 287 215 303 249
rect 337 215 381 249
rect 415 215 459 249
rect 493 215 537 249
rect 571 215 615 249
rect 287 199 615 215
rect 162 177 192 199
rect 287 177 317 199
rect 383 177 413 199
rect 479 177 509 199
rect 585 177 615 199
rect 90 21 120 47
rect 162 21 192 47
rect 287 21 317 47
rect 383 21 413 47
rect 479 21 509 47
rect 585 21 615 47
<< polycont >>
rect 53 215 87 249
rect 172 215 206 249
rect 303 215 337 249
rect 381 215 415 249
rect 459 215 493 249
rect 537 215 571 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 19 485 85 527
rect 19 451 35 485
rect 69 451 85 485
rect 19 417 85 451
rect 19 383 35 417
rect 69 383 85 417
rect 19 376 85 383
rect 131 477 167 493
rect 165 443 167 477
rect 131 409 167 443
rect 165 375 167 409
rect 218 489 284 527
rect 218 455 234 489
rect 268 455 284 489
rect 218 421 284 455
rect 218 387 234 421
rect 268 387 284 421
rect 336 477 374 493
rect 336 443 338 477
rect 372 443 374 477
rect 336 409 374 443
rect 131 350 167 375
rect 336 375 338 409
rect 372 375 374 409
rect 408 489 484 527
rect 408 455 434 489
rect 468 455 484 489
rect 408 421 484 455
rect 408 387 434 421
rect 468 387 484 421
rect 528 477 566 493
rect 528 443 530 477
rect 564 443 566 477
rect 528 409 566 443
rect 336 352 374 375
rect 528 375 530 409
rect 564 375 566 409
rect 600 489 676 527
rect 600 455 626 489
rect 660 455 676 489
rect 600 421 676 455
rect 600 387 626 421
rect 660 387 676 421
rect 528 353 566 375
rect 528 352 714 353
rect 25 249 87 323
rect 131 316 292 350
rect 250 271 292 316
rect 336 341 714 352
rect 336 307 530 341
rect 564 307 714 341
rect 25 215 53 249
rect 25 199 87 215
rect 121 249 216 265
rect 121 215 172 249
rect 206 215 216 249
rect 121 199 216 215
rect 250 249 587 271
rect 250 215 303 249
rect 337 215 381 249
rect 415 215 459 249
rect 493 215 537 249
rect 571 215 587 249
rect 250 204 587 215
rect 250 161 292 204
rect 658 169 714 307
rect 19 127 35 161
rect 69 127 292 161
rect 19 123 292 127
rect 336 153 530 169
rect 19 93 85 123
rect 336 119 338 153
rect 372 135 530 153
rect 564 135 714 169
rect 372 123 714 135
rect 372 119 374 123
rect 336 103 374 119
rect 19 59 35 93
rect 69 59 85 93
rect 528 101 566 123
rect 19 51 85 59
rect 211 55 227 89
rect 261 55 277 89
rect 211 17 277 55
rect 408 55 434 89
rect 468 55 484 89
rect 408 17 484 55
rect 528 67 530 101
rect 564 67 566 101
rect 528 51 566 67
rect 600 55 626 89
rect 660 55 676 89
rect 600 17 676 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel corelocali s 668 153 702 187 0 FreeSans 340 0 0 0 X
port 7 nsew
flabel corelocali s 131 221 165 255 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 29 289 63 323 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew
rlabel comment s 0 0 0 0 4 and2_4
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1495088
string GDS_START 1489050
<< end >>
