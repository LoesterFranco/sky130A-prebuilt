magic
tech sky130A
magscale 1 2
timestamp 1601050056
<< nwell >>
rect -38 332 710 704
<< pwell >>
rect 0 0 672 49
<< scpmos >>
rect 100 392 136 592
rect 184 392 220 592
rect 298 392 334 592
rect 412 392 448 592
rect 550 368 586 592
<< nmoslvt >>
rect 98 112 128 222
rect 184 112 214 222
rect 331 112 361 222
rect 449 112 479 222
rect 551 74 581 222
<< ndiff >>
rect 27 184 98 222
rect 27 150 53 184
rect 87 150 98 184
rect 27 112 98 150
rect 128 184 184 222
rect 128 150 139 184
rect 173 150 184 184
rect 128 112 184 150
rect 214 152 331 222
rect 214 118 255 152
rect 289 118 331 152
rect 214 112 331 118
rect 361 184 449 222
rect 361 150 388 184
rect 422 150 449 184
rect 361 112 449 150
rect 479 152 551 222
rect 479 118 506 152
rect 540 118 551 152
rect 479 112 551 118
rect 229 106 316 112
rect 494 74 551 112
rect 581 210 638 222
rect 581 176 592 210
rect 626 176 638 210
rect 581 120 638 176
rect 581 86 592 120
rect 626 86 638 120
rect 581 74 638 86
<< pdiff >>
rect 44 580 100 592
rect 44 546 56 580
rect 90 546 100 580
rect 44 510 100 546
rect 44 476 56 510
rect 90 476 100 510
rect 44 440 100 476
rect 44 406 56 440
rect 90 406 100 440
rect 44 392 100 406
rect 136 392 184 592
rect 220 392 298 592
rect 334 392 412 592
rect 448 580 550 592
rect 448 546 458 580
rect 492 546 550 580
rect 448 508 550 546
rect 448 474 458 508
rect 492 474 550 508
rect 448 392 550 474
rect 500 368 550 392
rect 586 580 642 592
rect 586 546 596 580
rect 630 546 642 580
rect 586 497 642 546
rect 586 463 596 497
rect 630 463 642 497
rect 586 414 642 463
rect 586 380 596 414
rect 630 380 642 414
rect 586 368 642 380
<< ndiffc >>
rect 53 150 87 184
rect 139 150 173 184
rect 255 118 289 152
rect 388 150 422 184
rect 506 118 540 152
rect 592 176 626 210
rect 592 86 626 120
<< pdiffc >>
rect 56 546 90 580
rect 56 476 90 510
rect 56 406 90 440
rect 458 546 492 580
rect 458 474 492 508
rect 596 546 630 580
rect 596 463 630 497
rect 596 380 630 414
<< poly >>
rect 100 592 136 618
rect 184 592 220 618
rect 298 592 334 618
rect 412 592 448 618
rect 550 592 586 618
rect 100 350 136 392
rect 184 350 220 392
rect 298 350 334 392
rect 64 334 130 350
rect 64 300 80 334
rect 114 300 130 334
rect 64 284 130 300
rect 184 334 250 350
rect 184 300 200 334
rect 234 300 250 334
rect 184 284 250 300
rect 298 334 364 350
rect 298 300 314 334
rect 348 300 364 334
rect 298 284 364 300
rect 412 336 448 392
rect 412 320 479 336
rect 550 326 586 368
rect 412 286 428 320
rect 462 286 479 320
rect 98 222 128 284
rect 184 222 214 284
rect 331 222 361 284
rect 412 270 479 286
rect 449 222 479 270
rect 521 310 587 326
rect 521 276 537 310
rect 571 276 587 310
rect 521 260 587 276
rect 551 222 581 260
rect 98 86 128 112
rect 184 86 214 112
rect 331 86 361 112
rect 449 86 479 112
rect 551 48 581 74
<< polycont >>
rect 80 300 114 334
rect 200 300 234 334
rect 314 300 348 334
rect 428 286 462 320
rect 537 276 571 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 40 580 106 596
rect 40 546 56 580
rect 90 546 106 580
rect 40 510 106 546
rect 40 476 56 510
rect 90 476 106 510
rect 40 440 106 476
rect 430 580 513 649
rect 430 546 458 580
rect 492 546 513 580
rect 430 508 513 546
rect 430 474 458 508
rect 492 474 513 508
rect 430 458 513 474
rect 580 580 655 596
rect 580 546 596 580
rect 630 546 655 580
rect 580 497 655 546
rect 580 463 596 497
rect 630 463 655 497
rect 40 406 56 440
rect 90 424 106 440
rect 90 406 546 424
rect 40 390 546 406
rect 25 334 130 356
rect 25 300 80 334
rect 114 300 130 334
rect 25 284 130 300
rect 184 334 259 356
rect 184 300 200 334
rect 234 300 259 334
rect 184 284 259 300
rect 298 334 364 356
rect 298 300 314 334
rect 348 300 364 334
rect 298 284 364 300
rect 409 320 478 356
rect 409 286 428 320
rect 462 286 478 320
rect 409 270 478 286
rect 512 326 546 390
rect 580 414 655 463
rect 580 380 596 414
rect 630 380 655 414
rect 580 364 655 380
rect 512 310 587 326
rect 512 276 537 310
rect 571 276 587 310
rect 512 260 587 276
rect 512 236 546 260
rect 23 184 89 226
rect 23 150 53 184
rect 87 150 89 184
rect 23 17 89 150
rect 123 202 546 236
rect 621 226 655 364
rect 592 210 655 226
rect 123 184 189 202
rect 123 150 139 184
rect 173 150 189 184
rect 372 184 438 202
rect 123 108 189 150
rect 225 152 320 168
rect 225 118 255 152
rect 289 118 320 152
rect 225 17 320 118
rect 372 150 388 184
rect 422 150 438 184
rect 626 176 655 210
rect 372 108 438 150
rect 490 152 556 168
rect 490 118 506 152
rect 540 118 556 152
rect 490 17 556 118
rect 592 120 655 176
rect 626 86 655 120
rect 592 70 655 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
rlabel comment s 0 0 0 0 4 or4_1
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 D
port 4 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 607 390 641 424 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 607 464 641 498 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 607 538 641 572 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 B
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 672 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 813974
string GDS_START 808088
<< end >>
