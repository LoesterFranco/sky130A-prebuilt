magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 518 704
<< pwell >>
rect 0 0 480 49
<< scnmos >>
rect 84 74 114 222
rect 266 74 296 222
rect 352 74 382 222
<< pmoshvt >>
rect 132 368 162 592
rect 216 368 246 592
rect 347 368 377 592
<< ndiff >>
rect 27 202 84 222
rect 27 168 39 202
rect 73 168 84 202
rect 27 120 84 168
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 84 266 222
rect 114 74 137 84
rect 129 50 137 74
rect 171 50 209 84
rect 243 74 266 84
rect 296 148 352 222
rect 296 114 307 148
rect 341 114 352 148
rect 296 74 352 114
rect 382 210 453 222
rect 382 176 407 210
rect 441 176 453 210
rect 382 120 453 176
rect 382 86 407 120
rect 441 86 453 120
rect 382 74 453 86
rect 243 50 251 74
rect 129 38 251 50
<< pdiff >>
rect 49 580 132 592
rect 49 546 77 580
rect 111 546 132 580
rect 49 497 132 546
rect 49 463 77 497
rect 111 463 132 497
rect 49 414 132 463
rect 49 380 77 414
rect 111 380 132 414
rect 49 368 132 380
rect 162 368 216 592
rect 246 580 347 592
rect 246 546 259 580
rect 293 546 347 580
rect 246 510 347 546
rect 246 476 259 510
rect 293 476 347 510
rect 246 440 347 476
rect 246 406 259 440
rect 293 406 347 440
rect 246 368 347 406
rect 377 580 436 592
rect 377 546 390 580
rect 424 546 436 580
rect 377 510 436 546
rect 377 476 390 510
rect 424 476 436 510
rect 377 440 436 476
rect 377 406 390 440
rect 424 406 436 440
rect 377 368 436 406
<< ndiffc >>
rect 39 168 73 202
rect 39 86 73 120
rect 137 50 171 84
rect 209 50 243 84
rect 307 114 341 148
rect 407 176 441 210
rect 407 86 441 120
<< pdiffc >>
rect 77 546 111 580
rect 77 463 111 497
rect 77 380 111 414
rect 259 546 293 580
rect 259 476 293 510
rect 259 406 293 440
rect 390 546 424 580
rect 390 476 424 510
rect 390 406 424 440
<< poly >>
rect 132 592 162 618
rect 216 592 246 618
rect 347 592 377 618
rect 132 353 162 368
rect 216 353 246 368
rect 347 353 377 368
rect 129 310 165 353
rect 45 294 165 310
rect 45 260 61 294
rect 95 260 165 294
rect 213 336 249 353
rect 344 336 380 353
rect 213 320 296 336
rect 213 286 229 320
rect 263 286 296 320
rect 213 270 296 286
rect 344 320 410 336
rect 344 286 360 320
rect 394 286 410 320
rect 344 270 410 286
rect 45 244 165 260
rect 84 222 114 244
rect 266 222 296 270
rect 352 222 382 270
rect 84 48 114 74
rect 266 48 296 74
rect 352 48 382 74
<< polycont >>
rect 61 260 95 294
rect 229 286 263 320
rect 360 286 394 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 61 580 111 649
rect 61 546 77 580
rect 61 497 111 546
rect 61 463 77 497
rect 61 414 111 463
rect 61 380 77 414
rect 61 364 111 380
rect 145 580 309 596
rect 145 546 259 580
rect 293 546 309 580
rect 145 510 309 546
rect 145 476 259 510
rect 293 476 309 510
rect 145 440 309 476
rect 145 406 259 440
rect 293 406 309 440
rect 145 390 309 406
rect 374 580 440 649
rect 374 546 390 580
rect 424 546 440 580
rect 374 510 440 546
rect 374 476 390 510
rect 424 476 440 510
rect 374 440 440 476
rect 374 406 390 440
rect 424 406 440 440
rect 374 390 440 406
rect 25 294 111 310
rect 25 260 61 294
rect 95 260 111 294
rect 25 236 111 260
rect 145 236 179 390
rect 213 320 279 356
rect 213 286 229 320
rect 263 286 279 320
rect 213 270 279 286
rect 313 320 455 356
rect 313 286 360 320
rect 394 286 455 320
rect 313 270 455 286
rect 145 210 457 236
rect 145 202 407 210
rect 23 168 39 202
rect 73 168 89 202
rect 391 176 407 202
rect 441 176 457 210
rect 23 148 357 168
rect 23 134 307 148
rect 23 120 84 134
rect 23 86 39 120
rect 73 86 84 120
rect 296 114 307 134
rect 341 114 357 148
rect 23 70 84 86
rect 121 84 259 100
rect 121 50 137 84
rect 171 50 209 84
rect 243 50 259 84
rect 296 70 357 114
rect 391 120 457 176
rect 391 86 407 120
rect 441 86 457 120
rect 391 70 457 86
rect 121 17 259 50
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< metal1 >>
rect 0 683 480 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 0 617 480 649
rect 0 17 480 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
rect 0 -49 480 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o21ai_1
flabel pwell s 0 0 480 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 0 617 480 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 480 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 480 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 223 464 257 498 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 223 538 257 572 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 A1
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 480 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1358702
string GDS_START 1353676
<< end >>
