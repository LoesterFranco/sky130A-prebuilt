magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1380 561
rect 129 359 171 527
rect 213 325 255 493
rect 289 359 339 527
rect 373 325 423 493
rect 457 359 507 527
rect 645 325 695 425
rect 813 325 863 425
rect 213 291 863 325
rect 981 359 1031 527
rect 1149 359 1199 527
rect 489 289 863 291
rect 17 215 111 257
rect 489 215 579 289
rect 1317 257 1362 491
rect 613 215 895 255
rect 929 215 1362 257
rect 45 17 79 179
rect 489 163 535 215
rect 284 129 535 163
rect 653 17 687 111
rect 821 17 855 111
rect 989 17 1023 111
rect 1157 17 1191 111
rect 0 -17 1380 17
<< obsli1 >>
rect 29 325 95 487
rect 555 459 947 493
rect 555 359 611 459
rect 729 359 779 459
rect 29 291 179 325
rect 897 325 947 459
rect 1065 325 1115 493
rect 1233 325 1283 493
rect 897 291 1283 325
rect 145 257 179 291
rect 145 215 455 257
rect 145 179 179 215
rect 113 58 179 179
rect 569 145 1291 181
rect 569 95 619 145
rect 216 61 619 95
rect 721 51 787 145
rect 889 51 955 145
rect 1057 51 1123 145
rect 1225 51 1291 145
<< metal1 >>
rect 0 496 1380 592
rect 0 -48 1380 48
<< labels >>
rlabel locali s 1317 257 1362 491 6 A1
port 1 nsew signal input
rlabel locali s 929 215 1362 257 6 A1
port 1 nsew signal input
rlabel locali s 613 215 895 255 6 A2
port 2 nsew signal input
rlabel locali s 17 215 111 257 6 B1_N
port 3 nsew signal input
rlabel locali s 813 325 863 425 6 Y
port 4 nsew signal output
rlabel locali s 645 325 695 425 6 Y
port 4 nsew signal output
rlabel locali s 489 289 863 291 6 Y
port 4 nsew signal output
rlabel locali s 489 215 579 289 6 Y
port 4 nsew signal output
rlabel locali s 489 163 535 215 6 Y
port 4 nsew signal output
rlabel locali s 373 325 423 493 6 Y
port 4 nsew signal output
rlabel locali s 284 129 535 163 6 Y
port 4 nsew signal output
rlabel locali s 213 325 255 493 6 Y
port 4 nsew signal output
rlabel locali s 213 291 863 325 6 Y
port 4 nsew signal output
rlabel locali s 1157 17 1191 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 989 17 1023 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 821 17 855 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 653 17 687 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 45 17 79 179 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 1380 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1380 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 1149 359 1199 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 981 359 1031 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 457 359 507 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 289 359 339 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 129 359 171 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 1380 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 1380 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1380 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1412390
string GDS_START 1401582
<< end >>
