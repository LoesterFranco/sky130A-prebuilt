magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 1326 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 80 47 110 177
rect 186 47 216 177
rect 282 47 312 177
rect 378 47 408 177
rect 472 47 502 177
rect 568 47 598 177
rect 664 47 694 177
rect 760 47 790 177
rect 866 47 896 177
rect 952 47 982 177
rect 1048 47 1078 177
rect 1144 47 1174 177
<< pmoshvt >>
rect 82 297 118 497
rect 178 297 214 497
rect 274 297 310 497
rect 370 297 406 497
rect 472 297 508 497
rect 570 297 606 497
rect 666 297 702 497
rect 762 297 798 497
rect 858 297 894 497
rect 954 297 990 497
rect 1050 297 1086 497
rect 1146 297 1182 497
<< ndiff >>
rect 27 161 80 177
rect 27 127 35 161
rect 69 127 80 161
rect 27 93 80 127
rect 27 59 35 93
rect 69 59 80 93
rect 27 47 80 59
rect 110 124 186 177
rect 110 90 131 124
rect 165 90 186 124
rect 110 47 186 90
rect 216 89 282 177
rect 216 55 227 89
rect 261 55 282 89
rect 216 47 282 55
rect 312 169 378 177
rect 312 135 323 169
rect 357 135 378 169
rect 312 101 378 135
rect 312 67 323 101
rect 357 67 378 101
rect 312 47 378 67
rect 408 89 472 177
rect 408 55 427 89
rect 461 55 472 89
rect 408 47 472 55
rect 502 101 568 177
rect 502 67 523 101
rect 557 67 568 101
rect 502 47 568 67
rect 598 169 664 177
rect 598 135 619 169
rect 653 135 664 169
rect 598 47 664 135
rect 694 101 760 177
rect 694 67 715 101
rect 749 67 760 101
rect 694 47 760 67
rect 790 169 866 177
rect 790 135 811 169
rect 845 135 866 169
rect 790 47 866 135
rect 896 157 952 177
rect 896 123 907 157
rect 941 123 952 157
rect 896 89 952 123
rect 896 55 907 89
rect 941 55 952 89
rect 896 47 952 55
rect 982 97 1048 177
rect 982 63 1003 97
rect 1037 63 1048 97
rect 982 47 1048 63
rect 1078 164 1144 177
rect 1078 130 1099 164
rect 1133 130 1144 164
rect 1078 96 1144 130
rect 1078 62 1099 96
rect 1133 62 1144 96
rect 1078 47 1144 62
rect 1174 161 1237 177
rect 1174 127 1195 161
rect 1229 127 1237 161
rect 1174 93 1237 127
rect 1174 59 1195 93
rect 1229 59 1237 93
rect 1174 47 1237 59
<< pdiff >>
rect 28 477 82 497
rect 28 443 36 477
rect 70 443 82 477
rect 28 409 82 443
rect 28 375 36 409
rect 70 375 82 409
rect 28 297 82 375
rect 118 387 178 497
rect 118 353 131 387
rect 165 353 178 387
rect 118 297 178 353
rect 214 489 274 497
rect 214 455 227 489
rect 261 455 274 489
rect 214 297 274 455
rect 310 395 370 497
rect 310 361 323 395
rect 357 361 370 395
rect 310 297 370 361
rect 406 477 472 497
rect 406 443 425 477
rect 459 443 472 477
rect 406 297 472 443
rect 508 489 570 497
rect 508 455 523 489
rect 557 455 570 489
rect 508 297 570 455
rect 606 477 666 497
rect 606 443 619 477
rect 653 443 666 477
rect 606 409 666 443
rect 606 375 619 409
rect 653 375 666 409
rect 606 297 666 375
rect 702 489 762 497
rect 702 455 715 489
rect 749 455 762 489
rect 702 297 762 455
rect 798 477 858 497
rect 798 443 811 477
rect 845 443 858 477
rect 798 409 858 443
rect 798 375 811 409
rect 845 375 858 409
rect 798 297 858 375
rect 894 489 954 497
rect 894 455 907 489
rect 941 455 954 489
rect 894 297 954 455
rect 990 477 1050 497
rect 990 443 1003 477
rect 1037 443 1050 477
rect 990 297 1050 443
rect 1086 489 1146 497
rect 1086 455 1099 489
rect 1133 455 1146 489
rect 1086 297 1146 455
rect 1182 477 1237 497
rect 1182 443 1195 477
rect 1229 443 1237 477
rect 1182 409 1237 443
rect 1182 375 1195 409
rect 1229 375 1237 409
rect 1182 297 1237 375
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 131 90 165 124
rect 227 55 261 89
rect 323 135 357 169
rect 323 67 357 101
rect 427 55 461 89
rect 523 67 557 101
rect 619 135 653 169
rect 715 67 749 101
rect 811 135 845 169
rect 907 123 941 157
rect 907 55 941 89
rect 1003 63 1037 97
rect 1099 130 1133 164
rect 1099 62 1133 96
rect 1195 127 1229 161
rect 1195 59 1229 93
<< pdiffc >>
rect 36 443 70 477
rect 36 375 70 409
rect 131 353 165 387
rect 227 455 261 489
rect 323 361 357 395
rect 425 443 459 477
rect 523 455 557 489
rect 619 443 653 477
rect 619 375 653 409
rect 715 455 749 489
rect 811 443 845 477
rect 811 375 845 409
rect 907 455 941 489
rect 1003 443 1037 477
rect 1099 455 1133 489
rect 1195 443 1229 477
rect 1195 375 1229 409
<< poly >>
rect 82 497 118 523
rect 178 497 214 523
rect 274 497 310 523
rect 370 497 406 523
rect 472 497 508 523
rect 570 497 606 523
rect 666 497 702 523
rect 762 497 798 523
rect 858 497 894 523
rect 954 497 990 523
rect 1050 497 1086 523
rect 1146 497 1182 523
rect 82 282 118 297
rect 178 282 214 297
rect 274 282 310 297
rect 370 282 406 297
rect 472 282 508 297
rect 570 282 606 297
rect 666 282 702 297
rect 762 282 798 297
rect 858 282 894 297
rect 954 282 990 297
rect 1050 282 1086 297
rect 1146 282 1182 297
rect 80 265 120 282
rect 176 265 216 282
rect 272 265 312 282
rect 368 265 408 282
rect 470 265 510 282
rect 22 249 408 265
rect 22 215 32 249
rect 66 215 100 249
rect 134 215 178 249
rect 212 215 256 249
rect 290 215 408 249
rect 22 199 408 215
rect 450 249 526 265
rect 450 215 466 249
rect 500 215 526 249
rect 450 199 526 215
rect 568 259 608 282
rect 664 259 704 282
rect 760 259 800 282
rect 856 259 896 282
rect 568 249 896 259
rect 568 215 592 249
rect 626 215 670 249
rect 704 215 748 249
rect 782 215 826 249
rect 860 215 896 249
rect 80 177 110 199
rect 186 177 216 199
rect 282 177 312 199
rect 378 177 408 199
rect 472 177 502 199
rect 568 198 896 215
rect 568 177 598 198
rect 664 177 694 198
rect 760 177 790 198
rect 866 177 896 198
rect 952 265 992 282
rect 1048 265 1088 282
rect 1144 265 1184 282
rect 952 249 1208 265
rect 952 215 1008 249
rect 1042 215 1076 249
rect 1110 215 1154 249
rect 1188 215 1208 249
rect 952 199 1208 215
rect 952 177 982 199
rect 1048 177 1078 199
rect 1144 177 1174 199
rect 80 21 110 47
rect 186 21 216 47
rect 282 21 312 47
rect 378 21 408 47
rect 472 21 502 47
rect 568 21 598 47
rect 664 21 694 47
rect 760 21 790 47
rect 866 21 896 47
rect 952 21 982 47
rect 1048 21 1078 47
rect 1144 21 1174 47
<< polycont >>
rect 32 215 66 249
rect 100 215 134 249
rect 178 215 212 249
rect 256 215 290 249
rect 466 215 500 249
rect 592 215 626 249
rect 670 215 704 249
rect 748 215 782 249
rect 826 215 860 249
rect 1008 215 1042 249
rect 1076 215 1110 249
rect 1154 215 1188 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 36 489 463 493
rect 36 477 227 489
rect 70 455 227 477
rect 261 477 463 489
rect 261 455 425 477
rect 70 443 425 455
rect 459 443 463 477
rect 497 489 573 527
rect 497 455 523 489
rect 557 455 573 489
rect 617 477 655 493
rect 36 409 75 443
rect 201 441 463 443
rect 70 375 75 409
rect 423 421 463 441
rect 617 443 619 477
rect 653 443 655 477
rect 689 489 765 527
rect 689 455 715 489
rect 749 455 765 489
rect 809 477 847 493
rect 617 421 655 443
rect 809 443 811 477
rect 845 443 847 477
rect 881 489 957 527
rect 881 455 907 489
rect 941 455 957 489
rect 1001 477 1037 493
rect 809 421 847 443
rect 1001 443 1003 477
rect 1073 489 1149 527
rect 1073 455 1099 489
rect 1133 455 1149 489
rect 1193 477 1245 493
rect 1001 421 1037 443
rect 1193 443 1195 477
rect 1229 443 1245 477
rect 1193 421 1245 443
rect 423 409 1245 421
rect 36 359 75 375
rect 126 395 379 407
rect 126 387 323 395
rect 126 353 131 387
rect 165 361 323 387
rect 357 361 379 395
rect 423 375 619 409
rect 653 375 811 409
rect 845 375 1195 409
rect 1229 375 1245 409
rect 165 353 379 361
rect 126 341 379 353
rect 126 317 416 341
rect 18 249 316 283
rect 18 215 32 249
rect 66 215 100 249
rect 134 215 178 249
rect 212 215 256 249
rect 290 215 316 249
rect 18 207 316 215
rect 18 199 80 207
rect 350 179 416 317
rect 450 296 1214 341
rect 450 249 529 296
rect 450 215 466 249
rect 500 215 529 249
rect 450 213 529 215
rect 563 249 880 262
rect 563 215 592 249
rect 626 215 670 249
rect 704 215 748 249
rect 782 215 826 249
rect 860 215 880 249
rect 935 249 1214 296
rect 935 215 1008 249
rect 1042 215 1076 249
rect 1110 215 1154 249
rect 1188 215 1214 249
rect 563 213 880 215
rect 350 173 861 179
rect 129 169 861 173
rect 18 127 35 161
rect 69 127 85 161
rect 18 93 85 127
rect 18 59 35 93
rect 69 59 85 93
rect 129 135 323 169
rect 357 139 619 169
rect 357 135 359 139
rect 495 135 619 139
rect 653 135 811 169
rect 845 135 861 169
rect 905 164 1149 181
rect 905 157 1099 164
rect 129 124 359 135
rect 129 90 131 124
rect 165 123 359 124
rect 165 90 167 123
rect 129 74 167 90
rect 321 101 359 123
rect 905 123 907 157
rect 941 147 1099 157
rect 941 123 957 147
rect 18 17 85 59
rect 201 55 227 89
rect 261 55 277 89
rect 201 17 277 55
rect 321 67 323 101
rect 357 67 359 101
rect 321 51 359 67
rect 397 89 463 105
rect 905 101 957 123
rect 1073 130 1099 147
rect 1133 130 1149 164
rect 397 55 427 89
rect 461 55 463 89
rect 397 17 463 55
rect 497 67 523 101
rect 557 67 715 101
rect 749 89 957 101
rect 749 67 907 89
rect 497 55 907 67
rect 941 55 957 89
rect 497 51 957 55
rect 1001 97 1039 113
rect 1001 63 1003 97
rect 1037 63 1039 97
rect 1001 17 1039 63
rect 1073 96 1149 130
rect 1073 62 1099 96
rect 1133 62 1149 96
rect 1073 51 1149 62
rect 1193 161 1245 177
rect 1193 127 1195 161
rect 1229 127 1245 161
rect 1193 93 1245 127
rect 1193 59 1195 93
rect 1229 59 1245 93
rect 1193 17 1245 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
flabel corelocali s 215 221 249 255 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 1059 306 1059 306 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 768 221 802 255 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 307 357 341 391 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 1288 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1214842
string GDS_START 1205838
<< end >>
