magic
tech sky130A
magscale 1 2
timestamp 1604502705
<< nwell >>
rect -38 332 1862 704
rect 291 312 459 332
<< pwell >>
rect 0 0 1824 49
<< scnmos >>
rect 84 112 114 222
rect 200 74 230 222
rect 420 74 450 222
rect 562 74 592 202
rect 640 74 670 202
rect 760 74 790 158
rect 838 74 868 158
rect 1036 74 1066 222
rect 1114 74 1144 222
rect 1232 74 1262 222
rect 1318 74 1348 222
rect 1418 74 1448 202
rect 1616 74 1646 222
rect 1710 74 1740 222
<< pmoshvt >>
rect 86 424 116 592
rect 222 424 252 592
rect 441 392 471 560
rect 565 392 595 592
rect 643 392 673 592
rect 753 508 783 592
rect 878 508 908 592
rect 1033 368 1063 592
rect 1125 368 1155 592
rect 1225 368 1255 592
rect 1315 368 1345 592
rect 1416 368 1446 568
rect 1618 368 1648 592
rect 1708 368 1738 592
<< ndiff >>
rect 27 180 84 222
rect 27 146 39 180
rect 73 146 84 180
rect 27 112 84 146
rect 114 202 200 222
rect 114 168 141 202
rect 175 168 200 202
rect 114 123 200 168
rect 114 112 141 123
rect 129 89 141 112
rect 175 89 200 123
rect 129 74 200 89
rect 230 202 287 222
rect 230 168 241 202
rect 275 168 287 202
rect 230 120 287 168
rect 230 86 241 120
rect 275 86 287 120
rect 230 74 287 86
rect 363 192 420 222
rect 363 158 375 192
rect 409 158 420 192
rect 363 120 420 158
rect 363 86 375 120
rect 409 86 420 120
rect 363 74 420 86
rect 450 202 500 222
rect 450 120 562 202
rect 450 86 496 120
rect 530 86 562 120
rect 450 74 562 86
rect 592 74 640 202
rect 670 158 720 202
rect 979 210 1036 222
rect 979 176 991 210
rect 1025 176 1036 210
rect 670 122 760 158
rect 670 88 698 122
rect 732 88 760 122
rect 670 74 760 88
rect 790 74 838 158
rect 868 123 925 158
rect 868 89 879 123
rect 913 89 925 123
rect 868 74 925 89
rect 979 120 1036 176
rect 979 86 991 120
rect 1025 86 1036 120
rect 979 74 1036 86
rect 1066 74 1114 222
rect 1144 199 1232 222
rect 1144 165 1155 199
rect 1189 165 1232 199
rect 1144 120 1232 165
rect 1144 86 1155 120
rect 1189 86 1232 120
rect 1144 74 1232 86
rect 1262 207 1318 222
rect 1262 173 1273 207
rect 1307 173 1318 207
rect 1262 74 1318 173
rect 1348 202 1398 222
rect 1348 194 1418 202
rect 1348 160 1359 194
rect 1393 160 1418 194
rect 1348 120 1418 160
rect 1348 86 1359 120
rect 1393 86 1418 120
rect 1348 74 1418 86
rect 1448 190 1505 202
rect 1448 156 1459 190
rect 1493 156 1505 190
rect 1448 120 1505 156
rect 1448 86 1459 120
rect 1493 86 1505 120
rect 1448 74 1505 86
rect 1559 194 1616 222
rect 1559 160 1571 194
rect 1605 160 1616 194
rect 1559 123 1616 160
rect 1559 89 1571 123
rect 1605 89 1616 123
rect 1559 74 1616 89
rect 1646 210 1710 222
rect 1646 176 1661 210
rect 1695 176 1710 210
rect 1646 74 1710 176
rect 1740 210 1797 222
rect 1740 176 1751 210
rect 1785 176 1797 210
rect 1740 123 1797 176
rect 1740 89 1751 123
rect 1785 89 1797 123
rect 1740 74 1797 89
<< pdiff >>
rect 489 614 547 626
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 470 86 546
rect 27 436 39 470
rect 73 436 86 470
rect 27 424 86 436
rect 116 559 222 592
rect 116 525 129 559
rect 163 525 222 559
rect 116 424 222 525
rect 252 475 311 592
rect 489 580 501 614
rect 535 592 547 614
rect 535 580 565 592
rect 489 560 565 580
rect 252 441 265 475
rect 299 441 311 475
rect 252 424 311 441
rect 365 394 441 560
rect 365 360 377 394
rect 411 392 441 394
rect 471 392 565 560
rect 595 392 643 592
rect 673 531 753 592
rect 673 497 687 531
rect 721 508 753 531
rect 783 508 878 592
rect 908 580 1033 592
rect 908 546 949 580
rect 983 546 1033 580
rect 908 508 1033 546
rect 721 497 735 508
rect 673 392 735 497
rect 411 360 423 392
rect 365 348 423 360
rect 980 368 1033 508
rect 1063 580 1125 592
rect 1063 546 1078 580
rect 1112 546 1125 580
rect 1063 497 1125 546
rect 1063 463 1078 497
rect 1112 463 1125 497
rect 1063 414 1125 463
rect 1063 380 1078 414
rect 1112 380 1125 414
rect 1063 368 1125 380
rect 1155 573 1225 592
rect 1155 539 1178 573
rect 1212 539 1225 573
rect 1155 368 1225 539
rect 1255 414 1315 592
rect 1255 380 1268 414
rect 1302 380 1315 414
rect 1255 368 1315 380
rect 1345 568 1398 592
rect 1559 580 1618 592
rect 1345 553 1416 568
rect 1345 519 1358 553
rect 1392 519 1416 553
rect 1345 368 1416 519
rect 1446 556 1505 568
rect 1446 522 1459 556
rect 1493 522 1505 556
rect 1446 485 1505 522
rect 1446 451 1459 485
rect 1493 451 1505 485
rect 1446 414 1505 451
rect 1446 380 1459 414
rect 1493 380 1505 414
rect 1446 368 1505 380
rect 1559 546 1571 580
rect 1605 546 1618 580
rect 1559 497 1618 546
rect 1559 463 1571 497
rect 1605 463 1618 497
rect 1559 414 1618 463
rect 1559 380 1571 414
rect 1605 380 1618 414
rect 1559 368 1618 380
rect 1648 580 1708 592
rect 1648 546 1661 580
rect 1695 546 1708 580
rect 1648 497 1708 546
rect 1648 463 1661 497
rect 1695 463 1708 497
rect 1648 414 1708 463
rect 1648 380 1661 414
rect 1695 380 1708 414
rect 1648 368 1708 380
rect 1738 580 1797 592
rect 1738 546 1751 580
rect 1785 546 1797 580
rect 1738 497 1797 546
rect 1738 463 1751 497
rect 1785 463 1797 497
rect 1738 414 1797 463
rect 1738 380 1751 414
rect 1785 380 1797 414
rect 1738 368 1797 380
<< ndiffc >>
rect 39 146 73 180
rect 141 168 175 202
rect 141 89 175 123
rect 241 168 275 202
rect 241 86 275 120
rect 375 158 409 192
rect 375 86 409 120
rect 496 86 530 120
rect 991 176 1025 210
rect 698 88 732 122
rect 879 89 913 123
rect 991 86 1025 120
rect 1155 165 1189 199
rect 1155 86 1189 120
rect 1273 173 1307 207
rect 1359 160 1393 194
rect 1359 86 1393 120
rect 1459 156 1493 190
rect 1459 86 1493 120
rect 1571 160 1605 194
rect 1571 89 1605 123
rect 1661 176 1695 210
rect 1751 176 1785 210
rect 1751 89 1785 123
<< pdiffc >>
rect 39 546 73 580
rect 39 436 73 470
rect 129 525 163 559
rect 501 580 535 614
rect 265 441 299 475
rect 377 360 411 394
rect 687 497 721 531
rect 949 546 983 580
rect 1078 546 1112 580
rect 1078 463 1112 497
rect 1078 380 1112 414
rect 1178 539 1212 573
rect 1268 380 1302 414
rect 1358 519 1392 553
rect 1459 522 1493 556
rect 1459 451 1493 485
rect 1459 380 1493 414
rect 1571 546 1605 580
rect 1571 463 1605 497
rect 1571 380 1605 414
rect 1661 546 1695 580
rect 1661 463 1695 497
rect 1661 380 1695 414
rect 1751 546 1785 580
rect 1751 463 1785 497
rect 1751 380 1785 414
<< poly >>
rect 86 592 116 618
rect 222 592 252 618
rect 441 560 471 586
rect 565 592 595 618
rect 643 592 673 618
rect 753 592 783 618
rect 878 592 908 618
rect 1033 592 1063 618
rect 1125 592 1155 618
rect 1225 592 1255 618
rect 1315 592 1345 618
rect 86 409 116 424
rect 222 409 252 424
rect 83 386 119 409
rect 219 386 255 409
rect 83 370 151 386
rect 83 336 101 370
rect 135 336 151 370
rect 83 302 151 336
rect 83 268 101 302
rect 135 268 151 302
rect 83 252 151 268
rect 193 370 259 386
rect 193 336 209 370
rect 243 336 259 370
rect 753 493 783 508
rect 878 493 908 508
rect 750 476 786 493
rect 750 460 833 476
rect 750 426 783 460
rect 817 426 833 460
rect 750 410 833 426
rect 875 473 911 493
rect 875 457 941 473
rect 875 423 891 457
rect 925 423 941 457
rect 875 407 941 423
rect 441 377 471 392
rect 565 377 595 392
rect 643 377 673 392
rect 193 302 259 336
rect 438 310 474 377
rect 562 360 598 377
rect 532 344 598 360
rect 532 310 548 344
rect 582 310 598 344
rect 640 368 676 377
rect 640 338 790 368
rect 193 268 209 302
rect 243 268 259 302
rect 193 252 259 268
rect 420 294 490 310
rect 532 294 598 310
rect 760 311 790 338
rect 760 295 826 311
rect 420 260 440 294
rect 474 260 490 294
rect 84 222 114 252
rect 200 222 230 252
rect 420 244 490 260
rect 420 222 450 244
rect 84 86 114 112
rect 562 202 592 294
rect 640 274 706 290
rect 640 240 656 274
rect 690 240 706 274
rect 640 224 706 240
rect 760 261 776 295
rect 810 261 826 295
rect 760 245 826 261
rect 640 202 670 224
rect 760 158 790 245
rect 875 203 905 407
rect 1416 568 1446 594
rect 1618 592 1648 618
rect 1708 592 1738 618
rect 1033 353 1063 368
rect 1125 353 1155 368
rect 1225 353 1255 368
rect 1315 353 1345 368
rect 1416 353 1446 368
rect 1618 353 1648 368
rect 1708 353 1738 368
rect 1030 336 1066 353
rect 947 320 1066 336
rect 947 286 963 320
rect 997 286 1066 320
rect 1122 310 1158 353
rect 947 270 1066 286
rect 1036 222 1066 270
rect 1114 294 1180 310
rect 1114 260 1130 294
rect 1164 260 1180 294
rect 1222 294 1258 353
rect 1312 330 1348 353
rect 1413 330 1449 353
rect 1312 314 1449 330
rect 1312 294 1341 314
rect 1222 280 1341 294
rect 1375 280 1449 314
rect 1615 322 1651 353
rect 1615 310 1646 322
rect 1222 264 1449 280
rect 1512 294 1646 310
rect 1114 244 1180 260
rect 1114 222 1144 244
rect 1232 222 1262 264
rect 1318 222 1348 264
rect 838 173 905 203
rect 838 158 868 173
rect 1418 202 1448 264
rect 1512 260 1528 294
rect 1562 260 1596 294
rect 1630 274 1646 294
rect 1705 274 1741 353
rect 1630 260 1740 274
rect 1512 244 1740 260
rect 1616 222 1646 244
rect 1710 222 1740 244
rect 200 48 230 74
rect 420 48 450 74
rect 562 48 592 74
rect 640 48 670 74
rect 760 48 790 74
rect 838 48 868 74
rect 1036 48 1066 74
rect 1114 48 1144 74
rect 1232 48 1262 74
rect 1318 48 1348 74
rect 1418 48 1448 74
rect 1616 48 1646 74
rect 1710 48 1740 74
<< polycont >>
rect 101 336 135 370
rect 101 268 135 302
rect 209 336 243 370
rect 783 426 817 460
rect 891 423 925 457
rect 548 310 582 344
rect 209 268 243 302
rect 440 260 474 294
rect 656 240 690 274
rect 776 261 810 295
rect 963 286 997 320
rect 1130 260 1164 294
rect 1341 280 1375 314
rect 1528 260 1562 294
rect 1596 260 1630 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 17 580 89 596
rect 17 546 39 580
rect 73 546 89 580
rect 17 470 89 546
rect 129 559 163 649
rect 485 614 551 649
rect 485 580 501 614
rect 535 580 551 614
rect 485 564 551 580
rect 602 581 833 615
rect 129 488 163 525
rect 197 530 393 564
rect 17 436 39 470
rect 73 454 89 470
rect 197 454 231 530
rect 359 496 566 530
rect 73 436 231 454
rect 17 420 231 436
rect 265 475 325 496
rect 299 462 325 475
rect 299 441 495 462
rect 265 428 495 441
rect 265 420 325 428
rect 17 218 51 420
rect 85 370 161 386
rect 85 336 101 370
rect 135 336 161 370
rect 85 302 161 336
rect 85 268 101 302
rect 135 268 161 302
rect 85 252 161 268
rect 195 370 257 386
rect 195 336 209 370
rect 243 336 257 370
rect 195 302 257 336
rect 195 268 209 302
rect 243 268 257 302
rect 195 252 257 268
rect 291 218 325 420
rect 17 180 89 218
rect 17 146 39 180
rect 73 146 89 180
rect 17 108 89 146
rect 125 202 191 218
rect 125 168 141 202
rect 175 168 191 202
rect 125 123 191 168
rect 125 89 141 123
rect 175 89 191 123
rect 125 17 191 89
rect 225 202 325 218
rect 225 168 241 202
rect 275 168 325 202
rect 225 120 325 168
rect 225 86 241 120
rect 275 86 325 120
rect 225 70 325 86
rect 359 360 377 394
rect 411 360 427 394
rect 359 344 427 360
rect 359 192 393 344
rect 461 310 495 428
rect 427 294 495 310
rect 532 360 566 496
rect 602 428 636 581
rect 670 531 733 547
rect 670 497 687 531
rect 721 497 733 531
rect 670 481 733 497
rect 602 394 665 428
rect 532 344 597 360
rect 532 310 548 344
rect 582 310 597 344
rect 532 294 597 310
rect 427 260 440 294
rect 474 260 495 294
rect 631 290 665 394
rect 699 376 733 481
rect 767 460 833 581
rect 905 580 1028 649
rect 905 546 949 580
rect 983 546 1028 580
rect 905 530 1028 546
rect 1062 580 1128 596
rect 1062 546 1078 580
rect 1112 546 1128 580
rect 1062 497 1128 546
rect 1162 573 1228 649
rect 1162 539 1178 573
rect 1212 539 1228 573
rect 1162 516 1228 539
rect 1342 553 1408 649
rect 1555 580 1605 649
rect 1342 519 1358 553
rect 1392 519 1408 553
rect 1342 516 1408 519
rect 1443 556 1509 572
rect 1443 522 1459 556
rect 1493 522 1509 556
rect 1062 470 1078 497
rect 767 426 783 460
rect 817 426 833 460
rect 767 410 833 426
rect 875 463 1078 470
rect 1112 482 1128 497
rect 1443 485 1509 522
rect 1112 463 1391 482
rect 875 457 1391 463
rect 875 423 891 457
rect 925 448 1391 457
rect 925 423 1128 448
rect 875 414 1128 423
rect 875 410 1078 414
rect 1046 380 1078 410
rect 1112 380 1128 414
rect 699 342 1012 376
rect 743 295 826 308
rect 631 274 706 290
rect 631 260 656 274
rect 427 240 656 260
rect 690 240 706 274
rect 427 226 706 240
rect 631 224 706 226
rect 743 261 776 295
rect 810 261 826 295
rect 743 245 826 261
rect 359 158 375 192
rect 409 190 425 192
rect 743 190 777 245
rect 860 211 894 342
rect 947 320 1012 342
rect 947 286 963 320
rect 997 286 1012 320
rect 947 270 1012 286
rect 1046 364 1128 380
rect 1252 380 1268 414
rect 1302 380 1318 414
rect 1252 364 1318 380
rect 1046 226 1080 364
rect 1114 294 1223 310
rect 1114 260 1130 294
rect 1164 260 1223 294
rect 1114 236 1223 260
rect 409 158 777 190
rect 359 156 777 158
rect 811 177 894 211
rect 975 210 1080 226
rect 359 120 425 156
rect 811 122 845 177
rect 975 176 991 210
rect 1025 176 1080 210
rect 1257 226 1291 364
rect 1357 330 1391 448
rect 1325 314 1391 330
rect 1325 280 1341 314
rect 1375 280 1391 314
rect 1325 264 1391 280
rect 1443 451 1459 485
rect 1493 451 1509 485
rect 1443 414 1509 451
rect 1443 380 1459 414
rect 1493 380 1509 414
rect 1443 310 1509 380
rect 1555 546 1571 580
rect 1555 497 1605 546
rect 1555 463 1571 497
rect 1555 414 1605 463
rect 1555 380 1571 414
rect 1555 364 1605 380
rect 1645 580 1715 596
rect 1645 546 1661 580
rect 1695 546 1715 580
rect 1645 497 1715 546
rect 1645 463 1661 497
rect 1695 463 1715 497
rect 1645 414 1715 463
rect 1645 380 1661 414
rect 1695 380 1715 414
rect 1645 364 1715 380
rect 1751 580 1801 649
rect 1785 546 1801 580
rect 1751 497 1801 546
rect 1785 463 1801 497
rect 1751 414 1801 463
rect 1785 380 1801 414
rect 1751 364 1801 380
rect 1443 294 1646 310
rect 1443 260 1528 294
rect 1562 260 1596 294
rect 1630 260 1646 294
rect 1443 244 1646 260
rect 1257 207 1323 226
rect 359 86 375 120
rect 409 86 425 120
rect 359 70 425 86
rect 459 86 496 120
rect 530 86 567 120
rect 459 17 567 86
rect 665 88 698 122
rect 732 88 845 122
rect 665 72 845 88
rect 879 123 929 143
rect 913 89 929 123
rect 879 17 929 89
rect 975 120 1080 176
rect 975 86 991 120
rect 1025 86 1080 120
rect 975 70 1080 86
rect 1139 199 1205 202
rect 1139 165 1155 199
rect 1189 165 1205 199
rect 1139 120 1205 165
rect 1257 173 1273 207
rect 1307 173 1323 207
rect 1257 154 1323 173
rect 1357 194 1409 210
rect 1357 160 1359 194
rect 1393 160 1409 194
rect 1139 86 1155 120
rect 1189 86 1205 120
rect 1139 17 1205 86
rect 1357 120 1409 160
rect 1357 86 1359 120
rect 1393 86 1409 120
rect 1357 17 1409 86
rect 1443 190 1509 244
rect 1681 210 1715 364
rect 1443 156 1459 190
rect 1493 156 1509 190
rect 1443 120 1509 156
rect 1443 86 1459 120
rect 1493 86 1509 120
rect 1443 70 1509 86
rect 1555 194 1607 210
rect 1555 160 1571 194
rect 1605 160 1607 194
rect 1641 176 1661 210
rect 1695 176 1715 210
rect 1749 210 1801 226
rect 1749 176 1751 210
rect 1785 176 1801 210
rect 1555 123 1607 160
rect 1555 89 1571 123
rect 1605 89 1607 123
rect 1555 17 1607 89
rect 1749 123 1801 176
rect 1749 89 1751 123
rect 1785 89 1801 123
rect 1749 17 1801 89
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
<< metal1 >>
rect 0 683 1824 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 0 617 1824 649
rect 0 17 1824 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
rect 0 -49 1824 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dlrbn_2
flabel pwell s 0 0 1824 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 1824 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 1824 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 1824 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 1 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew
flabel corelocali s 1183 242 1217 276 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew
flabel corelocali s 1279 168 1313 202 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 1663 390 1697 424 0 FreeSans 340 0 0 0 Q_N
port 9 nsew
flabel corelocali s 1663 464 1697 498 0 FreeSans 340 0 0 0 Q_N
port 9 nsew
flabel corelocali s 1663 538 1697 572 0 FreeSans 340 0 0 0 Q_N
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 1824 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2870226
string GDS_START 2856226
<< end >>
