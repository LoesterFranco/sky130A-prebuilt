magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1472 561
rect 29 291 79 527
rect 197 425 247 527
rect 533 425 685 527
rect 971 425 1021 527
rect 1063 391 1105 493
rect 1139 425 1189 527
rect 1063 357 1180 391
rect 1146 323 1180 357
rect 1223 323 1273 493
rect 1307 359 1357 527
rect 18 215 88 255
rect 205 289 549 323
rect 205 215 304 289
rect 338 215 449 255
rect 483 215 549 289
rect 601 289 955 323
rect 1146 289 1384 323
rect 601 215 721 289
rect 905 255 955 289
rect 755 215 871 255
rect 905 215 1007 255
rect 1315 181 1384 289
rect 629 17 677 109
rect 811 17 845 111
rect 979 17 1013 181
rect 1047 147 1384 181
rect 1047 145 1281 147
rect 1047 51 1113 145
rect 1147 17 1181 111
rect 1215 51 1281 145
rect 1315 17 1366 113
rect 0 -17 1472 17
<< obsli1 >>
rect 113 391 163 493
rect 281 459 499 493
rect 281 425 331 459
rect 449 425 499 459
rect 719 459 937 493
rect 719 425 769 459
rect 887 425 937 459
rect 365 391 415 425
rect 803 391 853 425
rect 113 357 1029 391
rect 113 289 169 357
rect 995 323 1029 357
rect 17 95 69 179
rect 122 173 169 289
rect 995 289 1075 323
rect 1041 255 1075 289
rect 1041 215 1281 255
rect 103 129 169 173
rect 203 95 237 181
rect 271 145 945 181
rect 271 143 777 145
rect 271 129 507 143
rect 17 51 591 95
rect 711 51 777 143
rect 879 51 945 145
<< metal1 >>
rect 0 496 1472 592
rect 0 -48 1472 48
<< labels >>
rlabel locali s 905 255 955 289 6 A1
port 1 nsew signal input
rlabel locali s 905 215 1007 255 6 A1
port 1 nsew signal input
rlabel locali s 601 289 955 323 6 A1
port 1 nsew signal input
rlabel locali s 601 215 721 289 6 A1
port 1 nsew signal input
rlabel locali s 755 215 871 255 6 A2
port 2 nsew signal input
rlabel locali s 483 215 549 289 6 B1
port 3 nsew signal input
rlabel locali s 205 289 549 323 6 B1
port 3 nsew signal input
rlabel locali s 205 215 304 289 6 B1
port 3 nsew signal input
rlabel locali s 338 215 449 255 6 B2
port 4 nsew signal input
rlabel locali s 18 215 88 255 6 C1
port 5 nsew signal input
rlabel locali s 1315 181 1384 289 6 X
port 6 nsew signal output
rlabel locali s 1223 323 1273 493 6 X
port 6 nsew signal output
rlabel locali s 1215 51 1281 145 6 X
port 6 nsew signal output
rlabel locali s 1146 323 1180 357 6 X
port 6 nsew signal output
rlabel locali s 1146 289 1384 323 6 X
port 6 nsew signal output
rlabel locali s 1063 391 1105 493 6 X
port 6 nsew signal output
rlabel locali s 1063 357 1180 391 6 X
port 6 nsew signal output
rlabel locali s 1047 147 1384 181 6 X
port 6 nsew signal output
rlabel locali s 1047 145 1281 147 6 X
port 6 nsew signal output
rlabel locali s 1047 51 1113 145 6 X
port 6 nsew signal output
rlabel locali s 1315 17 1366 113 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1147 17 1181 111 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 979 17 1013 181 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 811 17 845 111 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 629 17 677 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 1472 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1472 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1307 359 1357 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1139 425 1189 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 971 425 1021 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 533 425 685 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 197 425 247 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 29 291 79 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 1472 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 1472 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1472 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1438068
string GDS_START 1427258
<< end >>
