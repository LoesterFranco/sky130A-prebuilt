magic
tech sky130A
magscale 1 2
timestamp 1601050082
<< locali >>
rect 113 390 179 596
rect 313 390 379 596
rect 537 472 1181 506
rect 113 356 379 390
rect 537 356 571 472
rect 113 330 179 356
rect 25 296 179 330
rect 25 262 71 296
rect 25 228 203 262
rect 505 290 571 356
rect 1147 370 1181 472
rect 137 222 203 228
rect 785 254 851 356
rect 899 336 1181 370
rect 1215 356 1281 360
rect 899 290 965 336
rect 1215 316 1607 356
rect 1013 236 1147 302
rect 1215 226 1281 316
rect 1513 290 1607 316
rect 1369 224 1459 282
rect 137 188 403 222
rect 137 70 203 188
rect 337 70 403 188
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 23 364 73 649
rect 213 424 279 649
rect 417 390 483 649
rect 531 540 805 592
rect 839 540 905 649
rect 957 540 1249 596
rect 1361 546 1427 649
rect 1215 512 1249 540
rect 1543 512 1609 596
rect 1215 478 1609 512
rect 251 256 471 322
rect 646 404 1113 438
rect 646 384 715 404
rect 646 256 712 384
rect 1231 440 1335 444
rect 1231 394 1519 440
rect 1453 390 1519 394
rect 1553 390 1609 478
rect 437 222 712 256
rect 37 17 103 194
rect 660 220 712 222
rect 237 17 303 154
rect 448 17 514 188
rect 560 85 626 188
rect 660 186 912 220
rect 660 119 712 186
rect 746 85 812 152
rect 846 119 912 186
rect 946 192 1012 202
rect 946 190 1212 192
rect 1543 190 1609 206
rect 946 158 1609 190
rect 946 85 1012 158
rect 1146 156 1609 158
rect 560 51 1012 85
rect 1046 17 1112 124
rect 1146 70 1212 156
rect 1246 17 1312 122
rect 1348 70 1398 156
rect 1432 17 1509 120
rect 1543 70 1609 156
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
rlabel locali s 1369 224 1459 282 6 A1
port 1 nsew signal input
rlabel locali s 1513 290 1607 316 6 A2
port 2 nsew signal input
rlabel locali s 1215 356 1281 360 6 A2
port 2 nsew signal input
rlabel locali s 1215 316 1607 356 6 A2
port 2 nsew signal input
rlabel locali s 1215 226 1281 316 6 A2
port 2 nsew signal input
rlabel locali s 1013 236 1147 302 6 A3
port 3 nsew signal input
rlabel locali s 1147 370 1181 472 6 B1
port 4 nsew signal input
rlabel locali s 899 336 1181 370 6 B1
port 4 nsew signal input
rlabel locali s 899 290 965 336 6 B1
port 4 nsew signal input
rlabel locali s 537 472 1181 506 6 B1
port 4 nsew signal input
rlabel locali s 537 356 571 472 6 B1
port 4 nsew signal input
rlabel locali s 505 290 571 356 6 B1
port 4 nsew signal input
rlabel locali s 785 254 851 356 6 B2
port 5 nsew signal input
rlabel locali s 337 70 403 188 6 X
port 6 nsew signal output
rlabel locali s 313 390 379 596 6 X
port 6 nsew signal output
rlabel locali s 137 222 203 228 6 X
port 6 nsew signal output
rlabel locali s 137 188 403 222 6 X
port 6 nsew signal output
rlabel locali s 137 70 203 188 6 X
port 6 nsew signal output
rlabel locali s 113 390 179 596 6 X
port 6 nsew signal output
rlabel locali s 113 356 379 390 6 X
port 6 nsew signal output
rlabel locali s 113 330 179 356 6 X
port 6 nsew signal output
rlabel locali s 25 296 179 330 6 X
port 6 nsew signal output
rlabel locali s 25 262 71 296 6 X
port 6 nsew signal output
rlabel locali s 25 228 203 262 6 X
port 6 nsew signal output
rlabel metal1 s 0 -49 1632 49 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1632 715 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 875358
string GDS_START 862596
<< end >>
