magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 276 561
rect 17 333 69 527
rect 17 75 65 265
rect 103 258 169 493
rect 203 333 259 527
rect 103 152 259 258
rect 103 51 168 152
rect 202 17 259 118
rect 0 -17 276 17
<< metal1 >>
rect 0 496 276 592
rect 0 -48 276 48
<< labels >>
rlabel locali s 17 75 65 265 6 A
port 1 nsew signal input
rlabel locali s 103 258 169 493 6 Y
port 2 nsew signal output
rlabel locali s 103 152 259 258 6 Y
port 2 nsew signal output
rlabel locali s 103 51 168 152 6 Y
port 2 nsew signal output
rlabel locali s 202 17 259 118 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 0 -17 276 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 276 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 203 333 259 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 17 333 69 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 0 527 276 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 496 276 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 276 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3202140
string GDS_START 3198366
<< end >>
