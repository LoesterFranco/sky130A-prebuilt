magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 17 289 367 323
rect 17 215 125 289
rect 171 215 289 255
rect 333 249 367 289
rect 1165 391 1215 493
rect 1353 391 1403 493
rect 1165 357 1403 391
rect 1353 331 1403 357
rect 333 215 419 249
rect 755 289 1093 323
rect 755 265 801 289
rect 723 215 801 265
rect 841 215 983 255
rect 1017 215 1093 289
rect 1353 283 1535 331
rect 1462 181 1535 283
rect 1147 145 1535 181
rect 1147 55 1223 145
rect 1335 55 1411 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 27 391 77 493
rect 121 425 171 527
rect 215 391 265 493
rect 309 425 359 527
rect 403 459 641 493
rect 403 391 453 459
rect 591 427 641 459
rect 695 427 745 527
rect 789 459 1027 493
rect 789 427 839 459
rect 27 357 453 391
rect 411 291 453 357
rect 497 393 547 425
rect 883 393 933 425
rect 497 283 574 393
rect 687 357 933 393
rect 977 357 1027 459
rect 1071 359 1121 527
rect 1259 433 1309 527
rect 1447 365 1497 527
rect 687 333 721 357
rect 651 299 721 333
rect 497 181 539 283
rect 651 249 689 299
rect 573 215 689 249
rect 1127 249 1202 323
rect 1127 215 1418 249
rect 651 181 689 215
rect 35 17 69 179
rect 103 95 163 181
rect 197 147 555 181
rect 197 129 274 147
rect 103 51 367 95
rect 411 17 445 111
rect 479 51 555 147
rect 651 145 1035 181
rect 599 17 737 111
rect 771 51 847 145
rect 891 17 925 111
rect 959 51 1035 145
rect 1079 17 1113 179
rect 1267 17 1301 111
rect 1455 17 1489 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
<< metal1 >>
rect 0 561 1564 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 0 496 1564 527
rect 0 17 1564 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
rect 0 -48 1564 -17
<< obsm1 >>
rect 528 320 596 329
rect 1134 320 1192 329
rect 528 292 1192 320
rect 528 283 596 292
rect 1134 283 1192 292
<< labels >>
rlabel locali s 1017 215 1093 289 6 A1_N
port 1 nsew signal input
rlabel locali s 755 289 1093 323 6 A1_N
port 1 nsew signal input
rlabel locali s 755 265 801 289 6 A1_N
port 1 nsew signal input
rlabel locali s 723 215 801 265 6 A1_N
port 1 nsew signal input
rlabel locali s 841 215 983 255 6 A2_N
port 2 nsew signal input
rlabel locali s 333 249 367 289 6 B1
port 3 nsew signal input
rlabel locali s 333 215 419 249 6 B1
port 3 nsew signal input
rlabel locali s 17 289 367 323 6 B1
port 3 nsew signal input
rlabel locali s 17 215 125 289 6 B1
port 3 nsew signal input
rlabel locali s 171 215 289 255 6 B2
port 4 nsew signal input
rlabel locali s 1462 181 1535 283 6 X
port 5 nsew signal output
rlabel locali s 1353 391 1403 493 6 X
port 5 nsew signal output
rlabel locali s 1353 331 1403 357 6 X
port 5 nsew signal output
rlabel locali s 1353 283 1535 331 6 X
port 5 nsew signal output
rlabel locali s 1335 55 1411 145 6 X
port 5 nsew signal output
rlabel locali s 1165 391 1215 493 6 X
port 5 nsew signal output
rlabel locali s 1165 357 1403 391 6 X
port 5 nsew signal output
rlabel locali s 1147 145 1535 181 6 X
port 5 nsew signal output
rlabel locali s 1147 55 1223 145 6 X
port 5 nsew signal output
rlabel metal1 s 0 -48 1564 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 1564 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1564 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1332082
string GDS_START 1320070
<< end >>
