magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 1862 704
<< pwell >>
rect 0 0 1824 49
<< scnmos >>
rect 96 74 126 222
rect 350 74 380 222
rect 436 74 466 222
rect 522 74 552 222
rect 622 74 652 222
rect 708 74 738 222
rect 808 74 838 222
rect 894 74 924 222
rect 980 74 1010 222
rect 1066 74 1096 222
rect 1152 74 1182 222
rect 1238 74 1268 222
rect 1324 74 1354 222
rect 1424 74 1454 222
rect 1510 74 1540 222
rect 1596 74 1626 222
rect 1710 74 1740 222
<< pmoshvt >>
rect 96 368 126 592
rect 298 368 328 592
rect 398 368 428 592
rect 488 368 518 592
rect 588 368 618 592
rect 678 368 708 592
rect 778 368 808 592
rect 868 368 898 592
rect 978 368 1008 592
rect 1068 368 1098 592
rect 1158 368 1188 592
rect 1248 368 1278 592
rect 1348 368 1378 592
rect 1438 368 1468 592
rect 1528 368 1558 592
rect 1618 368 1648 592
rect 1708 368 1738 592
<< ndiff >>
rect 39 196 96 222
rect 39 162 51 196
rect 85 162 96 196
rect 39 120 96 162
rect 39 86 51 120
rect 85 86 96 120
rect 39 74 96 86
rect 126 210 183 222
rect 126 176 137 210
rect 171 176 183 210
rect 126 120 183 176
rect 126 86 137 120
rect 171 86 183 120
rect 126 74 183 86
rect 293 210 350 222
rect 293 176 305 210
rect 339 176 350 210
rect 293 120 350 176
rect 293 86 305 120
rect 339 86 350 120
rect 293 74 350 86
rect 380 210 436 222
rect 380 176 391 210
rect 425 176 436 210
rect 380 120 436 176
rect 380 86 391 120
rect 425 86 436 120
rect 380 74 436 86
rect 466 210 522 222
rect 466 176 477 210
rect 511 176 522 210
rect 466 120 522 176
rect 466 86 477 120
rect 511 86 522 120
rect 466 74 522 86
rect 552 210 622 222
rect 552 176 563 210
rect 597 176 622 210
rect 552 120 622 176
rect 552 86 563 120
rect 597 86 622 120
rect 552 74 622 86
rect 652 210 708 222
rect 652 176 663 210
rect 697 176 708 210
rect 652 120 708 176
rect 652 86 663 120
rect 697 86 708 120
rect 652 74 708 86
rect 738 210 808 222
rect 738 176 749 210
rect 783 176 808 210
rect 738 120 808 176
rect 738 86 749 120
rect 783 86 808 120
rect 738 74 808 86
rect 838 210 894 222
rect 838 176 849 210
rect 883 176 894 210
rect 838 120 894 176
rect 838 86 849 120
rect 883 86 894 120
rect 838 74 894 86
rect 924 192 980 222
rect 924 158 935 192
rect 969 158 980 192
rect 924 120 980 158
rect 924 86 935 120
rect 969 86 980 120
rect 924 74 980 86
rect 1010 210 1066 222
rect 1010 176 1021 210
rect 1055 176 1066 210
rect 1010 120 1066 176
rect 1010 86 1021 120
rect 1055 86 1066 120
rect 1010 74 1066 86
rect 1096 207 1152 222
rect 1096 173 1107 207
rect 1141 173 1152 207
rect 1096 74 1152 173
rect 1182 120 1238 222
rect 1182 86 1193 120
rect 1227 86 1238 120
rect 1182 74 1238 86
rect 1268 199 1324 222
rect 1268 165 1279 199
rect 1313 165 1324 199
rect 1268 74 1324 165
rect 1354 149 1424 222
rect 1354 115 1379 149
rect 1413 115 1424 149
rect 1354 74 1424 115
rect 1454 173 1510 222
rect 1454 139 1465 173
rect 1499 139 1510 173
rect 1454 74 1510 139
rect 1540 149 1596 222
rect 1540 115 1551 149
rect 1585 115 1596 149
rect 1540 74 1596 115
rect 1626 173 1710 222
rect 1626 139 1651 173
rect 1685 139 1710 173
rect 1626 74 1710 139
rect 1740 210 1797 222
rect 1740 176 1751 210
rect 1785 176 1797 210
rect 1740 120 1797 176
rect 1740 86 1751 120
rect 1785 86 1797 120
rect 1740 74 1797 86
<< pdiff >>
rect 27 580 96 592
rect 27 546 39 580
rect 73 546 96 580
rect 27 497 96 546
rect 27 463 39 497
rect 73 463 96 497
rect 27 414 96 463
rect 27 380 39 414
rect 73 380 96 414
rect 27 368 96 380
rect 126 580 185 592
rect 126 546 139 580
rect 173 546 185 580
rect 126 497 185 546
rect 126 463 139 497
rect 173 463 185 497
rect 126 414 185 463
rect 126 380 139 414
rect 173 380 185 414
rect 126 368 185 380
rect 239 580 298 592
rect 239 546 251 580
rect 285 546 298 580
rect 239 510 298 546
rect 239 476 251 510
rect 285 476 298 510
rect 239 440 298 476
rect 239 406 251 440
rect 285 406 298 440
rect 239 368 298 406
rect 328 580 398 592
rect 328 546 341 580
rect 375 546 398 580
rect 328 504 398 546
rect 328 470 341 504
rect 375 470 398 504
rect 328 435 398 470
rect 328 401 341 435
rect 375 401 398 435
rect 328 368 398 401
rect 428 580 488 592
rect 428 546 441 580
rect 475 546 488 580
rect 428 510 488 546
rect 428 476 441 510
rect 475 476 488 510
rect 428 440 488 476
rect 428 406 441 440
rect 475 406 488 440
rect 428 368 488 406
rect 518 580 588 592
rect 518 546 531 580
rect 565 546 588 580
rect 518 504 588 546
rect 518 470 531 504
rect 565 470 588 504
rect 518 435 588 470
rect 518 401 531 435
rect 565 401 588 435
rect 518 368 588 401
rect 618 580 678 592
rect 618 546 631 580
rect 665 546 678 580
rect 618 510 678 546
rect 618 476 631 510
rect 665 476 678 510
rect 618 440 678 476
rect 618 406 631 440
rect 665 406 678 440
rect 618 368 678 406
rect 708 580 778 592
rect 708 546 721 580
rect 755 546 778 580
rect 708 504 778 546
rect 708 470 721 504
rect 755 470 778 504
rect 708 435 778 470
rect 708 401 721 435
rect 755 401 778 435
rect 708 368 778 401
rect 808 580 868 592
rect 808 546 821 580
rect 855 546 868 580
rect 808 510 868 546
rect 808 476 821 510
rect 855 476 868 510
rect 808 440 868 476
rect 808 406 821 440
rect 855 406 868 440
rect 808 368 868 406
rect 898 580 978 592
rect 898 546 921 580
rect 955 546 978 580
rect 898 508 978 546
rect 898 474 921 508
rect 955 474 978 508
rect 898 368 978 474
rect 1008 580 1068 592
rect 1008 546 1021 580
rect 1055 546 1068 580
rect 1008 510 1068 546
rect 1008 476 1021 510
rect 1055 476 1068 510
rect 1008 440 1068 476
rect 1008 406 1021 440
rect 1055 406 1068 440
rect 1008 368 1068 406
rect 1098 531 1158 592
rect 1098 497 1111 531
rect 1145 497 1158 531
rect 1098 414 1158 497
rect 1098 380 1111 414
rect 1145 380 1158 414
rect 1098 368 1158 380
rect 1188 580 1248 592
rect 1188 546 1201 580
rect 1235 546 1248 580
rect 1188 508 1248 546
rect 1188 474 1201 508
rect 1235 474 1248 508
rect 1188 368 1248 474
rect 1278 540 1348 592
rect 1278 506 1301 540
rect 1335 506 1348 540
rect 1278 424 1348 506
rect 1278 390 1301 424
rect 1335 390 1348 424
rect 1278 368 1348 390
rect 1378 580 1438 592
rect 1378 546 1391 580
rect 1425 546 1438 580
rect 1378 508 1438 546
rect 1378 474 1391 508
rect 1425 474 1438 508
rect 1378 368 1438 474
rect 1468 540 1528 592
rect 1468 506 1481 540
rect 1515 506 1528 540
rect 1468 424 1528 506
rect 1468 390 1481 424
rect 1515 390 1528 424
rect 1468 368 1528 390
rect 1558 580 1618 592
rect 1558 546 1571 580
rect 1605 546 1618 580
rect 1558 508 1618 546
rect 1558 474 1571 508
rect 1605 474 1618 508
rect 1558 368 1618 474
rect 1648 540 1708 592
rect 1648 506 1661 540
rect 1695 506 1708 540
rect 1648 424 1708 506
rect 1648 390 1661 424
rect 1695 390 1708 424
rect 1648 368 1708 390
rect 1738 580 1797 592
rect 1738 546 1751 580
rect 1785 546 1797 580
rect 1738 510 1797 546
rect 1738 476 1751 510
rect 1785 476 1797 510
rect 1738 440 1797 476
rect 1738 406 1751 440
rect 1785 406 1797 440
rect 1738 368 1797 406
<< ndiffc >>
rect 51 162 85 196
rect 51 86 85 120
rect 137 176 171 210
rect 137 86 171 120
rect 305 176 339 210
rect 305 86 339 120
rect 391 176 425 210
rect 391 86 425 120
rect 477 176 511 210
rect 477 86 511 120
rect 563 176 597 210
rect 563 86 597 120
rect 663 176 697 210
rect 663 86 697 120
rect 749 176 783 210
rect 749 86 783 120
rect 849 176 883 210
rect 849 86 883 120
rect 935 158 969 192
rect 935 86 969 120
rect 1021 176 1055 210
rect 1021 86 1055 120
rect 1107 173 1141 207
rect 1193 86 1227 120
rect 1279 165 1313 199
rect 1379 115 1413 149
rect 1465 139 1499 173
rect 1551 115 1585 149
rect 1651 139 1685 173
rect 1751 176 1785 210
rect 1751 86 1785 120
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 139 546 173 580
rect 139 463 173 497
rect 139 380 173 414
rect 251 546 285 580
rect 251 476 285 510
rect 251 406 285 440
rect 341 546 375 580
rect 341 470 375 504
rect 341 401 375 435
rect 441 546 475 580
rect 441 476 475 510
rect 441 406 475 440
rect 531 546 565 580
rect 531 470 565 504
rect 531 401 565 435
rect 631 546 665 580
rect 631 476 665 510
rect 631 406 665 440
rect 721 546 755 580
rect 721 470 755 504
rect 721 401 755 435
rect 821 546 855 580
rect 821 476 855 510
rect 821 406 855 440
rect 921 546 955 580
rect 921 474 955 508
rect 1021 546 1055 580
rect 1021 476 1055 510
rect 1021 406 1055 440
rect 1111 497 1145 531
rect 1111 380 1145 414
rect 1201 546 1235 580
rect 1201 474 1235 508
rect 1301 506 1335 540
rect 1301 390 1335 424
rect 1391 546 1425 580
rect 1391 474 1425 508
rect 1481 506 1515 540
rect 1481 390 1515 424
rect 1571 546 1605 580
rect 1571 474 1605 508
rect 1661 506 1695 540
rect 1661 390 1695 424
rect 1751 546 1785 580
rect 1751 476 1785 510
rect 1751 406 1785 440
<< poly >>
rect 96 592 126 618
rect 298 592 328 618
rect 398 592 428 618
rect 488 592 518 618
rect 588 592 618 618
rect 678 592 708 618
rect 778 592 808 618
rect 868 592 898 618
rect 978 592 1008 618
rect 1068 592 1098 618
rect 1158 592 1188 618
rect 1248 592 1278 618
rect 1348 592 1378 618
rect 1438 592 1468 618
rect 1528 592 1558 618
rect 1618 592 1648 618
rect 1708 592 1738 618
rect 96 353 126 368
rect 298 353 328 368
rect 398 353 428 368
rect 488 353 518 368
rect 588 353 618 368
rect 678 353 708 368
rect 778 353 808 368
rect 868 353 898 368
rect 978 353 1008 368
rect 1068 353 1098 368
rect 1158 353 1188 368
rect 1248 353 1278 368
rect 1348 353 1378 368
rect 1438 353 1468 368
rect 1528 353 1558 368
rect 1618 353 1648 368
rect 1708 353 1738 368
rect 93 345 129 353
rect 295 345 331 353
rect 395 345 431 353
rect 485 345 521 353
rect 585 345 621 353
rect 675 345 711 353
rect 775 345 811 353
rect 865 345 901 353
rect 975 345 1011 353
rect 21 315 1011 345
rect 1065 336 1101 353
rect 1155 336 1191 353
rect 1245 336 1281 353
rect 1345 336 1381 353
rect 1435 336 1471 353
rect 1525 336 1561 353
rect 1615 336 1651 353
rect 1705 336 1741 353
rect 1065 320 1741 336
rect 21 310 129 315
rect 21 276 37 310
rect 71 276 129 310
rect 21 260 129 276
rect 1065 286 1215 320
rect 1249 286 1283 320
rect 1317 286 1351 320
rect 1385 286 1419 320
rect 1453 286 1487 320
rect 1521 286 1555 320
rect 1589 286 1623 320
rect 1657 286 1691 320
rect 1725 286 1741 320
rect 1065 270 1741 286
rect 96 222 126 260
rect 205 251 1010 267
rect 205 217 221 251
rect 255 237 1010 251
rect 255 217 271 237
rect 350 222 380 237
rect 436 222 466 237
rect 522 222 552 237
rect 622 222 652 237
rect 708 222 738 237
rect 808 222 838 237
rect 894 222 924 237
rect 980 222 1010 237
rect 1066 222 1096 270
rect 1152 222 1182 270
rect 1238 222 1268 270
rect 1324 222 1354 270
rect 1424 222 1454 270
rect 1510 222 1540 270
rect 1596 222 1626 270
rect 1710 222 1740 270
rect 205 183 271 217
rect 205 149 221 183
rect 255 149 271 183
rect 205 115 271 149
rect 205 81 221 115
rect 255 81 271 115
rect 96 48 126 74
rect 205 65 271 81
rect 350 48 380 74
rect 436 48 466 74
rect 522 48 552 74
rect 622 48 652 74
rect 708 48 738 74
rect 808 48 838 74
rect 894 48 924 74
rect 980 48 1010 74
rect 1066 48 1096 74
rect 1152 48 1182 74
rect 1238 48 1268 74
rect 1324 48 1354 74
rect 1424 48 1454 74
rect 1510 48 1540 74
rect 1596 48 1626 74
rect 1710 48 1740 74
<< polycont >>
rect 37 276 71 310
rect 1215 286 1249 320
rect 1283 286 1317 320
rect 1351 286 1385 320
rect 1419 286 1453 320
rect 1487 286 1521 320
rect 1555 286 1589 320
rect 1623 286 1657 320
rect 1691 286 1725 320
rect 221 217 255 251
rect 221 149 255 183
rect 221 81 255 115
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 23 580 89 649
rect 23 546 39 580
rect 73 546 89 580
rect 23 497 89 546
rect 23 463 39 497
rect 73 463 89 497
rect 23 414 89 463
rect 23 380 39 414
rect 73 380 89 414
rect 23 364 89 380
rect 123 580 189 596
rect 123 546 139 580
rect 173 546 189 580
rect 123 497 189 546
rect 123 463 139 497
rect 173 463 189 497
rect 123 414 189 463
rect 123 380 139 414
rect 173 380 189 414
rect 21 310 87 326
rect 21 276 37 310
rect 71 276 87 310
rect 21 236 87 276
rect 123 267 189 380
rect 235 580 285 596
rect 235 546 251 580
rect 235 510 285 546
rect 235 476 251 510
rect 235 440 285 476
rect 235 406 251 440
rect 235 367 285 406
rect 325 580 391 649
rect 325 546 341 580
rect 375 546 391 580
rect 325 504 391 546
rect 325 470 341 504
rect 375 470 391 504
rect 325 435 391 470
rect 325 401 341 435
rect 375 401 391 435
rect 425 580 475 596
rect 425 546 441 580
rect 425 510 475 546
rect 425 476 441 510
rect 425 440 475 476
rect 425 406 441 440
rect 425 367 475 406
rect 515 580 581 649
rect 515 546 531 580
rect 565 546 581 580
rect 515 504 581 546
rect 515 470 531 504
rect 565 470 581 504
rect 515 435 581 470
rect 515 401 531 435
rect 565 401 581 435
rect 615 580 665 596
rect 615 546 631 580
rect 615 510 665 546
rect 615 476 631 510
rect 615 440 665 476
rect 615 406 631 440
rect 615 367 665 406
rect 705 580 771 649
rect 705 546 721 580
rect 755 546 771 580
rect 705 504 771 546
rect 705 470 721 504
rect 755 470 771 504
rect 705 435 771 470
rect 705 401 721 435
rect 755 401 771 435
rect 805 580 871 596
rect 805 546 821 580
rect 855 546 871 580
rect 805 510 871 546
rect 805 476 821 510
rect 855 476 871 510
rect 805 440 871 476
rect 905 580 971 649
rect 905 546 921 580
rect 955 546 971 580
rect 905 508 971 546
rect 905 474 921 508
rect 955 474 971 508
rect 905 458 971 474
rect 1005 581 1801 615
rect 1005 580 1071 581
rect 1005 546 1021 580
rect 1055 546 1071 580
rect 1185 580 1251 581
rect 1005 510 1071 546
rect 1005 476 1021 510
rect 1055 476 1071 510
rect 805 406 821 440
rect 855 424 871 440
rect 1005 440 1071 476
rect 1005 424 1021 440
rect 855 406 1021 424
rect 1055 406 1071 440
rect 805 390 1071 406
rect 1111 531 1145 547
rect 1111 424 1145 497
rect 1185 546 1201 580
rect 1235 546 1251 580
rect 1391 580 1425 581
rect 1185 508 1251 546
rect 1185 474 1201 508
rect 1235 474 1251 508
rect 1185 458 1251 474
rect 1285 540 1351 547
rect 1285 506 1301 540
rect 1335 506 1351 540
rect 1285 424 1351 506
rect 1571 580 1605 581
rect 1391 508 1425 546
rect 1391 458 1425 474
rect 1465 540 1531 547
rect 1465 506 1481 540
rect 1515 506 1531 540
rect 1465 424 1531 506
rect 1751 580 1801 581
rect 1571 508 1605 546
rect 1571 458 1605 474
rect 1645 540 1711 547
rect 1645 506 1661 540
rect 1695 506 1711 540
rect 1645 424 1711 506
rect 1111 414 1301 424
rect 805 367 899 390
rect 235 333 899 367
rect 1145 390 1301 414
rect 1335 390 1481 424
rect 1515 390 1661 424
rect 1695 390 1711 424
rect 1785 546 1801 580
rect 1751 510 1801 546
rect 1785 476 1801 510
rect 1751 440 1801 476
rect 1785 406 1801 440
rect 1751 390 1801 406
rect 1111 356 1145 380
rect 985 310 1145 356
rect 305 276 883 294
rect 123 251 271 267
rect 123 226 221 251
rect 137 217 221 226
rect 255 217 271 251
rect 137 210 271 217
rect 35 196 101 198
rect 35 162 51 196
rect 85 162 101 196
rect 35 120 101 162
rect 35 86 51 120
rect 85 86 101 120
rect 35 17 101 86
rect 171 183 271 210
rect 171 176 221 183
rect 137 149 221 176
rect 255 149 271 183
rect 137 120 271 149
rect 171 115 271 120
rect 171 86 221 115
rect 137 81 221 86
rect 255 81 271 115
rect 137 65 271 81
rect 305 260 1055 276
rect 305 210 339 260
rect 305 120 339 176
rect 305 70 339 86
rect 375 210 425 226
rect 375 176 391 210
rect 375 120 425 176
rect 375 86 391 120
rect 375 17 425 86
rect 461 210 511 260
rect 461 176 477 210
rect 461 120 511 176
rect 461 86 477 120
rect 461 70 511 86
rect 547 210 613 226
rect 547 176 563 210
rect 597 176 613 210
rect 547 120 613 176
rect 547 86 563 120
rect 597 86 613 120
rect 547 17 613 86
rect 647 210 697 260
rect 833 242 1055 260
rect 647 176 663 210
rect 647 120 697 176
rect 647 86 663 120
rect 647 70 697 86
rect 733 210 799 226
rect 733 176 749 210
rect 783 176 799 210
rect 733 120 799 176
rect 733 86 749 120
rect 783 86 799 120
rect 733 17 799 86
rect 833 210 883 242
rect 833 176 849 210
rect 1021 210 1055 242
rect 833 120 883 176
rect 833 86 849 120
rect 833 70 883 86
rect 919 192 985 208
rect 919 158 935 192
rect 969 158 985 192
rect 919 120 985 158
rect 919 86 935 120
rect 969 86 985 120
rect 919 17 985 86
rect 1021 120 1055 176
rect 1091 226 1145 310
rect 1199 320 1799 356
rect 1199 286 1215 320
rect 1249 286 1283 320
rect 1317 286 1351 320
rect 1385 286 1419 320
rect 1453 286 1487 320
rect 1521 286 1555 320
rect 1589 286 1623 320
rect 1657 286 1691 320
rect 1725 286 1799 320
rect 1199 270 1799 286
rect 1263 226 1701 236
rect 1091 207 1701 226
rect 1091 173 1107 207
rect 1141 202 1701 207
rect 1141 199 1329 202
rect 1141 173 1279 199
rect 1091 165 1279 173
rect 1313 165 1329 199
rect 1465 173 1499 202
rect 1091 154 1329 165
rect 1363 149 1429 165
rect 1363 120 1379 149
rect 1055 86 1193 120
rect 1227 115 1379 120
rect 1413 115 1429 149
rect 1635 173 1701 202
rect 1465 123 1499 139
rect 1535 149 1601 165
rect 1227 86 1429 115
rect 1021 85 1429 86
rect 1535 115 1551 149
rect 1585 115 1601 149
rect 1635 139 1651 173
rect 1685 139 1701 173
rect 1635 123 1701 139
rect 1735 210 1801 226
rect 1735 176 1751 210
rect 1785 176 1801 210
rect 1535 85 1601 115
rect 1735 120 1801 176
rect 1735 86 1751 120
rect 1785 86 1801 120
rect 1735 85 1801 86
rect 1021 51 1801 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
<< metal1 >>
rect 0 683 1824 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 0 617 1824 649
rect 0 17 1824 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
rect 0 -49 1824 -17
<< labels >>
rlabel comment s 0 0 0 0 4 einvn_8
flabel pwell s 0 0 1824 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 0 617 1824 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 0 617 1824 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 1824 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 1375 316 1409 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 1471 316 1505 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 1567 316 1601 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 1663 316 1697 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 1759 316 1793 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 TE_B
port 2 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 Z
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 1824 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2110200
string GDS_START 2096102
<< end >>
