magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 920 561
rect 146 455 236 527
rect 349 455 415 527
rect 529 455 596 527
rect 701 455 767 527
rect 445 307 707 341
rect 204 145 247 268
rect 305 199 343 268
rect 654 169 707 307
rect 457 123 707 169
rect 743 123 799 341
rect 457 103 495 123
rect 356 17 422 89
rect 529 17 595 89
rect 629 51 667 123
rect 701 17 767 89
rect 0 -17 920 17
<< obsli1 >>
rect 30 299 102 433
rect 136 375 889 421
rect 30 161 74 299
rect 136 265 170 375
rect 256 305 411 339
rect 377 271 411 305
rect 108 199 170 265
rect 30 109 127 161
rect 377 204 620 271
rect 377 161 423 204
rect 284 123 423 161
rect 284 109 320 123
rect 30 71 320 109
rect 30 51 127 71
rect 833 85 889 375
<< metal1 >>
rect 0 496 920 592
rect 0 -48 920 48
<< labels >>
rlabel locali s 743 123 799 341 6 A_N
port 1 nsew signal input
rlabel locali s 204 145 247 268 6 B
port 2 nsew signal input
rlabel locali s 305 199 343 268 6 C
port 3 nsew signal input
rlabel locali s 654 169 707 307 6 X
port 4 nsew signal output
rlabel locali s 629 51 667 123 6 X
port 4 nsew signal output
rlabel locali s 457 123 707 169 6 X
port 4 nsew signal output
rlabel locali s 457 103 495 123 6 X
port 4 nsew signal output
rlabel locali s 445 307 707 341 6 X
port 4 nsew signal output
rlabel locali s 701 17 767 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 529 17 595 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 356 17 422 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 920 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 920 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 701 455 767 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 529 455 596 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 349 455 415 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 146 455 236 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 920 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 920 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 920 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3827886
string GDS_START 3821302
<< end >>
