magic
tech sky130A
magscale 1 2
timestamp 1599588218
<< nwell >>
rect -38 388 902 704
rect -38 332 274 388
rect 644 332 902 388
<< pwell >>
rect 0 0 864 49
<< scpmos >>
rect 83 424 119 592
rect 193 424 229 592
rect 299 424 335 592
rect 513 424 549 592
rect 613 424 649 592
rect 745 368 781 592
<< nmoslvt >>
rect 84 74 114 184
rect 323 124 353 252
rect 418 139 448 267
rect 496 139 526 267
rect 634 120 664 248
rect 750 100 780 248
<< ndiff >>
rect 27 146 84 184
rect 27 112 39 146
rect 73 112 84 146
rect 27 74 84 112
rect 114 120 167 184
rect 114 86 125 120
rect 159 86 167 120
rect 114 74 167 86
rect 368 252 418 267
rect 266 240 323 252
rect 266 206 278 240
rect 312 206 323 240
rect 266 170 323 206
rect 266 136 278 170
rect 312 136 323 170
rect 266 124 323 136
rect 353 139 418 252
rect 448 139 496 267
rect 526 248 576 267
rect 526 139 634 248
rect 353 124 403 139
rect 584 120 634 139
rect 664 192 750 248
rect 664 158 691 192
rect 725 158 750 192
rect 664 120 750 158
rect 679 100 750 120
rect 780 220 837 248
rect 780 186 791 220
rect 825 186 837 220
rect 780 146 837 186
rect 780 112 791 146
rect 825 112 837 146
rect 780 100 837 112
<< pdiff >>
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 470 83 546
rect 27 436 39 470
rect 73 436 83 470
rect 27 424 83 436
rect 119 584 193 592
rect 119 550 139 584
rect 173 550 193 584
rect 119 508 193 550
rect 119 474 139 508
rect 173 474 193 508
rect 119 424 193 474
rect 229 476 299 592
rect 229 442 242 476
rect 276 442 299 476
rect 229 424 299 442
rect 335 554 513 592
rect 335 520 345 554
rect 379 520 469 554
rect 503 520 513 554
rect 335 424 513 520
rect 549 580 613 592
rect 549 546 569 580
rect 603 546 613 580
rect 549 470 613 546
rect 549 436 569 470
rect 603 436 613 470
rect 549 424 613 436
rect 649 580 745 592
rect 649 546 683 580
rect 717 546 745 580
rect 649 470 745 546
rect 649 436 683 470
rect 717 436 745 470
rect 649 424 745 436
rect 695 368 745 424
rect 781 580 837 592
rect 781 546 791 580
rect 825 546 837 580
rect 781 500 837 546
rect 781 466 791 500
rect 825 466 837 500
rect 781 420 837 466
rect 781 386 791 420
rect 825 386 837 420
rect 781 368 837 386
<< ndiffc >>
rect 39 112 73 146
rect 125 86 159 120
rect 278 206 312 240
rect 278 136 312 170
rect 691 158 725 192
rect 791 186 825 220
rect 791 112 825 146
<< pdiffc >>
rect 39 546 73 580
rect 39 436 73 470
rect 139 550 173 584
rect 139 474 173 508
rect 242 442 276 476
rect 345 520 379 554
rect 469 520 503 554
rect 569 546 603 580
rect 569 436 603 470
rect 683 546 717 580
rect 683 436 717 470
rect 791 546 825 580
rect 791 466 825 500
rect 791 386 825 420
<< poly >>
rect 83 592 119 618
rect 193 592 229 618
rect 299 592 335 618
rect 513 592 549 618
rect 613 592 649 618
rect 745 592 781 618
rect 83 372 119 424
rect 193 376 229 424
rect 299 392 335 424
rect 299 376 448 392
rect 53 356 119 372
rect 53 322 69 356
rect 103 322 119 356
rect 53 288 119 322
rect 185 360 251 376
rect 185 326 201 360
rect 235 326 251 360
rect 299 342 329 376
rect 363 342 398 376
rect 432 342 448 376
rect 299 326 448 342
rect 185 310 251 326
rect 53 254 69 288
rect 103 254 119 288
rect 53 238 119 254
rect 84 184 114 238
rect 221 109 251 310
rect 323 252 353 278
rect 418 267 448 326
rect 513 312 549 424
rect 613 376 649 424
rect 496 282 549 312
rect 597 360 664 376
rect 597 326 613 360
rect 647 326 664 360
rect 745 336 781 368
rect 597 310 664 326
rect 496 267 526 282
rect 634 248 664 310
rect 712 320 781 336
rect 712 286 728 320
rect 762 286 781 320
rect 712 270 781 286
rect 750 248 780 270
rect 323 109 353 124
rect 418 113 448 139
rect 496 117 526 139
rect 221 79 353 109
rect 496 101 562 117
rect 84 48 114 74
rect 496 67 512 101
rect 546 67 562 101
rect 634 94 664 120
rect 750 74 780 100
rect 496 51 562 67
<< polycont >>
rect 69 322 103 356
rect 201 326 235 360
rect 329 342 363 376
rect 398 342 432 376
rect 69 254 103 288
rect 613 326 647 360
rect 728 286 762 320
rect 512 67 546 101
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 23 580 89 596
rect 23 546 39 580
rect 73 546 89 580
rect 23 470 89 546
rect 123 584 189 649
rect 123 550 139 584
rect 173 550 189 584
rect 123 508 189 550
rect 123 474 139 508
rect 173 474 189 508
rect 329 554 519 649
rect 329 520 345 554
rect 379 520 469 554
rect 503 520 519 554
rect 329 507 519 520
rect 553 580 619 596
rect 553 546 569 580
rect 603 546 619 580
rect 223 476 292 492
rect 23 436 39 470
rect 73 440 89 470
rect 223 442 242 476
rect 276 470 292 476
rect 553 470 619 546
rect 276 442 569 470
rect 73 436 189 440
rect 23 406 189 436
rect 223 436 569 442
rect 603 436 619 470
rect 223 426 619 436
rect 155 376 189 406
rect 519 420 619 426
rect 667 580 733 649
rect 667 546 683 580
rect 717 546 733 580
rect 667 470 733 546
rect 667 436 683 470
rect 717 436 733 470
rect 667 420 733 436
rect 775 580 846 596
rect 775 546 791 580
rect 825 546 846 580
rect 775 500 846 546
rect 775 466 791 500
rect 825 466 846 500
rect 775 420 846 466
rect 313 376 455 392
rect 25 356 119 372
rect 25 322 69 356
rect 103 322 119 356
rect 25 288 119 322
rect 25 254 69 288
rect 103 254 119 288
rect 25 238 119 254
rect 155 360 251 376
rect 155 326 201 360
rect 235 326 251 360
rect 155 310 251 326
rect 313 342 329 376
rect 363 342 398 376
rect 432 342 455 376
rect 313 310 455 342
rect 155 204 189 310
rect 519 276 553 420
rect 775 386 791 420
rect 825 386 846 420
rect 597 360 663 376
rect 775 370 846 386
rect 597 326 613 360
rect 647 326 663 360
rect 597 310 663 326
rect 707 320 778 336
rect 707 286 728 320
rect 762 286 778 320
rect 707 276 778 286
rect 23 170 189 204
rect 262 270 778 276
rect 262 242 741 270
rect 262 240 328 242
rect 262 206 278 240
rect 312 206 328 240
rect 812 236 846 370
rect 775 220 846 236
rect 262 170 328 206
rect 23 146 81 170
rect 23 112 39 146
rect 73 112 81 146
rect 262 136 278 170
rect 312 136 328 170
rect 23 70 81 112
rect 115 120 175 136
rect 262 120 328 136
rect 675 192 741 208
rect 675 158 691 192
rect 725 158 741 192
rect 115 86 125 120
rect 159 86 175 120
rect 115 17 175 86
rect 409 101 562 134
rect 409 67 512 101
rect 546 67 562 101
rect 409 51 562 67
rect 675 17 741 158
rect 775 186 791 220
rect 825 186 846 220
rect 775 146 846 186
rect 775 112 791 146
rect 825 112 846 146
rect 775 96 846 112
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
rlabel comment s 0 0 0 0 4 and4b_1
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 799 390 833 424 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 799 464 833 498 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 799 538 833 572 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 D
port 4 nsew
flabel corelocali s 415 94 449 128 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 511 94 545 128 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 B
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 864 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3273720
string GDS_START 3266026
<< end >>
