magic
tech sky130A
magscale 1 2
timestamp 1604502729
<< locali >>
rect 372 390 463 596
rect 21 236 87 302
rect 121 224 220 290
rect 372 236 406 390
rect 445 260 551 356
rect 585 260 651 356
rect 322 202 406 236
rect 322 70 372 202
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 28 379 94 649
rect 128 358 194 555
rect 228 395 338 649
rect 599 390 649 649
rect 128 324 338 358
rect 254 270 338 324
rect 254 190 288 270
rect 23 17 89 190
rect 187 70 288 190
rect 440 192 644 226
rect 440 168 474 192
rect 406 89 474 168
rect 508 17 542 158
rect 578 70 644 192
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel locali s 21 236 87 302 6 A1_N
port 1 nsew signal input
rlabel locali s 121 224 220 290 6 A2_N
port 2 nsew signal input
rlabel locali s 585 260 651 356 6 B1
port 3 nsew signal input
rlabel locali s 445 260 551 356 6 B2
port 4 nsew signal input
rlabel locali s 372 390 463 596 6 Y
port 5 nsew signal output
rlabel locali s 372 236 406 390 6 Y
port 5 nsew signal output
rlabel locali s 322 202 406 236 6 Y
port 5 nsew signal output
rlabel locali s 322 70 372 202 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -49 672 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 672 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1233306
string GDS_START 1226706
<< end >>
