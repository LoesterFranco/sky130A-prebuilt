magic
tech sky130A
magscale 1 2
timestamp 1601050088
<< locali >>
rect 123 378 189 596
rect 430 430 486 547
rect 610 430 666 547
rect 430 378 666 430
rect 123 344 666 378
rect 25 236 229 310
rect 295 202 361 344
rect 409 236 632 310
rect 125 168 361 202
rect 125 119 159 168
rect 295 119 361 168
rect 879 236 1223 310
rect 1273 236 1607 310
rect 1657 236 1991 310
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 23 364 89 649
rect 223 412 289 649
rect 335 581 1141 615
rect 335 412 396 581
rect 520 464 576 581
rect 700 360 761 581
rect 795 378 861 547
rect 895 412 961 581
rect 995 378 1041 547
rect 1075 412 1141 581
rect 1187 581 1603 615
rect 1187 578 1433 581
rect 1187 412 1253 578
rect 1287 378 1333 544
rect 1367 412 1433 578
rect 1467 378 1513 547
rect 795 344 1513 378
rect 1547 378 1603 581
rect 1637 412 1703 649
rect 1737 378 1803 600
rect 1837 412 1903 649
rect 1937 378 1993 600
rect 1547 344 1993 378
rect 666 260 838 294
rect 666 202 700 260
rect 23 85 89 202
rect 195 85 261 134
rect 395 168 700 202
rect 395 85 461 168
rect 23 51 461 85
rect 495 17 598 120
rect 632 70 700 168
rect 734 17 768 226
rect 804 202 838 260
rect 804 168 1993 202
rect 804 70 870 168
rect 904 17 970 134
rect 1006 70 1056 168
rect 1090 17 1156 134
rect 1192 70 1242 168
rect 1276 17 1342 134
rect 1378 70 1412 168
rect 1448 17 1514 134
rect 1557 70 1607 168
rect 1641 17 1707 134
rect 1741 70 1807 168
rect 1841 17 1907 134
rect 1943 70 1993 168
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
rlabel locali s 1657 236 1991 310 6 A1
port 1 nsew signal input
rlabel locali s 1273 236 1607 310 6 A2
port 2 nsew signal input
rlabel locali s 879 236 1223 310 6 A3
port 3 nsew signal input
rlabel locali s 409 236 632 310 6 A4
port 4 nsew signal input
rlabel locali s 25 236 229 310 6 B1
port 5 nsew signal input
rlabel locali s 610 430 666 547 6 Y
port 6 nsew signal output
rlabel locali s 430 430 486 547 6 Y
port 6 nsew signal output
rlabel locali s 430 378 666 430 6 Y
port 6 nsew signal output
rlabel locali s 295 202 361 344 6 Y
port 6 nsew signal output
rlabel locali s 295 119 361 168 6 Y
port 6 nsew signal output
rlabel locali s 125 168 361 202 6 Y
port 6 nsew signal output
rlabel locali s 125 119 159 168 6 Y
port 6 nsew signal output
rlabel locali s 123 378 189 596 6 Y
port 6 nsew signal output
rlabel locali s 123 344 666 378 6 Y
port 6 nsew signal output
rlabel metal1 s 0 -49 2016 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 617 2016 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2016 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 793602
string GDS_START 777448
<< end >>
