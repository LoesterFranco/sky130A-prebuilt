magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 552 561
rect 17 269 71 489
rect 194 375 260 527
rect 294 325 359 493
rect 17 199 107 269
rect 237 291 359 325
rect 454 307 529 527
rect 237 165 271 291
rect 305 215 405 257
rect 439 215 535 257
rect 17 17 72 165
rect 223 129 271 165
rect 223 51 257 129
rect 399 17 433 111
rect 0 -17 552 17
<< obsli1 >>
rect 105 341 160 442
rect 105 307 203 341
rect 144 199 203 307
rect 144 165 178 199
rect 116 131 178 165
rect 116 99 154 131
rect 314 147 533 181
rect 314 97 348 147
rect 298 51 364 97
rect 467 54 533 147
<< metal1 >>
rect 0 496 552 592
rect 0 -48 552 48
<< labels >>
rlabel locali s 439 215 535 257 6 A1
port 1 nsew signal input
rlabel locali s 305 215 405 257 6 A2
port 2 nsew signal input
rlabel locali s 17 269 71 489 6 B1_N
port 3 nsew signal input
rlabel locali s 17 199 107 269 6 B1_N
port 3 nsew signal input
rlabel locali s 294 325 359 493 6 Y
port 4 nsew signal output
rlabel locali s 237 291 359 325 6 Y
port 4 nsew signal output
rlabel locali s 237 165 271 291 6 Y
port 4 nsew signal output
rlabel locali s 223 129 271 165 6 Y
port 4 nsew signal output
rlabel locali s 223 51 257 129 6 Y
port 4 nsew signal output
rlabel locali s 399 17 433 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 17 17 72 165 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 552 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 552 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 454 307 529 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 194 375 260 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 552 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 552 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 552 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1394410
string GDS_START 1388898
<< end >>
