magic
tech sky130A
magscale 1 2
timestamp 1604502697
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 79 93 109 177
rect 267 47 297 177
rect 351 47 381 177
rect 435 47 465 177
rect 529 47 559 177
<< pmoshvt >>
rect 81 297 117 381
rect 189 297 225 497
rect 295 297 331 497
rect 425 297 461 497
rect 521 297 557 497
<< ndiff >>
rect 27 152 79 177
rect 27 118 35 152
rect 69 118 79 152
rect 27 93 79 118
rect 109 139 161 177
rect 109 105 119 139
rect 153 105 161 139
rect 109 93 161 105
rect 215 93 267 177
rect 215 59 223 93
rect 257 59 267 93
rect 215 47 267 59
rect 297 161 351 177
rect 297 127 307 161
rect 341 127 351 161
rect 297 47 351 127
rect 381 161 435 177
rect 381 127 391 161
rect 425 127 435 161
rect 381 93 435 127
rect 381 59 391 93
rect 425 59 435 93
rect 381 47 435 59
rect 465 89 529 177
rect 465 55 485 89
rect 519 55 529 89
rect 465 47 529 55
rect 559 161 611 177
rect 559 127 569 161
rect 603 127 611 161
rect 559 93 611 127
rect 559 59 569 93
rect 603 59 611 93
rect 559 47 611 59
<< pdiff >>
rect 135 485 189 497
rect 135 451 143 485
rect 177 451 189 485
rect 135 417 189 451
rect 135 383 143 417
rect 177 383 189 417
rect 135 381 189 383
rect 27 356 81 381
rect 27 322 35 356
rect 69 322 81 356
rect 27 297 81 322
rect 117 297 189 381
rect 225 485 295 497
rect 225 451 243 485
rect 277 451 295 485
rect 225 417 295 451
rect 225 383 243 417
rect 277 383 295 417
rect 225 297 295 383
rect 331 485 425 497
rect 331 451 367 485
rect 401 451 425 485
rect 331 297 425 451
rect 461 485 521 497
rect 461 451 473 485
rect 507 451 521 485
rect 461 417 521 451
rect 461 383 473 417
rect 507 383 521 417
rect 461 349 521 383
rect 461 315 473 349
rect 507 315 521 349
rect 461 297 521 315
rect 557 485 614 497
rect 557 451 569 485
rect 603 451 614 485
rect 557 417 614 451
rect 557 383 569 417
rect 603 383 614 417
rect 557 297 614 383
<< ndiffc >>
rect 35 118 69 152
rect 119 105 153 139
rect 223 59 257 93
rect 307 127 341 161
rect 391 127 425 161
rect 391 59 425 93
rect 485 55 519 89
rect 569 127 603 161
rect 569 59 603 93
<< pdiffc >>
rect 143 451 177 485
rect 143 383 177 417
rect 35 322 69 356
rect 243 451 277 485
rect 243 383 277 417
rect 367 451 401 485
rect 473 451 507 485
rect 473 383 507 417
rect 473 315 507 349
rect 569 451 603 485
rect 569 383 603 417
<< poly >>
rect 189 497 225 523
rect 295 497 331 523
rect 425 497 461 523
rect 521 497 557 523
rect 81 381 117 407
rect 81 282 117 297
rect 189 282 225 297
rect 295 282 331 297
rect 425 282 461 297
rect 521 282 557 297
rect 79 265 119 282
rect 79 249 145 265
rect 79 215 91 249
rect 125 215 145 249
rect 79 199 145 215
rect 187 259 227 282
rect 293 259 333 282
rect 423 259 463 282
rect 519 259 559 282
rect 187 249 381 259
rect 187 215 204 249
rect 238 215 381 249
rect 187 205 381 215
rect 423 249 559 259
rect 423 215 439 249
rect 473 215 507 249
rect 541 215 559 249
rect 423 205 559 215
rect 79 177 109 199
rect 267 177 297 205
rect 351 177 381 205
rect 435 177 465 205
rect 529 177 559 205
rect 79 67 109 93
rect 267 21 297 47
rect 351 21 381 47
rect 435 21 465 47
rect 529 21 559 47
<< polycont >>
rect 91 215 125 249
rect 204 215 238 249
rect 439 215 473 249
rect 507 215 541 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 126 485 177 527
rect 126 451 143 485
rect 126 417 177 451
rect 126 383 143 417
rect 22 356 82 372
rect 126 367 177 383
rect 227 485 293 493
rect 227 451 243 485
rect 277 451 293 485
rect 227 417 293 451
rect 345 485 420 527
rect 345 451 367 485
rect 401 451 420 485
rect 345 435 420 451
rect 457 485 523 493
rect 457 451 473 485
rect 507 451 523 485
rect 227 383 243 417
rect 277 401 293 417
rect 457 417 523 451
rect 457 401 473 417
rect 277 383 473 401
rect 507 383 523 417
rect 227 367 523 383
rect 569 485 603 527
rect 569 417 603 451
rect 569 367 603 383
rect 22 322 35 356
rect 69 333 82 356
rect 69 322 238 333
rect 22 299 238 322
rect 22 168 56 299
rect 91 249 170 265
rect 125 215 170 249
rect 91 199 170 215
rect 204 249 238 299
rect 204 199 238 215
rect 22 152 69 168
rect 291 161 357 367
rect 468 349 523 367
rect 468 315 473 349
rect 507 315 523 349
rect 468 299 523 315
rect 581 255 619 331
rect 422 249 619 255
rect 422 215 439 249
rect 473 215 507 249
rect 541 215 619 249
rect 22 118 35 152
rect 22 102 69 118
rect 119 139 153 155
rect 291 127 307 161
rect 341 127 357 161
rect 391 161 619 181
rect 425 139 569 161
rect 425 127 441 139
rect 119 17 153 105
rect 391 93 441 127
rect 553 127 569 139
rect 603 127 619 161
rect 207 59 223 93
rect 257 59 391 93
rect 425 59 441 93
rect 207 51 441 59
rect 485 89 519 105
rect 485 17 519 55
rect 553 93 619 127
rect 553 59 569 93
rect 603 59 619 93
rect 553 51 619 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel corelocali s 581 221 615 255 0 FreeSans 250 0 0 0 B
port 2 nsew
flabel corelocali s 486 221 520 255 0 FreeSans 250 0 0 0 B
port 2 nsew
flabel corelocali s 310 153 344 187 0 FreeSans 250 0 0 0 Y
port 7 nsew
flabel corelocali s 305 221 339 255 0 FreeSans 250 0 0 0 Y
port 7 nsew
flabel corelocali s 305 289 339 323 0 FreeSans 250 0 0 0 Y
port 7 nsew
flabel corelocali s 305 357 339 391 0 FreeSans 250 0 0 0 Y
port 7 nsew
flabel corelocali s 132 221 166 255 0 FreeSans 250 0 0 0 A_N
port 1 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew
rlabel comment s 0 0 0 0 4 nand2b_2
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2228600
string GDS_START 2222406
<< end >>
