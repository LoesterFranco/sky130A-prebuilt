magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 109 70 173 493
rect 445 215 568 265
rect 1427 289 1553 323
rect 1427 199 1471 289
rect 1611 215 1739 265
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 17 298 75 527
rect 17 17 75 147
rect 209 443 286 527
rect 322 447 636 481
rect 787 447 853 527
rect 940 455 1599 489
rect 1691 455 1758 527
rect 322 409 366 447
rect 940 413 974 455
rect 209 375 366 409
rect 434 379 974 413
rect 209 173 253 375
rect 299 307 636 341
rect 209 139 343 173
rect 207 17 265 105
rect 299 85 343 139
rect 377 119 411 307
rect 602 265 636 307
rect 680 305 757 339
rect 701 275 757 305
rect 602 199 667 265
rect 471 159 547 181
rect 701 159 735 275
rect 791 241 825 379
rect 871 289 975 343
rect 471 125 735 159
rect 769 207 825 241
rect 769 91 803 207
rect 536 85 633 91
rect 299 51 633 85
rect 677 57 803 91
rect 837 17 871 173
rect 917 83 975 289
rect 1011 119 1045 421
rect 1079 178 1113 455
rect 1838 421 1897 493
rect 1159 323 1242 409
rect 1359 387 1897 421
rect 1159 289 1325 323
rect 1162 199 1247 254
rect 1079 165 1131 178
rect 1079 144 1171 165
rect 1087 131 1171 144
rect 1011 97 1053 119
rect 1011 53 1093 97
rect 1137 64 1171 131
rect 1205 126 1247 199
rect 1291 85 1325 289
rect 1359 119 1393 387
rect 1790 375 1897 387
rect 1597 299 1807 341
rect 1773 265 1807 299
rect 1505 189 1567 255
rect 1773 199 1829 265
rect 1505 146 1546 189
rect 1773 181 1807 199
rect 1613 150 1807 181
rect 1605 147 1807 150
rect 1427 85 1530 93
rect 1291 51 1530 85
rect 1605 59 1663 147
rect 1863 117 1897 375
rect 1707 17 1741 113
rect 1837 51 1897 117
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< obsm1 >>
rect 711 320 769 329
rect 1201 320 1259 329
rect 711 292 1259 320
rect 711 283 769 292
rect 1201 283 1259 292
rect 905 184 963 193
rect 1201 184 1259 193
rect 1497 184 1555 193
rect 905 156 1555 184
rect 905 147 963 156
rect 1201 147 1259 156
rect 1497 147 1555 156
rect 1007 116 1065 125
rect 1599 116 1657 125
rect 1007 88 1657 116
rect 1007 79 1065 88
rect 1599 79 1657 88
<< labels >>
rlabel locali s 1611 215 1739 265 6 A
port 1 nsew signal input
rlabel locali s 1427 289 1553 323 6 B
port 2 nsew signal input
rlabel locali s 1427 199 1471 289 6 B
port 2 nsew signal input
rlabel locali s 445 215 568 265 6 C
port 3 nsew signal input
rlabel locali s 109 70 173 493 6 X
port 4 nsew signal output
rlabel metal1 s 0 -48 1932 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 1932 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1932 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 735940
string GDS_START 723148
<< end >>
