magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 1510 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 89 47 119 131
rect 183 47 213 131
rect 381 47 411 131
rect 475 47 505 131
rect 593 47 623 119
rect 679 47 709 119
rect 774 47 804 131
rect 982 47 1012 177
rect 1079 47 1109 177
rect 1173 47 1203 177
rect 1267 47 1297 177
rect 1361 47 1391 177
<< pmoshvt >>
rect 81 363 117 491
rect 175 363 211 491
rect 373 369 409 497
rect 467 369 503 497
rect 573 413 609 497
rect 667 413 703 497
rect 776 413 812 497
rect 974 297 1010 497
rect 1071 297 1107 497
rect 1165 297 1201 497
rect 1259 297 1295 497
rect 1353 297 1389 497
<< ndiff >>
rect 27 119 89 131
rect 27 85 35 119
rect 69 85 89 119
rect 27 47 89 85
rect 119 93 183 131
rect 119 59 129 93
rect 163 59 183 93
rect 119 47 183 59
rect 213 119 265 131
rect 213 85 223 119
rect 257 85 265 119
rect 213 47 265 85
rect 319 119 381 131
rect 319 85 327 119
rect 361 85 381 119
rect 319 47 381 85
rect 411 89 475 131
rect 411 55 421 89
rect 455 55 475 89
rect 411 47 475 55
rect 505 119 555 131
rect 920 133 982 177
rect 724 119 774 131
rect 505 47 593 119
rect 623 107 679 119
rect 623 73 634 107
rect 668 73 679 107
rect 623 47 679 73
rect 709 47 774 119
rect 804 106 866 131
rect 804 72 824 106
rect 858 72 866 106
rect 804 47 866 72
rect 920 99 934 133
rect 968 99 982 133
rect 920 47 982 99
rect 1012 127 1079 177
rect 1012 93 1025 127
rect 1059 93 1079 127
rect 1012 47 1079 93
rect 1109 133 1173 177
rect 1109 99 1119 133
rect 1153 99 1173 133
rect 1109 47 1173 99
rect 1203 127 1267 177
rect 1203 93 1213 127
rect 1247 93 1267 127
rect 1203 47 1267 93
rect 1297 127 1361 177
rect 1297 93 1307 127
rect 1341 93 1361 127
rect 1297 47 1361 93
rect 1391 127 1443 177
rect 1391 93 1401 127
rect 1435 93 1443 127
rect 1391 47 1443 93
<< pdiff >>
rect 27 477 81 491
rect 27 443 35 477
rect 69 443 81 477
rect 27 409 81 443
rect 27 375 35 409
rect 69 375 81 409
rect 27 363 81 375
rect 117 461 175 491
rect 117 427 129 461
rect 163 427 175 461
rect 117 363 175 427
rect 211 477 265 491
rect 211 443 223 477
rect 257 443 265 477
rect 211 409 265 443
rect 211 375 223 409
rect 257 375 265 409
rect 211 363 265 375
rect 319 483 373 497
rect 319 449 327 483
rect 361 449 373 483
rect 319 415 373 449
rect 319 381 327 415
rect 361 381 373 415
rect 319 369 373 381
rect 409 485 467 497
rect 409 451 421 485
rect 455 451 467 485
rect 409 417 467 451
rect 409 383 421 417
rect 455 383 467 417
rect 409 369 467 383
rect 503 413 573 497
rect 609 485 667 497
rect 609 451 621 485
rect 655 451 667 485
rect 609 413 667 451
rect 703 413 776 497
rect 812 477 866 497
rect 812 443 824 477
rect 858 443 866 477
rect 812 413 866 443
rect 920 471 974 497
rect 920 437 928 471
rect 962 437 974 471
rect 503 369 555 413
rect 920 368 974 437
rect 920 334 928 368
rect 962 334 974 368
rect 920 297 974 334
rect 1010 484 1071 497
rect 1010 450 1025 484
rect 1059 450 1071 484
rect 1010 364 1071 450
rect 1010 330 1025 364
rect 1059 330 1071 364
rect 1010 297 1071 330
rect 1107 475 1165 497
rect 1107 441 1119 475
rect 1153 441 1165 475
rect 1107 384 1165 441
rect 1107 350 1119 384
rect 1153 350 1165 384
rect 1107 297 1165 350
rect 1201 475 1259 497
rect 1201 441 1213 475
rect 1247 441 1259 475
rect 1201 384 1259 441
rect 1201 350 1213 384
rect 1247 350 1259 384
rect 1201 297 1259 350
rect 1295 475 1353 497
rect 1295 441 1307 475
rect 1341 441 1353 475
rect 1295 384 1353 441
rect 1295 350 1307 384
rect 1341 350 1353 384
rect 1295 297 1353 350
rect 1389 475 1443 497
rect 1389 441 1401 475
rect 1435 441 1443 475
rect 1389 384 1443 441
rect 1389 350 1401 384
rect 1435 350 1443 384
rect 1389 297 1443 350
<< ndiffc >>
rect 35 85 69 119
rect 129 59 163 93
rect 223 85 257 119
rect 327 85 361 119
rect 421 55 455 89
rect 634 73 668 107
rect 824 72 858 106
rect 934 99 968 133
rect 1025 93 1059 127
rect 1119 99 1153 133
rect 1213 93 1247 127
rect 1307 93 1341 127
rect 1401 93 1435 127
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 129 427 163 461
rect 223 443 257 477
rect 223 375 257 409
rect 327 449 361 483
rect 327 381 361 415
rect 421 451 455 485
rect 421 383 455 417
rect 621 451 655 485
rect 824 443 858 477
rect 928 437 962 471
rect 928 334 962 368
rect 1025 450 1059 484
rect 1025 330 1059 364
rect 1119 441 1153 475
rect 1119 350 1153 384
rect 1213 441 1247 475
rect 1213 350 1247 384
rect 1307 441 1341 475
rect 1307 350 1341 384
rect 1401 441 1435 475
rect 1401 350 1435 384
<< poly >>
rect 81 491 117 517
rect 175 491 211 517
rect 373 497 409 523
rect 467 497 503 523
rect 573 497 609 523
rect 667 497 703 523
rect 776 497 812 523
rect 974 497 1010 523
rect 1071 497 1107 523
rect 1165 497 1201 523
rect 1259 497 1295 523
rect 1353 497 1389 523
rect 573 398 609 413
rect 667 398 703 413
rect 776 398 812 413
rect 81 348 117 363
rect 175 348 211 363
rect 373 354 409 369
rect 467 354 503 369
rect 46 318 119 348
rect 46 280 76 318
rect 21 264 76 280
rect 173 274 213 348
rect 21 230 32 264
rect 66 230 76 264
rect 21 214 76 230
rect 128 264 213 274
rect 128 230 144 264
rect 178 230 213 264
rect 371 241 411 354
rect 128 220 213 230
rect 46 176 76 214
rect 46 146 119 176
rect 89 131 119 146
rect 183 131 213 220
rect 318 225 411 241
rect 318 191 328 225
rect 362 191 411 225
rect 465 219 505 354
rect 571 337 611 398
rect 665 375 705 398
rect 547 321 611 337
rect 663 365 729 375
rect 663 331 679 365
rect 713 331 729 365
rect 663 321 729 331
rect 774 373 814 398
rect 774 357 872 373
rect 774 323 828 357
rect 862 323 872 357
rect 547 287 557 321
rect 591 287 611 321
rect 547 279 611 287
rect 774 307 872 323
rect 547 271 709 279
rect 571 249 709 271
rect 318 175 411 191
rect 381 131 411 175
rect 454 203 518 219
rect 454 169 464 203
rect 498 169 518 203
rect 454 153 518 169
rect 573 191 637 207
rect 573 157 583 191
rect 617 157 637 191
rect 475 131 505 153
rect 573 141 637 157
rect 593 119 623 141
rect 679 119 709 249
rect 774 131 804 307
rect 974 282 1010 297
rect 1071 282 1107 297
rect 1165 282 1201 297
rect 1259 282 1295 297
rect 1353 282 1389 297
rect 972 265 1012 282
rect 1069 265 1109 282
rect 1163 265 1203 282
rect 1257 265 1297 282
rect 1351 265 1391 282
rect 856 249 1012 265
rect 856 215 866 249
rect 900 215 1012 249
rect 856 199 1012 215
rect 1054 249 1391 265
rect 1054 215 1064 249
rect 1098 215 1391 249
rect 1054 199 1391 215
rect 982 177 1012 199
rect 1079 177 1109 199
rect 1173 177 1203 199
rect 1267 177 1297 199
rect 1361 177 1391 199
rect 89 21 119 47
rect 183 21 213 47
rect 381 21 411 47
rect 475 21 505 47
rect 593 21 623 47
rect 679 21 709 47
rect 774 21 804 47
rect 982 21 1012 47
rect 1079 21 1109 47
rect 1173 21 1203 47
rect 1267 21 1297 47
rect 1361 21 1391 47
<< polycont >>
rect 32 230 66 264
rect 144 230 178 264
rect 328 191 362 225
rect 679 331 713 365
rect 828 323 862 357
rect 557 287 591 321
rect 464 169 498 203
rect 583 157 617 191
rect 866 215 900 249
rect 1064 215 1098 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 35 477 69 493
rect 35 409 69 443
rect 103 461 179 527
rect 103 427 129 461
rect 163 427 179 461
rect 223 477 257 493
rect 421 485 484 527
rect 223 409 257 443
rect 69 375 178 393
rect 35 359 178 375
rect 17 264 66 325
rect 17 230 32 264
rect 17 197 66 230
rect 132 314 178 359
rect 166 280 178 314
rect 132 264 178 280
rect 132 230 144 264
rect 132 161 178 230
rect 35 127 178 161
rect 35 119 69 127
rect 223 119 257 354
rect 311 449 327 483
rect 361 449 377 483
rect 311 415 377 449
rect 311 381 327 415
rect 361 381 377 415
rect 311 333 377 381
rect 455 451 484 485
rect 605 451 621 485
rect 655 451 790 485
rect 421 417 484 451
rect 455 383 484 417
rect 421 367 484 383
rect 534 388 591 401
rect 568 354 591 388
rect 311 299 458 333
rect 295 225 378 265
rect 295 191 328 225
rect 362 191 378 225
rect 424 219 458 299
rect 534 321 591 354
rect 534 287 557 321
rect 534 271 591 287
rect 635 365 713 399
rect 635 331 679 365
rect 635 314 713 331
rect 669 283 713 314
rect 424 203 508 219
rect 635 207 669 280
rect 424 169 464 203
rect 498 169 508 203
rect 424 157 508 169
rect 35 69 69 85
rect 103 59 129 93
rect 163 59 179 93
rect 223 69 257 85
rect 327 153 508 157
rect 583 191 669 207
rect 617 157 669 191
rect 327 123 458 153
rect 583 141 669 157
rect 756 265 790 451
rect 824 477 858 527
rect 824 427 858 443
rect 928 471 972 487
rect 962 437 972 471
rect 928 373 972 437
rect 828 368 972 373
rect 828 357 928 368
rect 862 334 928 357
rect 962 334 972 368
rect 862 323 972 334
rect 828 307 972 323
rect 934 265 972 307
rect 1018 484 1075 527
rect 1018 450 1025 484
rect 1059 450 1075 484
rect 1018 364 1075 450
rect 1018 330 1025 364
rect 1059 330 1075 364
rect 1018 299 1075 330
rect 1119 475 1179 491
rect 1153 441 1179 475
rect 1119 384 1179 441
rect 1153 350 1179 384
rect 1119 299 1179 350
rect 1213 475 1263 527
rect 1247 441 1263 475
rect 1213 384 1263 441
rect 1247 350 1263 384
rect 1213 299 1263 350
rect 1307 475 1361 491
rect 1341 441 1361 475
rect 1307 384 1361 441
rect 1341 350 1361 384
rect 1142 265 1179 299
rect 1307 265 1361 350
rect 1401 475 1435 527
rect 1401 384 1435 441
rect 1401 299 1435 350
rect 756 249 900 265
rect 756 215 866 249
rect 756 199 900 215
rect 934 249 1098 265
rect 934 215 1064 249
rect 934 199 1098 215
rect 1142 199 1447 265
rect 327 119 361 123
rect 756 107 790 199
rect 934 133 972 199
rect 1142 149 1179 199
rect 327 69 361 85
rect 103 17 179 59
rect 395 55 421 89
rect 455 55 471 89
rect 618 73 634 107
rect 668 73 790 107
rect 824 106 858 122
rect 395 17 471 55
rect 968 99 972 133
rect 934 83 972 99
rect 1018 127 1075 143
rect 1018 93 1025 127
rect 1059 93 1075 127
rect 824 17 858 72
rect 1018 17 1075 93
rect 1119 133 1179 149
rect 1153 99 1179 133
rect 1119 83 1179 99
rect 1213 127 1263 165
rect 1247 93 1263 127
rect 1213 17 1263 93
rect 1307 127 1361 199
rect 1341 93 1361 127
rect 1307 77 1361 93
rect 1401 127 1435 143
rect 1401 17 1435 93
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 132 280 166 314
rect 223 375 257 388
rect 223 354 257 375
rect 534 354 568 388
rect 635 280 669 314
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 211 388 269 394
rect 522 388 580 394
rect 211 354 223 388
rect 257 360 534 388
rect 257 354 269 360
rect 211 348 269 354
rect 522 354 534 360
rect 568 354 580 388
rect 522 348 580 354
rect 120 314 682 320
rect 120 280 132 314
rect 166 292 635 314
rect 166 280 178 292
rect 120 274 178 280
rect 623 280 635 292
rect 669 280 682 314
rect 623 274 682 280
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< labels >>
flabel corelocali s 305 221 339 255 0 FreeSans 200 0 0 0 D
port 1 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 200 0 0 0 GATE_N
port 2 nsew
flabel corelocali s 1129 357 1163 391 0 FreeSans 200 0 0 0 Q
port 7 nsew
flabel corelocali s 30 289 64 323 0 FreeSans 200 0 0 0 GATE_N
port 2 nsew
flabel corelocali s 1129 425 1163 459 0 FreeSans 200 0 0 0 Q
port 7 nsew
flabel corelocali s 1129 85 1163 119 0 FreeSans 200 0 0 0 Q
port 7 nsew
flabel corelocali s 1407 221 1441 255 0 FreeSans 200 0 0 0 Q
port 7 nsew
flabel corelocali s 1229 221 1263 255 0 FreeSans 200 0 0 0 Q
port 7 nsew
flabel corelocali s 1320 221 1354 255 0 FreeSans 200 0 0 0 Q
port 7 nsew
flabel corelocali s 1319 357 1353 391 0 FreeSans 200 0 0 0 Q
port 7 nsew
flabel corelocali s 1319 425 1353 459 0 FreeSans 200 0 0 0 Q
port 7 nsew
flabel corelocali s 1319 153 1353 187 0 FreeSans 200 0 0 0 Q
port 7 nsew
flabel corelocali s 1319 85 1353 119 0 FreeSans 200 0 0 0 Q
port 7 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew
rlabel comment s 0 0 0 0 4 dlxtn_4
<< properties >>
string FIXED_BBOX 0 0 1472 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1960880
string GDS_START 1948756
<< end >>
