magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 2117 333 2183 493
rect 2305 333 2371 493
rect 2493 333 2559 493
rect 2681 333 2747 493
rect 2869 333 2935 493
rect 3057 333 3123 493
rect 3245 333 3311 493
rect 3433 333 3499 493
rect 2117 299 3499 333
rect 113 215 383 265
rect 585 215 855 265
rect 1621 215 1891 265
rect 3417 181 3499 299
rect 2117 145 3499 181
rect 2117 51 2183 145
rect 2305 51 2371 145
rect 2493 51 2559 145
rect 2681 51 2747 145
rect 2869 51 2935 145
rect 3057 51 3123 145
rect 3245 51 3311 145
rect 3433 51 3499 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3157 561
rect 3191 527 3249 561
rect 3283 527 3341 561
rect 3375 527 3433 561
rect 3467 527 3525 561
rect 3559 527 3617 561
rect 3651 527 3680 561
rect 19 459 461 493
rect 19 85 79 459
rect 113 333 179 425
rect 213 367 267 459
rect 301 333 367 425
rect 113 299 367 333
rect 401 299 461 459
rect 505 299 559 527
rect 593 333 659 493
rect 693 367 747 527
rect 781 333 847 493
rect 593 299 847 333
rect 881 299 935 527
rect 969 265 1035 493
rect 1069 299 1123 527
rect 1157 333 1223 493
rect 1257 367 1311 527
rect 1345 333 1411 493
rect 1157 299 1411 333
rect 1445 299 1499 527
rect 1543 459 1985 493
rect 1543 299 1603 459
rect 1637 333 1703 425
rect 1737 367 1791 459
rect 1825 333 1891 425
rect 1637 299 1891 333
rect 1925 265 1985 459
rect 2029 299 2083 527
rect 2217 367 2271 527
rect 2405 367 2459 527
rect 2593 367 2647 527
rect 2781 367 2835 527
rect 2969 367 3023 527
rect 3157 367 3211 527
rect 3345 367 3399 527
rect 3533 299 3587 527
rect 969 215 1419 265
rect 1925 215 3373 265
rect 113 145 847 181
rect 113 119 179 145
rect 301 119 367 145
rect 213 85 267 109
rect 401 85 461 110
rect 19 51 461 85
rect 505 17 559 110
rect 593 51 659 145
rect 693 17 747 109
rect 781 51 847 145
rect 881 17 935 181
rect 969 51 1035 215
rect 1069 17 1123 181
rect 1157 145 1891 181
rect 1157 51 1223 145
rect 1257 17 1311 109
rect 1345 51 1411 145
rect 1637 119 1703 145
rect 1825 119 1891 145
rect 1445 17 1499 110
rect 1543 85 1603 110
rect 1737 85 1791 109
rect 1925 85 1985 215
rect 1543 51 1985 85
rect 2029 17 2083 181
rect 2217 17 2271 109
rect 2405 17 2459 109
rect 2593 17 2647 109
rect 2781 17 2835 110
rect 2969 17 3023 109
rect 3157 17 3211 109
rect 3345 17 3399 109
rect 3533 17 3587 181
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3341 17
rect 3375 -17 3433 17
rect 3467 -17 3525 17
rect 3559 -17 3617 17
rect 3651 -17 3680 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 2881 527 2915 561
rect 2973 527 3007 561
rect 3065 527 3099 561
rect 3157 527 3191 561
rect 3249 527 3283 561
rect 3341 527 3375 561
rect 3433 527 3467 561
rect 3525 527 3559 561
rect 3617 527 3651 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
rect 2881 -17 2915 17
rect 2973 -17 3007 17
rect 3065 -17 3099 17
rect 3157 -17 3191 17
rect 3249 -17 3283 17
rect 3341 -17 3375 17
rect 3433 -17 3467 17
rect 3525 -17 3559 17
rect 3617 -17 3651 17
<< metal1 >>
rect 0 561 3680 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3157 561
rect 3191 527 3249 561
rect 3283 527 3341 561
rect 3375 527 3433 561
rect 3467 527 3525 561
rect 3559 527 3617 561
rect 3651 527 3680 561
rect 0 496 3680 527
rect 0 17 3680 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3341 17
rect 3375 -17 3433 17
rect 3467 -17 3525 17
rect 3559 -17 3617 17
rect 3651 -17 3680 17
rect 0 -48 3680 -17
<< obsm1 >>
rect 597 456 655 465
rect 785 456 843 465
rect 597 428 1532 456
rect 597 419 655 428
rect 785 419 843 428
rect 117 388 175 397
rect 305 388 363 397
rect 1161 388 1219 397
rect 1349 388 1407 397
rect 117 360 1407 388
rect 1504 388 1532 428
rect 1641 388 1699 397
rect 1829 388 1887 397
rect 1504 360 1887 388
rect 117 351 175 360
rect 305 351 363 360
rect 1161 351 1219 360
rect 1349 351 1407 360
rect 1641 351 1699 360
rect 1829 351 1887 360
rect 23 116 81 125
rect 1923 116 1981 125
rect 23 88 1981 116
rect 23 79 81 88
rect 1923 79 1981 88
<< labels >>
rlabel locali s 1621 215 1891 265 6 A0
port 1 nsew signal input
rlabel locali s 113 215 383 265 6 A1
port 2 nsew signal input
rlabel locali s 585 215 855 265 6 S
port 3 nsew signal input
rlabel locali s 3433 333 3499 493 6 X
port 4 nsew signal output
rlabel locali s 3433 51 3499 145 6 X
port 4 nsew signal output
rlabel locali s 3417 181 3499 299 6 X
port 4 nsew signal output
rlabel locali s 3245 333 3311 493 6 X
port 4 nsew signal output
rlabel locali s 3245 51 3311 145 6 X
port 4 nsew signal output
rlabel locali s 3057 333 3123 493 6 X
port 4 nsew signal output
rlabel locali s 3057 51 3123 145 6 X
port 4 nsew signal output
rlabel locali s 2869 333 2935 493 6 X
port 4 nsew signal output
rlabel locali s 2869 51 2935 145 6 X
port 4 nsew signal output
rlabel locali s 2681 333 2747 493 6 X
port 4 nsew signal output
rlabel locali s 2681 51 2747 145 6 X
port 4 nsew signal output
rlabel locali s 2493 333 2559 493 6 X
port 4 nsew signal output
rlabel locali s 2493 51 2559 145 6 X
port 4 nsew signal output
rlabel locali s 2305 333 2371 493 6 X
port 4 nsew signal output
rlabel locali s 2305 51 2371 145 6 X
port 4 nsew signal output
rlabel locali s 2117 333 2183 493 6 X
port 4 nsew signal output
rlabel locali s 2117 299 3499 333 6 X
port 4 nsew signal output
rlabel locali s 2117 145 3499 181 6 X
port 4 nsew signal output
rlabel locali s 2117 51 2183 145 6 X
port 4 nsew signal output
rlabel metal1 s 0 -48 3680 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 3680 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 3680 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3430384
string GDS_START 3403082
<< end >>
