magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 617 415 655 493
rect 617 381 807 415
rect 17 199 72 265
rect 186 199 262 265
rect 301 199 389 265
rect 433 199 535 265
rect 753 157 807 381
rect 589 123 807 157
rect 589 51 665 123
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 18 353 71 493
rect 105 387 181 527
rect 225 353 364 493
rect 475 387 571 527
rect 689 451 765 527
rect 18 347 364 353
rect 18 302 605 347
rect 106 165 152 302
rect 571 265 605 302
rect 571 199 713 265
rect 19 85 152 165
rect 186 127 475 165
rect 19 51 86 85
rect 307 17 374 93
rect 508 17 555 105
rect 709 17 775 89
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
rlabel locali s 433 199 535 265 6 A1
port 1 nsew signal input
rlabel locali s 301 199 389 265 6 A2
port 2 nsew signal input
rlabel locali s 186 199 262 265 6 B1
port 3 nsew signal input
rlabel locali s 17 199 72 265 6 C1
port 4 nsew signal input
rlabel locali s 753 157 807 381 6 X
port 5 nsew signal output
rlabel locali s 617 415 655 493 6 X
port 5 nsew signal output
rlabel locali s 617 381 807 415 6 X
port 5 nsew signal output
rlabel locali s 589 123 807 157 6 X
port 5 nsew signal output
rlabel locali s 589 51 665 123 6 X
port 5 nsew signal output
rlabel metal1 s 0 -48 828 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 828 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2574944
string GDS_START 2568348
<< end >>
