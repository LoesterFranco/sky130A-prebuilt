magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 93 47 123 177
rect 323 47 353 177
rect 417 47 447 177
rect 529 47 559 177
rect 613 47 643 177
<< pmoshvt >>
rect 85 297 121 497
rect 315 297 351 497
rect 403 297 439 497
rect 533 297 569 497
rect 615 297 651 497
<< ndiff >>
rect 27 136 93 177
rect 27 102 35 136
rect 69 102 93 136
rect 27 47 93 102
rect 123 95 175 177
rect 123 61 133 95
rect 167 61 175 95
rect 123 47 175 61
rect 261 163 323 177
rect 261 129 269 163
rect 303 129 323 163
rect 261 47 323 129
rect 353 95 417 177
rect 353 61 363 95
rect 397 61 417 95
rect 353 47 417 61
rect 447 149 529 177
rect 447 115 457 149
rect 491 115 529 149
rect 447 47 529 115
rect 559 89 613 177
rect 559 55 569 89
rect 603 55 613 89
rect 559 47 613 55
rect 643 163 705 177
rect 643 129 663 163
rect 697 129 705 163
rect 643 95 705 129
rect 643 61 663 95
rect 697 61 705 95
rect 643 47 705 61
<< pdiff >>
rect 27 477 85 497
rect 27 443 39 477
rect 73 443 85 477
rect 27 409 85 443
rect 27 375 39 409
rect 73 375 85 409
rect 27 341 85 375
rect 27 307 39 341
rect 73 307 85 341
rect 27 297 85 307
rect 121 477 315 497
rect 121 443 136 477
rect 170 443 266 477
rect 300 443 315 477
rect 121 409 315 443
rect 121 375 136 409
rect 170 375 266 409
rect 300 375 315 409
rect 121 297 315 375
rect 351 297 403 497
rect 439 485 533 497
rect 439 451 451 485
rect 485 451 533 485
rect 439 417 533 451
rect 439 383 451 417
rect 485 383 533 417
rect 439 349 533 383
rect 439 315 451 349
rect 485 315 533 349
rect 439 297 533 315
rect 569 297 615 497
rect 651 485 705 497
rect 651 451 663 485
rect 697 451 705 485
rect 651 417 705 451
rect 651 383 663 417
rect 697 383 705 417
rect 651 349 705 383
rect 651 315 663 349
rect 697 315 705 349
rect 651 297 705 315
<< ndiffc >>
rect 35 102 69 136
rect 133 61 167 95
rect 269 129 303 163
rect 363 61 397 95
rect 457 115 491 149
rect 569 55 603 89
rect 663 129 697 163
rect 663 61 697 95
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 136 443 170 477
rect 266 443 300 477
rect 136 375 170 409
rect 266 375 300 409
rect 451 451 485 485
rect 451 383 485 417
rect 451 315 485 349
rect 663 451 697 485
rect 663 383 697 417
rect 663 315 697 349
<< poly >>
rect 85 497 121 523
rect 315 497 351 523
rect 403 497 439 523
rect 533 497 569 523
rect 615 497 651 523
rect 85 282 121 297
rect 315 282 351 297
rect 403 282 439 297
rect 533 282 569 297
rect 615 282 651 297
rect 83 265 123 282
rect 313 265 353 282
rect 49 249 123 265
rect 49 215 59 249
rect 93 215 123 249
rect 49 199 123 215
rect 275 249 353 265
rect 275 215 285 249
rect 319 215 353 249
rect 275 199 353 215
rect 401 265 441 282
rect 531 265 571 282
rect 401 249 465 265
rect 401 215 411 249
rect 445 215 465 249
rect 401 199 465 215
rect 507 249 571 265
rect 507 215 517 249
rect 551 215 571 249
rect 507 199 571 215
rect 613 265 653 282
rect 613 249 708 265
rect 613 215 658 249
rect 692 215 708 249
rect 613 199 708 215
rect 93 177 123 199
rect 323 177 353 199
rect 417 177 447 199
rect 529 177 559 199
rect 613 177 643 199
rect 93 21 123 47
rect 323 21 353 47
rect 417 21 447 47
rect 529 21 559 47
rect 613 21 643 47
<< polycont >>
rect 59 215 93 249
rect 285 215 319 249
rect 411 215 445 249
rect 517 215 551 249
rect 658 215 692 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 17 477 73 493
rect 17 443 39 477
rect 17 409 73 443
rect 17 375 39 409
rect 120 477 316 527
rect 120 443 136 477
rect 170 443 266 477
rect 300 443 316 477
rect 120 409 316 443
rect 120 375 136 409
rect 170 375 266 409
rect 300 375 316 409
rect 380 485 501 493
rect 380 451 451 485
rect 485 451 501 485
rect 663 485 715 527
rect 380 436 501 451
rect 380 417 493 436
rect 380 383 451 417
rect 485 383 493 417
rect 17 341 73 375
rect 380 349 493 383
rect 380 341 451 349
rect 17 307 39 341
rect 73 315 451 341
rect 485 315 493 349
rect 571 323 625 481
rect 73 307 493 315
rect 17 299 493 307
rect 17 249 93 265
rect 17 215 59 249
rect 17 199 93 215
rect 135 165 169 299
rect 527 289 625 323
rect 697 451 715 485
rect 663 417 715 451
rect 697 383 715 417
rect 663 349 715 383
rect 697 315 715 349
rect 663 291 715 315
rect 203 249 319 265
rect 203 215 285 249
rect 203 199 319 215
rect 363 249 465 265
rect 527 249 579 289
rect 363 215 411 249
rect 445 215 465 249
rect 501 215 517 249
rect 551 215 579 249
rect 613 249 715 255
rect 613 215 658 249
rect 692 215 715 249
rect 363 199 465 215
rect 489 165 715 173
rect 17 136 169 165
rect 17 102 35 136
rect 69 129 169 136
rect 250 163 715 165
rect 250 129 269 163
rect 303 149 663 163
rect 303 129 457 149
rect 17 73 69 102
rect 491 139 663 149
rect 491 115 512 139
rect 103 61 133 95
rect 167 61 363 95
rect 397 61 413 95
rect 457 56 512 115
rect 637 129 663 139
rect 697 129 715 163
rect 569 89 603 105
rect 637 95 715 129
rect 637 61 663 95
rect 697 61 715 95
rect 637 56 715 61
rect 569 17 603 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel corelocali s 582 357 616 391 0 FreeSans 400 0 0 0 A2
port 2 nsew
flabel corelocali s 400 425 434 459 0 FreeSans 400 0 0 0 Y
port 10 nsew
flabel corelocali s 214 221 248 255 0 FreeSans 400 0 0 0 B1
port 3 nsew
flabel corelocali s 29 221 63 255 0 FreeSans 400 0 0 0 C1
port 5 nsew
flabel corelocali s 669 221 703 255 0 FreeSans 400 0 0 0 A1
port 1 nsew
flabel corelocali s 400 357 434 391 0 FreeSans 400 0 0 0 Y
port 10 nsew
flabel corelocali s 396 238 396 238 0 FreeSans 400 0 0 0 B2
port 4 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew
rlabel comment s 0 0 0 0 4 o221ai_1
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 835850
string GDS_START 829290
<< end >>
