magic
tech sky130A
magscale 1 2
timestamp 1599588209
<< nwell >>
rect -38 332 902 704
<< pwell >>
rect 0 0 864 49
<< scpmos >>
rect 86 368 116 592
rect 176 368 206 592
rect 266 368 296 592
rect 360 368 390 592
rect 467 409 497 577
rect 562 409 592 577
rect 657 409 687 577
rect 747 409 777 577
<< nmoslvt >>
rect 84 99 114 247
rect 170 99 200 247
rect 256 99 286 247
rect 372 99 402 247
rect 474 119 504 247
rect 565 119 595 247
rect 660 119 690 247
rect 750 119 780 247
<< ndiff >>
rect 27 235 84 247
rect 27 201 39 235
rect 73 201 84 235
rect 27 145 84 201
rect 27 111 39 145
rect 73 111 84 145
rect 27 99 84 111
rect 114 235 170 247
rect 114 201 125 235
rect 159 201 170 235
rect 114 145 170 201
rect 114 111 125 145
rect 159 111 170 145
rect 114 99 170 111
rect 200 151 256 247
rect 200 117 211 151
rect 245 117 256 151
rect 200 99 256 117
rect 286 219 372 247
rect 286 185 311 219
rect 345 185 372 219
rect 286 145 372 185
rect 286 111 311 145
rect 345 111 372 145
rect 286 99 372 111
rect 402 235 474 247
rect 402 201 413 235
rect 447 201 474 235
rect 402 157 474 201
rect 402 123 413 157
rect 447 123 474 157
rect 402 119 474 123
rect 504 229 565 247
rect 504 195 515 229
rect 549 195 565 229
rect 504 161 565 195
rect 504 127 515 161
rect 549 127 565 161
rect 504 119 565 127
rect 595 239 660 247
rect 595 205 615 239
rect 649 205 660 239
rect 595 161 660 205
rect 595 127 615 161
rect 649 127 660 161
rect 595 119 660 127
rect 690 168 750 247
rect 690 134 701 168
rect 735 134 750 168
rect 690 119 750 134
rect 780 235 837 247
rect 780 201 791 235
rect 825 201 837 235
rect 780 165 837 201
rect 780 131 791 165
rect 825 131 837 165
rect 780 119 837 131
rect 402 99 459 119
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 497 86 546
rect 27 463 39 497
rect 73 463 86 497
rect 27 414 86 463
rect 27 380 39 414
rect 73 380 86 414
rect 27 368 86 380
rect 116 580 176 592
rect 116 546 129 580
rect 163 546 176 580
rect 116 499 176 546
rect 116 465 129 499
rect 163 465 176 499
rect 116 419 176 465
rect 116 385 129 419
rect 163 385 176 419
rect 116 368 176 385
rect 206 580 266 592
rect 206 546 219 580
rect 253 546 266 580
rect 206 487 266 546
rect 206 453 219 487
rect 253 453 266 487
rect 206 368 266 453
rect 296 580 360 592
rect 296 546 309 580
rect 343 546 360 580
rect 296 499 360 546
rect 296 465 309 499
rect 343 465 360 499
rect 296 419 360 465
rect 296 385 309 419
rect 343 385 360 419
rect 296 368 360 385
rect 390 580 449 592
rect 390 546 403 580
rect 437 577 449 580
rect 437 546 467 577
rect 390 508 467 546
rect 390 474 403 508
rect 437 474 467 508
rect 390 409 467 474
rect 497 565 562 577
rect 497 531 510 565
rect 544 531 562 565
rect 497 455 562 531
rect 497 421 510 455
rect 544 421 562 455
rect 497 409 562 421
rect 592 568 657 577
rect 592 534 610 568
rect 644 534 657 568
rect 592 500 657 534
rect 592 466 610 500
rect 644 466 657 500
rect 592 409 657 466
rect 687 565 747 577
rect 687 531 700 565
rect 734 531 747 565
rect 687 455 747 531
rect 687 421 700 455
rect 734 421 747 455
rect 687 409 747 421
rect 777 565 836 577
rect 777 531 790 565
rect 824 531 836 565
rect 777 455 836 531
rect 777 421 790 455
rect 824 421 836 455
rect 777 409 836 421
rect 390 368 443 409
<< ndiffc >>
rect 39 201 73 235
rect 39 111 73 145
rect 125 201 159 235
rect 125 111 159 145
rect 211 117 245 151
rect 311 185 345 219
rect 311 111 345 145
rect 413 201 447 235
rect 413 123 447 157
rect 515 195 549 229
rect 515 127 549 161
rect 615 205 649 239
rect 615 127 649 161
rect 701 134 735 168
rect 791 201 825 235
rect 791 131 825 165
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 129 546 163 580
rect 129 465 163 499
rect 129 385 163 419
rect 219 546 253 580
rect 219 453 253 487
rect 309 546 343 580
rect 309 465 343 499
rect 309 385 343 419
rect 403 546 437 580
rect 403 474 437 508
rect 510 531 544 565
rect 510 421 544 455
rect 610 534 644 568
rect 610 466 644 500
rect 700 531 734 565
rect 700 421 734 455
rect 790 531 824 565
rect 790 421 824 455
<< poly >>
rect 86 592 116 618
rect 176 592 206 618
rect 266 592 296 618
rect 360 592 390 618
rect 467 577 497 603
rect 562 577 592 603
rect 657 577 687 603
rect 747 577 777 603
rect 467 394 497 409
rect 562 394 592 409
rect 657 394 687 409
rect 747 394 777 409
rect 86 353 116 368
rect 176 353 206 368
rect 266 353 296 368
rect 360 353 390 368
rect 83 335 119 353
rect 173 335 209 353
rect 263 335 299 353
rect 357 335 393 353
rect 464 335 500 394
rect 559 383 595 394
rect 654 383 690 394
rect 559 340 690 383
rect 83 319 403 335
rect 83 285 217 319
rect 251 285 285 319
rect 319 285 353 319
rect 387 285 403 319
rect 83 269 403 285
rect 451 319 517 335
rect 451 285 467 319
rect 501 285 517 319
rect 559 306 601 340
rect 635 306 690 340
rect 559 290 690 306
rect 451 269 517 285
rect 84 247 114 269
rect 170 247 200 269
rect 256 247 286 269
rect 372 247 402 269
rect 474 247 504 269
rect 565 247 595 290
rect 660 247 690 290
rect 744 262 780 394
rect 750 247 780 262
rect 84 73 114 99
rect 170 73 200 99
rect 256 73 286 99
rect 372 73 402 99
rect 474 51 504 119
rect 565 93 595 119
rect 660 93 690 119
rect 750 51 780 119
rect 474 21 780 51
<< polycont >>
rect 217 285 251 319
rect 285 285 319 319
rect 353 285 387 319
rect 467 285 501 319
rect 601 306 635 340
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 23 580 73 649
rect 23 546 39 580
rect 23 497 73 546
rect 23 463 39 497
rect 23 414 73 463
rect 23 380 39 414
rect 23 364 73 380
rect 109 580 163 596
rect 109 546 129 580
rect 109 499 163 546
rect 109 465 129 499
rect 109 419 163 465
rect 203 580 253 649
rect 203 546 219 580
rect 203 487 253 546
rect 203 453 219 487
rect 203 437 253 453
rect 293 580 343 596
rect 293 546 309 580
rect 293 499 343 546
rect 293 465 309 499
rect 109 385 129 419
rect 293 419 343 465
rect 387 580 453 649
rect 387 546 403 580
rect 437 546 453 580
rect 387 508 453 546
rect 387 474 403 508
rect 437 474 453 508
rect 387 458 453 474
rect 494 565 560 581
rect 494 531 510 565
rect 544 531 560 565
rect 494 455 560 531
rect 594 568 660 649
rect 594 534 610 568
rect 644 534 660 568
rect 594 500 660 534
rect 594 466 610 500
rect 644 466 660 500
rect 594 458 660 466
rect 700 565 734 581
rect 494 424 510 455
rect 293 403 309 419
rect 163 385 309 403
rect 109 369 343 385
rect 377 421 510 424
rect 544 424 560 455
rect 700 455 734 531
rect 544 421 700 424
rect 377 390 734 421
rect 774 565 840 649
rect 774 531 790 565
rect 824 531 840 565
rect 774 455 840 531
rect 774 421 790 455
rect 824 421 840 455
rect 774 405 840 421
rect 109 310 167 369
rect 377 335 411 390
rect 201 319 411 335
rect 23 235 73 251
rect 23 201 39 235
rect 23 145 73 201
rect 23 111 39 145
rect 23 17 73 111
rect 109 235 159 310
rect 201 285 217 319
rect 251 285 285 319
rect 319 285 353 319
rect 387 285 411 319
rect 201 269 411 285
rect 451 319 551 356
rect 451 285 467 319
rect 501 285 551 319
rect 585 340 651 356
rect 585 306 601 340
rect 635 306 651 340
rect 585 290 651 306
rect 451 269 551 285
rect 700 256 734 390
rect 599 239 734 256
rect 109 201 125 235
rect 159 219 345 235
rect 159 201 311 219
rect 109 145 159 201
rect 295 185 311 201
rect 109 111 125 145
rect 109 95 159 111
rect 195 151 261 167
rect 195 117 211 151
rect 245 117 261 151
rect 195 17 261 117
rect 295 145 345 185
rect 295 111 311 145
rect 295 95 345 111
rect 397 201 413 235
rect 447 201 463 235
rect 397 157 463 201
rect 397 123 413 157
rect 447 123 463 157
rect 397 17 463 123
rect 499 229 565 235
rect 499 195 515 229
rect 549 195 565 229
rect 499 161 565 195
rect 499 127 515 161
rect 549 127 565 161
rect 499 85 565 127
rect 599 205 615 239
rect 649 222 734 239
rect 775 235 841 251
rect 649 205 665 222
rect 599 161 665 205
rect 775 201 791 235
rect 825 201 841 235
rect 599 127 615 161
rect 649 127 665 161
rect 599 119 665 127
rect 701 168 735 188
rect 701 85 735 134
rect 499 51 735 85
rect 775 165 841 201
rect 775 131 791 165
rect 825 131 841 165
rect 775 17 841 131
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel comment s 0 0 0 0 4 and2_4
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 X
port 7 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 B
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 864 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3204348
string GDS_START 3196774
<< end >>
