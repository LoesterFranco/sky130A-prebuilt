magic
tech sky130A
magscale 1 2
timestamp 1599588244
<< locali >>
rect 107 364 179 596
rect 107 226 141 364
rect 283 270 359 356
rect 397 270 463 356
rect 505 270 571 356
rect 619 270 743 356
rect 107 192 210 226
rect 144 70 210 192
rect 871 236 937 578
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 23 364 73 649
rect 213 458 320 649
rect 535 424 622 576
rect 763 458 829 649
rect 213 390 837 424
rect 23 158 73 228
rect 213 330 247 390
rect 175 264 247 330
rect 23 17 108 158
rect 244 17 310 226
rect 344 202 610 236
rect 803 209 837 390
rect 344 70 410 202
rect 444 17 510 168
rect 544 104 610 202
rect 644 143 837 209
rect 871 104 923 202
rect 544 70 923 104
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
rlabel locali s 283 270 359 356 6 A1
port 1 nsew signal input
rlabel locali s 397 270 463 356 6 A2
port 2 nsew signal input
rlabel locali s 505 270 571 356 6 A3
port 3 nsew signal input
rlabel locali s 871 236 937 578 6 B1
port 4 nsew signal input
rlabel locali s 619 270 743 356 6 B2
port 5 nsew signal input
rlabel locali s 144 70 210 192 6 X
port 6 nsew signal output
rlabel locali s 107 364 179 596 6 X
port 6 nsew signal output
rlabel locali s 107 226 141 364 6 X
port 6 nsew signal output
rlabel locali s 107 192 210 226 6 X
port 6 nsew signal output
rlabel metal1 s 0 -49 960 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 8 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 9 nsew power bidirectional
rlabel metal1 s 0 617 960 715 6 VPWR
port 10 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 665538
string GDS_START 657422
<< end >>
