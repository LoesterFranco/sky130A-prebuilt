magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 1694 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 102 47 132 177
rect 196 47 226 177
rect 290 47 320 177
rect 384 47 414 177
rect 478 47 508 177
rect 572 47 602 177
rect 666 47 696 177
rect 760 47 790 177
rect 854 47 884 177
rect 948 47 978 177
rect 1042 47 1072 177
rect 1136 47 1166 177
rect 1230 47 1260 177
rect 1324 47 1354 177
rect 1418 47 1448 177
rect 1512 47 1542 177
<< pmoshvt >>
rect 94 297 130 497
rect 188 297 224 497
rect 282 297 318 497
rect 376 297 412 497
rect 470 297 506 497
rect 564 297 600 497
rect 658 297 694 497
rect 752 297 788 497
rect 846 297 882 497
rect 940 297 976 497
rect 1034 297 1070 497
rect 1128 297 1164 497
rect 1222 297 1258 497
rect 1316 297 1352 497
rect 1410 297 1446 497
rect 1504 297 1540 497
<< ndiff >>
rect 40 161 102 177
rect 40 127 48 161
rect 82 127 102 161
rect 40 93 102 127
rect 40 59 48 93
rect 82 59 102 93
rect 40 47 102 59
rect 132 161 196 177
rect 132 127 142 161
rect 176 127 196 161
rect 132 93 196 127
rect 132 59 142 93
rect 176 59 196 93
rect 132 47 196 59
rect 226 93 290 177
rect 226 59 236 93
rect 270 59 290 93
rect 226 47 290 59
rect 320 161 384 177
rect 320 127 330 161
rect 364 127 384 161
rect 320 93 384 127
rect 320 59 330 93
rect 364 59 384 93
rect 320 47 384 59
rect 414 93 478 177
rect 414 59 424 93
rect 458 59 478 93
rect 414 47 478 59
rect 508 161 572 177
rect 508 127 518 161
rect 552 127 572 161
rect 508 93 572 127
rect 508 59 518 93
rect 552 59 572 93
rect 508 47 572 59
rect 602 93 666 177
rect 602 59 612 93
rect 646 59 666 93
rect 602 47 666 59
rect 696 161 760 177
rect 696 127 706 161
rect 740 127 760 161
rect 696 93 760 127
rect 696 59 706 93
rect 740 59 760 93
rect 696 47 760 59
rect 790 93 854 177
rect 790 59 800 93
rect 834 59 854 93
rect 790 47 854 59
rect 884 161 948 177
rect 884 127 894 161
rect 928 127 948 161
rect 884 93 948 127
rect 884 59 894 93
rect 928 59 948 93
rect 884 47 948 59
rect 978 93 1042 177
rect 978 59 988 93
rect 1022 59 1042 93
rect 978 47 1042 59
rect 1072 161 1136 177
rect 1072 127 1082 161
rect 1116 127 1136 161
rect 1072 93 1136 127
rect 1072 59 1082 93
rect 1116 59 1136 93
rect 1072 47 1136 59
rect 1166 93 1230 177
rect 1166 59 1176 93
rect 1210 59 1230 93
rect 1166 47 1230 59
rect 1260 161 1324 177
rect 1260 127 1270 161
rect 1304 127 1324 161
rect 1260 93 1324 127
rect 1260 59 1270 93
rect 1304 59 1324 93
rect 1260 47 1324 59
rect 1354 93 1418 177
rect 1354 59 1364 93
rect 1398 59 1418 93
rect 1354 47 1418 59
rect 1448 161 1512 177
rect 1448 127 1458 161
rect 1492 127 1512 161
rect 1448 93 1512 127
rect 1448 59 1458 93
rect 1492 59 1512 93
rect 1448 47 1512 59
rect 1542 161 1594 177
rect 1542 127 1552 161
rect 1586 127 1594 161
rect 1542 93 1594 127
rect 1542 59 1552 93
rect 1586 59 1594 93
rect 1542 47 1594 59
<< pdiff >>
rect 40 485 94 497
rect 40 451 48 485
rect 82 451 94 485
rect 40 417 94 451
rect 40 383 48 417
rect 82 383 94 417
rect 40 347 94 383
rect 40 313 48 347
rect 82 313 94 347
rect 40 297 94 313
rect 130 485 188 497
rect 130 451 142 485
rect 176 451 188 485
rect 130 417 188 451
rect 130 383 142 417
rect 176 383 188 417
rect 130 347 188 383
rect 130 313 142 347
rect 176 313 188 347
rect 130 297 188 313
rect 224 485 282 497
rect 224 451 236 485
rect 270 451 282 485
rect 224 417 282 451
rect 224 383 236 417
rect 270 383 282 417
rect 224 297 282 383
rect 318 485 376 497
rect 318 451 330 485
rect 364 451 376 485
rect 318 417 376 451
rect 318 383 330 417
rect 364 383 376 417
rect 318 347 376 383
rect 318 313 330 347
rect 364 313 376 347
rect 318 297 376 313
rect 412 485 470 497
rect 412 451 424 485
rect 458 451 470 485
rect 412 417 470 451
rect 412 383 424 417
rect 458 383 470 417
rect 412 297 470 383
rect 506 485 564 497
rect 506 451 518 485
rect 552 451 564 485
rect 506 417 564 451
rect 506 383 518 417
rect 552 383 564 417
rect 506 347 564 383
rect 506 313 518 347
rect 552 313 564 347
rect 506 297 564 313
rect 600 485 658 497
rect 600 451 612 485
rect 646 451 658 485
rect 600 417 658 451
rect 600 383 612 417
rect 646 383 658 417
rect 600 297 658 383
rect 694 485 752 497
rect 694 451 706 485
rect 740 451 752 485
rect 694 417 752 451
rect 694 383 706 417
rect 740 383 752 417
rect 694 347 752 383
rect 694 313 706 347
rect 740 313 752 347
rect 694 297 752 313
rect 788 485 846 497
rect 788 451 800 485
rect 834 451 846 485
rect 788 417 846 451
rect 788 383 800 417
rect 834 383 846 417
rect 788 297 846 383
rect 882 485 940 497
rect 882 451 894 485
rect 928 451 940 485
rect 882 417 940 451
rect 882 383 894 417
rect 928 383 940 417
rect 882 347 940 383
rect 882 313 894 347
rect 928 313 940 347
rect 882 297 940 313
rect 976 485 1034 497
rect 976 451 988 485
rect 1022 451 1034 485
rect 976 417 1034 451
rect 976 383 988 417
rect 1022 383 1034 417
rect 976 297 1034 383
rect 1070 485 1128 497
rect 1070 451 1082 485
rect 1116 451 1128 485
rect 1070 417 1128 451
rect 1070 383 1082 417
rect 1116 383 1128 417
rect 1070 347 1128 383
rect 1070 313 1082 347
rect 1116 313 1128 347
rect 1070 297 1128 313
rect 1164 485 1222 497
rect 1164 451 1176 485
rect 1210 451 1222 485
rect 1164 417 1222 451
rect 1164 383 1176 417
rect 1210 383 1222 417
rect 1164 297 1222 383
rect 1258 485 1316 497
rect 1258 451 1270 485
rect 1304 451 1316 485
rect 1258 417 1316 451
rect 1258 383 1270 417
rect 1304 383 1316 417
rect 1258 347 1316 383
rect 1258 313 1270 347
rect 1304 313 1316 347
rect 1258 297 1316 313
rect 1352 485 1410 497
rect 1352 451 1364 485
rect 1398 451 1410 485
rect 1352 417 1410 451
rect 1352 383 1364 417
rect 1398 383 1410 417
rect 1352 297 1410 383
rect 1446 485 1504 497
rect 1446 451 1458 485
rect 1492 451 1504 485
rect 1446 417 1504 451
rect 1446 383 1458 417
rect 1492 383 1504 417
rect 1446 347 1504 383
rect 1446 313 1458 347
rect 1492 313 1504 347
rect 1446 297 1504 313
rect 1540 485 1594 497
rect 1540 451 1552 485
rect 1586 451 1594 485
rect 1540 417 1594 451
rect 1540 383 1552 417
rect 1586 383 1594 417
rect 1540 297 1594 383
<< ndiffc >>
rect 48 127 82 161
rect 48 59 82 93
rect 142 127 176 161
rect 142 59 176 93
rect 236 59 270 93
rect 330 127 364 161
rect 330 59 364 93
rect 424 59 458 93
rect 518 127 552 161
rect 518 59 552 93
rect 612 59 646 93
rect 706 127 740 161
rect 706 59 740 93
rect 800 59 834 93
rect 894 127 928 161
rect 894 59 928 93
rect 988 59 1022 93
rect 1082 127 1116 161
rect 1082 59 1116 93
rect 1176 59 1210 93
rect 1270 127 1304 161
rect 1270 59 1304 93
rect 1364 59 1398 93
rect 1458 127 1492 161
rect 1458 59 1492 93
rect 1552 127 1586 161
rect 1552 59 1586 93
<< pdiffc >>
rect 48 451 82 485
rect 48 383 82 417
rect 48 313 82 347
rect 142 451 176 485
rect 142 383 176 417
rect 142 313 176 347
rect 236 451 270 485
rect 236 383 270 417
rect 330 451 364 485
rect 330 383 364 417
rect 330 313 364 347
rect 424 451 458 485
rect 424 383 458 417
rect 518 451 552 485
rect 518 383 552 417
rect 518 313 552 347
rect 612 451 646 485
rect 612 383 646 417
rect 706 451 740 485
rect 706 383 740 417
rect 706 313 740 347
rect 800 451 834 485
rect 800 383 834 417
rect 894 451 928 485
rect 894 383 928 417
rect 894 313 928 347
rect 988 451 1022 485
rect 988 383 1022 417
rect 1082 451 1116 485
rect 1082 383 1116 417
rect 1082 313 1116 347
rect 1176 451 1210 485
rect 1176 383 1210 417
rect 1270 451 1304 485
rect 1270 383 1304 417
rect 1270 313 1304 347
rect 1364 451 1398 485
rect 1364 383 1398 417
rect 1458 451 1492 485
rect 1458 383 1492 417
rect 1458 313 1492 347
rect 1552 451 1586 485
rect 1552 383 1586 417
<< poly >>
rect 94 497 130 523
rect 188 497 224 523
rect 282 497 318 523
rect 376 497 412 523
rect 470 497 506 523
rect 564 497 600 523
rect 658 497 694 523
rect 752 497 788 523
rect 846 497 882 523
rect 940 497 976 523
rect 1034 497 1070 523
rect 1128 497 1164 523
rect 1222 497 1258 523
rect 1316 497 1352 523
rect 1410 497 1446 523
rect 1504 497 1540 523
rect 94 282 130 297
rect 188 282 224 297
rect 282 282 318 297
rect 376 282 412 297
rect 470 282 506 297
rect 564 282 600 297
rect 658 282 694 297
rect 752 282 788 297
rect 846 282 882 297
rect 940 282 976 297
rect 1034 282 1070 297
rect 1128 282 1164 297
rect 1222 282 1258 297
rect 1316 282 1352 297
rect 1410 282 1446 297
rect 1504 282 1540 297
rect 92 265 132 282
rect 186 265 226 282
rect 280 265 320 282
rect 374 265 414 282
rect 468 265 508 282
rect 562 265 602 282
rect 656 265 696 282
rect 750 265 790 282
rect 844 265 884 282
rect 938 265 978 282
rect 1032 265 1072 282
rect 1126 265 1166 282
rect 1220 265 1260 282
rect 1314 265 1354 282
rect 1408 265 1448 282
rect 1502 265 1542 282
rect 26 249 1542 265
rect 26 215 42 249
rect 76 215 236 249
rect 270 215 424 249
rect 458 215 613 249
rect 647 215 800 249
rect 834 215 988 249
rect 1022 215 1175 249
rect 1209 215 1542 249
rect 26 199 1542 215
rect 102 177 132 199
rect 196 177 226 199
rect 290 177 320 199
rect 384 177 414 199
rect 478 177 508 199
rect 572 177 602 199
rect 666 177 696 199
rect 760 177 790 199
rect 854 177 884 199
rect 948 177 978 199
rect 1042 177 1072 199
rect 1136 177 1166 199
rect 1230 177 1260 199
rect 1324 177 1354 199
rect 1418 177 1448 199
rect 1512 177 1542 199
rect 102 21 132 47
rect 196 21 226 47
rect 290 21 320 47
rect 384 21 414 47
rect 478 21 508 47
rect 572 21 602 47
rect 666 21 696 47
rect 760 21 790 47
rect 854 21 884 47
rect 948 21 978 47
rect 1042 21 1072 47
rect 1136 21 1166 47
rect 1230 21 1260 47
rect 1324 21 1354 47
rect 1418 21 1448 47
rect 1512 21 1542 47
<< polycont >>
rect 42 215 76 249
rect 236 215 270 249
rect 424 215 458 249
rect 613 215 647 249
rect 800 215 834 249
rect 988 215 1022 249
rect 1175 215 1209 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 40 485 82 527
rect 40 451 48 485
rect 40 417 82 451
rect 40 383 48 417
rect 40 347 82 383
rect 40 313 48 347
rect 40 297 82 313
rect 116 485 192 493
rect 116 451 142 485
rect 176 451 192 485
rect 116 417 192 451
rect 116 383 142 417
rect 176 383 192 417
rect 116 347 192 383
rect 236 485 270 527
rect 236 417 270 451
rect 236 367 270 383
rect 304 485 380 493
rect 304 451 330 485
rect 364 451 380 485
rect 304 417 380 451
rect 304 383 330 417
rect 364 383 380 417
rect 116 313 142 347
rect 176 333 192 347
rect 304 347 380 383
rect 424 485 458 527
rect 424 417 458 451
rect 424 367 458 383
rect 492 485 568 493
rect 492 451 518 485
rect 552 451 568 485
rect 492 417 568 451
rect 492 383 518 417
rect 552 383 568 417
rect 304 333 330 347
rect 176 313 330 333
rect 364 333 380 347
rect 492 347 568 383
rect 612 485 646 527
rect 612 417 646 451
rect 612 367 646 383
rect 680 485 756 493
rect 680 451 706 485
rect 740 451 756 485
rect 680 417 756 451
rect 680 383 706 417
rect 740 383 756 417
rect 492 333 518 347
rect 364 313 518 333
rect 552 333 568 347
rect 680 347 756 383
rect 800 485 834 527
rect 800 417 834 451
rect 800 367 834 383
rect 868 485 944 493
rect 868 451 894 485
rect 928 451 944 485
rect 868 417 944 451
rect 868 383 894 417
rect 928 383 944 417
rect 680 333 706 347
rect 552 313 706 333
rect 740 333 756 347
rect 868 347 944 383
rect 988 485 1022 527
rect 988 417 1022 451
rect 988 367 1022 383
rect 1056 485 1132 493
rect 1056 451 1082 485
rect 1116 451 1132 485
rect 1056 417 1132 451
rect 1056 383 1082 417
rect 1116 383 1132 417
rect 868 333 894 347
rect 740 313 894 333
rect 928 333 944 347
rect 1056 347 1132 383
rect 1176 485 1210 527
rect 1176 417 1210 451
rect 1176 367 1210 383
rect 1244 485 1320 493
rect 1244 451 1270 485
rect 1304 451 1320 485
rect 1244 417 1320 451
rect 1244 383 1270 417
rect 1304 383 1320 417
rect 1056 333 1082 347
rect 928 313 1082 333
rect 1116 333 1132 347
rect 1244 347 1320 383
rect 1364 485 1398 527
rect 1364 417 1398 451
rect 1364 367 1398 383
rect 1432 485 1508 493
rect 1432 451 1458 485
rect 1492 451 1508 485
rect 1432 417 1508 451
rect 1432 383 1458 417
rect 1492 383 1508 417
rect 1244 333 1270 347
rect 1116 313 1270 333
rect 1304 333 1320 347
rect 1432 347 1508 383
rect 1552 485 1594 527
rect 1586 451 1594 485
rect 1552 417 1594 451
rect 1586 383 1594 417
rect 1552 367 1594 383
rect 1432 333 1458 347
rect 1304 313 1458 333
rect 1492 313 1508 347
rect 116 299 1508 313
rect 17 249 1225 263
rect 17 215 42 249
rect 76 215 236 249
rect 270 215 424 249
rect 458 215 613 249
rect 647 215 800 249
rect 834 215 988 249
rect 1022 215 1175 249
rect 1209 215 1225 249
rect 1403 181 1508 299
rect 36 161 82 177
rect 36 127 48 161
rect 36 93 82 127
rect 36 59 48 93
rect 36 17 82 59
rect 116 161 1508 181
rect 116 127 142 161
rect 176 143 330 161
rect 176 127 192 143
rect 116 93 192 127
rect 304 127 330 143
rect 364 143 518 161
rect 364 127 380 143
rect 116 59 142 93
rect 176 59 192 93
rect 116 51 192 59
rect 236 93 270 109
rect 236 17 270 59
rect 304 93 380 127
rect 492 127 518 143
rect 552 143 706 161
rect 552 127 568 143
rect 304 59 330 93
rect 364 59 380 93
rect 304 51 380 59
rect 424 93 458 109
rect 424 17 458 59
rect 492 93 568 127
rect 680 127 706 143
rect 740 143 894 161
rect 740 127 756 143
rect 492 59 518 93
rect 552 59 568 93
rect 492 51 568 59
rect 612 93 646 109
rect 612 17 646 59
rect 680 93 756 127
rect 868 127 894 143
rect 928 143 1082 161
rect 928 127 944 143
rect 680 59 706 93
rect 740 59 756 93
rect 680 51 756 59
rect 800 93 834 109
rect 800 17 834 59
rect 868 93 944 127
rect 1056 127 1082 143
rect 1116 143 1270 161
rect 1116 127 1132 143
rect 868 59 894 93
rect 928 59 944 93
rect 868 51 944 59
rect 988 93 1022 109
rect 988 17 1022 59
rect 1056 93 1132 127
rect 1244 127 1270 143
rect 1304 143 1458 161
rect 1304 127 1320 143
rect 1056 59 1082 93
rect 1116 59 1132 93
rect 1056 51 1132 59
rect 1176 93 1210 109
rect 1176 17 1210 59
rect 1244 93 1320 127
rect 1432 127 1458 143
rect 1492 127 1508 161
rect 1244 59 1270 93
rect 1304 59 1320 93
rect 1244 51 1320 59
rect 1364 93 1398 109
rect 1364 17 1398 59
rect 1432 93 1508 127
rect 1432 59 1458 93
rect 1492 59 1508 93
rect 1432 51 1508 59
rect 1552 161 1594 177
rect 1586 127 1594 161
rect 1552 93 1594 127
rect 1586 59 1594 93
rect 1552 17 1594 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
<< metal1 >>
rect 0 561 1656 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 0 496 1656 527
rect 0 17 1656 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
rect 0 -48 1656 -17
<< labels >>
flabel corelocali s 1467 221 1501 255 0 FreeSans 340 0 0 0 Y
port 6 nsew
flabel corelocali s 1467 153 1501 187 0 FreeSans 340 0 0 0 Y
port 6 nsew
flabel corelocali s 29 221 63 255 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 233 221 267 255 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 437 221 471 255 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 641 221 675 255 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 845 221 879 255 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 947 221 981 255 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew
rlabel comment s 0 0 0 0 4 inv_16
<< properties >>
string FIXED_BBOX 0 0 1656 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2097992
string GDS_START 2085580
<< end >>
