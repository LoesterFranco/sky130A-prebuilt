magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 19 195 89 325
rect 376 157 443 337
rect 549 271 630 337
rect 667 157 701 223
rect 745 207 819 331
rect 376 123 701 157
rect 1986 309 2094 479
rect 2046 164 2094 309
rect 1986 61 2094 164
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 36 393 70 493
rect 104 427 180 527
rect 36 382 179 393
rect 36 359 133 382
rect 167 348 179 382
rect 133 161 179 348
rect 35 127 179 161
rect 223 178 269 493
rect 223 144 231 178
rect 265 144 269 178
rect 35 69 69 127
rect 103 17 179 93
rect 223 69 269 144
rect 307 415 362 489
rect 396 449 472 527
rect 579 449 778 483
rect 307 372 708 415
rect 307 89 341 372
rect 477 225 511 372
rect 666 271 708 372
rect 744 399 778 449
rect 822 433 856 527
rect 913 413 960 488
rect 1009 438 1246 472
rect 913 399 947 413
rect 744 365 947 399
rect 1077 382 1175 402
rect 477 191 543 225
rect 913 173 947 365
rect 745 139 947 173
rect 981 207 1039 381
rect 1077 348 1133 382
rect 1167 348 1175 382
rect 1077 331 1175 348
rect 1209 315 1246 438
rect 1280 367 1314 527
rect 1209 297 1337 315
rect 1141 263 1337 297
rect 981 178 1107 207
rect 981 144 1031 178
rect 1065 144 1107 178
rect 981 141 1107 144
rect 745 89 779 139
rect 913 107 947 139
rect 1141 107 1175 263
rect 1371 219 1412 493
rect 1450 433 1657 467
rect 1446 382 1494 393
rect 1446 348 1448 382
rect 1482 348 1494 382
rect 1446 249 1494 348
rect 1209 153 1412 219
rect 1547 207 1589 381
rect 307 55 381 89
rect 415 17 481 89
rect 614 55 779 89
rect 823 17 863 105
rect 913 73 983 107
rect 1027 73 1175 107
rect 1245 17 1319 117
rect 1355 107 1412 153
rect 1450 178 1589 207
rect 1450 144 1462 178
rect 1496 144 1589 178
rect 1450 141 1589 144
rect 1623 265 1657 433
rect 1693 427 1754 527
rect 1824 381 1881 491
rect 1691 315 1881 381
rect 1918 325 1952 527
rect 1844 265 1881 315
rect 1623 199 1810 265
rect 1844 199 2006 265
rect 1623 107 1657 199
rect 1844 165 1880 199
rect 1355 73 1452 107
rect 1491 73 1657 107
rect 1691 17 1754 123
rect 1808 60 1880 165
rect 1918 17 1952 139
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 133 348 167 382
rect 231 144 265 178
rect 1133 348 1167 382
rect 1031 144 1065 178
rect 1448 348 1482 382
rect 1462 144 1496 178
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
<< metal1 >>
rect 0 561 2116 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 0 496 2116 527
rect 0 17 2116 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
rect 0 -48 2116 -17
<< obsm1 >>
rect 121 382 1494 388
rect 121 348 133 382
rect 167 360 1133 382
rect 167 348 179 360
rect 121 342 179 348
rect 1111 348 1133 360
rect 1167 360 1448 382
rect 1167 348 1179 360
rect 1111 342 1179 348
rect 1426 348 1448 360
rect 1482 348 1494 382
rect 1426 342 1494 348
rect 219 178 1508 184
rect 219 144 231 178
rect 265 156 1031 178
rect 265 144 277 156
rect 219 138 277 144
rect 1009 144 1031 156
rect 1065 156 1462 178
rect 1065 144 1077 156
rect 1009 138 1077 144
rect 1446 144 1462 156
rect 1496 144 1508 178
rect 1446 138 1508 144
<< labels >>
rlabel locali s 19 195 89 325 6 CLK
port 1 nsew signal input
rlabel locali s 549 271 630 337 6 D
port 2 nsew signal input
rlabel locali s 2046 164 2094 309 6 Q
port 3 nsew signal output
rlabel locali s 1986 309 2094 479 6 Q
port 3 nsew signal output
rlabel locali s 1986 61 2094 164 6 Q
port 3 nsew signal output
rlabel locali s 745 207 819 331 6 SCD
port 4 nsew signal input
rlabel locali s 667 157 701 223 6 SCE
port 5 nsew signal input
rlabel locali s 376 157 443 337 6 SCE
port 5 nsew signal input
rlabel locali s 376 123 701 157 6 SCE
port 5 nsew signal input
rlabel metal1 s 0 -48 2116 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 2116 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2116 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 336706
string GDS_START 321576
<< end >>
