magic
tech sky130A
magscale 1 2
timestamp 1599588218
<< nwell >>
rect -38 332 1766 704
rect 307 312 1416 332
rect 1005 306 1416 312
<< pwell >>
rect 0 0 1728 49
<< scpmos >>
rect 83 424 119 592
rect 235 424 271 592
rect 454 392 490 560
rect 578 392 614 592
rect 662 392 698 592
rect 769 508 805 592
rect 906 508 942 592
rect 1091 342 1127 566
rect 1183 342 1219 566
rect 1289 342 1325 566
rect 1501 384 1537 552
rect 1609 368 1645 592
<< nmoslvt >>
rect 85 112 115 222
rect 201 74 231 222
rect 430 74 460 222
rect 578 74 608 202
rect 656 74 686 202
rect 811 118 841 202
rect 889 118 919 202
rect 1103 74 1133 222
rect 1181 74 1211 222
rect 1289 74 1319 222
rect 1507 112 1537 222
rect 1610 74 1640 222
<< ndiff >>
rect 28 180 85 222
rect 28 146 40 180
rect 74 146 85 180
rect 28 112 85 146
rect 115 202 201 222
rect 115 168 142 202
rect 176 168 201 202
rect 115 120 201 168
rect 115 112 142 120
rect 130 86 142 112
rect 176 86 201 120
rect 130 74 201 86
rect 231 202 288 222
rect 231 168 242 202
rect 276 168 288 202
rect 231 120 288 168
rect 231 86 242 120
rect 276 86 288 120
rect 231 74 288 86
rect 373 192 430 222
rect 373 158 385 192
rect 419 158 430 192
rect 373 120 430 158
rect 373 86 385 120
rect 419 86 430 120
rect 373 74 430 86
rect 460 202 510 222
rect 460 120 578 202
rect 460 86 509 120
rect 543 86 578 120
rect 460 74 578 86
rect 608 74 656 202
rect 686 122 811 202
rect 686 88 727 122
rect 761 118 811 122
rect 841 118 889 202
rect 919 177 992 202
rect 919 143 946 177
rect 980 143 992 177
rect 919 118 992 143
rect 1046 194 1103 222
rect 1046 160 1058 194
rect 1092 160 1103 194
rect 1046 120 1103 160
rect 761 88 796 118
rect 686 74 796 88
rect 1046 86 1058 120
rect 1092 86 1103 120
rect 1046 74 1103 86
rect 1133 74 1181 222
rect 1211 197 1289 222
rect 1211 163 1222 197
rect 1256 163 1289 197
rect 1211 116 1289 163
rect 1211 82 1222 116
rect 1256 82 1289 116
rect 1211 74 1289 82
rect 1319 210 1376 222
rect 1319 176 1330 210
rect 1364 176 1376 210
rect 1319 120 1376 176
rect 1319 86 1330 120
rect 1364 86 1376 120
rect 1437 184 1507 222
rect 1437 150 1462 184
rect 1496 150 1507 184
rect 1437 112 1507 150
rect 1537 210 1610 222
rect 1537 176 1565 210
rect 1599 176 1610 210
rect 1537 116 1610 176
rect 1537 112 1565 116
rect 1319 74 1376 86
rect 1552 82 1565 112
rect 1599 82 1610 116
rect 1552 74 1610 82
rect 1640 210 1697 222
rect 1640 176 1651 210
rect 1685 176 1697 210
rect 1640 120 1697 176
rect 1640 86 1651 120
rect 1685 86 1697 120
rect 1640 74 1697 86
<< pdiff >>
rect 505 614 563 626
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 470 83 546
rect 27 436 39 470
rect 73 436 83 470
rect 27 424 83 436
rect 119 584 235 592
rect 119 550 129 584
rect 163 550 235 584
rect 119 516 235 550
rect 119 482 129 516
rect 163 482 235 516
rect 119 424 235 482
rect 271 483 327 592
rect 505 580 517 614
rect 551 592 563 614
rect 551 580 578 592
rect 505 560 578 580
rect 271 449 281 483
rect 315 449 327 483
rect 271 424 327 449
rect 381 394 454 560
rect 381 360 393 394
rect 427 392 454 394
rect 490 392 578 560
rect 614 392 662 592
rect 698 531 769 592
rect 698 497 708 531
rect 742 508 769 531
rect 805 508 906 592
rect 942 566 992 592
rect 1557 580 1609 592
rect 942 554 1091 566
rect 942 520 952 554
rect 986 520 1039 554
rect 1073 520 1091 554
rect 942 508 1091 520
rect 742 497 754 508
rect 698 392 754 497
rect 427 360 439 392
rect 381 348 439 360
rect 1041 342 1091 508
rect 1127 554 1183 566
rect 1127 520 1139 554
rect 1173 520 1183 554
rect 1127 474 1183 520
rect 1127 440 1139 474
rect 1173 440 1183 474
rect 1127 394 1183 440
rect 1127 360 1139 394
rect 1173 360 1183 394
rect 1127 342 1183 360
rect 1219 547 1289 566
rect 1219 513 1239 547
rect 1273 513 1289 547
rect 1219 446 1289 513
rect 1219 412 1239 446
rect 1273 412 1289 446
rect 1219 342 1289 412
rect 1325 554 1380 566
rect 1325 520 1338 554
rect 1372 520 1380 554
rect 1557 552 1565 580
rect 1325 472 1380 520
rect 1325 438 1338 472
rect 1372 438 1380 472
rect 1325 394 1380 438
rect 1325 360 1338 394
rect 1372 360 1380 394
rect 1449 540 1501 552
rect 1449 506 1457 540
rect 1491 506 1501 540
rect 1449 430 1501 506
rect 1449 396 1457 430
rect 1491 396 1501 430
rect 1449 384 1501 396
rect 1537 546 1565 552
rect 1599 546 1609 580
rect 1537 497 1609 546
rect 1537 463 1565 497
rect 1599 463 1609 497
rect 1537 414 1609 463
rect 1537 384 1565 414
rect 1325 342 1380 360
rect 1557 380 1565 384
rect 1599 380 1609 414
rect 1557 368 1609 380
rect 1645 580 1701 592
rect 1645 546 1655 580
rect 1689 546 1701 580
rect 1645 497 1701 546
rect 1645 463 1655 497
rect 1689 463 1701 497
rect 1645 414 1701 463
rect 1645 380 1655 414
rect 1689 380 1701 414
rect 1645 368 1701 380
<< ndiffc >>
rect 40 146 74 180
rect 142 168 176 202
rect 142 86 176 120
rect 242 168 276 202
rect 242 86 276 120
rect 385 158 419 192
rect 385 86 419 120
rect 509 86 543 120
rect 727 88 761 122
rect 946 143 980 177
rect 1058 160 1092 194
rect 1058 86 1092 120
rect 1222 163 1256 197
rect 1222 82 1256 116
rect 1330 176 1364 210
rect 1330 86 1364 120
rect 1462 150 1496 184
rect 1565 176 1599 210
rect 1565 82 1599 116
rect 1651 176 1685 210
rect 1651 86 1685 120
<< pdiffc >>
rect 39 546 73 580
rect 39 436 73 470
rect 129 550 163 584
rect 129 482 163 516
rect 517 580 551 614
rect 281 449 315 483
rect 393 360 427 394
rect 708 497 742 531
rect 952 520 986 554
rect 1039 520 1073 554
rect 1139 520 1173 554
rect 1139 440 1173 474
rect 1139 360 1173 394
rect 1239 513 1273 547
rect 1239 412 1273 446
rect 1338 520 1372 554
rect 1338 438 1372 472
rect 1338 360 1372 394
rect 1457 506 1491 540
rect 1457 396 1491 430
rect 1565 546 1599 580
rect 1565 463 1599 497
rect 1565 380 1599 414
rect 1655 546 1689 580
rect 1655 463 1689 497
rect 1655 380 1689 414
<< poly >>
rect 83 592 119 618
rect 235 592 271 618
rect 454 560 490 586
rect 578 592 614 618
rect 662 592 698 618
rect 769 592 805 618
rect 906 592 942 618
rect 1609 592 1645 618
rect 83 386 119 424
rect 235 386 271 424
rect 83 370 153 386
rect 83 336 103 370
rect 137 336 153 370
rect 83 302 153 336
rect 83 268 103 302
rect 137 268 153 302
rect 83 252 153 268
rect 201 370 271 386
rect 201 336 217 370
rect 251 336 271 370
rect 1091 566 1127 592
rect 1183 566 1219 592
rect 1289 566 1325 592
rect 769 476 805 508
rect 769 460 858 476
rect 769 426 808 460
rect 842 426 858 460
rect 769 410 858 426
rect 906 458 942 508
rect 906 442 972 458
rect 906 408 922 442
rect 956 408 972 442
rect 906 392 972 408
rect 201 302 271 336
rect 454 310 490 392
rect 578 360 614 392
rect 548 344 614 360
rect 548 310 564 344
rect 598 310 614 344
rect 662 368 698 392
rect 906 368 936 392
rect 662 338 805 368
rect 201 268 217 302
rect 251 268 271 302
rect 201 252 271 268
rect 430 294 503 310
rect 548 294 614 310
rect 430 260 453 294
rect 487 260 503 294
rect 85 222 115 252
rect 201 222 231 252
rect 430 244 503 260
rect 430 222 460 244
rect 85 86 115 112
rect 578 202 608 294
rect 775 290 805 338
rect 889 338 936 368
rect 1501 552 1537 578
rect 1501 352 1537 384
rect 656 274 722 290
rect 656 240 672 274
rect 706 240 722 274
rect 656 224 722 240
rect 775 274 841 290
rect 775 240 791 274
rect 825 240 841 274
rect 775 224 841 240
rect 656 202 686 224
rect 811 202 841 224
rect 889 202 919 338
rect 1091 310 1127 342
rect 1183 310 1219 342
rect 1289 316 1325 342
rect 1455 316 1537 352
rect 1609 326 1645 368
rect 968 294 1127 310
rect 968 260 984 294
rect 1018 274 1127 294
rect 1175 294 1241 310
rect 1018 260 1133 274
rect 968 244 1133 260
rect 1175 260 1191 294
rect 1225 260 1241 294
rect 1175 244 1241 260
rect 1289 294 1537 316
rect 1289 260 1312 294
rect 1346 260 1537 294
rect 1579 310 1645 326
rect 1579 276 1595 310
rect 1629 276 1645 310
rect 1579 260 1645 276
rect 1289 244 1537 260
rect 1103 222 1133 244
rect 1181 222 1211 244
rect 1289 222 1319 244
rect 1507 222 1537 244
rect 1610 222 1640 260
rect 811 92 841 118
rect 889 92 919 118
rect 1507 86 1537 112
rect 201 48 231 74
rect 430 48 460 74
rect 578 48 608 74
rect 656 48 686 74
rect 1103 48 1133 74
rect 1181 48 1211 74
rect 1289 48 1319 74
rect 1610 48 1640 74
<< polycont >>
rect 103 336 137 370
rect 103 268 137 302
rect 217 336 251 370
rect 808 426 842 460
rect 922 408 956 442
rect 564 310 598 344
rect 217 268 251 302
rect 453 260 487 294
rect 672 240 706 274
rect 791 240 825 274
rect 984 260 1018 294
rect 1191 260 1225 294
rect 1312 260 1346 294
rect 1595 276 1629 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 19 580 73 596
rect 19 546 39 580
rect 19 470 73 546
rect 113 584 179 649
rect 113 550 129 584
rect 163 550 179 584
rect 501 614 567 649
rect 501 580 517 614
rect 551 580 567 614
rect 624 581 858 615
rect 113 516 179 550
rect 113 482 129 516
rect 163 482 179 516
rect 213 546 403 580
rect 19 436 39 470
rect 213 448 247 546
rect 369 512 582 546
rect 73 436 247 448
rect 19 414 247 436
rect 281 483 335 512
rect 315 478 335 483
rect 315 449 511 478
rect 281 444 511 449
rect 281 420 335 444
rect 19 218 53 414
rect 87 370 167 380
rect 87 336 103 370
rect 137 336 167 370
rect 87 302 167 336
rect 87 268 103 302
rect 137 268 167 302
rect 87 252 167 268
rect 201 370 267 380
rect 201 336 217 370
rect 251 336 267 370
rect 201 302 267 336
rect 201 268 217 302
rect 251 268 267 302
rect 201 252 267 268
rect 301 218 335 420
rect 19 180 90 218
rect 19 146 40 180
rect 74 146 90 180
rect 19 108 90 146
rect 126 202 192 218
rect 126 168 142 202
rect 176 168 192 202
rect 126 120 192 168
rect 126 86 142 120
rect 176 86 192 120
rect 126 17 192 86
rect 226 202 335 218
rect 226 168 242 202
rect 276 168 335 202
rect 226 120 335 168
rect 226 86 242 120
rect 276 86 335 120
rect 226 70 335 86
rect 369 394 443 410
rect 369 360 393 394
rect 427 360 443 394
rect 369 344 443 360
rect 369 192 403 344
rect 477 310 511 444
rect 437 294 511 310
rect 548 360 582 512
rect 624 428 658 581
rect 692 531 758 547
rect 692 497 708 531
rect 742 497 758 531
rect 692 481 758 497
rect 624 394 690 428
rect 548 344 614 360
rect 548 310 564 344
rect 598 310 614 344
rect 548 294 614 310
rect 437 260 453 294
rect 487 260 511 294
rect 656 290 690 394
rect 724 358 758 481
rect 792 460 858 581
rect 936 554 1089 649
rect 936 520 952 554
rect 986 520 1039 554
rect 1073 520 1089 554
rect 936 504 1089 520
rect 1123 554 1189 570
rect 1123 520 1139 554
rect 1173 520 1189 554
rect 792 426 808 460
rect 842 426 858 460
rect 1123 474 1189 520
rect 1123 458 1139 474
rect 792 410 858 426
rect 906 442 1139 458
rect 906 408 922 442
rect 956 440 1139 442
rect 1173 440 1189 474
rect 956 408 1189 440
rect 1223 547 1289 649
rect 1549 580 1602 649
rect 1223 513 1239 547
rect 1273 513 1289 547
rect 1223 446 1289 513
rect 1223 412 1239 446
rect 1273 412 1289 446
rect 1338 554 1423 570
rect 1372 520 1423 554
rect 1338 472 1423 520
rect 1372 438 1423 472
rect 906 394 1189 408
rect 906 392 1139 394
rect 1058 360 1139 392
rect 1173 378 1189 394
rect 1338 394 1423 438
rect 1173 360 1304 378
rect 724 324 945 358
rect 875 310 945 324
rect 1058 344 1304 360
rect 1372 360 1423 394
rect 1338 344 1423 360
rect 875 294 1024 310
rect 656 274 722 290
rect 656 260 672 274
rect 437 240 672 260
rect 706 240 722 274
rect 437 226 722 240
rect 656 224 722 226
rect 775 274 841 290
rect 775 240 791 274
rect 825 240 841 274
rect 369 158 385 192
rect 419 190 435 192
rect 775 190 841 240
rect 419 158 841 190
rect 369 156 841 158
rect 875 260 984 294
rect 1018 260 1024 294
rect 875 244 1024 260
rect 369 120 435 156
rect 875 122 909 244
rect 1058 210 1092 344
rect 1270 310 1304 344
rect 1175 294 1236 310
rect 1175 260 1191 294
rect 1225 260 1236 294
rect 1175 236 1236 260
rect 1270 294 1355 310
rect 1270 260 1312 294
rect 1346 260 1355 294
rect 1270 244 1355 260
rect 1389 210 1423 344
rect 369 86 385 120
rect 419 86 435 120
rect 369 70 435 86
rect 469 86 509 120
rect 543 86 583 120
rect 469 17 583 86
rect 681 88 727 122
rect 761 88 909 122
rect 681 72 909 88
rect 946 177 996 206
rect 980 143 996 177
rect 946 17 996 143
rect 1042 194 1092 210
rect 1042 160 1058 194
rect 1042 120 1092 160
rect 1042 86 1058 120
rect 1042 70 1092 86
rect 1206 197 1272 202
rect 1206 163 1222 197
rect 1256 163 1272 197
rect 1206 116 1272 163
rect 1206 82 1222 116
rect 1256 82 1272 116
rect 1206 17 1272 82
rect 1313 176 1330 210
rect 1364 176 1423 210
rect 1313 120 1423 176
rect 1313 86 1330 120
rect 1364 86 1423 120
rect 1457 540 1507 556
rect 1491 506 1507 540
rect 1457 430 1507 506
rect 1491 396 1507 430
rect 1457 326 1507 396
rect 1549 546 1565 580
rect 1599 546 1602 580
rect 1549 497 1602 546
rect 1549 463 1565 497
rect 1599 463 1602 497
rect 1549 414 1602 463
rect 1549 380 1565 414
rect 1599 380 1602 414
rect 1549 364 1602 380
rect 1639 580 1706 596
rect 1639 546 1655 580
rect 1689 546 1706 580
rect 1639 497 1706 546
rect 1639 463 1655 497
rect 1689 463 1706 497
rect 1639 414 1706 463
rect 1639 380 1655 414
rect 1689 380 1706 414
rect 1639 364 1706 380
rect 1457 310 1638 326
rect 1457 276 1595 310
rect 1629 276 1638 310
rect 1457 260 1638 276
rect 1457 184 1512 260
rect 1672 226 1706 364
rect 1457 150 1462 184
rect 1496 150 1512 184
rect 1457 108 1512 150
rect 1549 210 1615 226
rect 1549 176 1565 210
rect 1599 176 1615 210
rect 1549 116 1615 176
rect 1313 70 1423 86
rect 1549 82 1565 116
rect 1599 82 1615 116
rect 1549 17 1615 82
rect 1649 210 1706 226
rect 1649 176 1651 210
rect 1685 176 1706 210
rect 1649 120 1706 176
rect 1649 86 1651 120
rect 1685 86 1706 120
rect 1649 70 1706 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
<< metal1 >>
rect 0 683 1728 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 0 617 1728 649
rect 0 17 1728 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
rect 0 -49 1728 -17
<< labels >>
flabel pwell s 0 0 1728 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 0 617 1728 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
rlabel comment s 0 0 0 0 4 dlrbn_1
flabel metal1 s 0 617 1728 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 1728 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 1663 390 1697 424 0 FreeSans 340 0 0 0 Q_N
port 9 nsew
flabel corelocali s 1663 464 1697 498 0 FreeSans 340 0 0 0 Q_N
port 9 nsew
flabel corelocali s 1663 538 1697 572 0 FreeSans 340 0 0 0 Q_N
port 9 nsew
flabel corelocali s 1375 94 1409 128 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 1375 168 1409 202 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 1375 390 1409 424 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 1375 464 1409 498 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew
flabel corelocali s 1183 242 1217 276 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 1728 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 2979232
string GDS_START 2966006
<< end >>
