magic
tech sky130A
magscale 1 2
timestamp 1604502705
<< nwell >>
rect -38 332 1478 704
<< pwell >>
rect 0 0 1440 49
<< scnmos >>
rect 162 74 192 222
rect 248 74 278 222
rect 334 74 364 222
rect 420 74 450 222
rect 556 94 586 222
rect 642 94 672 222
rect 872 74 902 222
rect 1062 74 1092 202
rect 1148 74 1178 202
rect 1234 74 1264 202
rect 1328 74 1358 202
<< pmoshvt >>
rect 175 368 205 592
rect 265 368 295 592
rect 355 368 385 592
rect 445 368 475 592
rect 553 368 583 592
rect 631 368 661 592
rect 875 392 905 592
rect 965 392 995 592
rect 1055 392 1085 592
rect 1145 392 1175 592
rect 1235 392 1265 592
rect 1325 392 1355 592
<< ndiff >>
rect 109 142 162 222
rect 109 108 117 142
rect 151 108 162 142
rect 109 74 162 108
rect 192 210 248 222
rect 192 176 203 210
rect 237 176 248 210
rect 192 120 248 176
rect 192 86 203 120
rect 237 86 248 120
rect 192 74 248 86
rect 278 142 334 222
rect 278 108 289 142
rect 323 108 334 142
rect 278 74 334 108
rect 364 210 420 222
rect 364 176 375 210
rect 409 176 420 210
rect 364 120 420 176
rect 364 86 375 120
rect 409 86 420 120
rect 364 74 420 86
rect 450 152 556 222
rect 450 118 461 152
rect 495 118 556 152
rect 450 94 556 118
rect 586 178 642 222
rect 586 144 597 178
rect 631 144 642 178
rect 586 94 642 144
rect 672 152 872 222
rect 672 118 740 152
rect 774 118 827 152
rect 861 118 872 152
rect 672 94 872 118
rect 450 74 503 94
rect 819 74 872 94
rect 902 210 955 222
rect 902 176 913 210
rect 947 176 955 210
rect 902 120 955 176
rect 902 86 913 120
rect 947 86 955 120
rect 902 74 955 86
rect 1009 189 1062 202
rect 1009 155 1017 189
rect 1051 155 1062 189
rect 1009 74 1062 155
rect 1092 120 1148 202
rect 1092 86 1103 120
rect 1137 86 1148 120
rect 1092 74 1148 86
rect 1178 190 1234 202
rect 1178 156 1189 190
rect 1223 156 1234 190
rect 1178 120 1234 156
rect 1178 86 1189 120
rect 1223 86 1234 120
rect 1178 74 1234 86
rect 1264 127 1328 202
rect 1264 93 1279 127
rect 1313 93 1328 127
rect 1264 74 1328 93
rect 1358 190 1411 202
rect 1358 156 1369 190
rect 1403 156 1411 190
rect 1358 120 1411 156
rect 1358 86 1369 120
rect 1403 86 1411 120
rect 1358 74 1411 86
<< pdiff >>
rect 120 580 175 592
rect 120 546 128 580
rect 162 546 175 580
rect 120 478 175 546
rect 120 444 128 478
rect 162 444 175 478
rect 120 368 175 444
rect 205 580 265 592
rect 205 546 218 580
rect 252 546 265 580
rect 205 497 265 546
rect 205 463 218 497
rect 252 463 265 497
rect 205 414 265 463
rect 205 380 218 414
rect 252 380 265 414
rect 205 368 265 380
rect 295 580 355 592
rect 295 546 308 580
rect 342 546 355 580
rect 295 478 355 546
rect 295 444 308 478
rect 342 444 355 478
rect 295 368 355 444
rect 385 580 445 592
rect 385 546 398 580
rect 432 546 445 580
rect 385 497 445 546
rect 385 463 398 497
rect 432 463 445 497
rect 385 414 445 463
rect 385 380 398 414
rect 432 380 445 414
rect 385 368 445 380
rect 475 580 553 592
rect 475 546 502 580
rect 536 546 553 580
rect 475 510 553 546
rect 475 476 502 510
rect 536 476 553 510
rect 475 440 553 476
rect 475 406 502 440
rect 536 406 553 440
rect 475 368 553 406
rect 583 368 631 592
rect 661 580 716 592
rect 661 546 674 580
rect 708 546 716 580
rect 661 510 716 546
rect 661 476 674 510
rect 708 476 716 510
rect 661 440 716 476
rect 661 406 674 440
rect 708 406 716 440
rect 661 368 716 406
rect 820 580 875 592
rect 820 546 828 580
rect 862 546 875 580
rect 820 508 875 546
rect 820 474 828 508
rect 862 474 875 508
rect 820 392 875 474
rect 905 531 965 592
rect 905 497 918 531
rect 952 497 965 531
rect 905 438 965 497
rect 905 404 918 438
rect 952 404 965 438
rect 905 392 965 404
rect 995 580 1055 592
rect 995 546 1008 580
rect 1042 546 1055 580
rect 995 510 1055 546
rect 995 476 1008 510
rect 1042 476 1055 510
rect 995 440 1055 476
rect 995 406 1008 440
rect 1042 406 1055 440
rect 995 392 1055 406
rect 1085 580 1145 592
rect 1085 546 1098 580
rect 1132 546 1145 580
rect 1085 508 1145 546
rect 1085 474 1098 508
rect 1132 474 1145 508
rect 1085 392 1145 474
rect 1175 580 1235 592
rect 1175 546 1188 580
rect 1222 546 1235 580
rect 1175 510 1235 546
rect 1175 476 1188 510
rect 1222 476 1235 510
rect 1175 440 1235 476
rect 1175 406 1188 440
rect 1222 406 1235 440
rect 1175 392 1235 406
rect 1265 580 1325 592
rect 1265 546 1278 580
rect 1312 546 1325 580
rect 1265 508 1325 546
rect 1265 474 1278 508
rect 1312 474 1325 508
rect 1265 392 1325 474
rect 1355 580 1410 592
rect 1355 546 1368 580
rect 1402 546 1410 580
rect 1355 510 1410 546
rect 1355 476 1368 510
rect 1402 476 1410 510
rect 1355 440 1410 476
rect 1355 406 1368 440
rect 1402 406 1410 440
rect 1355 392 1410 406
<< ndiffc >>
rect 117 108 151 142
rect 203 176 237 210
rect 203 86 237 120
rect 289 108 323 142
rect 375 176 409 210
rect 375 86 409 120
rect 461 118 495 152
rect 597 144 631 178
rect 740 118 774 152
rect 827 118 861 152
rect 913 176 947 210
rect 913 86 947 120
rect 1017 155 1051 189
rect 1103 86 1137 120
rect 1189 156 1223 190
rect 1189 86 1223 120
rect 1279 93 1313 127
rect 1369 156 1403 190
rect 1369 86 1403 120
<< pdiffc >>
rect 128 546 162 580
rect 128 444 162 478
rect 218 546 252 580
rect 218 463 252 497
rect 218 380 252 414
rect 308 546 342 580
rect 308 444 342 478
rect 398 546 432 580
rect 398 463 432 497
rect 398 380 432 414
rect 502 546 536 580
rect 502 476 536 510
rect 502 406 536 440
rect 674 546 708 580
rect 674 476 708 510
rect 674 406 708 440
rect 828 546 862 580
rect 828 474 862 508
rect 918 497 952 531
rect 918 404 952 438
rect 1008 546 1042 580
rect 1008 476 1042 510
rect 1008 406 1042 440
rect 1098 546 1132 580
rect 1098 474 1132 508
rect 1188 546 1222 580
rect 1188 476 1222 510
rect 1188 406 1222 440
rect 1278 546 1312 580
rect 1278 474 1312 508
rect 1368 546 1402 580
rect 1368 476 1402 510
rect 1368 406 1402 440
<< poly >>
rect 175 592 205 618
rect 265 592 295 618
rect 355 592 385 618
rect 445 592 475 618
rect 553 592 583 618
rect 631 592 661 618
rect 875 592 905 618
rect 965 592 995 618
rect 1055 592 1085 618
rect 1145 592 1175 618
rect 1235 592 1265 618
rect 1325 592 1355 618
rect 875 377 905 392
rect 965 377 995 392
rect 1055 377 1085 392
rect 1145 377 1175 392
rect 1235 377 1265 392
rect 1325 377 1355 392
rect 175 353 205 368
rect 265 353 295 368
rect 355 353 385 368
rect 445 353 475 368
rect 553 353 583 368
rect 631 353 661 368
rect 872 360 908 377
rect 962 360 998 377
rect 172 326 208 353
rect 262 326 298 353
rect 352 326 388 353
rect 442 326 478 353
rect 550 336 586 353
rect 162 310 478 326
rect 162 276 223 310
rect 257 276 291 310
rect 325 276 359 310
rect 393 276 427 310
rect 461 276 478 310
rect 162 260 478 276
rect 520 320 586 336
rect 520 286 536 320
rect 570 286 586 320
rect 520 270 586 286
rect 628 336 664 353
rect 764 344 998 360
rect 628 320 722 336
rect 628 286 672 320
rect 706 286 722 320
rect 764 310 780 344
rect 814 330 998 344
rect 814 310 830 330
rect 764 294 830 310
rect 628 270 722 286
rect 162 222 192 260
rect 248 222 278 260
rect 334 222 364 260
rect 420 222 450 260
rect 556 222 586 270
rect 642 222 672 270
rect 872 222 902 330
rect 1052 318 1088 377
rect 1142 318 1178 377
rect 1052 302 1178 318
rect 1052 268 1097 302
rect 1131 268 1178 302
rect 1052 252 1178 268
rect 1232 318 1268 377
rect 1322 318 1358 377
rect 1232 302 1358 318
rect 1232 268 1289 302
rect 1323 268 1358 302
rect 1232 252 1358 268
rect 162 48 192 74
rect 248 48 278 74
rect 334 48 364 74
rect 420 48 450 74
rect 556 68 586 94
rect 642 68 672 94
rect 1062 202 1092 252
rect 1148 202 1178 252
rect 1234 202 1264 252
rect 1328 202 1358 252
rect 872 48 902 74
rect 1062 48 1092 74
rect 1148 48 1178 74
rect 1234 48 1264 74
rect 1328 48 1358 74
<< polycont >>
rect 223 276 257 310
rect 291 276 325 310
rect 359 276 393 310
rect 427 276 461 310
rect 536 286 570 320
rect 672 286 706 320
rect 780 310 814 344
rect 1097 268 1131 302
rect 1289 268 1323 302
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 112 580 162 649
rect 112 546 128 580
rect 112 478 162 546
rect 112 444 128 478
rect 112 428 162 444
rect 202 580 268 596
rect 202 546 218 580
rect 252 546 268 580
rect 202 497 268 546
rect 202 463 218 497
rect 252 463 268 497
rect 202 414 268 463
rect 308 580 342 649
rect 308 478 342 546
rect 308 428 342 444
rect 382 580 448 596
rect 382 546 398 580
rect 432 546 448 580
rect 382 497 448 546
rect 382 463 398 497
rect 432 463 448 497
rect 202 394 218 414
rect 133 380 218 394
rect 252 394 268 414
rect 382 414 448 463
rect 382 394 398 414
rect 252 380 398 394
rect 432 380 448 414
rect 482 580 556 649
rect 482 546 502 580
rect 536 546 556 580
rect 482 510 556 546
rect 482 476 502 510
rect 536 476 556 510
rect 482 440 556 476
rect 482 406 502 440
rect 536 406 556 440
rect 658 580 724 596
rect 658 546 674 580
rect 708 546 724 580
rect 658 510 724 546
rect 658 476 674 510
rect 708 476 724 510
rect 658 440 724 476
rect 812 581 1042 615
rect 812 580 878 581
rect 812 546 828 580
rect 862 546 878 580
rect 992 580 1042 581
rect 812 508 878 546
rect 812 474 828 508
rect 862 474 878 508
rect 812 458 878 474
rect 913 531 952 547
rect 913 497 918 531
rect 658 424 674 440
rect 482 390 556 406
rect 604 406 674 424
rect 708 424 724 440
rect 913 438 952 497
rect 708 406 830 424
rect 604 390 830 406
rect 133 360 448 380
rect 133 356 167 360
rect 25 226 167 356
rect 207 310 477 326
rect 207 276 223 310
rect 257 276 291 310
rect 325 276 359 310
rect 393 276 427 310
rect 461 276 477 310
rect 207 260 477 276
rect 511 320 570 356
rect 511 286 536 320
rect 511 270 570 286
rect 443 236 477 260
rect 25 210 409 226
rect 25 192 203 210
rect 187 176 203 192
rect 237 192 375 210
rect 101 142 151 158
rect 101 108 117 142
rect 101 17 151 108
rect 187 120 237 176
rect 359 176 375 192
rect 443 202 563 236
rect 604 226 638 390
rect 672 320 737 356
rect 706 286 737 320
rect 771 344 830 390
rect 771 310 780 344
rect 814 310 830 344
rect 771 294 830 310
rect 913 404 918 438
rect 672 270 737 286
rect 913 236 952 404
rect 992 546 1008 580
rect 992 510 1042 546
rect 992 476 1008 510
rect 992 440 1042 476
rect 1082 580 1132 649
rect 1082 546 1098 580
rect 1082 508 1132 546
rect 1082 474 1098 508
rect 1082 458 1132 474
rect 1172 580 1238 596
rect 1172 546 1188 580
rect 1222 546 1238 580
rect 1172 510 1238 546
rect 1172 476 1188 510
rect 1222 476 1238 510
rect 992 406 1008 440
rect 1172 440 1238 476
rect 1278 580 1312 649
rect 1278 508 1312 546
rect 1278 458 1312 474
rect 1352 580 1418 596
rect 1352 546 1368 580
rect 1402 546 1418 580
rect 1352 510 1418 546
rect 1352 476 1368 510
rect 1402 476 1418 510
rect 1172 424 1188 440
rect 1042 406 1188 424
rect 1222 424 1238 440
rect 1352 440 1418 476
rect 1352 424 1368 440
rect 1222 406 1368 424
rect 1402 406 1418 440
rect 992 390 1418 406
rect 1081 302 1223 356
rect 1081 268 1097 302
rect 1131 268 1223 302
rect 1081 252 1223 268
rect 1273 302 1415 356
rect 1273 268 1289 302
rect 1323 268 1415 302
rect 1273 252 1415 268
rect 187 86 203 120
rect 187 70 237 86
rect 273 142 323 158
rect 273 108 289 142
rect 273 17 323 108
rect 359 120 409 176
rect 359 86 375 120
rect 359 70 409 86
rect 445 152 495 168
rect 445 118 461 152
rect 445 17 495 118
rect 529 85 563 202
rect 597 178 638 226
rect 631 144 638 178
rect 597 119 638 144
rect 672 210 963 236
rect 672 202 913 210
rect 672 85 706 202
rect 947 176 963 210
rect 529 51 706 85
rect 740 152 877 168
rect 774 118 827 152
rect 861 118 877 152
rect 740 17 877 118
rect 913 120 963 176
rect 1001 190 1419 218
rect 1001 189 1189 190
rect 1001 155 1017 189
rect 1051 156 1189 189
rect 1223 184 1369 190
rect 1051 155 1223 156
rect 1001 154 1223 155
rect 1189 120 1223 154
rect 1403 156 1419 190
rect 947 86 1103 120
rect 1137 86 1153 120
rect 913 70 1153 86
rect 1189 70 1223 86
rect 1259 127 1333 150
rect 1259 93 1279 127
rect 1313 93 1333 127
rect 1259 70 1333 93
rect 1369 120 1419 156
rect 1403 86 1419 120
rect 1369 70 1419 86
rect 1299 17 1333 70
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 683 1440 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 0 617 1440 649
rect 0 17 1440 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -49 1440 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a2bb2o_4
flabel pwell s 0 0 1440 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 1440 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 1440 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 1440 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 127 242 161 276 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 1087 316 1121 350 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 1183 316 1217 350 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 1279 316 1313 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 1375 316 1409 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 A2_N
port 2 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 A1_N
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 1440 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3651272
string GDS_START 3639722
<< end >>
