magic
tech sky130A
magscale 1 2
timestamp 1599588238
<< locali >>
rect 95 196 161 398
rect 263 236 359 310
rect 2137 210 2187 596
rect 2100 70 2187 210
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 21 480 71 596
rect 111 514 177 649
rect 308 514 374 649
rect 414 581 751 615
rect 414 480 464 581
rect 21 446 352 480
rect 498 459 582 547
rect 616 459 683 547
rect 498 446 532 459
rect 21 162 55 446
rect 318 412 532 446
rect 195 378 284 412
rect 195 344 463 378
rect 195 202 229 344
rect 397 252 463 344
rect 21 70 73 162
rect 109 17 159 162
rect 195 70 287 202
rect 323 17 357 202
rect 393 85 459 218
rect 497 185 532 412
rect 566 287 615 421
rect 497 119 547 185
rect 581 85 615 287
rect 393 51 615 85
rect 649 204 683 459
rect 717 451 751 581
rect 790 485 846 649
rect 880 581 1073 615
rect 880 451 914 581
rect 717 417 914 451
rect 948 464 1005 547
rect 1039 498 1073 581
rect 1107 532 1157 649
rect 1295 525 1520 596
rect 1554 530 1588 649
rect 1039 464 1195 498
rect 717 287 751 417
rect 948 383 982 464
rect 811 349 982 383
rect 1016 424 1127 430
rect 1016 390 1087 424
rect 1121 390 1127 424
rect 1016 364 1127 390
rect 1161 377 1195 464
rect 1295 410 1362 525
rect 1486 496 1520 525
rect 1628 496 1694 586
rect 1733 530 1783 649
rect 1823 530 1889 596
rect 811 337 877 349
rect 1161 343 1281 377
rect 961 303 1213 309
rect 785 269 1213 303
rect 785 204 819 269
rect 961 243 1213 269
rect 1247 290 1281 343
rect 1315 360 1362 410
rect 1396 428 1452 471
rect 1486 462 1821 496
rect 1396 394 1465 428
rect 1315 326 1397 360
rect 649 170 819 204
rect 853 206 925 235
rect 1247 224 1329 290
rect 853 172 1002 206
rect 649 83 715 170
rect 813 17 891 136
rect 925 114 1002 172
rect 1124 17 1190 206
rect 1247 85 1281 224
rect 1363 185 1397 326
rect 1315 119 1397 185
rect 1431 85 1465 394
rect 1637 424 1703 428
rect 1637 390 1663 424
rect 1697 390 1703 424
rect 1499 192 1546 311
rect 1637 226 1703 390
rect 1755 274 1821 462
rect 1855 240 1889 530
rect 1818 206 1889 240
rect 1927 310 1993 575
rect 2031 364 2097 649
rect 1927 244 2103 310
rect 1818 192 1852 206
rect 1499 158 1852 192
rect 1927 172 1964 244
rect 1247 51 1465 85
rect 1574 17 1752 120
rect 1786 70 1852 158
rect 1898 70 1964 172
rect 2000 17 2066 206
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 1087 390 1121 424
rect 1663 390 1697 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
<< metal1 >>
rect 0 683 2208 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 0 617 2208 649
rect 1075 424 1133 430
rect 1075 390 1087 424
rect 1121 421 1133 424
rect 1651 424 1709 430
rect 1651 421 1663 424
rect 1121 393 1663 421
rect 1121 390 1133 393
rect 1075 384 1133 390
rect 1651 390 1663 393
rect 1697 390 1709 424
rect 1651 384 1709 390
rect 0 17 2208 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
rect 0 -49 2208 -17
<< labels >>
rlabel locali s 95 196 161 398 6 D
port 1 nsew signal input
rlabel locali s 2137 210 2187 596 6 Q
port 2 nsew signal output
rlabel locali s 2100 70 2187 210 6 Q
port 2 nsew signal output
rlabel metal1 s 1651 421 1709 430 6 SET_B
port 3 nsew signal input
rlabel metal1 s 1651 384 1709 393 6 SET_B
port 3 nsew signal input
rlabel metal1 s 1075 421 1133 430 6 SET_B
port 3 nsew signal input
rlabel metal1 s 1075 393 1709 421 6 SET_B
port 3 nsew signal input
rlabel metal1 s 1075 384 1133 393 6 SET_B
port 3 nsew signal input
rlabel locali s 263 236 359 310 6 CLK
port 4 nsew clock input
rlabel metal1 s 0 -49 2208 49 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 617 2208 715 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2208 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2749860
string GDS_START 2732446
<< end >>
