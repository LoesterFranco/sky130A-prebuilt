magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 336 352 374 493
rect 528 353 566 493
rect 528 352 714 353
rect 25 199 87 323
rect 336 307 714 352
rect 121 199 216 265
rect 658 169 714 307
rect 336 123 714 169
rect 336 103 374 123
rect 528 51 566 123
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 19 376 85 527
rect 131 350 167 493
rect 218 387 284 527
rect 408 387 484 527
rect 600 387 676 527
rect 131 316 292 350
rect 250 271 292 316
rect 250 204 587 271
rect 250 161 292 204
rect 19 123 292 161
rect 19 51 85 123
rect 211 17 277 89
rect 408 17 484 89
rect 600 17 676 89
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel locali s 25 199 87 323 6 A
port 1 nsew signal input
rlabel locali s 121 199 216 265 6 B
port 2 nsew signal input
rlabel locali s 658 169 714 307 6 X
port 3 nsew signal output
rlabel locali s 528 353 566 493 6 X
port 3 nsew signal output
rlabel locali s 528 352 714 353 6 X
port 3 nsew signal output
rlabel locali s 528 51 566 123 6 X
port 3 nsew signal output
rlabel locali s 336 352 374 493 6 X
port 3 nsew signal output
rlabel locali s 336 307 714 352 6 X
port 3 nsew signal output
rlabel locali s 336 123 714 169 6 X
port 3 nsew signal output
rlabel locali s 336 103 374 123 6 X
port 3 nsew signal output
rlabel metal1 s 0 -48 736 48 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 496 736 592 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1495088
string GDS_START 1489050
<< end >>
