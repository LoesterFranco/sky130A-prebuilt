magic
tech sky130A
magscale 1 2
timestamp 1601050088
<< locali >>
rect 85 290 161 356
rect 195 236 257 310
rect 1259 394 1293 596
rect 1259 360 1415 394
rect 1087 236 1157 310
rect 1369 226 1415 360
rect 1230 192 1415 226
rect 1645 364 1717 596
rect 1683 226 1717 364
rect 1230 70 1296 192
rect 1649 70 1717 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 17 506 89 564
rect 130 540 196 649
rect 466 540 539 649
rect 595 581 807 615
rect 17 472 561 506
rect 17 390 89 472
rect 17 226 51 390
rect 237 388 325 438
rect 359 388 441 438
rect 291 334 325 388
rect 291 268 373 334
rect 17 108 89 226
rect 291 202 325 268
rect 407 260 441 388
rect 497 294 561 472
rect 595 296 629 581
rect 663 364 697 547
rect 741 410 807 581
rect 885 530 1013 649
rect 1047 464 1113 596
rect 849 398 1113 464
rect 1147 412 1213 649
rect 1019 378 1113 398
rect 1333 428 1399 649
rect 663 330 985 364
rect 595 260 677 296
rect 407 234 677 260
rect 125 17 191 202
rect 225 150 325 202
rect 359 226 677 234
rect 359 184 441 226
rect 714 192 748 330
rect 921 270 985 330
rect 1019 344 1225 378
rect 1019 226 1053 344
rect 1191 326 1225 344
rect 1191 260 1330 326
rect 636 158 748 192
rect 225 116 596 150
rect 225 70 325 116
rect 562 102 596 116
rect 461 17 528 82
rect 562 51 779 102
rect 846 17 912 212
rect 958 70 1053 226
rect 1122 17 1188 202
rect 1449 326 1511 572
rect 1545 364 1611 649
rect 1751 364 1801 649
rect 1449 260 1649 326
rect 1449 226 1511 260
rect 1330 17 1396 158
rect 1449 90 1515 226
rect 1549 17 1615 226
rect 1751 17 1801 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
<< metal1 >>
rect 0 683 1824 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 0 617 1824 649
rect 0 17 1824 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
rect 0 -49 1824 -17
<< labels >>
rlabel locali s 85 290 161 356 6 D
port 1 nsew signal input
rlabel locali s 1369 226 1415 360 6 Q
port 2 nsew signal output
rlabel locali s 1259 394 1293 596 6 Q
port 2 nsew signal output
rlabel locali s 1259 360 1415 394 6 Q
port 2 nsew signal output
rlabel locali s 1230 192 1415 226 6 Q
port 2 nsew signal output
rlabel locali s 1230 70 1296 192 6 Q
port 2 nsew signal output
rlabel locali s 1683 226 1717 364 6 Q_N
port 3 nsew signal output
rlabel locali s 1649 70 1717 226 6 Q_N
port 3 nsew signal output
rlabel locali s 1645 364 1717 596 6 Q_N
port 3 nsew signal output
rlabel locali s 1087 236 1157 310 6 RESET_B
port 4 nsew signal input
rlabel locali s 195 236 257 310 6 GATE
port 5 nsew clock input
rlabel metal1 s 0 -49 1824 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 1824 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1824 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3048910
string GDS_START 3035568
<< end >>
