magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 1670 704
<< pwell >>
rect 0 0 1632 49
<< scnmos >>
rect 84 74 114 222
rect 208 74 238 222
rect 474 119 504 203
rect 606 125 636 209
rect 701 101 731 185
rect 773 101 803 185
rect 909 75 939 185
rect 1011 98 1041 208
rect 1138 124 1168 208
rect 1221 124 1251 208
rect 1419 74 1449 184
rect 1518 74 1548 222
<< pmoshvt >>
rect 86 368 116 592
rect 176 368 206 592
rect 424 503 454 587
rect 531 463 561 547
rect 638 503 668 587
rect 716 503 746 587
rect 840 424 870 592
rect 981 424 1011 592
rect 1088 508 1118 592
rect 1213 508 1243 592
rect 1415 368 1445 536
rect 1516 368 1546 592
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 131 208 222
rect 114 97 125 131
rect 159 97 208 131
rect 114 74 208 97
rect 238 189 307 222
rect 238 155 261 189
rect 295 155 307 189
rect 238 74 307 155
rect 519 248 591 260
rect 519 214 538 248
rect 572 214 591 248
rect 519 209 591 214
rect 519 203 606 209
rect 401 119 474 203
rect 504 125 606 203
rect 636 185 686 209
rect 954 185 1011 208
rect 636 173 701 185
rect 636 139 648 173
rect 682 139 701 173
rect 636 125 701 139
rect 504 119 554 125
rect 401 112 459 119
rect 401 78 413 112
rect 447 78 459 112
rect 651 101 701 125
rect 731 101 773 185
rect 803 101 909 185
rect 401 66 459 78
rect 818 88 909 101
rect 818 54 830 88
rect 864 75 909 88
rect 939 182 1011 185
rect 939 148 966 182
rect 1000 148 1011 182
rect 939 98 1011 148
rect 1041 180 1138 208
rect 1041 146 1072 180
rect 1106 146 1138 180
rect 1041 124 1138 146
rect 1168 124 1221 208
rect 1251 183 1308 208
rect 1468 184 1518 222
rect 1251 149 1262 183
rect 1296 149 1308 183
rect 1251 124 1308 149
rect 1362 146 1419 184
rect 1041 98 1091 124
rect 939 75 989 98
rect 864 54 876 75
rect 818 42 876 54
rect 1362 112 1374 146
rect 1408 112 1419 146
rect 1362 74 1419 112
rect 1449 120 1518 184
rect 1449 86 1466 120
rect 1500 86 1518 120
rect 1449 74 1518 86
rect 1548 210 1605 222
rect 1548 176 1559 210
rect 1593 176 1605 210
rect 1548 120 1605 176
rect 1548 86 1559 120
rect 1593 86 1605 120
rect 1548 74 1605 86
<< pdiff >>
rect 319 627 378 639
rect 319 593 331 627
rect 365 593 378 627
rect 764 627 822 639
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 510 86 546
rect 27 476 39 510
rect 73 476 86 510
rect 27 440 86 476
rect 27 406 39 440
rect 73 406 86 440
rect 27 368 86 406
rect 116 580 176 592
rect 116 546 129 580
rect 163 546 176 580
rect 116 508 176 546
rect 116 474 129 508
rect 163 474 176 508
rect 116 368 176 474
rect 206 580 265 592
rect 206 546 219 580
rect 253 546 265 580
rect 206 497 265 546
rect 319 587 378 593
rect 764 593 776 627
rect 810 593 822 627
rect 764 592 822 593
rect 764 587 840 592
rect 319 503 424 587
rect 454 547 507 587
rect 585 547 638 587
rect 454 509 531 547
rect 454 503 484 509
rect 206 463 219 497
rect 253 463 265 497
rect 206 414 265 463
rect 206 380 219 414
rect 253 380 265 414
rect 472 475 484 503
rect 518 475 531 509
rect 472 463 531 475
rect 561 509 638 547
rect 561 475 574 509
rect 608 503 638 509
rect 668 503 716 587
rect 746 503 840 587
rect 608 475 620 503
rect 561 463 620 475
rect 206 368 265 380
rect 787 424 840 503
rect 870 475 981 592
rect 870 441 885 475
rect 919 441 981 475
rect 870 424 981 441
rect 1011 513 1088 592
rect 1011 479 1024 513
rect 1058 508 1088 513
rect 1118 508 1213 592
rect 1243 567 1302 592
rect 1243 533 1256 567
rect 1290 533 1302 567
rect 1463 536 1516 592
rect 1243 508 1302 533
rect 1356 524 1415 536
rect 1058 479 1070 508
rect 1011 424 1070 479
rect 1356 490 1368 524
rect 1402 490 1415 524
rect 1356 414 1415 490
rect 1356 380 1368 414
rect 1402 380 1415 414
rect 1356 368 1415 380
rect 1445 524 1516 536
rect 1445 490 1458 524
rect 1492 490 1516 524
rect 1445 444 1516 490
rect 1445 410 1458 444
rect 1492 410 1516 444
rect 1445 368 1516 410
rect 1546 580 1605 592
rect 1546 546 1559 580
rect 1593 546 1605 580
rect 1546 512 1605 546
rect 1546 478 1559 512
rect 1593 478 1605 512
rect 1546 444 1605 478
rect 1546 410 1559 444
rect 1593 410 1605 444
rect 1546 368 1605 410
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 125 97 159 131
rect 261 155 295 189
rect 538 214 572 248
rect 648 139 682 173
rect 413 78 447 112
rect 830 54 864 88
rect 966 148 1000 182
rect 1072 146 1106 180
rect 1262 149 1296 183
rect 1374 112 1408 146
rect 1466 86 1500 120
rect 1559 176 1593 210
rect 1559 86 1593 120
<< pdiffc >>
rect 331 593 365 627
rect 39 546 73 580
rect 39 476 73 510
rect 39 406 73 440
rect 129 546 163 580
rect 129 474 163 508
rect 219 546 253 580
rect 776 593 810 627
rect 219 463 253 497
rect 219 380 253 414
rect 484 475 518 509
rect 574 475 608 509
rect 885 441 919 475
rect 1024 479 1058 513
rect 1256 533 1290 567
rect 1368 490 1402 524
rect 1368 380 1402 414
rect 1458 490 1492 524
rect 1458 410 1492 444
rect 1559 546 1593 580
rect 1559 478 1593 512
rect 1559 410 1593 444
<< poly >>
rect 86 592 116 618
rect 176 592 206 618
rect 424 587 454 613
rect 638 587 668 613
rect 716 587 746 613
rect 840 592 870 618
rect 981 592 1011 618
rect 1088 592 1118 618
rect 1213 592 1243 618
rect 1516 592 1546 618
rect 531 547 561 573
rect 424 488 454 503
rect 421 471 457 488
rect 374 455 457 471
rect 638 488 668 503
rect 716 488 746 503
rect 374 421 390 455
rect 424 421 457 455
rect 531 448 561 463
rect 374 405 457 421
rect 86 353 116 368
rect 176 353 206 368
rect 528 363 564 448
rect 635 416 671 488
rect 713 458 752 488
rect 83 326 119 353
rect 35 310 119 326
rect 173 310 209 353
rect 286 333 564 363
rect 606 400 680 416
rect 606 366 630 400
rect 664 366 680 400
rect 606 350 680 366
rect 286 320 352 333
rect 35 276 51 310
rect 85 276 119 310
rect 35 260 119 276
rect 161 294 238 310
rect 161 260 177 294
rect 211 260 238 294
rect 286 286 302 320
rect 336 286 352 320
rect 286 270 352 286
rect 84 222 114 260
rect 161 244 238 260
rect 208 222 238 244
rect 84 48 114 74
rect 208 48 238 74
rect 322 51 352 270
rect 394 275 460 291
rect 394 241 410 275
rect 444 255 460 275
rect 444 241 504 255
rect 394 225 504 241
rect 474 203 504 225
rect 606 209 636 350
rect 722 283 752 458
rect 1415 536 1445 562
rect 1088 493 1118 508
rect 1213 493 1243 508
rect 1085 476 1121 493
rect 1085 460 1168 476
rect 1085 426 1118 460
rect 1152 426 1168 460
rect 840 409 870 424
rect 981 409 1011 424
rect 1085 410 1168 426
rect 1210 448 1246 493
rect 1210 432 1276 448
rect 837 391 873 409
rect 794 375 873 391
rect 794 341 810 375
rect 844 355 873 375
rect 978 368 1014 409
rect 1210 398 1226 432
rect 1260 398 1276 432
rect 844 341 930 355
rect 794 325 930 341
rect 978 338 1168 368
rect 900 290 930 325
rect 722 267 852 283
rect 722 253 802 267
rect 773 233 802 253
rect 836 233 852 267
rect 900 260 939 290
rect 773 217 852 233
rect 701 185 731 211
rect 773 185 803 217
rect 909 185 939 260
rect 1011 280 1096 296
rect 1011 246 1046 280
rect 1080 246 1096 280
rect 1011 230 1096 246
rect 1011 208 1041 230
rect 1138 208 1168 338
rect 1210 364 1276 398
rect 1210 330 1226 364
rect 1260 330 1276 364
rect 1415 353 1445 368
rect 1516 353 1546 368
rect 1210 314 1276 330
rect 1221 208 1251 314
rect 1412 304 1448 353
rect 1513 336 1549 353
rect 1375 288 1448 304
rect 1375 254 1391 288
rect 1425 268 1448 288
rect 1491 320 1557 336
rect 1491 286 1507 320
rect 1541 286 1557 320
rect 1491 270 1557 286
rect 1425 254 1449 268
rect 1375 238 1449 254
rect 474 93 504 119
rect 606 99 636 125
rect 701 51 731 101
rect 773 75 803 101
rect 322 21 731 51
rect 1419 184 1449 238
rect 1518 222 1548 270
rect 1138 102 1168 124
rect 909 49 939 75
rect 1011 72 1041 98
rect 1113 86 1179 102
rect 1221 98 1251 124
rect 1113 52 1129 86
rect 1163 52 1179 86
rect 1113 36 1179 52
rect 1419 48 1449 74
rect 1518 48 1548 74
<< polycont >>
rect 390 421 424 455
rect 630 366 664 400
rect 51 276 85 310
rect 177 260 211 294
rect 302 286 336 320
rect 410 241 444 275
rect 1118 426 1152 460
rect 810 341 844 375
rect 1226 398 1260 432
rect 802 233 836 267
rect 1046 246 1080 280
rect 1226 330 1260 364
rect 1391 254 1425 288
rect 1507 286 1541 320
rect 1129 52 1163 86
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 23 580 89 596
rect 23 546 39 580
rect 73 546 89 580
rect 23 510 89 546
rect 23 476 39 510
rect 73 476 89 510
rect 23 440 89 476
rect 129 580 163 649
rect 315 627 382 649
rect 129 508 163 546
rect 129 458 163 474
rect 203 580 269 596
rect 315 593 331 627
rect 365 593 382 627
rect 760 627 826 649
rect 760 593 776 627
rect 810 593 826 627
rect 203 546 219 580
rect 253 559 269 580
rect 416 559 692 593
rect 956 581 1168 615
rect 956 559 990 581
rect 253 546 450 559
rect 203 525 450 546
rect 658 525 990 559
rect 203 497 295 525
rect 203 463 219 497
rect 253 463 295 497
rect 484 509 518 525
rect 23 406 39 440
rect 73 424 89 440
rect 73 406 169 424
rect 23 390 169 406
rect 25 310 101 356
rect 25 276 51 310
rect 85 276 101 310
rect 25 260 101 276
rect 135 310 169 390
rect 203 414 295 463
rect 203 380 219 414
rect 253 380 295 414
rect 374 455 450 471
rect 374 421 390 455
rect 424 421 450 455
rect 374 405 450 421
rect 203 364 295 380
rect 261 336 295 364
rect 261 320 352 336
rect 135 294 227 310
rect 135 260 177 294
rect 211 260 227 294
rect 135 226 227 260
rect 23 210 227 226
rect 23 176 39 210
rect 73 192 227 210
rect 23 120 73 176
rect 23 86 39 120
rect 23 70 73 86
rect 109 131 159 158
rect 109 97 125 131
rect 109 17 159 97
rect 193 85 227 192
rect 261 286 302 320
rect 336 286 352 320
rect 261 270 352 286
rect 394 275 450 405
rect 261 189 295 270
rect 394 241 410 275
rect 444 241 450 275
rect 394 225 450 241
rect 484 248 518 475
rect 552 509 624 525
rect 552 475 574 509
rect 608 491 624 509
rect 608 475 828 491
rect 552 457 828 475
rect 552 316 586 457
rect 620 400 752 416
rect 620 366 630 400
rect 664 366 752 400
rect 620 350 752 366
rect 552 282 684 316
rect 484 214 538 248
rect 572 214 595 248
rect 261 119 295 155
rect 329 146 531 180
rect 329 85 363 146
rect 193 51 363 85
rect 397 78 413 112
rect 447 78 463 112
rect 397 17 463 78
rect 497 89 531 146
rect 631 173 684 282
rect 631 139 648 173
rect 682 139 684 173
rect 631 123 684 139
rect 718 172 752 350
rect 794 391 828 457
rect 867 475 922 491
rect 867 441 885 475
rect 919 441 922 475
rect 867 425 922 441
rect 794 375 854 391
rect 794 341 810 375
rect 844 341 854 375
rect 794 325 854 341
rect 786 267 852 283
rect 786 233 802 267
rect 836 240 852 267
rect 888 240 922 425
rect 956 308 990 525
rect 1024 513 1058 547
rect 1024 376 1058 479
rect 1102 460 1168 581
rect 1240 567 1306 649
rect 1240 533 1256 567
rect 1290 533 1306 567
rect 1240 504 1306 533
rect 1352 524 1402 540
rect 1102 426 1118 460
rect 1152 426 1168 460
rect 1352 490 1368 524
rect 1102 410 1168 426
rect 1210 432 1276 448
rect 1210 398 1226 432
rect 1260 398 1276 432
rect 1024 342 1164 376
rect 956 280 1096 308
rect 956 274 1046 280
rect 1034 246 1046 274
rect 1080 246 1096 280
rect 836 233 1000 240
rect 786 206 1000 233
rect 1034 230 1096 246
rect 1130 280 1164 342
rect 1210 372 1276 398
rect 1352 414 1402 490
rect 1352 380 1368 414
rect 1442 524 1508 649
rect 1442 490 1458 524
rect 1492 490 1508 524
rect 1442 444 1508 490
rect 1442 410 1458 444
rect 1492 410 1508 444
rect 1442 406 1508 410
rect 1543 580 1615 596
rect 1543 546 1559 580
rect 1593 546 1615 580
rect 1543 512 1615 546
rect 1543 478 1559 512
rect 1593 478 1615 512
rect 1543 444 1615 478
rect 1543 410 1559 444
rect 1593 410 1615 444
rect 1543 406 1615 410
rect 1352 372 1402 380
rect 1210 364 1547 372
rect 1210 330 1226 364
rect 1260 338 1547 364
rect 1260 330 1276 338
rect 1210 314 1276 330
rect 1475 320 1547 338
rect 1375 288 1441 304
rect 1375 280 1391 288
rect 1130 254 1391 280
rect 1425 254 1441 288
rect 1130 246 1441 254
rect 966 182 1000 206
rect 1130 196 1164 246
rect 1375 238 1441 246
rect 1475 286 1507 320
rect 1541 286 1547 320
rect 1475 270 1547 286
rect 718 138 932 172
rect 718 89 752 138
rect 497 55 752 89
rect 814 88 864 104
rect 814 54 830 88
rect 814 17 864 54
rect 898 85 932 138
rect 966 119 1000 148
rect 1044 180 1164 196
rect 1044 146 1072 180
rect 1106 146 1164 180
rect 1246 183 1312 212
rect 1475 204 1509 270
rect 1581 226 1615 406
rect 1246 149 1262 183
rect 1296 149 1312 183
rect 1113 86 1179 102
rect 1113 85 1129 86
rect 898 52 1129 85
rect 1163 52 1179 86
rect 898 51 1179 52
rect 1246 17 1312 149
rect 1358 170 1509 204
rect 1543 210 1615 226
rect 1543 176 1559 210
rect 1593 176 1615 210
rect 1358 146 1408 170
rect 1358 112 1374 146
rect 1358 70 1408 112
rect 1444 120 1507 136
rect 1444 86 1466 120
rect 1500 86 1507 120
rect 1444 17 1507 86
rect 1543 120 1615 176
rect 1543 86 1559 120
rect 1593 86 1615 120
rect 1543 70 1615 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dfxtp_1
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 1567 94 1601 128 0 FreeSans 340 0 0 0 Q
port 7 nsew
flabel corelocali s 1567 168 1601 202 0 FreeSans 340 0 0 0 Q
port 7 nsew
flabel corelocali s 415 390 449 424 0 FreeSans 340 0 0 0 D
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 1632 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2664938
string GDS_START 2652306
<< end >>
