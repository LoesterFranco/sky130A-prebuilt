magic
tech sky130A
magscale 1 2
timestamp 1601050082
<< locali >>
rect 25 258 110 392
rect 159 326 260 430
rect 1442 364 1513 596
rect 1067 236 1133 310
rect 1479 226 1513 364
rect 1459 70 1525 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 21 426 87 649
rect 189 498 255 596
rect 297 532 363 649
rect 510 498 560 551
rect 189 464 560 498
rect 294 278 328 464
rect 144 244 328 278
rect 362 343 468 430
rect 510 377 560 464
rect 600 447 672 539
rect 362 309 604 343
rect 144 224 178 244
rect 23 17 73 224
rect 109 142 178 224
rect 362 210 396 309
rect 538 277 604 309
rect 638 283 672 447
rect 798 419 848 649
rect 888 478 965 584
rect 1102 512 1168 649
rect 888 444 1201 478
rect 888 385 965 444
rect 706 351 965 385
rect 706 317 772 351
rect 831 283 897 317
rect 313 176 396 210
rect 430 240 496 272
rect 638 249 897 283
rect 430 206 543 240
rect 109 108 475 142
rect 211 17 277 74
rect 425 70 475 108
rect 509 85 543 206
rect 638 169 672 249
rect 931 215 965 351
rect 577 119 672 169
rect 706 181 876 215
rect 706 85 740 181
rect 509 51 740 85
rect 774 17 808 147
rect 842 85 876 181
rect 910 119 965 215
rect 999 344 1062 410
rect 999 202 1033 344
rect 1167 326 1201 444
rect 1235 394 1301 578
rect 1342 428 1408 649
rect 1235 360 1408 394
rect 1548 364 1598 649
rect 1374 326 1408 360
rect 1167 260 1306 326
rect 1374 260 1445 326
rect 1374 226 1408 260
rect 999 85 1072 202
rect 842 51 1072 85
rect 1106 17 1172 202
rect 1265 192 1408 226
rect 1265 70 1331 192
rect 1373 17 1423 158
rect 1561 17 1611 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
rlabel locali s 159 326 260 430 6 GATE
port 1 nsew signal input
rlabel locali s 1479 226 1513 364 6 GCLK
port 2 nsew signal output
rlabel locali s 1459 70 1525 226 6 GCLK
port 2 nsew signal output
rlabel locali s 1442 364 1513 596 6 GCLK
port 2 nsew signal output
rlabel locali s 25 258 110 392 6 SCE
port 3 nsew signal input
rlabel locali s 1067 236 1133 310 6 CLK
port 4 nsew clock input
rlabel metal1 s 0 -49 1632 49 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1632 715 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 433364
string GDS_START 420868
<< end >>
