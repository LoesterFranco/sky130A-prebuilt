magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 130 517 467 524
rect 25 490 467 517
rect 25 483 164 490
rect 25 326 71 483
rect 25 260 96 326
rect 275 289 359 356
rect 433 336 467 490
rect 601 446 658 596
rect 893 446 939 547
rect 601 412 939 446
rect 393 270 467 336
rect 601 226 658 412
rect 739 356 1019 378
rect 739 344 1099 356
rect 739 270 805 344
rect 869 236 935 310
rect 985 270 1099 344
rect 600 119 658 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 23 551 89 649
rect 237 558 303 649
rect 344 449 399 456
rect 130 390 399 449
rect 130 255 196 390
rect 501 364 567 649
rect 692 480 758 649
rect 793 581 1039 615
rect 793 480 859 581
rect 973 412 1039 581
rect 501 260 567 326
rect 130 236 281 255
rect 501 236 535 260
rect 130 221 535 236
rect 1079 390 1129 649
rect 29 17 95 206
rect 231 202 535 221
rect 129 85 195 187
rect 231 121 281 202
rect 316 85 382 165
rect 129 51 382 85
rect 416 17 468 165
rect 514 85 564 165
rect 692 202 758 226
rect 1063 202 1129 226
rect 692 168 1129 202
rect 692 85 758 168
rect 894 154 1129 168
rect 514 51 758 85
rect 792 17 858 134
rect 894 70 938 154
rect 974 17 1043 120
rect 1079 70 1129 154
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
rlabel locali s 433 336 467 490 6 A1_N
port 1 nsew signal input
rlabel locali s 393 270 467 336 6 A1_N
port 1 nsew signal input
rlabel locali s 130 517 467 524 6 A1_N
port 1 nsew signal input
rlabel locali s 25 490 467 517 6 A1_N
port 1 nsew signal input
rlabel locali s 25 483 164 490 6 A1_N
port 1 nsew signal input
rlabel locali s 25 326 71 483 6 A1_N
port 1 nsew signal input
rlabel locali s 25 260 96 326 6 A1_N
port 1 nsew signal input
rlabel locali s 275 289 359 356 6 A2_N
port 2 nsew signal input
rlabel locali s 985 270 1099 344 6 B1
port 3 nsew signal input
rlabel locali s 739 356 1019 378 6 B1
port 3 nsew signal input
rlabel locali s 739 344 1099 356 6 B1
port 3 nsew signal input
rlabel locali s 739 270 805 344 6 B1
port 3 nsew signal input
rlabel locali s 869 236 935 310 6 B2
port 4 nsew signal input
rlabel locali s 893 446 939 547 6 Y
port 5 nsew signal output
rlabel locali s 601 446 658 596 6 Y
port 5 nsew signal output
rlabel locali s 601 412 939 446 6 Y
port 5 nsew signal output
rlabel locali s 601 226 658 412 6 Y
port 5 nsew signal output
rlabel locali s 600 119 658 226 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -49 1152 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 1152 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1283472
string GDS_START 1273612
<< end >>
