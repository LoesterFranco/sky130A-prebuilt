magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 301 333 377 493
rect 489 333 568 493
rect 680 333 756 493
rect 868 333 944 493
rect 301 289 944 333
rect 22 215 88 255
rect 515 181 568 289
rect 681 215 1078 255
rect 301 127 568 181
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 18 333 85 493
rect 129 367 267 527
rect 18 289 166 333
rect 204 289 267 367
rect 421 367 455 527
rect 612 367 646 527
rect 800 367 834 527
rect 994 299 1060 527
rect 132 255 166 289
rect 132 215 471 255
rect 132 181 166 215
rect 18 143 166 181
rect 18 51 85 143
rect 129 17 168 109
rect 217 93 267 181
rect 612 143 1060 181
rect 612 93 662 143
rect 217 51 662 93
rect 706 17 740 109
rect 774 51 850 143
rect 894 17 942 109
rect 994 51 1060 143
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
rlabel locali s 22 215 88 255 6 A_N
port 1 nsew signal input
rlabel locali s 681 215 1078 255 6 B
port 2 nsew signal input
rlabel locali s 868 333 944 493 6 Y
port 3 nsew signal output
rlabel locali s 680 333 756 493 6 Y
port 3 nsew signal output
rlabel locali s 515 181 568 289 6 Y
port 3 nsew signal output
rlabel locali s 489 333 568 493 6 Y
port 3 nsew signal output
rlabel locali s 301 333 377 493 6 Y
port 3 nsew signal output
rlabel locali s 301 289 944 333 6 Y
port 3 nsew signal output
rlabel locali s 301 127 568 181 6 Y
port 3 nsew signal output
rlabel metal1 s 0 -48 1104 48 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 496 1104 592 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1104 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2238036
string GDS_START 2228660
<< end >>
