magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 828 561
rect 27 324 78 492
rect 113 363 179 527
rect 27 51 93 324
rect 303 258 344 493
rect 258 210 344 258
rect 378 210 444 493
rect 480 199 536 493
rect 665 367 708 527
rect 581 199 658 265
rect 702 205 802 258
rect 597 169 658 199
rect 127 17 262 94
rect 417 17 486 97
rect 597 57 708 169
rect 743 17 791 152
rect 0 -17 828 17
<< obsli1 >>
rect 227 329 269 492
rect 139 293 269 329
rect 139 165 183 293
rect 572 333 629 492
rect 744 333 798 492
rect 572 299 798 333
rect 139 131 561 165
rect 139 130 383 131
rect 317 52 383 130
rect 520 52 561 131
<< metal1 >>
rect 0 496 828 592
rect 0 -48 828 48
<< labels >>
rlabel locali s 597 169 658 199 6 A1
port 1 nsew signal input
rlabel locali s 597 57 708 169 6 A1
port 1 nsew signal input
rlabel locali s 581 199 658 265 6 A1
port 1 nsew signal input
rlabel locali s 702 205 802 258 6 A2
port 2 nsew signal input
rlabel locali s 480 199 536 493 6 B1
port 3 nsew signal input
rlabel locali s 378 210 444 493 6 C1
port 4 nsew signal input
rlabel locali s 303 258 344 493 6 D1
port 5 nsew signal input
rlabel locali s 258 210 344 258 6 D1
port 5 nsew signal input
rlabel locali s 27 324 78 492 6 X
port 6 nsew signal output
rlabel locali s 27 51 93 324 6 X
port 6 nsew signal output
rlabel locali s 743 17 791 152 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 417 17 486 97 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 127 17 262 94 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 828 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 828 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 665 367 708 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 113 363 179 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 828 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 828 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3867694
string GDS_START 3859002
<< end >>
