magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 368 561
rect 114 447 198 527
rect 232 425 351 493
rect 17 199 130 345
rect 232 119 266 425
rect 300 153 351 391
rect 106 17 198 97
rect 232 51 351 119
rect 0 -17 368 17
<< obsli1 >>
rect 17 413 80 493
rect 17 379 198 413
rect 164 165 198 379
rect 17 131 198 165
rect 17 51 72 131
<< metal1 >>
rect 0 496 368 592
rect 0 -48 368 48
<< labels >>
rlabel locali s 300 153 351 391 6 A
port 1 nsew signal input
rlabel locali s 17 199 130 345 6 TE_B
port 2 nsew signal input
rlabel locali s 232 425 351 493 6 Z
port 3 nsew signal output
rlabel locali s 232 119 266 425 6 Z
port 3 nsew signal output
rlabel locali s 232 51 351 119 6 Z
port 3 nsew signal output
rlabel locali s 106 17 198 97 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 368 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 368 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 114 447 198 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 368 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 368 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 368 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2888674
string GDS_START 2884432
<< end >>
