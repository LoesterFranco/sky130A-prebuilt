magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 10434 827
<< pwell >>
rect 29 1071 63 1105
rect 2513 1071 2547 1105
rect 2605 1071 2639 1105
rect 5089 1071 5123 1105
rect 5273 1071 5307 1105
rect 7757 1071 7791 1105
rect 7849 1071 7883 1105
rect 10333 1071 10367 1105
rect 29 -17 63 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 5089 -17 5123 17
rect 5273 -17 5307 17
rect 7757 -17 7791 17
rect 7849 -17 7883 17
rect 10333 -17 10367 17
<< scnmos >>
rect 89 911 119 1041
rect 173 911 203 1041
rect 277 911 307 1041
rect 361 911 391 1041
rect 549 918 579 1022
rect 633 918 663 1022
rect 717 918 747 1022
rect 801 918 831 1022
rect 1060 957 1090 1041
rect 1144 957 1174 1041
rect 1402 957 1432 1041
rect 1486 957 1516 1041
rect 1745 918 1775 1022
rect 1829 918 1859 1022
rect 1913 918 1943 1022
rect 1997 918 2027 1022
rect 2185 911 2215 1041
rect 2269 911 2299 1041
rect 2373 911 2403 1041
rect 2457 911 2487 1041
rect 2665 911 2695 1041
rect 2749 911 2779 1041
rect 2853 911 2883 1041
rect 2937 911 2967 1041
rect 3125 918 3155 1022
rect 3209 918 3239 1022
rect 3293 918 3323 1022
rect 3377 918 3407 1022
rect 3636 957 3666 1041
rect 3720 957 3750 1041
rect 3978 957 4008 1041
rect 4062 957 4092 1041
rect 4321 918 4351 1022
rect 4405 918 4435 1022
rect 4489 918 4519 1022
rect 4573 918 4603 1022
rect 4761 911 4791 1041
rect 4845 911 4875 1041
rect 4949 911 4979 1041
rect 5033 911 5063 1041
rect 5333 911 5363 1041
rect 5417 911 5447 1041
rect 5521 911 5551 1041
rect 5605 911 5635 1041
rect 5793 918 5823 1022
rect 5877 918 5907 1022
rect 5961 918 5991 1022
rect 6045 918 6075 1022
rect 6304 957 6334 1041
rect 6388 957 6418 1041
rect 6646 957 6676 1041
rect 6730 957 6760 1041
rect 6989 918 7019 1022
rect 7073 918 7103 1022
rect 7157 918 7187 1022
rect 7241 918 7271 1022
rect 7429 911 7459 1041
rect 7513 911 7543 1041
rect 7617 911 7647 1041
rect 7701 911 7731 1041
rect 7909 911 7939 1041
rect 7993 911 8023 1041
rect 8097 911 8127 1041
rect 8181 911 8211 1041
rect 8369 918 8399 1022
rect 8453 918 8483 1022
rect 8537 918 8567 1022
rect 8621 918 8651 1022
rect 8880 957 8910 1041
rect 8964 957 8994 1041
rect 9222 957 9252 1041
rect 9306 957 9336 1041
rect 9565 918 9595 1022
rect 9649 918 9679 1022
rect 9733 918 9763 1022
rect 9817 918 9847 1022
rect 10005 911 10035 1041
rect 10089 911 10119 1041
rect 10193 911 10223 1041
rect 10277 911 10307 1041
rect 89 47 119 177
rect 173 47 203 177
rect 277 47 307 177
rect 361 47 391 177
rect 549 66 579 170
rect 633 66 663 170
rect 717 66 747 170
rect 801 66 831 170
rect 1060 47 1090 131
rect 1144 47 1174 131
rect 1402 47 1432 131
rect 1486 47 1516 131
rect 1745 66 1775 170
rect 1829 66 1859 170
rect 1913 66 1943 170
rect 1997 66 2027 170
rect 2185 47 2215 177
rect 2269 47 2299 177
rect 2373 47 2403 177
rect 2457 47 2487 177
rect 2665 47 2695 177
rect 2749 47 2779 177
rect 2853 47 2883 177
rect 2937 47 2967 177
rect 3125 66 3155 170
rect 3209 66 3239 170
rect 3293 66 3323 170
rect 3377 66 3407 170
rect 3636 47 3666 131
rect 3720 47 3750 131
rect 3978 47 4008 131
rect 4062 47 4092 131
rect 4321 66 4351 170
rect 4405 66 4435 170
rect 4489 66 4519 170
rect 4573 66 4603 170
rect 4761 47 4791 177
rect 4845 47 4875 177
rect 4949 47 4979 177
rect 5033 47 5063 177
rect 5333 47 5363 177
rect 5417 47 5447 177
rect 5521 47 5551 177
rect 5605 47 5635 177
rect 5793 66 5823 170
rect 5877 66 5907 170
rect 5961 66 5991 170
rect 6045 66 6075 170
rect 6304 47 6334 131
rect 6388 47 6418 131
rect 6646 47 6676 131
rect 6730 47 6760 131
rect 6989 66 7019 170
rect 7073 66 7103 170
rect 7157 66 7187 170
rect 7241 66 7271 170
rect 7429 47 7459 177
rect 7513 47 7543 177
rect 7617 47 7647 177
rect 7701 47 7731 177
rect 7909 47 7939 177
rect 7993 47 8023 177
rect 8097 47 8127 177
rect 8181 47 8211 177
rect 8369 66 8399 170
rect 8453 66 8483 170
rect 8537 66 8567 170
rect 8621 66 8651 170
rect 8880 47 8910 131
rect 8964 47 8994 131
rect 9222 47 9252 131
rect 9306 47 9336 131
rect 9565 66 9595 170
rect 9649 66 9679 170
rect 9733 66 9763 170
rect 9817 66 9847 170
rect 10005 47 10035 177
rect 10089 47 10119 177
rect 10193 47 10223 177
rect 10277 47 10307 177
<< pmoshvt >>
rect 81 591 117 791
rect 175 591 211 791
rect 269 591 305 791
rect 363 591 399 791
rect 561 613 597 777
rect 655 613 691 777
rect 749 613 785 777
rect 843 613 879 777
rect 1052 599 1088 763
rect 1146 599 1182 763
rect 1394 599 1430 763
rect 1488 599 1524 763
rect 1697 613 1733 777
rect 1791 613 1827 777
rect 1885 613 1921 777
rect 1979 613 2015 777
rect 2177 591 2213 791
rect 2271 591 2307 791
rect 2365 591 2401 791
rect 2459 591 2495 791
rect 2657 591 2693 791
rect 2751 591 2787 791
rect 2845 591 2881 791
rect 2939 591 2975 791
rect 3137 613 3173 777
rect 3231 613 3267 777
rect 3325 613 3361 777
rect 3419 613 3455 777
rect 3628 599 3664 763
rect 3722 599 3758 763
rect 3970 599 4006 763
rect 4064 599 4100 763
rect 4273 613 4309 777
rect 4367 613 4403 777
rect 4461 613 4497 777
rect 4555 613 4591 777
rect 4753 591 4789 791
rect 4847 591 4883 791
rect 4941 591 4977 791
rect 5035 591 5071 791
rect 5325 591 5361 791
rect 5419 591 5455 791
rect 5513 591 5549 791
rect 5607 591 5643 791
rect 5805 613 5841 777
rect 5899 613 5935 777
rect 5993 613 6029 777
rect 6087 613 6123 777
rect 6296 599 6332 763
rect 6390 599 6426 763
rect 6638 599 6674 763
rect 6732 599 6768 763
rect 6941 613 6977 777
rect 7035 613 7071 777
rect 7129 613 7165 777
rect 7223 613 7259 777
rect 7421 591 7457 791
rect 7515 591 7551 791
rect 7609 591 7645 791
rect 7703 591 7739 791
rect 7901 591 7937 791
rect 7995 591 8031 791
rect 8089 591 8125 791
rect 8183 591 8219 791
rect 8381 613 8417 777
rect 8475 613 8511 777
rect 8569 613 8605 777
rect 8663 613 8699 777
rect 8872 599 8908 763
rect 8966 599 9002 763
rect 9214 599 9250 763
rect 9308 599 9344 763
rect 9517 613 9553 777
rect 9611 613 9647 777
rect 9705 613 9741 777
rect 9799 613 9835 777
rect 9997 591 10033 791
rect 10091 591 10127 791
rect 10185 591 10221 791
rect 10279 591 10315 791
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 561 311 597 475
rect 655 311 691 475
rect 749 311 785 475
rect 843 311 879 475
rect 1052 325 1088 489
rect 1146 325 1182 489
rect 1394 325 1430 489
rect 1488 325 1524 489
rect 1697 311 1733 475
rect 1791 311 1827 475
rect 1885 311 1921 475
rect 1979 311 2015 475
rect 2177 297 2213 497
rect 2271 297 2307 497
rect 2365 297 2401 497
rect 2459 297 2495 497
rect 2657 297 2693 497
rect 2751 297 2787 497
rect 2845 297 2881 497
rect 2939 297 2975 497
rect 3137 311 3173 475
rect 3231 311 3267 475
rect 3325 311 3361 475
rect 3419 311 3455 475
rect 3628 325 3664 489
rect 3722 325 3758 489
rect 3970 325 4006 489
rect 4064 325 4100 489
rect 4273 311 4309 475
rect 4367 311 4403 475
rect 4461 311 4497 475
rect 4555 311 4591 475
rect 4753 297 4789 497
rect 4847 297 4883 497
rect 4941 297 4977 497
rect 5035 297 5071 497
rect 5325 297 5361 497
rect 5419 297 5455 497
rect 5513 297 5549 497
rect 5607 297 5643 497
rect 5805 311 5841 475
rect 5899 311 5935 475
rect 5993 311 6029 475
rect 6087 311 6123 475
rect 6296 325 6332 489
rect 6390 325 6426 489
rect 6638 325 6674 489
rect 6732 325 6768 489
rect 6941 311 6977 475
rect 7035 311 7071 475
rect 7129 311 7165 475
rect 7223 311 7259 475
rect 7421 297 7457 497
rect 7515 297 7551 497
rect 7609 297 7645 497
rect 7703 297 7739 497
rect 7901 297 7937 497
rect 7995 297 8031 497
rect 8089 297 8125 497
rect 8183 297 8219 497
rect 8381 311 8417 475
rect 8475 311 8511 475
rect 8569 311 8605 475
rect 8663 311 8699 475
rect 8872 325 8908 489
rect 8966 325 9002 489
rect 9214 325 9250 489
rect 9308 325 9344 489
rect 9517 311 9553 475
rect 9611 311 9647 475
rect 9705 311 9741 475
rect 9799 311 9835 475
rect 9997 297 10033 497
rect 10091 297 10127 497
rect 10185 297 10221 497
rect 10279 297 10315 497
<< ndiff >>
rect 27 1029 89 1041
rect 27 995 45 1029
rect 79 995 89 1029
rect 27 961 89 995
rect 27 927 45 961
rect 79 927 89 961
rect 27 911 89 927
rect 119 1029 173 1041
rect 119 995 129 1029
rect 163 995 173 1029
rect 119 961 173 995
rect 119 927 129 961
rect 163 927 173 961
rect 119 911 173 927
rect 203 1029 277 1041
rect 203 995 223 1029
rect 257 995 277 1029
rect 203 911 277 995
rect 307 1029 361 1041
rect 307 995 317 1029
rect 351 995 361 1029
rect 307 961 361 995
rect 307 927 317 961
rect 351 927 361 961
rect 307 911 361 927
rect 391 1029 443 1041
rect 391 995 401 1029
rect 435 995 443 1029
rect 391 911 443 995
rect 497 987 549 1022
rect 497 953 505 987
rect 539 953 549 987
rect 497 918 549 953
rect 579 969 633 1022
rect 579 935 589 969
rect 623 935 633 969
rect 579 918 633 935
rect 663 987 717 1022
rect 663 953 673 987
rect 707 953 717 987
rect 663 918 717 953
rect 747 969 801 1022
rect 747 935 757 969
rect 791 935 801 969
rect 747 918 801 935
rect 831 987 883 1022
rect 831 953 841 987
rect 875 953 883 987
rect 831 918 883 953
rect 1008 1016 1060 1041
rect 1008 982 1016 1016
rect 1050 982 1060 1016
rect 1008 957 1060 982
rect 1090 1016 1144 1041
rect 1090 982 1100 1016
rect 1134 982 1144 1016
rect 1090 957 1144 982
rect 1174 1016 1226 1041
rect 1174 982 1184 1016
rect 1218 982 1226 1016
rect 1174 957 1226 982
rect 1350 1016 1402 1041
rect 1350 982 1358 1016
rect 1392 982 1402 1016
rect 1350 957 1402 982
rect 1432 1016 1486 1041
rect 1432 982 1442 1016
rect 1476 982 1486 1016
rect 1432 957 1486 982
rect 1516 1016 1568 1041
rect 1516 982 1526 1016
rect 1560 982 1568 1016
rect 1516 957 1568 982
rect 2133 1029 2185 1041
rect 1693 987 1745 1022
rect 1693 953 1701 987
rect 1735 953 1745 987
rect 1693 918 1745 953
rect 1775 969 1829 1022
rect 1775 935 1785 969
rect 1819 935 1829 969
rect 1775 918 1829 935
rect 1859 987 1913 1022
rect 1859 953 1869 987
rect 1903 953 1913 987
rect 1859 918 1913 953
rect 1943 969 1997 1022
rect 1943 935 1953 969
rect 1987 935 1997 969
rect 1943 918 1997 935
rect 2027 987 2079 1022
rect 2027 953 2037 987
rect 2071 953 2079 987
rect 2027 918 2079 953
rect 2133 995 2141 1029
rect 2175 995 2185 1029
rect 2133 911 2185 995
rect 2215 1029 2269 1041
rect 2215 995 2225 1029
rect 2259 995 2269 1029
rect 2215 961 2269 995
rect 2215 927 2225 961
rect 2259 927 2269 961
rect 2215 911 2269 927
rect 2299 1029 2373 1041
rect 2299 995 2319 1029
rect 2353 995 2373 1029
rect 2299 911 2373 995
rect 2403 1029 2457 1041
rect 2403 995 2413 1029
rect 2447 995 2457 1029
rect 2403 961 2457 995
rect 2403 927 2413 961
rect 2447 927 2457 961
rect 2403 911 2457 927
rect 2487 1029 2549 1041
rect 2487 995 2497 1029
rect 2531 995 2549 1029
rect 2487 961 2549 995
rect 2487 927 2497 961
rect 2531 927 2549 961
rect 2487 911 2549 927
rect 2603 1029 2665 1041
rect 2603 995 2621 1029
rect 2655 995 2665 1029
rect 2603 961 2665 995
rect 2603 927 2621 961
rect 2655 927 2665 961
rect 2603 911 2665 927
rect 2695 1029 2749 1041
rect 2695 995 2705 1029
rect 2739 995 2749 1029
rect 2695 961 2749 995
rect 2695 927 2705 961
rect 2739 927 2749 961
rect 2695 911 2749 927
rect 2779 1029 2853 1041
rect 2779 995 2799 1029
rect 2833 995 2853 1029
rect 2779 911 2853 995
rect 2883 1029 2937 1041
rect 2883 995 2893 1029
rect 2927 995 2937 1029
rect 2883 961 2937 995
rect 2883 927 2893 961
rect 2927 927 2937 961
rect 2883 911 2937 927
rect 2967 1029 3019 1041
rect 2967 995 2977 1029
rect 3011 995 3019 1029
rect 2967 911 3019 995
rect 3073 987 3125 1022
rect 3073 953 3081 987
rect 3115 953 3125 987
rect 3073 918 3125 953
rect 3155 969 3209 1022
rect 3155 935 3165 969
rect 3199 935 3209 969
rect 3155 918 3209 935
rect 3239 987 3293 1022
rect 3239 953 3249 987
rect 3283 953 3293 987
rect 3239 918 3293 953
rect 3323 969 3377 1022
rect 3323 935 3333 969
rect 3367 935 3377 969
rect 3323 918 3377 935
rect 3407 987 3459 1022
rect 3407 953 3417 987
rect 3451 953 3459 987
rect 3407 918 3459 953
rect 3584 1016 3636 1041
rect 3584 982 3592 1016
rect 3626 982 3636 1016
rect 3584 957 3636 982
rect 3666 1016 3720 1041
rect 3666 982 3676 1016
rect 3710 982 3720 1016
rect 3666 957 3720 982
rect 3750 1016 3802 1041
rect 3750 982 3760 1016
rect 3794 982 3802 1016
rect 3750 957 3802 982
rect 3926 1016 3978 1041
rect 3926 982 3934 1016
rect 3968 982 3978 1016
rect 3926 957 3978 982
rect 4008 1016 4062 1041
rect 4008 982 4018 1016
rect 4052 982 4062 1016
rect 4008 957 4062 982
rect 4092 1016 4144 1041
rect 4092 982 4102 1016
rect 4136 982 4144 1016
rect 4092 957 4144 982
rect 4709 1029 4761 1041
rect 4269 987 4321 1022
rect 4269 953 4277 987
rect 4311 953 4321 987
rect 4269 918 4321 953
rect 4351 969 4405 1022
rect 4351 935 4361 969
rect 4395 935 4405 969
rect 4351 918 4405 935
rect 4435 987 4489 1022
rect 4435 953 4445 987
rect 4479 953 4489 987
rect 4435 918 4489 953
rect 4519 969 4573 1022
rect 4519 935 4529 969
rect 4563 935 4573 969
rect 4519 918 4573 935
rect 4603 987 4655 1022
rect 4603 953 4613 987
rect 4647 953 4655 987
rect 4603 918 4655 953
rect 4709 995 4717 1029
rect 4751 995 4761 1029
rect 4709 911 4761 995
rect 4791 1029 4845 1041
rect 4791 995 4801 1029
rect 4835 995 4845 1029
rect 4791 961 4845 995
rect 4791 927 4801 961
rect 4835 927 4845 961
rect 4791 911 4845 927
rect 4875 1029 4949 1041
rect 4875 995 4895 1029
rect 4929 995 4949 1029
rect 4875 911 4949 995
rect 4979 1029 5033 1041
rect 4979 995 4989 1029
rect 5023 995 5033 1029
rect 4979 961 5033 995
rect 4979 927 4989 961
rect 5023 927 5033 961
rect 4979 911 5033 927
rect 5063 1029 5125 1041
rect 5063 995 5073 1029
rect 5107 995 5125 1029
rect 5271 1029 5333 1041
rect 5063 961 5125 995
rect 5063 927 5073 961
rect 5107 927 5125 961
rect 5063 911 5125 927
rect 5271 995 5289 1029
rect 5323 995 5333 1029
rect 5271 961 5333 995
rect 5271 927 5289 961
rect 5323 927 5333 961
rect 5271 911 5333 927
rect 5363 1029 5417 1041
rect 5363 995 5373 1029
rect 5407 995 5417 1029
rect 5363 961 5417 995
rect 5363 927 5373 961
rect 5407 927 5417 961
rect 5363 911 5417 927
rect 5447 1029 5521 1041
rect 5447 995 5467 1029
rect 5501 995 5521 1029
rect 5447 911 5521 995
rect 5551 1029 5605 1041
rect 5551 995 5561 1029
rect 5595 995 5605 1029
rect 5551 961 5605 995
rect 5551 927 5561 961
rect 5595 927 5605 961
rect 5551 911 5605 927
rect 5635 1029 5687 1041
rect 5635 995 5645 1029
rect 5679 995 5687 1029
rect 5635 911 5687 995
rect 5741 987 5793 1022
rect 5741 953 5749 987
rect 5783 953 5793 987
rect 5741 918 5793 953
rect 5823 969 5877 1022
rect 5823 935 5833 969
rect 5867 935 5877 969
rect 5823 918 5877 935
rect 5907 987 5961 1022
rect 5907 953 5917 987
rect 5951 953 5961 987
rect 5907 918 5961 953
rect 5991 969 6045 1022
rect 5991 935 6001 969
rect 6035 935 6045 969
rect 5991 918 6045 935
rect 6075 987 6127 1022
rect 6075 953 6085 987
rect 6119 953 6127 987
rect 6075 918 6127 953
rect 6252 1016 6304 1041
rect 6252 982 6260 1016
rect 6294 982 6304 1016
rect 6252 957 6304 982
rect 6334 1016 6388 1041
rect 6334 982 6344 1016
rect 6378 982 6388 1016
rect 6334 957 6388 982
rect 6418 1016 6470 1041
rect 6418 982 6428 1016
rect 6462 982 6470 1016
rect 6418 957 6470 982
rect 6594 1016 6646 1041
rect 6594 982 6602 1016
rect 6636 982 6646 1016
rect 6594 957 6646 982
rect 6676 1016 6730 1041
rect 6676 982 6686 1016
rect 6720 982 6730 1016
rect 6676 957 6730 982
rect 6760 1016 6812 1041
rect 6760 982 6770 1016
rect 6804 982 6812 1016
rect 6760 957 6812 982
rect 7377 1029 7429 1041
rect 6937 987 6989 1022
rect 6937 953 6945 987
rect 6979 953 6989 987
rect 6937 918 6989 953
rect 7019 969 7073 1022
rect 7019 935 7029 969
rect 7063 935 7073 969
rect 7019 918 7073 935
rect 7103 987 7157 1022
rect 7103 953 7113 987
rect 7147 953 7157 987
rect 7103 918 7157 953
rect 7187 969 7241 1022
rect 7187 935 7197 969
rect 7231 935 7241 969
rect 7187 918 7241 935
rect 7271 987 7323 1022
rect 7271 953 7281 987
rect 7315 953 7323 987
rect 7271 918 7323 953
rect 7377 995 7385 1029
rect 7419 995 7429 1029
rect 7377 911 7429 995
rect 7459 1029 7513 1041
rect 7459 995 7469 1029
rect 7503 995 7513 1029
rect 7459 961 7513 995
rect 7459 927 7469 961
rect 7503 927 7513 961
rect 7459 911 7513 927
rect 7543 1029 7617 1041
rect 7543 995 7563 1029
rect 7597 995 7617 1029
rect 7543 911 7617 995
rect 7647 1029 7701 1041
rect 7647 995 7657 1029
rect 7691 995 7701 1029
rect 7647 961 7701 995
rect 7647 927 7657 961
rect 7691 927 7701 961
rect 7647 911 7701 927
rect 7731 1029 7793 1041
rect 7731 995 7741 1029
rect 7775 995 7793 1029
rect 7731 961 7793 995
rect 7731 927 7741 961
rect 7775 927 7793 961
rect 7731 911 7793 927
rect 7847 1029 7909 1041
rect 7847 995 7865 1029
rect 7899 995 7909 1029
rect 7847 961 7909 995
rect 7847 927 7865 961
rect 7899 927 7909 961
rect 7847 911 7909 927
rect 7939 1029 7993 1041
rect 7939 995 7949 1029
rect 7983 995 7993 1029
rect 7939 961 7993 995
rect 7939 927 7949 961
rect 7983 927 7993 961
rect 7939 911 7993 927
rect 8023 1029 8097 1041
rect 8023 995 8043 1029
rect 8077 995 8097 1029
rect 8023 911 8097 995
rect 8127 1029 8181 1041
rect 8127 995 8137 1029
rect 8171 995 8181 1029
rect 8127 961 8181 995
rect 8127 927 8137 961
rect 8171 927 8181 961
rect 8127 911 8181 927
rect 8211 1029 8263 1041
rect 8211 995 8221 1029
rect 8255 995 8263 1029
rect 8211 911 8263 995
rect 8317 987 8369 1022
rect 8317 953 8325 987
rect 8359 953 8369 987
rect 8317 918 8369 953
rect 8399 969 8453 1022
rect 8399 935 8409 969
rect 8443 935 8453 969
rect 8399 918 8453 935
rect 8483 987 8537 1022
rect 8483 953 8493 987
rect 8527 953 8537 987
rect 8483 918 8537 953
rect 8567 969 8621 1022
rect 8567 935 8577 969
rect 8611 935 8621 969
rect 8567 918 8621 935
rect 8651 987 8703 1022
rect 8651 953 8661 987
rect 8695 953 8703 987
rect 8651 918 8703 953
rect 8828 1016 8880 1041
rect 8828 982 8836 1016
rect 8870 982 8880 1016
rect 8828 957 8880 982
rect 8910 1016 8964 1041
rect 8910 982 8920 1016
rect 8954 982 8964 1016
rect 8910 957 8964 982
rect 8994 1016 9046 1041
rect 8994 982 9004 1016
rect 9038 982 9046 1016
rect 8994 957 9046 982
rect 9170 1016 9222 1041
rect 9170 982 9178 1016
rect 9212 982 9222 1016
rect 9170 957 9222 982
rect 9252 1016 9306 1041
rect 9252 982 9262 1016
rect 9296 982 9306 1016
rect 9252 957 9306 982
rect 9336 1016 9388 1041
rect 9336 982 9346 1016
rect 9380 982 9388 1016
rect 9336 957 9388 982
rect 9953 1029 10005 1041
rect 9513 987 9565 1022
rect 9513 953 9521 987
rect 9555 953 9565 987
rect 9513 918 9565 953
rect 9595 969 9649 1022
rect 9595 935 9605 969
rect 9639 935 9649 969
rect 9595 918 9649 935
rect 9679 987 9733 1022
rect 9679 953 9689 987
rect 9723 953 9733 987
rect 9679 918 9733 953
rect 9763 969 9817 1022
rect 9763 935 9773 969
rect 9807 935 9817 969
rect 9763 918 9817 935
rect 9847 987 9899 1022
rect 9847 953 9857 987
rect 9891 953 9899 987
rect 9847 918 9899 953
rect 9953 995 9961 1029
rect 9995 995 10005 1029
rect 9953 911 10005 995
rect 10035 1029 10089 1041
rect 10035 995 10045 1029
rect 10079 995 10089 1029
rect 10035 961 10089 995
rect 10035 927 10045 961
rect 10079 927 10089 961
rect 10035 911 10089 927
rect 10119 1029 10193 1041
rect 10119 995 10139 1029
rect 10173 995 10193 1029
rect 10119 911 10193 995
rect 10223 1029 10277 1041
rect 10223 995 10233 1029
rect 10267 995 10277 1029
rect 10223 961 10277 995
rect 10223 927 10233 961
rect 10267 927 10277 961
rect 10223 911 10277 927
rect 10307 1029 10369 1041
rect 10307 995 10317 1029
rect 10351 995 10369 1029
rect 10307 961 10369 995
rect 10307 927 10317 961
rect 10351 927 10369 961
rect 10307 911 10369 927
rect 27 161 89 177
rect 27 127 45 161
rect 79 127 89 161
rect 27 93 89 127
rect 27 59 45 93
rect 79 59 89 93
rect 27 47 89 59
rect 119 161 173 177
rect 119 127 129 161
rect 163 127 173 161
rect 119 93 173 127
rect 119 59 129 93
rect 163 59 173 93
rect 119 47 173 59
rect 203 93 277 177
rect 203 59 223 93
rect 257 59 277 93
rect 203 47 277 59
rect 307 161 361 177
rect 307 127 317 161
rect 351 127 361 161
rect 307 93 361 127
rect 307 59 317 93
rect 351 59 361 93
rect 307 47 361 59
rect 391 93 443 177
rect 391 59 401 93
rect 435 59 443 93
rect 497 135 549 170
rect 497 101 505 135
rect 539 101 549 135
rect 497 66 549 101
rect 579 153 633 170
rect 579 119 589 153
rect 623 119 633 153
rect 579 66 633 119
rect 663 135 717 170
rect 663 101 673 135
rect 707 101 717 135
rect 663 66 717 101
rect 747 153 801 170
rect 747 119 757 153
rect 791 119 801 153
rect 747 66 801 119
rect 831 135 883 170
rect 831 101 841 135
rect 875 101 883 135
rect 831 66 883 101
rect 391 47 443 59
rect 1008 106 1060 131
rect 1008 72 1016 106
rect 1050 72 1060 106
rect 1008 47 1060 72
rect 1090 106 1144 131
rect 1090 72 1100 106
rect 1134 72 1144 106
rect 1090 47 1144 72
rect 1174 106 1226 131
rect 1174 72 1184 106
rect 1218 72 1226 106
rect 1174 47 1226 72
rect 1350 106 1402 131
rect 1350 72 1358 106
rect 1392 72 1402 106
rect 1350 47 1402 72
rect 1432 106 1486 131
rect 1432 72 1442 106
rect 1476 72 1486 106
rect 1432 47 1486 72
rect 1516 106 1568 131
rect 1516 72 1526 106
rect 1560 72 1568 106
rect 1516 47 1568 72
rect 1693 135 1745 170
rect 1693 101 1701 135
rect 1735 101 1745 135
rect 1693 66 1745 101
rect 1775 153 1829 170
rect 1775 119 1785 153
rect 1819 119 1829 153
rect 1775 66 1829 119
rect 1859 135 1913 170
rect 1859 101 1869 135
rect 1903 101 1913 135
rect 1859 66 1913 101
rect 1943 153 1997 170
rect 1943 119 1953 153
rect 1987 119 1997 153
rect 1943 66 1997 119
rect 2027 135 2079 170
rect 2027 101 2037 135
rect 2071 101 2079 135
rect 2027 66 2079 101
rect 2133 93 2185 177
rect 2133 59 2141 93
rect 2175 59 2185 93
rect 2133 47 2185 59
rect 2215 161 2269 177
rect 2215 127 2225 161
rect 2259 127 2269 161
rect 2215 93 2269 127
rect 2215 59 2225 93
rect 2259 59 2269 93
rect 2215 47 2269 59
rect 2299 93 2373 177
rect 2299 59 2319 93
rect 2353 59 2373 93
rect 2299 47 2373 59
rect 2403 161 2457 177
rect 2403 127 2413 161
rect 2447 127 2457 161
rect 2403 93 2457 127
rect 2403 59 2413 93
rect 2447 59 2457 93
rect 2403 47 2457 59
rect 2487 161 2549 177
rect 2487 127 2497 161
rect 2531 127 2549 161
rect 2487 93 2549 127
rect 2487 59 2497 93
rect 2531 59 2549 93
rect 2487 47 2549 59
rect 2603 161 2665 177
rect 2603 127 2621 161
rect 2655 127 2665 161
rect 2603 93 2665 127
rect 2603 59 2621 93
rect 2655 59 2665 93
rect 2603 47 2665 59
rect 2695 161 2749 177
rect 2695 127 2705 161
rect 2739 127 2749 161
rect 2695 93 2749 127
rect 2695 59 2705 93
rect 2739 59 2749 93
rect 2695 47 2749 59
rect 2779 93 2853 177
rect 2779 59 2799 93
rect 2833 59 2853 93
rect 2779 47 2853 59
rect 2883 161 2937 177
rect 2883 127 2893 161
rect 2927 127 2937 161
rect 2883 93 2937 127
rect 2883 59 2893 93
rect 2927 59 2937 93
rect 2883 47 2937 59
rect 2967 93 3019 177
rect 2967 59 2977 93
rect 3011 59 3019 93
rect 3073 135 3125 170
rect 3073 101 3081 135
rect 3115 101 3125 135
rect 3073 66 3125 101
rect 3155 153 3209 170
rect 3155 119 3165 153
rect 3199 119 3209 153
rect 3155 66 3209 119
rect 3239 135 3293 170
rect 3239 101 3249 135
rect 3283 101 3293 135
rect 3239 66 3293 101
rect 3323 153 3377 170
rect 3323 119 3333 153
rect 3367 119 3377 153
rect 3323 66 3377 119
rect 3407 135 3459 170
rect 3407 101 3417 135
rect 3451 101 3459 135
rect 3407 66 3459 101
rect 2967 47 3019 59
rect 3584 106 3636 131
rect 3584 72 3592 106
rect 3626 72 3636 106
rect 3584 47 3636 72
rect 3666 106 3720 131
rect 3666 72 3676 106
rect 3710 72 3720 106
rect 3666 47 3720 72
rect 3750 106 3802 131
rect 3750 72 3760 106
rect 3794 72 3802 106
rect 3750 47 3802 72
rect 3926 106 3978 131
rect 3926 72 3934 106
rect 3968 72 3978 106
rect 3926 47 3978 72
rect 4008 106 4062 131
rect 4008 72 4018 106
rect 4052 72 4062 106
rect 4008 47 4062 72
rect 4092 106 4144 131
rect 4092 72 4102 106
rect 4136 72 4144 106
rect 4092 47 4144 72
rect 4269 135 4321 170
rect 4269 101 4277 135
rect 4311 101 4321 135
rect 4269 66 4321 101
rect 4351 153 4405 170
rect 4351 119 4361 153
rect 4395 119 4405 153
rect 4351 66 4405 119
rect 4435 135 4489 170
rect 4435 101 4445 135
rect 4479 101 4489 135
rect 4435 66 4489 101
rect 4519 153 4573 170
rect 4519 119 4529 153
rect 4563 119 4573 153
rect 4519 66 4573 119
rect 4603 135 4655 170
rect 4603 101 4613 135
rect 4647 101 4655 135
rect 4603 66 4655 101
rect 4709 93 4761 177
rect 4709 59 4717 93
rect 4751 59 4761 93
rect 4709 47 4761 59
rect 4791 161 4845 177
rect 4791 127 4801 161
rect 4835 127 4845 161
rect 4791 93 4845 127
rect 4791 59 4801 93
rect 4835 59 4845 93
rect 4791 47 4845 59
rect 4875 93 4949 177
rect 4875 59 4895 93
rect 4929 59 4949 93
rect 4875 47 4949 59
rect 4979 161 5033 177
rect 4979 127 4989 161
rect 5023 127 5033 161
rect 4979 93 5033 127
rect 4979 59 4989 93
rect 5023 59 5033 93
rect 4979 47 5033 59
rect 5063 161 5125 177
rect 5063 127 5073 161
rect 5107 127 5125 161
rect 5063 93 5125 127
rect 5063 59 5073 93
rect 5107 59 5125 93
rect 5271 161 5333 177
rect 5271 127 5289 161
rect 5323 127 5333 161
rect 5271 93 5333 127
rect 5063 47 5125 59
rect 5271 59 5289 93
rect 5323 59 5333 93
rect 5271 47 5333 59
rect 5363 161 5417 177
rect 5363 127 5373 161
rect 5407 127 5417 161
rect 5363 93 5417 127
rect 5363 59 5373 93
rect 5407 59 5417 93
rect 5363 47 5417 59
rect 5447 93 5521 177
rect 5447 59 5467 93
rect 5501 59 5521 93
rect 5447 47 5521 59
rect 5551 161 5605 177
rect 5551 127 5561 161
rect 5595 127 5605 161
rect 5551 93 5605 127
rect 5551 59 5561 93
rect 5595 59 5605 93
rect 5551 47 5605 59
rect 5635 93 5687 177
rect 5635 59 5645 93
rect 5679 59 5687 93
rect 5741 135 5793 170
rect 5741 101 5749 135
rect 5783 101 5793 135
rect 5741 66 5793 101
rect 5823 153 5877 170
rect 5823 119 5833 153
rect 5867 119 5877 153
rect 5823 66 5877 119
rect 5907 135 5961 170
rect 5907 101 5917 135
rect 5951 101 5961 135
rect 5907 66 5961 101
rect 5991 153 6045 170
rect 5991 119 6001 153
rect 6035 119 6045 153
rect 5991 66 6045 119
rect 6075 135 6127 170
rect 6075 101 6085 135
rect 6119 101 6127 135
rect 6075 66 6127 101
rect 5635 47 5687 59
rect 6252 106 6304 131
rect 6252 72 6260 106
rect 6294 72 6304 106
rect 6252 47 6304 72
rect 6334 106 6388 131
rect 6334 72 6344 106
rect 6378 72 6388 106
rect 6334 47 6388 72
rect 6418 106 6470 131
rect 6418 72 6428 106
rect 6462 72 6470 106
rect 6418 47 6470 72
rect 6594 106 6646 131
rect 6594 72 6602 106
rect 6636 72 6646 106
rect 6594 47 6646 72
rect 6676 106 6730 131
rect 6676 72 6686 106
rect 6720 72 6730 106
rect 6676 47 6730 72
rect 6760 106 6812 131
rect 6760 72 6770 106
rect 6804 72 6812 106
rect 6760 47 6812 72
rect 6937 135 6989 170
rect 6937 101 6945 135
rect 6979 101 6989 135
rect 6937 66 6989 101
rect 7019 153 7073 170
rect 7019 119 7029 153
rect 7063 119 7073 153
rect 7019 66 7073 119
rect 7103 135 7157 170
rect 7103 101 7113 135
rect 7147 101 7157 135
rect 7103 66 7157 101
rect 7187 153 7241 170
rect 7187 119 7197 153
rect 7231 119 7241 153
rect 7187 66 7241 119
rect 7271 135 7323 170
rect 7271 101 7281 135
rect 7315 101 7323 135
rect 7271 66 7323 101
rect 7377 93 7429 177
rect 7377 59 7385 93
rect 7419 59 7429 93
rect 7377 47 7429 59
rect 7459 161 7513 177
rect 7459 127 7469 161
rect 7503 127 7513 161
rect 7459 93 7513 127
rect 7459 59 7469 93
rect 7503 59 7513 93
rect 7459 47 7513 59
rect 7543 93 7617 177
rect 7543 59 7563 93
rect 7597 59 7617 93
rect 7543 47 7617 59
rect 7647 161 7701 177
rect 7647 127 7657 161
rect 7691 127 7701 161
rect 7647 93 7701 127
rect 7647 59 7657 93
rect 7691 59 7701 93
rect 7647 47 7701 59
rect 7731 161 7793 177
rect 7731 127 7741 161
rect 7775 127 7793 161
rect 7731 93 7793 127
rect 7731 59 7741 93
rect 7775 59 7793 93
rect 7731 47 7793 59
rect 7847 161 7909 177
rect 7847 127 7865 161
rect 7899 127 7909 161
rect 7847 93 7909 127
rect 7847 59 7865 93
rect 7899 59 7909 93
rect 7847 47 7909 59
rect 7939 161 7993 177
rect 7939 127 7949 161
rect 7983 127 7993 161
rect 7939 93 7993 127
rect 7939 59 7949 93
rect 7983 59 7993 93
rect 7939 47 7993 59
rect 8023 93 8097 177
rect 8023 59 8043 93
rect 8077 59 8097 93
rect 8023 47 8097 59
rect 8127 161 8181 177
rect 8127 127 8137 161
rect 8171 127 8181 161
rect 8127 93 8181 127
rect 8127 59 8137 93
rect 8171 59 8181 93
rect 8127 47 8181 59
rect 8211 93 8263 177
rect 8211 59 8221 93
rect 8255 59 8263 93
rect 8317 135 8369 170
rect 8317 101 8325 135
rect 8359 101 8369 135
rect 8317 66 8369 101
rect 8399 153 8453 170
rect 8399 119 8409 153
rect 8443 119 8453 153
rect 8399 66 8453 119
rect 8483 135 8537 170
rect 8483 101 8493 135
rect 8527 101 8537 135
rect 8483 66 8537 101
rect 8567 153 8621 170
rect 8567 119 8577 153
rect 8611 119 8621 153
rect 8567 66 8621 119
rect 8651 135 8703 170
rect 8651 101 8661 135
rect 8695 101 8703 135
rect 8651 66 8703 101
rect 8211 47 8263 59
rect 8828 106 8880 131
rect 8828 72 8836 106
rect 8870 72 8880 106
rect 8828 47 8880 72
rect 8910 106 8964 131
rect 8910 72 8920 106
rect 8954 72 8964 106
rect 8910 47 8964 72
rect 8994 106 9046 131
rect 8994 72 9004 106
rect 9038 72 9046 106
rect 8994 47 9046 72
rect 9170 106 9222 131
rect 9170 72 9178 106
rect 9212 72 9222 106
rect 9170 47 9222 72
rect 9252 106 9306 131
rect 9252 72 9262 106
rect 9296 72 9306 106
rect 9252 47 9306 72
rect 9336 106 9388 131
rect 9336 72 9346 106
rect 9380 72 9388 106
rect 9336 47 9388 72
rect 9513 135 9565 170
rect 9513 101 9521 135
rect 9555 101 9565 135
rect 9513 66 9565 101
rect 9595 153 9649 170
rect 9595 119 9605 153
rect 9639 119 9649 153
rect 9595 66 9649 119
rect 9679 135 9733 170
rect 9679 101 9689 135
rect 9723 101 9733 135
rect 9679 66 9733 101
rect 9763 153 9817 170
rect 9763 119 9773 153
rect 9807 119 9817 153
rect 9763 66 9817 119
rect 9847 135 9899 170
rect 9847 101 9857 135
rect 9891 101 9899 135
rect 9847 66 9899 101
rect 9953 93 10005 177
rect 9953 59 9961 93
rect 9995 59 10005 93
rect 9953 47 10005 59
rect 10035 161 10089 177
rect 10035 127 10045 161
rect 10079 127 10089 161
rect 10035 93 10089 127
rect 10035 59 10045 93
rect 10079 59 10089 93
rect 10035 47 10089 59
rect 10119 93 10193 177
rect 10119 59 10139 93
rect 10173 59 10193 93
rect 10119 47 10193 59
rect 10223 161 10277 177
rect 10223 127 10233 161
rect 10267 127 10277 161
rect 10223 93 10277 127
rect 10223 59 10233 93
rect 10267 59 10277 93
rect 10223 47 10277 59
rect 10307 161 10369 177
rect 10307 127 10317 161
rect 10351 127 10369 161
rect 10307 93 10369 127
rect 10307 59 10317 93
rect 10351 59 10369 93
rect 10307 47 10369 59
<< pdiff >>
rect 27 773 81 791
rect 27 739 35 773
rect 69 739 81 773
rect 27 705 81 739
rect 27 671 35 705
rect 69 671 81 705
rect 27 637 81 671
rect 27 603 35 637
rect 69 603 81 637
rect 27 591 81 603
rect 117 773 175 791
rect 117 739 129 773
rect 163 739 175 773
rect 117 705 175 739
rect 117 671 129 705
rect 163 671 175 705
rect 117 637 175 671
rect 117 603 129 637
rect 163 603 175 637
rect 117 591 175 603
rect 211 705 269 791
rect 211 671 223 705
rect 257 671 269 705
rect 211 637 269 671
rect 211 603 223 637
rect 257 603 269 637
rect 211 591 269 603
rect 305 773 363 791
rect 305 739 317 773
rect 351 739 363 773
rect 305 705 363 739
rect 305 671 317 705
rect 351 671 363 705
rect 305 637 363 671
rect 305 603 317 637
rect 351 603 363 637
rect 305 591 363 603
rect 399 705 453 791
rect 399 671 411 705
rect 445 671 453 705
rect 399 637 453 671
rect 399 603 411 637
rect 445 603 453 637
rect 507 765 561 777
rect 507 731 515 765
rect 549 731 561 765
rect 507 659 561 731
rect 507 625 515 659
rect 549 625 561 659
rect 507 613 561 625
rect 597 765 655 777
rect 597 731 609 765
rect 643 731 655 765
rect 597 659 655 731
rect 597 625 609 659
rect 643 625 655 659
rect 597 613 655 625
rect 691 765 749 777
rect 691 731 703 765
rect 737 731 749 765
rect 691 659 749 731
rect 691 625 703 659
rect 737 625 749 659
rect 691 613 749 625
rect 785 765 843 777
rect 785 731 797 765
rect 831 731 843 765
rect 785 659 843 731
rect 785 625 797 659
rect 831 625 843 659
rect 785 613 843 625
rect 879 759 933 777
rect 879 725 891 759
rect 925 725 933 759
rect 879 659 933 725
rect 879 625 891 659
rect 925 625 933 659
rect 879 613 933 625
rect 998 751 1052 763
rect 998 717 1006 751
rect 1040 717 1052 751
rect 998 645 1052 717
rect 399 591 453 603
rect 998 611 1006 645
rect 1040 611 1052 645
rect 998 599 1052 611
rect 1088 751 1146 763
rect 1088 717 1100 751
rect 1134 717 1146 751
rect 1088 645 1146 717
rect 1088 611 1100 645
rect 1134 611 1146 645
rect 1088 599 1146 611
rect 1182 751 1236 763
rect 1182 717 1194 751
rect 1228 717 1236 751
rect 1182 645 1236 717
rect 1182 611 1194 645
rect 1228 611 1236 645
rect 1182 599 1236 611
rect 1340 751 1394 763
rect 1340 717 1348 751
rect 1382 717 1394 751
rect 1340 645 1394 717
rect 1340 611 1348 645
rect 1382 611 1394 645
rect 1340 599 1394 611
rect 1430 751 1488 763
rect 1430 717 1442 751
rect 1476 717 1488 751
rect 1430 645 1488 717
rect 1430 611 1442 645
rect 1476 611 1488 645
rect 1430 599 1488 611
rect 1524 751 1578 763
rect 1524 717 1536 751
rect 1570 717 1578 751
rect 1524 645 1578 717
rect 1524 611 1536 645
rect 1570 611 1578 645
rect 1643 759 1697 777
rect 1643 725 1651 759
rect 1685 725 1697 759
rect 1643 659 1697 725
rect 1643 625 1651 659
rect 1685 625 1697 659
rect 1643 613 1697 625
rect 1733 765 1791 777
rect 1733 731 1745 765
rect 1779 731 1791 765
rect 1733 659 1791 731
rect 1733 625 1745 659
rect 1779 625 1791 659
rect 1733 613 1791 625
rect 1827 765 1885 777
rect 1827 731 1839 765
rect 1873 731 1885 765
rect 1827 659 1885 731
rect 1827 625 1839 659
rect 1873 625 1885 659
rect 1827 613 1885 625
rect 1921 765 1979 777
rect 1921 731 1933 765
rect 1967 731 1979 765
rect 1921 659 1979 731
rect 1921 625 1933 659
rect 1967 625 1979 659
rect 1921 613 1979 625
rect 2015 765 2069 777
rect 2015 731 2027 765
rect 2061 731 2069 765
rect 2015 659 2069 731
rect 2015 625 2027 659
rect 2061 625 2069 659
rect 2015 613 2069 625
rect 2123 705 2177 791
rect 2123 671 2131 705
rect 2165 671 2177 705
rect 2123 637 2177 671
rect 1524 599 1578 611
rect 2123 603 2131 637
rect 2165 603 2177 637
rect 2123 591 2177 603
rect 2213 773 2271 791
rect 2213 739 2225 773
rect 2259 739 2271 773
rect 2213 705 2271 739
rect 2213 671 2225 705
rect 2259 671 2271 705
rect 2213 637 2271 671
rect 2213 603 2225 637
rect 2259 603 2271 637
rect 2213 591 2271 603
rect 2307 705 2365 791
rect 2307 671 2319 705
rect 2353 671 2365 705
rect 2307 637 2365 671
rect 2307 603 2319 637
rect 2353 603 2365 637
rect 2307 591 2365 603
rect 2401 773 2459 791
rect 2401 739 2413 773
rect 2447 739 2459 773
rect 2401 705 2459 739
rect 2401 671 2413 705
rect 2447 671 2459 705
rect 2401 637 2459 671
rect 2401 603 2413 637
rect 2447 603 2459 637
rect 2401 591 2459 603
rect 2495 773 2549 791
rect 2495 739 2507 773
rect 2541 739 2549 773
rect 2495 705 2549 739
rect 2495 671 2507 705
rect 2541 671 2549 705
rect 2495 637 2549 671
rect 2495 603 2507 637
rect 2541 603 2549 637
rect 2495 591 2549 603
rect 2603 773 2657 791
rect 2603 739 2611 773
rect 2645 739 2657 773
rect 2603 705 2657 739
rect 2603 671 2611 705
rect 2645 671 2657 705
rect 2603 637 2657 671
rect 2603 603 2611 637
rect 2645 603 2657 637
rect 2603 591 2657 603
rect 2693 773 2751 791
rect 2693 739 2705 773
rect 2739 739 2751 773
rect 2693 705 2751 739
rect 2693 671 2705 705
rect 2739 671 2751 705
rect 2693 637 2751 671
rect 2693 603 2705 637
rect 2739 603 2751 637
rect 2693 591 2751 603
rect 2787 705 2845 791
rect 2787 671 2799 705
rect 2833 671 2845 705
rect 2787 637 2845 671
rect 2787 603 2799 637
rect 2833 603 2845 637
rect 2787 591 2845 603
rect 2881 773 2939 791
rect 2881 739 2893 773
rect 2927 739 2939 773
rect 2881 705 2939 739
rect 2881 671 2893 705
rect 2927 671 2939 705
rect 2881 637 2939 671
rect 2881 603 2893 637
rect 2927 603 2939 637
rect 2881 591 2939 603
rect 2975 705 3029 791
rect 2975 671 2987 705
rect 3021 671 3029 705
rect 2975 637 3029 671
rect 2975 603 2987 637
rect 3021 603 3029 637
rect 3083 765 3137 777
rect 3083 731 3091 765
rect 3125 731 3137 765
rect 3083 659 3137 731
rect 3083 625 3091 659
rect 3125 625 3137 659
rect 3083 613 3137 625
rect 3173 765 3231 777
rect 3173 731 3185 765
rect 3219 731 3231 765
rect 3173 659 3231 731
rect 3173 625 3185 659
rect 3219 625 3231 659
rect 3173 613 3231 625
rect 3267 765 3325 777
rect 3267 731 3279 765
rect 3313 731 3325 765
rect 3267 659 3325 731
rect 3267 625 3279 659
rect 3313 625 3325 659
rect 3267 613 3325 625
rect 3361 765 3419 777
rect 3361 731 3373 765
rect 3407 731 3419 765
rect 3361 659 3419 731
rect 3361 625 3373 659
rect 3407 625 3419 659
rect 3361 613 3419 625
rect 3455 759 3509 777
rect 3455 725 3467 759
rect 3501 725 3509 759
rect 3455 659 3509 725
rect 3455 625 3467 659
rect 3501 625 3509 659
rect 3455 613 3509 625
rect 3574 751 3628 763
rect 3574 717 3582 751
rect 3616 717 3628 751
rect 3574 645 3628 717
rect 2975 591 3029 603
rect 3574 611 3582 645
rect 3616 611 3628 645
rect 3574 599 3628 611
rect 3664 751 3722 763
rect 3664 717 3676 751
rect 3710 717 3722 751
rect 3664 645 3722 717
rect 3664 611 3676 645
rect 3710 611 3722 645
rect 3664 599 3722 611
rect 3758 751 3812 763
rect 3758 717 3770 751
rect 3804 717 3812 751
rect 3758 645 3812 717
rect 3758 611 3770 645
rect 3804 611 3812 645
rect 3758 599 3812 611
rect 3916 751 3970 763
rect 3916 717 3924 751
rect 3958 717 3970 751
rect 3916 645 3970 717
rect 3916 611 3924 645
rect 3958 611 3970 645
rect 3916 599 3970 611
rect 4006 751 4064 763
rect 4006 717 4018 751
rect 4052 717 4064 751
rect 4006 645 4064 717
rect 4006 611 4018 645
rect 4052 611 4064 645
rect 4006 599 4064 611
rect 4100 751 4154 763
rect 4100 717 4112 751
rect 4146 717 4154 751
rect 4100 645 4154 717
rect 4100 611 4112 645
rect 4146 611 4154 645
rect 4219 759 4273 777
rect 4219 725 4227 759
rect 4261 725 4273 759
rect 4219 659 4273 725
rect 4219 625 4227 659
rect 4261 625 4273 659
rect 4219 613 4273 625
rect 4309 765 4367 777
rect 4309 731 4321 765
rect 4355 731 4367 765
rect 4309 659 4367 731
rect 4309 625 4321 659
rect 4355 625 4367 659
rect 4309 613 4367 625
rect 4403 765 4461 777
rect 4403 731 4415 765
rect 4449 731 4461 765
rect 4403 659 4461 731
rect 4403 625 4415 659
rect 4449 625 4461 659
rect 4403 613 4461 625
rect 4497 765 4555 777
rect 4497 731 4509 765
rect 4543 731 4555 765
rect 4497 659 4555 731
rect 4497 625 4509 659
rect 4543 625 4555 659
rect 4497 613 4555 625
rect 4591 765 4645 777
rect 4591 731 4603 765
rect 4637 731 4645 765
rect 4591 659 4645 731
rect 4591 625 4603 659
rect 4637 625 4645 659
rect 4591 613 4645 625
rect 4699 705 4753 791
rect 4699 671 4707 705
rect 4741 671 4753 705
rect 4699 637 4753 671
rect 4100 599 4154 611
rect 4699 603 4707 637
rect 4741 603 4753 637
rect 4699 591 4753 603
rect 4789 773 4847 791
rect 4789 739 4801 773
rect 4835 739 4847 773
rect 4789 705 4847 739
rect 4789 671 4801 705
rect 4835 671 4847 705
rect 4789 637 4847 671
rect 4789 603 4801 637
rect 4835 603 4847 637
rect 4789 591 4847 603
rect 4883 705 4941 791
rect 4883 671 4895 705
rect 4929 671 4941 705
rect 4883 637 4941 671
rect 4883 603 4895 637
rect 4929 603 4941 637
rect 4883 591 4941 603
rect 4977 773 5035 791
rect 4977 739 4989 773
rect 5023 739 5035 773
rect 4977 705 5035 739
rect 4977 671 4989 705
rect 5023 671 5035 705
rect 4977 637 5035 671
rect 4977 603 4989 637
rect 5023 603 5035 637
rect 4977 591 5035 603
rect 5071 773 5125 791
rect 5071 739 5083 773
rect 5117 739 5125 773
rect 5071 705 5125 739
rect 5071 671 5083 705
rect 5117 671 5125 705
rect 5071 637 5125 671
rect 5071 603 5083 637
rect 5117 603 5125 637
rect 5271 773 5325 791
rect 5271 739 5279 773
rect 5313 739 5325 773
rect 5271 705 5325 739
rect 5271 671 5279 705
rect 5313 671 5325 705
rect 5271 637 5325 671
rect 5071 591 5125 603
rect 5271 603 5279 637
rect 5313 603 5325 637
rect 5271 591 5325 603
rect 5361 773 5419 791
rect 5361 739 5373 773
rect 5407 739 5419 773
rect 5361 705 5419 739
rect 5361 671 5373 705
rect 5407 671 5419 705
rect 5361 637 5419 671
rect 5361 603 5373 637
rect 5407 603 5419 637
rect 5361 591 5419 603
rect 5455 705 5513 791
rect 5455 671 5467 705
rect 5501 671 5513 705
rect 5455 637 5513 671
rect 5455 603 5467 637
rect 5501 603 5513 637
rect 5455 591 5513 603
rect 5549 773 5607 791
rect 5549 739 5561 773
rect 5595 739 5607 773
rect 5549 705 5607 739
rect 5549 671 5561 705
rect 5595 671 5607 705
rect 5549 637 5607 671
rect 5549 603 5561 637
rect 5595 603 5607 637
rect 5549 591 5607 603
rect 5643 705 5697 791
rect 5643 671 5655 705
rect 5689 671 5697 705
rect 5643 637 5697 671
rect 5643 603 5655 637
rect 5689 603 5697 637
rect 5751 765 5805 777
rect 5751 731 5759 765
rect 5793 731 5805 765
rect 5751 659 5805 731
rect 5751 625 5759 659
rect 5793 625 5805 659
rect 5751 613 5805 625
rect 5841 765 5899 777
rect 5841 731 5853 765
rect 5887 731 5899 765
rect 5841 659 5899 731
rect 5841 625 5853 659
rect 5887 625 5899 659
rect 5841 613 5899 625
rect 5935 765 5993 777
rect 5935 731 5947 765
rect 5981 731 5993 765
rect 5935 659 5993 731
rect 5935 625 5947 659
rect 5981 625 5993 659
rect 5935 613 5993 625
rect 6029 765 6087 777
rect 6029 731 6041 765
rect 6075 731 6087 765
rect 6029 659 6087 731
rect 6029 625 6041 659
rect 6075 625 6087 659
rect 6029 613 6087 625
rect 6123 759 6177 777
rect 6123 725 6135 759
rect 6169 725 6177 759
rect 6123 659 6177 725
rect 6123 625 6135 659
rect 6169 625 6177 659
rect 6123 613 6177 625
rect 6242 751 6296 763
rect 6242 717 6250 751
rect 6284 717 6296 751
rect 6242 645 6296 717
rect 5643 591 5697 603
rect 6242 611 6250 645
rect 6284 611 6296 645
rect 6242 599 6296 611
rect 6332 751 6390 763
rect 6332 717 6344 751
rect 6378 717 6390 751
rect 6332 645 6390 717
rect 6332 611 6344 645
rect 6378 611 6390 645
rect 6332 599 6390 611
rect 6426 751 6480 763
rect 6426 717 6438 751
rect 6472 717 6480 751
rect 6426 645 6480 717
rect 6426 611 6438 645
rect 6472 611 6480 645
rect 6426 599 6480 611
rect 6584 751 6638 763
rect 6584 717 6592 751
rect 6626 717 6638 751
rect 6584 645 6638 717
rect 6584 611 6592 645
rect 6626 611 6638 645
rect 6584 599 6638 611
rect 6674 751 6732 763
rect 6674 717 6686 751
rect 6720 717 6732 751
rect 6674 645 6732 717
rect 6674 611 6686 645
rect 6720 611 6732 645
rect 6674 599 6732 611
rect 6768 751 6822 763
rect 6768 717 6780 751
rect 6814 717 6822 751
rect 6768 645 6822 717
rect 6768 611 6780 645
rect 6814 611 6822 645
rect 6887 759 6941 777
rect 6887 725 6895 759
rect 6929 725 6941 759
rect 6887 659 6941 725
rect 6887 625 6895 659
rect 6929 625 6941 659
rect 6887 613 6941 625
rect 6977 765 7035 777
rect 6977 731 6989 765
rect 7023 731 7035 765
rect 6977 659 7035 731
rect 6977 625 6989 659
rect 7023 625 7035 659
rect 6977 613 7035 625
rect 7071 765 7129 777
rect 7071 731 7083 765
rect 7117 731 7129 765
rect 7071 659 7129 731
rect 7071 625 7083 659
rect 7117 625 7129 659
rect 7071 613 7129 625
rect 7165 765 7223 777
rect 7165 731 7177 765
rect 7211 731 7223 765
rect 7165 659 7223 731
rect 7165 625 7177 659
rect 7211 625 7223 659
rect 7165 613 7223 625
rect 7259 765 7313 777
rect 7259 731 7271 765
rect 7305 731 7313 765
rect 7259 659 7313 731
rect 7259 625 7271 659
rect 7305 625 7313 659
rect 7259 613 7313 625
rect 7367 705 7421 791
rect 7367 671 7375 705
rect 7409 671 7421 705
rect 7367 637 7421 671
rect 6768 599 6822 611
rect 7367 603 7375 637
rect 7409 603 7421 637
rect 7367 591 7421 603
rect 7457 773 7515 791
rect 7457 739 7469 773
rect 7503 739 7515 773
rect 7457 705 7515 739
rect 7457 671 7469 705
rect 7503 671 7515 705
rect 7457 637 7515 671
rect 7457 603 7469 637
rect 7503 603 7515 637
rect 7457 591 7515 603
rect 7551 705 7609 791
rect 7551 671 7563 705
rect 7597 671 7609 705
rect 7551 637 7609 671
rect 7551 603 7563 637
rect 7597 603 7609 637
rect 7551 591 7609 603
rect 7645 773 7703 791
rect 7645 739 7657 773
rect 7691 739 7703 773
rect 7645 705 7703 739
rect 7645 671 7657 705
rect 7691 671 7703 705
rect 7645 637 7703 671
rect 7645 603 7657 637
rect 7691 603 7703 637
rect 7645 591 7703 603
rect 7739 773 7793 791
rect 7739 739 7751 773
rect 7785 739 7793 773
rect 7739 705 7793 739
rect 7739 671 7751 705
rect 7785 671 7793 705
rect 7739 637 7793 671
rect 7739 603 7751 637
rect 7785 603 7793 637
rect 7739 591 7793 603
rect 7847 773 7901 791
rect 7847 739 7855 773
rect 7889 739 7901 773
rect 7847 705 7901 739
rect 7847 671 7855 705
rect 7889 671 7901 705
rect 7847 637 7901 671
rect 7847 603 7855 637
rect 7889 603 7901 637
rect 7847 591 7901 603
rect 7937 773 7995 791
rect 7937 739 7949 773
rect 7983 739 7995 773
rect 7937 705 7995 739
rect 7937 671 7949 705
rect 7983 671 7995 705
rect 7937 637 7995 671
rect 7937 603 7949 637
rect 7983 603 7995 637
rect 7937 591 7995 603
rect 8031 705 8089 791
rect 8031 671 8043 705
rect 8077 671 8089 705
rect 8031 637 8089 671
rect 8031 603 8043 637
rect 8077 603 8089 637
rect 8031 591 8089 603
rect 8125 773 8183 791
rect 8125 739 8137 773
rect 8171 739 8183 773
rect 8125 705 8183 739
rect 8125 671 8137 705
rect 8171 671 8183 705
rect 8125 637 8183 671
rect 8125 603 8137 637
rect 8171 603 8183 637
rect 8125 591 8183 603
rect 8219 705 8273 791
rect 8219 671 8231 705
rect 8265 671 8273 705
rect 8219 637 8273 671
rect 8219 603 8231 637
rect 8265 603 8273 637
rect 8327 765 8381 777
rect 8327 731 8335 765
rect 8369 731 8381 765
rect 8327 659 8381 731
rect 8327 625 8335 659
rect 8369 625 8381 659
rect 8327 613 8381 625
rect 8417 765 8475 777
rect 8417 731 8429 765
rect 8463 731 8475 765
rect 8417 659 8475 731
rect 8417 625 8429 659
rect 8463 625 8475 659
rect 8417 613 8475 625
rect 8511 765 8569 777
rect 8511 731 8523 765
rect 8557 731 8569 765
rect 8511 659 8569 731
rect 8511 625 8523 659
rect 8557 625 8569 659
rect 8511 613 8569 625
rect 8605 765 8663 777
rect 8605 731 8617 765
rect 8651 731 8663 765
rect 8605 659 8663 731
rect 8605 625 8617 659
rect 8651 625 8663 659
rect 8605 613 8663 625
rect 8699 759 8753 777
rect 8699 725 8711 759
rect 8745 725 8753 759
rect 8699 659 8753 725
rect 8699 625 8711 659
rect 8745 625 8753 659
rect 8699 613 8753 625
rect 8818 751 8872 763
rect 8818 717 8826 751
rect 8860 717 8872 751
rect 8818 645 8872 717
rect 8219 591 8273 603
rect 8818 611 8826 645
rect 8860 611 8872 645
rect 8818 599 8872 611
rect 8908 751 8966 763
rect 8908 717 8920 751
rect 8954 717 8966 751
rect 8908 645 8966 717
rect 8908 611 8920 645
rect 8954 611 8966 645
rect 8908 599 8966 611
rect 9002 751 9056 763
rect 9002 717 9014 751
rect 9048 717 9056 751
rect 9002 645 9056 717
rect 9002 611 9014 645
rect 9048 611 9056 645
rect 9002 599 9056 611
rect 9160 751 9214 763
rect 9160 717 9168 751
rect 9202 717 9214 751
rect 9160 645 9214 717
rect 9160 611 9168 645
rect 9202 611 9214 645
rect 9160 599 9214 611
rect 9250 751 9308 763
rect 9250 717 9262 751
rect 9296 717 9308 751
rect 9250 645 9308 717
rect 9250 611 9262 645
rect 9296 611 9308 645
rect 9250 599 9308 611
rect 9344 751 9398 763
rect 9344 717 9356 751
rect 9390 717 9398 751
rect 9344 645 9398 717
rect 9344 611 9356 645
rect 9390 611 9398 645
rect 9463 759 9517 777
rect 9463 725 9471 759
rect 9505 725 9517 759
rect 9463 659 9517 725
rect 9463 625 9471 659
rect 9505 625 9517 659
rect 9463 613 9517 625
rect 9553 765 9611 777
rect 9553 731 9565 765
rect 9599 731 9611 765
rect 9553 659 9611 731
rect 9553 625 9565 659
rect 9599 625 9611 659
rect 9553 613 9611 625
rect 9647 765 9705 777
rect 9647 731 9659 765
rect 9693 731 9705 765
rect 9647 659 9705 731
rect 9647 625 9659 659
rect 9693 625 9705 659
rect 9647 613 9705 625
rect 9741 765 9799 777
rect 9741 731 9753 765
rect 9787 731 9799 765
rect 9741 659 9799 731
rect 9741 625 9753 659
rect 9787 625 9799 659
rect 9741 613 9799 625
rect 9835 765 9889 777
rect 9835 731 9847 765
rect 9881 731 9889 765
rect 9835 659 9889 731
rect 9835 625 9847 659
rect 9881 625 9889 659
rect 9835 613 9889 625
rect 9943 705 9997 791
rect 9943 671 9951 705
rect 9985 671 9997 705
rect 9943 637 9997 671
rect 9344 599 9398 611
rect 9943 603 9951 637
rect 9985 603 9997 637
rect 9943 591 9997 603
rect 10033 773 10091 791
rect 10033 739 10045 773
rect 10079 739 10091 773
rect 10033 705 10091 739
rect 10033 671 10045 705
rect 10079 671 10091 705
rect 10033 637 10091 671
rect 10033 603 10045 637
rect 10079 603 10091 637
rect 10033 591 10091 603
rect 10127 705 10185 791
rect 10127 671 10139 705
rect 10173 671 10185 705
rect 10127 637 10185 671
rect 10127 603 10139 637
rect 10173 603 10185 637
rect 10127 591 10185 603
rect 10221 773 10279 791
rect 10221 739 10233 773
rect 10267 739 10279 773
rect 10221 705 10279 739
rect 10221 671 10233 705
rect 10267 671 10279 705
rect 10221 637 10279 671
rect 10221 603 10233 637
rect 10267 603 10279 637
rect 10221 591 10279 603
rect 10315 773 10369 791
rect 10315 739 10327 773
rect 10361 739 10369 773
rect 10315 705 10369 739
rect 10315 671 10327 705
rect 10361 671 10369 705
rect 10315 637 10369 671
rect 10315 603 10327 637
rect 10361 603 10369 637
rect 10315 591 10369 603
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 485 175 497
rect 117 451 129 485
rect 163 451 175 485
rect 117 417 175 451
rect 117 383 129 417
rect 163 383 175 417
rect 117 349 175 383
rect 117 315 129 349
rect 163 315 175 349
rect 117 297 175 315
rect 211 485 269 497
rect 211 451 223 485
rect 257 451 269 485
rect 211 417 269 451
rect 211 383 223 417
rect 257 383 269 417
rect 211 297 269 383
rect 305 485 363 497
rect 305 451 317 485
rect 351 451 363 485
rect 305 417 363 451
rect 305 383 317 417
rect 351 383 363 417
rect 305 349 363 383
rect 305 315 317 349
rect 351 315 363 349
rect 305 297 363 315
rect 399 485 453 497
rect 399 451 411 485
rect 445 451 453 485
rect 998 477 1052 489
rect 399 417 453 451
rect 399 383 411 417
rect 445 383 453 417
rect 399 297 453 383
rect 507 463 561 475
rect 507 429 515 463
rect 549 429 561 463
rect 507 357 561 429
rect 507 323 515 357
rect 549 323 561 357
rect 507 311 561 323
rect 597 463 655 475
rect 597 429 609 463
rect 643 429 655 463
rect 597 357 655 429
rect 597 323 609 357
rect 643 323 655 357
rect 597 311 655 323
rect 691 463 749 475
rect 691 429 703 463
rect 737 429 749 463
rect 691 357 749 429
rect 691 323 703 357
rect 737 323 749 357
rect 691 311 749 323
rect 785 463 843 475
rect 785 429 797 463
rect 831 429 843 463
rect 785 357 843 429
rect 785 323 797 357
rect 831 323 843 357
rect 785 311 843 323
rect 879 463 933 475
rect 879 429 891 463
rect 925 429 933 463
rect 879 363 933 429
rect 879 329 891 363
rect 925 329 933 363
rect 879 311 933 329
rect 998 443 1006 477
rect 1040 443 1052 477
rect 998 371 1052 443
rect 998 337 1006 371
rect 1040 337 1052 371
rect 998 325 1052 337
rect 1088 477 1146 489
rect 1088 443 1100 477
rect 1134 443 1146 477
rect 1088 371 1146 443
rect 1088 337 1100 371
rect 1134 337 1146 371
rect 1088 325 1146 337
rect 1182 477 1236 489
rect 1182 443 1194 477
rect 1228 443 1236 477
rect 1182 371 1236 443
rect 1182 337 1194 371
rect 1228 337 1236 371
rect 1182 325 1236 337
rect 1340 477 1394 489
rect 1340 443 1348 477
rect 1382 443 1394 477
rect 1340 371 1394 443
rect 1340 337 1348 371
rect 1382 337 1394 371
rect 1340 325 1394 337
rect 1430 477 1488 489
rect 1430 443 1442 477
rect 1476 443 1488 477
rect 1430 371 1488 443
rect 1430 337 1442 371
rect 1476 337 1488 371
rect 1430 325 1488 337
rect 1524 477 1578 489
rect 1524 443 1536 477
rect 1570 443 1578 477
rect 2123 485 2177 497
rect 1524 371 1578 443
rect 1524 337 1536 371
rect 1570 337 1578 371
rect 1524 325 1578 337
rect 1643 463 1697 475
rect 1643 429 1651 463
rect 1685 429 1697 463
rect 1643 363 1697 429
rect 1643 329 1651 363
rect 1685 329 1697 363
rect 1643 311 1697 329
rect 1733 463 1791 475
rect 1733 429 1745 463
rect 1779 429 1791 463
rect 1733 357 1791 429
rect 1733 323 1745 357
rect 1779 323 1791 357
rect 1733 311 1791 323
rect 1827 463 1885 475
rect 1827 429 1839 463
rect 1873 429 1885 463
rect 1827 357 1885 429
rect 1827 323 1839 357
rect 1873 323 1885 357
rect 1827 311 1885 323
rect 1921 463 1979 475
rect 1921 429 1933 463
rect 1967 429 1979 463
rect 1921 357 1979 429
rect 1921 323 1933 357
rect 1967 323 1979 357
rect 1921 311 1979 323
rect 2015 463 2069 475
rect 2015 429 2027 463
rect 2061 429 2069 463
rect 2015 357 2069 429
rect 2015 323 2027 357
rect 2061 323 2069 357
rect 2015 311 2069 323
rect 2123 451 2131 485
rect 2165 451 2177 485
rect 2123 417 2177 451
rect 2123 383 2131 417
rect 2165 383 2177 417
rect 2123 297 2177 383
rect 2213 485 2271 497
rect 2213 451 2225 485
rect 2259 451 2271 485
rect 2213 417 2271 451
rect 2213 383 2225 417
rect 2259 383 2271 417
rect 2213 349 2271 383
rect 2213 315 2225 349
rect 2259 315 2271 349
rect 2213 297 2271 315
rect 2307 485 2365 497
rect 2307 451 2319 485
rect 2353 451 2365 485
rect 2307 417 2365 451
rect 2307 383 2319 417
rect 2353 383 2365 417
rect 2307 297 2365 383
rect 2401 485 2459 497
rect 2401 451 2413 485
rect 2447 451 2459 485
rect 2401 417 2459 451
rect 2401 383 2413 417
rect 2447 383 2459 417
rect 2401 349 2459 383
rect 2401 315 2413 349
rect 2447 315 2459 349
rect 2401 297 2459 315
rect 2495 485 2549 497
rect 2495 451 2507 485
rect 2541 451 2549 485
rect 2495 417 2549 451
rect 2495 383 2507 417
rect 2541 383 2549 417
rect 2495 349 2549 383
rect 2495 315 2507 349
rect 2541 315 2549 349
rect 2495 297 2549 315
rect 2603 485 2657 497
rect 2603 451 2611 485
rect 2645 451 2657 485
rect 2603 417 2657 451
rect 2603 383 2611 417
rect 2645 383 2657 417
rect 2603 349 2657 383
rect 2603 315 2611 349
rect 2645 315 2657 349
rect 2603 297 2657 315
rect 2693 485 2751 497
rect 2693 451 2705 485
rect 2739 451 2751 485
rect 2693 417 2751 451
rect 2693 383 2705 417
rect 2739 383 2751 417
rect 2693 349 2751 383
rect 2693 315 2705 349
rect 2739 315 2751 349
rect 2693 297 2751 315
rect 2787 485 2845 497
rect 2787 451 2799 485
rect 2833 451 2845 485
rect 2787 417 2845 451
rect 2787 383 2799 417
rect 2833 383 2845 417
rect 2787 297 2845 383
rect 2881 485 2939 497
rect 2881 451 2893 485
rect 2927 451 2939 485
rect 2881 417 2939 451
rect 2881 383 2893 417
rect 2927 383 2939 417
rect 2881 349 2939 383
rect 2881 315 2893 349
rect 2927 315 2939 349
rect 2881 297 2939 315
rect 2975 485 3029 497
rect 2975 451 2987 485
rect 3021 451 3029 485
rect 3574 477 3628 489
rect 2975 417 3029 451
rect 2975 383 2987 417
rect 3021 383 3029 417
rect 2975 297 3029 383
rect 3083 463 3137 475
rect 3083 429 3091 463
rect 3125 429 3137 463
rect 3083 357 3137 429
rect 3083 323 3091 357
rect 3125 323 3137 357
rect 3083 311 3137 323
rect 3173 463 3231 475
rect 3173 429 3185 463
rect 3219 429 3231 463
rect 3173 357 3231 429
rect 3173 323 3185 357
rect 3219 323 3231 357
rect 3173 311 3231 323
rect 3267 463 3325 475
rect 3267 429 3279 463
rect 3313 429 3325 463
rect 3267 357 3325 429
rect 3267 323 3279 357
rect 3313 323 3325 357
rect 3267 311 3325 323
rect 3361 463 3419 475
rect 3361 429 3373 463
rect 3407 429 3419 463
rect 3361 357 3419 429
rect 3361 323 3373 357
rect 3407 323 3419 357
rect 3361 311 3419 323
rect 3455 463 3509 475
rect 3455 429 3467 463
rect 3501 429 3509 463
rect 3455 363 3509 429
rect 3455 329 3467 363
rect 3501 329 3509 363
rect 3455 311 3509 329
rect 3574 443 3582 477
rect 3616 443 3628 477
rect 3574 371 3628 443
rect 3574 337 3582 371
rect 3616 337 3628 371
rect 3574 325 3628 337
rect 3664 477 3722 489
rect 3664 443 3676 477
rect 3710 443 3722 477
rect 3664 371 3722 443
rect 3664 337 3676 371
rect 3710 337 3722 371
rect 3664 325 3722 337
rect 3758 477 3812 489
rect 3758 443 3770 477
rect 3804 443 3812 477
rect 3758 371 3812 443
rect 3758 337 3770 371
rect 3804 337 3812 371
rect 3758 325 3812 337
rect 3916 477 3970 489
rect 3916 443 3924 477
rect 3958 443 3970 477
rect 3916 371 3970 443
rect 3916 337 3924 371
rect 3958 337 3970 371
rect 3916 325 3970 337
rect 4006 477 4064 489
rect 4006 443 4018 477
rect 4052 443 4064 477
rect 4006 371 4064 443
rect 4006 337 4018 371
rect 4052 337 4064 371
rect 4006 325 4064 337
rect 4100 477 4154 489
rect 4100 443 4112 477
rect 4146 443 4154 477
rect 4699 485 4753 497
rect 4100 371 4154 443
rect 4100 337 4112 371
rect 4146 337 4154 371
rect 4100 325 4154 337
rect 4219 463 4273 475
rect 4219 429 4227 463
rect 4261 429 4273 463
rect 4219 363 4273 429
rect 4219 329 4227 363
rect 4261 329 4273 363
rect 4219 311 4273 329
rect 4309 463 4367 475
rect 4309 429 4321 463
rect 4355 429 4367 463
rect 4309 357 4367 429
rect 4309 323 4321 357
rect 4355 323 4367 357
rect 4309 311 4367 323
rect 4403 463 4461 475
rect 4403 429 4415 463
rect 4449 429 4461 463
rect 4403 357 4461 429
rect 4403 323 4415 357
rect 4449 323 4461 357
rect 4403 311 4461 323
rect 4497 463 4555 475
rect 4497 429 4509 463
rect 4543 429 4555 463
rect 4497 357 4555 429
rect 4497 323 4509 357
rect 4543 323 4555 357
rect 4497 311 4555 323
rect 4591 463 4645 475
rect 4591 429 4603 463
rect 4637 429 4645 463
rect 4591 357 4645 429
rect 4591 323 4603 357
rect 4637 323 4645 357
rect 4591 311 4645 323
rect 4699 451 4707 485
rect 4741 451 4753 485
rect 4699 417 4753 451
rect 4699 383 4707 417
rect 4741 383 4753 417
rect 4699 297 4753 383
rect 4789 485 4847 497
rect 4789 451 4801 485
rect 4835 451 4847 485
rect 4789 417 4847 451
rect 4789 383 4801 417
rect 4835 383 4847 417
rect 4789 349 4847 383
rect 4789 315 4801 349
rect 4835 315 4847 349
rect 4789 297 4847 315
rect 4883 485 4941 497
rect 4883 451 4895 485
rect 4929 451 4941 485
rect 4883 417 4941 451
rect 4883 383 4895 417
rect 4929 383 4941 417
rect 4883 297 4941 383
rect 4977 485 5035 497
rect 4977 451 4989 485
rect 5023 451 5035 485
rect 4977 417 5035 451
rect 4977 383 4989 417
rect 5023 383 5035 417
rect 4977 349 5035 383
rect 4977 315 4989 349
rect 5023 315 5035 349
rect 4977 297 5035 315
rect 5071 485 5125 497
rect 5071 451 5083 485
rect 5117 451 5125 485
rect 5271 485 5325 497
rect 5071 417 5125 451
rect 5071 383 5083 417
rect 5117 383 5125 417
rect 5071 349 5125 383
rect 5071 315 5083 349
rect 5117 315 5125 349
rect 5071 297 5125 315
rect 5271 451 5279 485
rect 5313 451 5325 485
rect 5271 417 5325 451
rect 5271 383 5279 417
rect 5313 383 5325 417
rect 5271 349 5325 383
rect 5271 315 5279 349
rect 5313 315 5325 349
rect 5271 297 5325 315
rect 5361 485 5419 497
rect 5361 451 5373 485
rect 5407 451 5419 485
rect 5361 417 5419 451
rect 5361 383 5373 417
rect 5407 383 5419 417
rect 5361 349 5419 383
rect 5361 315 5373 349
rect 5407 315 5419 349
rect 5361 297 5419 315
rect 5455 485 5513 497
rect 5455 451 5467 485
rect 5501 451 5513 485
rect 5455 417 5513 451
rect 5455 383 5467 417
rect 5501 383 5513 417
rect 5455 297 5513 383
rect 5549 485 5607 497
rect 5549 451 5561 485
rect 5595 451 5607 485
rect 5549 417 5607 451
rect 5549 383 5561 417
rect 5595 383 5607 417
rect 5549 349 5607 383
rect 5549 315 5561 349
rect 5595 315 5607 349
rect 5549 297 5607 315
rect 5643 485 5697 497
rect 5643 451 5655 485
rect 5689 451 5697 485
rect 6242 477 6296 489
rect 5643 417 5697 451
rect 5643 383 5655 417
rect 5689 383 5697 417
rect 5643 297 5697 383
rect 5751 463 5805 475
rect 5751 429 5759 463
rect 5793 429 5805 463
rect 5751 357 5805 429
rect 5751 323 5759 357
rect 5793 323 5805 357
rect 5751 311 5805 323
rect 5841 463 5899 475
rect 5841 429 5853 463
rect 5887 429 5899 463
rect 5841 357 5899 429
rect 5841 323 5853 357
rect 5887 323 5899 357
rect 5841 311 5899 323
rect 5935 463 5993 475
rect 5935 429 5947 463
rect 5981 429 5993 463
rect 5935 357 5993 429
rect 5935 323 5947 357
rect 5981 323 5993 357
rect 5935 311 5993 323
rect 6029 463 6087 475
rect 6029 429 6041 463
rect 6075 429 6087 463
rect 6029 357 6087 429
rect 6029 323 6041 357
rect 6075 323 6087 357
rect 6029 311 6087 323
rect 6123 463 6177 475
rect 6123 429 6135 463
rect 6169 429 6177 463
rect 6123 363 6177 429
rect 6123 329 6135 363
rect 6169 329 6177 363
rect 6123 311 6177 329
rect 6242 443 6250 477
rect 6284 443 6296 477
rect 6242 371 6296 443
rect 6242 337 6250 371
rect 6284 337 6296 371
rect 6242 325 6296 337
rect 6332 477 6390 489
rect 6332 443 6344 477
rect 6378 443 6390 477
rect 6332 371 6390 443
rect 6332 337 6344 371
rect 6378 337 6390 371
rect 6332 325 6390 337
rect 6426 477 6480 489
rect 6426 443 6438 477
rect 6472 443 6480 477
rect 6426 371 6480 443
rect 6426 337 6438 371
rect 6472 337 6480 371
rect 6426 325 6480 337
rect 6584 477 6638 489
rect 6584 443 6592 477
rect 6626 443 6638 477
rect 6584 371 6638 443
rect 6584 337 6592 371
rect 6626 337 6638 371
rect 6584 325 6638 337
rect 6674 477 6732 489
rect 6674 443 6686 477
rect 6720 443 6732 477
rect 6674 371 6732 443
rect 6674 337 6686 371
rect 6720 337 6732 371
rect 6674 325 6732 337
rect 6768 477 6822 489
rect 6768 443 6780 477
rect 6814 443 6822 477
rect 7367 485 7421 497
rect 6768 371 6822 443
rect 6768 337 6780 371
rect 6814 337 6822 371
rect 6768 325 6822 337
rect 6887 463 6941 475
rect 6887 429 6895 463
rect 6929 429 6941 463
rect 6887 363 6941 429
rect 6887 329 6895 363
rect 6929 329 6941 363
rect 6887 311 6941 329
rect 6977 463 7035 475
rect 6977 429 6989 463
rect 7023 429 7035 463
rect 6977 357 7035 429
rect 6977 323 6989 357
rect 7023 323 7035 357
rect 6977 311 7035 323
rect 7071 463 7129 475
rect 7071 429 7083 463
rect 7117 429 7129 463
rect 7071 357 7129 429
rect 7071 323 7083 357
rect 7117 323 7129 357
rect 7071 311 7129 323
rect 7165 463 7223 475
rect 7165 429 7177 463
rect 7211 429 7223 463
rect 7165 357 7223 429
rect 7165 323 7177 357
rect 7211 323 7223 357
rect 7165 311 7223 323
rect 7259 463 7313 475
rect 7259 429 7271 463
rect 7305 429 7313 463
rect 7259 357 7313 429
rect 7259 323 7271 357
rect 7305 323 7313 357
rect 7259 311 7313 323
rect 7367 451 7375 485
rect 7409 451 7421 485
rect 7367 417 7421 451
rect 7367 383 7375 417
rect 7409 383 7421 417
rect 7367 297 7421 383
rect 7457 485 7515 497
rect 7457 451 7469 485
rect 7503 451 7515 485
rect 7457 417 7515 451
rect 7457 383 7469 417
rect 7503 383 7515 417
rect 7457 349 7515 383
rect 7457 315 7469 349
rect 7503 315 7515 349
rect 7457 297 7515 315
rect 7551 485 7609 497
rect 7551 451 7563 485
rect 7597 451 7609 485
rect 7551 417 7609 451
rect 7551 383 7563 417
rect 7597 383 7609 417
rect 7551 297 7609 383
rect 7645 485 7703 497
rect 7645 451 7657 485
rect 7691 451 7703 485
rect 7645 417 7703 451
rect 7645 383 7657 417
rect 7691 383 7703 417
rect 7645 349 7703 383
rect 7645 315 7657 349
rect 7691 315 7703 349
rect 7645 297 7703 315
rect 7739 485 7793 497
rect 7739 451 7751 485
rect 7785 451 7793 485
rect 7739 417 7793 451
rect 7739 383 7751 417
rect 7785 383 7793 417
rect 7739 349 7793 383
rect 7739 315 7751 349
rect 7785 315 7793 349
rect 7739 297 7793 315
rect 7847 485 7901 497
rect 7847 451 7855 485
rect 7889 451 7901 485
rect 7847 417 7901 451
rect 7847 383 7855 417
rect 7889 383 7901 417
rect 7847 349 7901 383
rect 7847 315 7855 349
rect 7889 315 7901 349
rect 7847 297 7901 315
rect 7937 485 7995 497
rect 7937 451 7949 485
rect 7983 451 7995 485
rect 7937 417 7995 451
rect 7937 383 7949 417
rect 7983 383 7995 417
rect 7937 349 7995 383
rect 7937 315 7949 349
rect 7983 315 7995 349
rect 7937 297 7995 315
rect 8031 485 8089 497
rect 8031 451 8043 485
rect 8077 451 8089 485
rect 8031 417 8089 451
rect 8031 383 8043 417
rect 8077 383 8089 417
rect 8031 297 8089 383
rect 8125 485 8183 497
rect 8125 451 8137 485
rect 8171 451 8183 485
rect 8125 417 8183 451
rect 8125 383 8137 417
rect 8171 383 8183 417
rect 8125 349 8183 383
rect 8125 315 8137 349
rect 8171 315 8183 349
rect 8125 297 8183 315
rect 8219 485 8273 497
rect 8219 451 8231 485
rect 8265 451 8273 485
rect 8818 477 8872 489
rect 8219 417 8273 451
rect 8219 383 8231 417
rect 8265 383 8273 417
rect 8219 297 8273 383
rect 8327 463 8381 475
rect 8327 429 8335 463
rect 8369 429 8381 463
rect 8327 357 8381 429
rect 8327 323 8335 357
rect 8369 323 8381 357
rect 8327 311 8381 323
rect 8417 463 8475 475
rect 8417 429 8429 463
rect 8463 429 8475 463
rect 8417 357 8475 429
rect 8417 323 8429 357
rect 8463 323 8475 357
rect 8417 311 8475 323
rect 8511 463 8569 475
rect 8511 429 8523 463
rect 8557 429 8569 463
rect 8511 357 8569 429
rect 8511 323 8523 357
rect 8557 323 8569 357
rect 8511 311 8569 323
rect 8605 463 8663 475
rect 8605 429 8617 463
rect 8651 429 8663 463
rect 8605 357 8663 429
rect 8605 323 8617 357
rect 8651 323 8663 357
rect 8605 311 8663 323
rect 8699 463 8753 475
rect 8699 429 8711 463
rect 8745 429 8753 463
rect 8699 363 8753 429
rect 8699 329 8711 363
rect 8745 329 8753 363
rect 8699 311 8753 329
rect 8818 443 8826 477
rect 8860 443 8872 477
rect 8818 371 8872 443
rect 8818 337 8826 371
rect 8860 337 8872 371
rect 8818 325 8872 337
rect 8908 477 8966 489
rect 8908 443 8920 477
rect 8954 443 8966 477
rect 8908 371 8966 443
rect 8908 337 8920 371
rect 8954 337 8966 371
rect 8908 325 8966 337
rect 9002 477 9056 489
rect 9002 443 9014 477
rect 9048 443 9056 477
rect 9002 371 9056 443
rect 9002 337 9014 371
rect 9048 337 9056 371
rect 9002 325 9056 337
rect 9160 477 9214 489
rect 9160 443 9168 477
rect 9202 443 9214 477
rect 9160 371 9214 443
rect 9160 337 9168 371
rect 9202 337 9214 371
rect 9160 325 9214 337
rect 9250 477 9308 489
rect 9250 443 9262 477
rect 9296 443 9308 477
rect 9250 371 9308 443
rect 9250 337 9262 371
rect 9296 337 9308 371
rect 9250 325 9308 337
rect 9344 477 9398 489
rect 9344 443 9356 477
rect 9390 443 9398 477
rect 9943 485 9997 497
rect 9344 371 9398 443
rect 9344 337 9356 371
rect 9390 337 9398 371
rect 9344 325 9398 337
rect 9463 463 9517 475
rect 9463 429 9471 463
rect 9505 429 9517 463
rect 9463 363 9517 429
rect 9463 329 9471 363
rect 9505 329 9517 363
rect 9463 311 9517 329
rect 9553 463 9611 475
rect 9553 429 9565 463
rect 9599 429 9611 463
rect 9553 357 9611 429
rect 9553 323 9565 357
rect 9599 323 9611 357
rect 9553 311 9611 323
rect 9647 463 9705 475
rect 9647 429 9659 463
rect 9693 429 9705 463
rect 9647 357 9705 429
rect 9647 323 9659 357
rect 9693 323 9705 357
rect 9647 311 9705 323
rect 9741 463 9799 475
rect 9741 429 9753 463
rect 9787 429 9799 463
rect 9741 357 9799 429
rect 9741 323 9753 357
rect 9787 323 9799 357
rect 9741 311 9799 323
rect 9835 463 9889 475
rect 9835 429 9847 463
rect 9881 429 9889 463
rect 9835 357 9889 429
rect 9835 323 9847 357
rect 9881 323 9889 357
rect 9835 311 9889 323
rect 9943 451 9951 485
rect 9985 451 9997 485
rect 9943 417 9997 451
rect 9943 383 9951 417
rect 9985 383 9997 417
rect 9943 297 9997 383
rect 10033 485 10091 497
rect 10033 451 10045 485
rect 10079 451 10091 485
rect 10033 417 10091 451
rect 10033 383 10045 417
rect 10079 383 10091 417
rect 10033 349 10091 383
rect 10033 315 10045 349
rect 10079 315 10091 349
rect 10033 297 10091 315
rect 10127 485 10185 497
rect 10127 451 10139 485
rect 10173 451 10185 485
rect 10127 417 10185 451
rect 10127 383 10139 417
rect 10173 383 10185 417
rect 10127 297 10185 383
rect 10221 485 10279 497
rect 10221 451 10233 485
rect 10267 451 10279 485
rect 10221 417 10279 451
rect 10221 383 10233 417
rect 10267 383 10279 417
rect 10221 349 10279 383
rect 10221 315 10233 349
rect 10267 315 10279 349
rect 10221 297 10279 315
rect 10315 485 10369 497
rect 10315 451 10327 485
rect 10361 451 10369 485
rect 10315 417 10369 451
rect 10315 383 10327 417
rect 10361 383 10369 417
rect 10315 349 10369 383
rect 10315 315 10327 349
rect 10361 315 10369 349
rect 10315 297 10369 315
<< ndiffc >>
rect 45 995 79 1029
rect 45 927 79 961
rect 129 995 163 1029
rect 129 927 163 961
rect 223 995 257 1029
rect 317 995 351 1029
rect 317 927 351 961
rect 401 995 435 1029
rect 505 953 539 987
rect 589 935 623 969
rect 673 953 707 987
rect 757 935 791 969
rect 841 953 875 987
rect 1016 982 1050 1016
rect 1100 982 1134 1016
rect 1184 982 1218 1016
rect 1358 982 1392 1016
rect 1442 982 1476 1016
rect 1526 982 1560 1016
rect 1701 953 1735 987
rect 1785 935 1819 969
rect 1869 953 1903 987
rect 1953 935 1987 969
rect 2037 953 2071 987
rect 2141 995 2175 1029
rect 2225 995 2259 1029
rect 2225 927 2259 961
rect 2319 995 2353 1029
rect 2413 995 2447 1029
rect 2413 927 2447 961
rect 2497 995 2531 1029
rect 2497 927 2531 961
rect 2621 995 2655 1029
rect 2621 927 2655 961
rect 2705 995 2739 1029
rect 2705 927 2739 961
rect 2799 995 2833 1029
rect 2893 995 2927 1029
rect 2893 927 2927 961
rect 2977 995 3011 1029
rect 3081 953 3115 987
rect 3165 935 3199 969
rect 3249 953 3283 987
rect 3333 935 3367 969
rect 3417 953 3451 987
rect 3592 982 3626 1016
rect 3676 982 3710 1016
rect 3760 982 3794 1016
rect 3934 982 3968 1016
rect 4018 982 4052 1016
rect 4102 982 4136 1016
rect 4277 953 4311 987
rect 4361 935 4395 969
rect 4445 953 4479 987
rect 4529 935 4563 969
rect 4613 953 4647 987
rect 4717 995 4751 1029
rect 4801 995 4835 1029
rect 4801 927 4835 961
rect 4895 995 4929 1029
rect 4989 995 5023 1029
rect 4989 927 5023 961
rect 5073 995 5107 1029
rect 5073 927 5107 961
rect 5289 995 5323 1029
rect 5289 927 5323 961
rect 5373 995 5407 1029
rect 5373 927 5407 961
rect 5467 995 5501 1029
rect 5561 995 5595 1029
rect 5561 927 5595 961
rect 5645 995 5679 1029
rect 5749 953 5783 987
rect 5833 935 5867 969
rect 5917 953 5951 987
rect 6001 935 6035 969
rect 6085 953 6119 987
rect 6260 982 6294 1016
rect 6344 982 6378 1016
rect 6428 982 6462 1016
rect 6602 982 6636 1016
rect 6686 982 6720 1016
rect 6770 982 6804 1016
rect 6945 953 6979 987
rect 7029 935 7063 969
rect 7113 953 7147 987
rect 7197 935 7231 969
rect 7281 953 7315 987
rect 7385 995 7419 1029
rect 7469 995 7503 1029
rect 7469 927 7503 961
rect 7563 995 7597 1029
rect 7657 995 7691 1029
rect 7657 927 7691 961
rect 7741 995 7775 1029
rect 7741 927 7775 961
rect 7865 995 7899 1029
rect 7865 927 7899 961
rect 7949 995 7983 1029
rect 7949 927 7983 961
rect 8043 995 8077 1029
rect 8137 995 8171 1029
rect 8137 927 8171 961
rect 8221 995 8255 1029
rect 8325 953 8359 987
rect 8409 935 8443 969
rect 8493 953 8527 987
rect 8577 935 8611 969
rect 8661 953 8695 987
rect 8836 982 8870 1016
rect 8920 982 8954 1016
rect 9004 982 9038 1016
rect 9178 982 9212 1016
rect 9262 982 9296 1016
rect 9346 982 9380 1016
rect 9521 953 9555 987
rect 9605 935 9639 969
rect 9689 953 9723 987
rect 9773 935 9807 969
rect 9857 953 9891 987
rect 9961 995 9995 1029
rect 10045 995 10079 1029
rect 10045 927 10079 961
rect 10139 995 10173 1029
rect 10233 995 10267 1029
rect 10233 927 10267 961
rect 10317 995 10351 1029
rect 10317 927 10351 961
rect 45 127 79 161
rect 45 59 79 93
rect 129 127 163 161
rect 129 59 163 93
rect 223 59 257 93
rect 317 127 351 161
rect 317 59 351 93
rect 401 59 435 93
rect 505 101 539 135
rect 589 119 623 153
rect 673 101 707 135
rect 757 119 791 153
rect 841 101 875 135
rect 1016 72 1050 106
rect 1100 72 1134 106
rect 1184 72 1218 106
rect 1358 72 1392 106
rect 1442 72 1476 106
rect 1526 72 1560 106
rect 1701 101 1735 135
rect 1785 119 1819 153
rect 1869 101 1903 135
rect 1953 119 1987 153
rect 2037 101 2071 135
rect 2141 59 2175 93
rect 2225 127 2259 161
rect 2225 59 2259 93
rect 2319 59 2353 93
rect 2413 127 2447 161
rect 2413 59 2447 93
rect 2497 127 2531 161
rect 2497 59 2531 93
rect 2621 127 2655 161
rect 2621 59 2655 93
rect 2705 127 2739 161
rect 2705 59 2739 93
rect 2799 59 2833 93
rect 2893 127 2927 161
rect 2893 59 2927 93
rect 2977 59 3011 93
rect 3081 101 3115 135
rect 3165 119 3199 153
rect 3249 101 3283 135
rect 3333 119 3367 153
rect 3417 101 3451 135
rect 3592 72 3626 106
rect 3676 72 3710 106
rect 3760 72 3794 106
rect 3934 72 3968 106
rect 4018 72 4052 106
rect 4102 72 4136 106
rect 4277 101 4311 135
rect 4361 119 4395 153
rect 4445 101 4479 135
rect 4529 119 4563 153
rect 4613 101 4647 135
rect 4717 59 4751 93
rect 4801 127 4835 161
rect 4801 59 4835 93
rect 4895 59 4929 93
rect 4989 127 5023 161
rect 4989 59 5023 93
rect 5073 127 5107 161
rect 5073 59 5107 93
rect 5289 127 5323 161
rect 5289 59 5323 93
rect 5373 127 5407 161
rect 5373 59 5407 93
rect 5467 59 5501 93
rect 5561 127 5595 161
rect 5561 59 5595 93
rect 5645 59 5679 93
rect 5749 101 5783 135
rect 5833 119 5867 153
rect 5917 101 5951 135
rect 6001 119 6035 153
rect 6085 101 6119 135
rect 6260 72 6294 106
rect 6344 72 6378 106
rect 6428 72 6462 106
rect 6602 72 6636 106
rect 6686 72 6720 106
rect 6770 72 6804 106
rect 6945 101 6979 135
rect 7029 119 7063 153
rect 7113 101 7147 135
rect 7197 119 7231 153
rect 7281 101 7315 135
rect 7385 59 7419 93
rect 7469 127 7503 161
rect 7469 59 7503 93
rect 7563 59 7597 93
rect 7657 127 7691 161
rect 7657 59 7691 93
rect 7741 127 7775 161
rect 7741 59 7775 93
rect 7865 127 7899 161
rect 7865 59 7899 93
rect 7949 127 7983 161
rect 7949 59 7983 93
rect 8043 59 8077 93
rect 8137 127 8171 161
rect 8137 59 8171 93
rect 8221 59 8255 93
rect 8325 101 8359 135
rect 8409 119 8443 153
rect 8493 101 8527 135
rect 8577 119 8611 153
rect 8661 101 8695 135
rect 8836 72 8870 106
rect 8920 72 8954 106
rect 9004 72 9038 106
rect 9178 72 9212 106
rect 9262 72 9296 106
rect 9346 72 9380 106
rect 9521 101 9555 135
rect 9605 119 9639 153
rect 9689 101 9723 135
rect 9773 119 9807 153
rect 9857 101 9891 135
rect 9961 59 9995 93
rect 10045 127 10079 161
rect 10045 59 10079 93
rect 10139 59 10173 93
rect 10233 127 10267 161
rect 10233 59 10267 93
rect 10317 127 10351 161
rect 10317 59 10351 93
<< pdiffc >>
rect 35 739 69 773
rect 35 671 69 705
rect 35 603 69 637
rect 129 739 163 773
rect 129 671 163 705
rect 129 603 163 637
rect 223 671 257 705
rect 223 603 257 637
rect 317 739 351 773
rect 317 671 351 705
rect 317 603 351 637
rect 411 671 445 705
rect 411 603 445 637
rect 515 731 549 765
rect 515 625 549 659
rect 609 731 643 765
rect 609 625 643 659
rect 703 731 737 765
rect 703 625 737 659
rect 797 731 831 765
rect 797 625 831 659
rect 891 725 925 759
rect 891 625 925 659
rect 1006 717 1040 751
rect 1006 611 1040 645
rect 1100 717 1134 751
rect 1100 611 1134 645
rect 1194 717 1228 751
rect 1194 611 1228 645
rect 1348 717 1382 751
rect 1348 611 1382 645
rect 1442 717 1476 751
rect 1442 611 1476 645
rect 1536 717 1570 751
rect 1536 611 1570 645
rect 1651 725 1685 759
rect 1651 625 1685 659
rect 1745 731 1779 765
rect 1745 625 1779 659
rect 1839 731 1873 765
rect 1839 625 1873 659
rect 1933 731 1967 765
rect 1933 625 1967 659
rect 2027 731 2061 765
rect 2027 625 2061 659
rect 2131 671 2165 705
rect 2131 603 2165 637
rect 2225 739 2259 773
rect 2225 671 2259 705
rect 2225 603 2259 637
rect 2319 671 2353 705
rect 2319 603 2353 637
rect 2413 739 2447 773
rect 2413 671 2447 705
rect 2413 603 2447 637
rect 2507 739 2541 773
rect 2507 671 2541 705
rect 2507 603 2541 637
rect 2611 739 2645 773
rect 2611 671 2645 705
rect 2611 603 2645 637
rect 2705 739 2739 773
rect 2705 671 2739 705
rect 2705 603 2739 637
rect 2799 671 2833 705
rect 2799 603 2833 637
rect 2893 739 2927 773
rect 2893 671 2927 705
rect 2893 603 2927 637
rect 2987 671 3021 705
rect 2987 603 3021 637
rect 3091 731 3125 765
rect 3091 625 3125 659
rect 3185 731 3219 765
rect 3185 625 3219 659
rect 3279 731 3313 765
rect 3279 625 3313 659
rect 3373 731 3407 765
rect 3373 625 3407 659
rect 3467 725 3501 759
rect 3467 625 3501 659
rect 3582 717 3616 751
rect 3582 611 3616 645
rect 3676 717 3710 751
rect 3676 611 3710 645
rect 3770 717 3804 751
rect 3770 611 3804 645
rect 3924 717 3958 751
rect 3924 611 3958 645
rect 4018 717 4052 751
rect 4018 611 4052 645
rect 4112 717 4146 751
rect 4112 611 4146 645
rect 4227 725 4261 759
rect 4227 625 4261 659
rect 4321 731 4355 765
rect 4321 625 4355 659
rect 4415 731 4449 765
rect 4415 625 4449 659
rect 4509 731 4543 765
rect 4509 625 4543 659
rect 4603 731 4637 765
rect 4603 625 4637 659
rect 4707 671 4741 705
rect 4707 603 4741 637
rect 4801 739 4835 773
rect 4801 671 4835 705
rect 4801 603 4835 637
rect 4895 671 4929 705
rect 4895 603 4929 637
rect 4989 739 5023 773
rect 4989 671 5023 705
rect 4989 603 5023 637
rect 5083 739 5117 773
rect 5083 671 5117 705
rect 5083 603 5117 637
rect 5279 739 5313 773
rect 5279 671 5313 705
rect 5279 603 5313 637
rect 5373 739 5407 773
rect 5373 671 5407 705
rect 5373 603 5407 637
rect 5467 671 5501 705
rect 5467 603 5501 637
rect 5561 739 5595 773
rect 5561 671 5595 705
rect 5561 603 5595 637
rect 5655 671 5689 705
rect 5655 603 5689 637
rect 5759 731 5793 765
rect 5759 625 5793 659
rect 5853 731 5887 765
rect 5853 625 5887 659
rect 5947 731 5981 765
rect 5947 625 5981 659
rect 6041 731 6075 765
rect 6041 625 6075 659
rect 6135 725 6169 759
rect 6135 625 6169 659
rect 6250 717 6284 751
rect 6250 611 6284 645
rect 6344 717 6378 751
rect 6344 611 6378 645
rect 6438 717 6472 751
rect 6438 611 6472 645
rect 6592 717 6626 751
rect 6592 611 6626 645
rect 6686 717 6720 751
rect 6686 611 6720 645
rect 6780 717 6814 751
rect 6780 611 6814 645
rect 6895 725 6929 759
rect 6895 625 6929 659
rect 6989 731 7023 765
rect 6989 625 7023 659
rect 7083 731 7117 765
rect 7083 625 7117 659
rect 7177 731 7211 765
rect 7177 625 7211 659
rect 7271 731 7305 765
rect 7271 625 7305 659
rect 7375 671 7409 705
rect 7375 603 7409 637
rect 7469 739 7503 773
rect 7469 671 7503 705
rect 7469 603 7503 637
rect 7563 671 7597 705
rect 7563 603 7597 637
rect 7657 739 7691 773
rect 7657 671 7691 705
rect 7657 603 7691 637
rect 7751 739 7785 773
rect 7751 671 7785 705
rect 7751 603 7785 637
rect 7855 739 7889 773
rect 7855 671 7889 705
rect 7855 603 7889 637
rect 7949 739 7983 773
rect 7949 671 7983 705
rect 7949 603 7983 637
rect 8043 671 8077 705
rect 8043 603 8077 637
rect 8137 739 8171 773
rect 8137 671 8171 705
rect 8137 603 8171 637
rect 8231 671 8265 705
rect 8231 603 8265 637
rect 8335 731 8369 765
rect 8335 625 8369 659
rect 8429 731 8463 765
rect 8429 625 8463 659
rect 8523 731 8557 765
rect 8523 625 8557 659
rect 8617 731 8651 765
rect 8617 625 8651 659
rect 8711 725 8745 759
rect 8711 625 8745 659
rect 8826 717 8860 751
rect 8826 611 8860 645
rect 8920 717 8954 751
rect 8920 611 8954 645
rect 9014 717 9048 751
rect 9014 611 9048 645
rect 9168 717 9202 751
rect 9168 611 9202 645
rect 9262 717 9296 751
rect 9262 611 9296 645
rect 9356 717 9390 751
rect 9356 611 9390 645
rect 9471 725 9505 759
rect 9471 625 9505 659
rect 9565 731 9599 765
rect 9565 625 9599 659
rect 9659 731 9693 765
rect 9659 625 9693 659
rect 9753 731 9787 765
rect 9753 625 9787 659
rect 9847 731 9881 765
rect 9847 625 9881 659
rect 9951 671 9985 705
rect 9951 603 9985 637
rect 10045 739 10079 773
rect 10045 671 10079 705
rect 10045 603 10079 637
rect 10139 671 10173 705
rect 10139 603 10173 637
rect 10233 739 10267 773
rect 10233 671 10267 705
rect 10233 603 10267 637
rect 10327 739 10361 773
rect 10327 671 10361 705
rect 10327 603 10361 637
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 451 163 485
rect 129 383 163 417
rect 129 315 163 349
rect 223 451 257 485
rect 223 383 257 417
rect 317 451 351 485
rect 317 383 351 417
rect 317 315 351 349
rect 411 451 445 485
rect 411 383 445 417
rect 515 429 549 463
rect 515 323 549 357
rect 609 429 643 463
rect 609 323 643 357
rect 703 429 737 463
rect 703 323 737 357
rect 797 429 831 463
rect 797 323 831 357
rect 891 429 925 463
rect 891 329 925 363
rect 1006 443 1040 477
rect 1006 337 1040 371
rect 1100 443 1134 477
rect 1100 337 1134 371
rect 1194 443 1228 477
rect 1194 337 1228 371
rect 1348 443 1382 477
rect 1348 337 1382 371
rect 1442 443 1476 477
rect 1442 337 1476 371
rect 1536 443 1570 477
rect 1536 337 1570 371
rect 1651 429 1685 463
rect 1651 329 1685 363
rect 1745 429 1779 463
rect 1745 323 1779 357
rect 1839 429 1873 463
rect 1839 323 1873 357
rect 1933 429 1967 463
rect 1933 323 1967 357
rect 2027 429 2061 463
rect 2027 323 2061 357
rect 2131 451 2165 485
rect 2131 383 2165 417
rect 2225 451 2259 485
rect 2225 383 2259 417
rect 2225 315 2259 349
rect 2319 451 2353 485
rect 2319 383 2353 417
rect 2413 451 2447 485
rect 2413 383 2447 417
rect 2413 315 2447 349
rect 2507 451 2541 485
rect 2507 383 2541 417
rect 2507 315 2541 349
rect 2611 451 2645 485
rect 2611 383 2645 417
rect 2611 315 2645 349
rect 2705 451 2739 485
rect 2705 383 2739 417
rect 2705 315 2739 349
rect 2799 451 2833 485
rect 2799 383 2833 417
rect 2893 451 2927 485
rect 2893 383 2927 417
rect 2893 315 2927 349
rect 2987 451 3021 485
rect 2987 383 3021 417
rect 3091 429 3125 463
rect 3091 323 3125 357
rect 3185 429 3219 463
rect 3185 323 3219 357
rect 3279 429 3313 463
rect 3279 323 3313 357
rect 3373 429 3407 463
rect 3373 323 3407 357
rect 3467 429 3501 463
rect 3467 329 3501 363
rect 3582 443 3616 477
rect 3582 337 3616 371
rect 3676 443 3710 477
rect 3676 337 3710 371
rect 3770 443 3804 477
rect 3770 337 3804 371
rect 3924 443 3958 477
rect 3924 337 3958 371
rect 4018 443 4052 477
rect 4018 337 4052 371
rect 4112 443 4146 477
rect 4112 337 4146 371
rect 4227 429 4261 463
rect 4227 329 4261 363
rect 4321 429 4355 463
rect 4321 323 4355 357
rect 4415 429 4449 463
rect 4415 323 4449 357
rect 4509 429 4543 463
rect 4509 323 4543 357
rect 4603 429 4637 463
rect 4603 323 4637 357
rect 4707 451 4741 485
rect 4707 383 4741 417
rect 4801 451 4835 485
rect 4801 383 4835 417
rect 4801 315 4835 349
rect 4895 451 4929 485
rect 4895 383 4929 417
rect 4989 451 5023 485
rect 4989 383 5023 417
rect 4989 315 5023 349
rect 5083 451 5117 485
rect 5083 383 5117 417
rect 5083 315 5117 349
rect 5279 451 5313 485
rect 5279 383 5313 417
rect 5279 315 5313 349
rect 5373 451 5407 485
rect 5373 383 5407 417
rect 5373 315 5407 349
rect 5467 451 5501 485
rect 5467 383 5501 417
rect 5561 451 5595 485
rect 5561 383 5595 417
rect 5561 315 5595 349
rect 5655 451 5689 485
rect 5655 383 5689 417
rect 5759 429 5793 463
rect 5759 323 5793 357
rect 5853 429 5887 463
rect 5853 323 5887 357
rect 5947 429 5981 463
rect 5947 323 5981 357
rect 6041 429 6075 463
rect 6041 323 6075 357
rect 6135 429 6169 463
rect 6135 329 6169 363
rect 6250 443 6284 477
rect 6250 337 6284 371
rect 6344 443 6378 477
rect 6344 337 6378 371
rect 6438 443 6472 477
rect 6438 337 6472 371
rect 6592 443 6626 477
rect 6592 337 6626 371
rect 6686 443 6720 477
rect 6686 337 6720 371
rect 6780 443 6814 477
rect 6780 337 6814 371
rect 6895 429 6929 463
rect 6895 329 6929 363
rect 6989 429 7023 463
rect 6989 323 7023 357
rect 7083 429 7117 463
rect 7083 323 7117 357
rect 7177 429 7211 463
rect 7177 323 7211 357
rect 7271 429 7305 463
rect 7271 323 7305 357
rect 7375 451 7409 485
rect 7375 383 7409 417
rect 7469 451 7503 485
rect 7469 383 7503 417
rect 7469 315 7503 349
rect 7563 451 7597 485
rect 7563 383 7597 417
rect 7657 451 7691 485
rect 7657 383 7691 417
rect 7657 315 7691 349
rect 7751 451 7785 485
rect 7751 383 7785 417
rect 7751 315 7785 349
rect 7855 451 7889 485
rect 7855 383 7889 417
rect 7855 315 7889 349
rect 7949 451 7983 485
rect 7949 383 7983 417
rect 7949 315 7983 349
rect 8043 451 8077 485
rect 8043 383 8077 417
rect 8137 451 8171 485
rect 8137 383 8171 417
rect 8137 315 8171 349
rect 8231 451 8265 485
rect 8231 383 8265 417
rect 8335 429 8369 463
rect 8335 323 8369 357
rect 8429 429 8463 463
rect 8429 323 8463 357
rect 8523 429 8557 463
rect 8523 323 8557 357
rect 8617 429 8651 463
rect 8617 323 8651 357
rect 8711 429 8745 463
rect 8711 329 8745 363
rect 8826 443 8860 477
rect 8826 337 8860 371
rect 8920 443 8954 477
rect 8920 337 8954 371
rect 9014 443 9048 477
rect 9014 337 9048 371
rect 9168 443 9202 477
rect 9168 337 9202 371
rect 9262 443 9296 477
rect 9262 337 9296 371
rect 9356 443 9390 477
rect 9356 337 9390 371
rect 9471 429 9505 463
rect 9471 329 9505 363
rect 9565 429 9599 463
rect 9565 323 9599 357
rect 9659 429 9693 463
rect 9659 323 9693 357
rect 9753 429 9787 463
rect 9753 323 9787 357
rect 9847 429 9881 463
rect 9847 323 9881 357
rect 9951 451 9985 485
rect 9951 383 9985 417
rect 10045 451 10079 485
rect 10045 383 10079 417
rect 10045 315 10079 349
rect 10139 451 10173 485
rect 10139 383 10173 417
rect 10233 451 10267 485
rect 10233 383 10267 417
rect 10233 315 10267 349
rect 10327 451 10361 485
rect 10327 383 10361 417
rect 10327 315 10361 349
<< psubdiff >>
rect 5181 977 5215 1024
rect 5181 919 5215 943
rect 5181 145 5215 169
rect 5181 64 5215 111
<< nsubdiff >>
rect 5181 759 5215 783
rect 5181 675 5215 725
rect 5181 608 5215 641
rect 5181 447 5215 480
rect 5181 363 5215 413
rect 5181 305 5215 329
<< psubdiffcont >>
rect 5181 943 5215 977
rect 5181 111 5215 145
<< nsubdiffcont >>
rect 5181 725 5215 759
rect 5181 641 5215 675
rect 5181 413 5215 447
rect 5181 329 5215 363
<< poly >>
rect 89 1041 119 1069
rect 173 1041 203 1067
rect 277 1041 307 1069
rect 361 1041 391 1067
rect 549 1037 983 1067
rect 1060 1041 1090 1067
rect 1144 1041 1174 1067
rect 1402 1041 1432 1067
rect 1486 1041 1516 1067
rect 549 1022 579 1037
rect 633 1022 663 1037
rect 717 1022 747 1037
rect 801 1022 831 1037
rect 953 941 983 1037
rect 1593 1037 2027 1067
rect 2185 1041 2215 1067
rect 2269 1041 2299 1069
rect 2373 1041 2403 1067
rect 2457 1041 2487 1069
rect 2665 1041 2695 1069
rect 2749 1041 2779 1067
rect 2853 1041 2883 1069
rect 2937 1041 2967 1067
rect 1060 941 1090 957
rect 1144 941 1174 957
rect 89 883 119 911
rect 173 883 203 911
rect 277 883 307 911
rect 361 883 391 911
rect 549 892 579 918
rect 633 892 663 918
rect 717 892 747 918
rect 801 892 831 918
rect 953 911 1174 941
rect 79 873 401 883
rect 79 839 103 873
rect 137 839 171 873
rect 205 839 239 873
rect 273 839 307 873
rect 341 839 401 873
rect 79 829 401 839
rect 874 859 1008 869
rect 81 791 117 829
rect 175 791 211 829
rect 269 791 305 829
rect 363 791 399 829
rect 874 825 890 859
rect 924 825 958 859
rect 992 825 1008 859
rect 874 823 1008 825
rect 559 815 1008 823
rect 559 793 925 815
rect 561 777 597 793
rect 655 777 691 793
rect 749 777 785 793
rect 843 777 879 793
rect 1050 778 1090 911
rect 1144 889 1174 911
rect 1402 941 1432 957
rect 1486 941 1516 957
rect 1593 941 1623 1037
rect 1745 1022 1775 1037
rect 1829 1022 1859 1037
rect 1913 1022 1943 1037
rect 1997 1022 2027 1037
rect 1402 911 1623 941
rect 1402 889 1432 911
rect 1144 873 1267 889
rect 1144 839 1155 873
rect 1189 839 1223 873
rect 1257 839 1267 873
rect 1144 823 1267 839
rect 1309 873 1432 889
rect 1309 839 1319 873
rect 1353 839 1387 873
rect 1421 839 1432 873
rect 1309 823 1432 839
rect 1144 778 1184 823
rect 1392 778 1432 823
rect 1486 778 1526 911
rect 1745 892 1775 918
rect 1829 892 1859 918
rect 1913 892 1943 918
rect 1997 892 2027 918
rect 3125 1037 3559 1067
rect 3636 1041 3666 1067
rect 3720 1041 3750 1067
rect 3978 1041 4008 1067
rect 4062 1041 4092 1067
rect 3125 1022 3155 1037
rect 3209 1022 3239 1037
rect 3293 1022 3323 1037
rect 3377 1022 3407 1037
rect 3529 941 3559 1037
rect 4169 1037 4603 1067
rect 4761 1041 4791 1067
rect 4845 1041 4875 1069
rect 4949 1041 4979 1067
rect 5033 1041 5063 1069
rect 5333 1041 5363 1069
rect 5417 1041 5447 1067
rect 5521 1041 5551 1069
rect 5605 1041 5635 1067
rect 3636 941 3666 957
rect 3720 941 3750 957
rect 2185 883 2215 911
rect 2269 883 2299 911
rect 2373 883 2403 911
rect 2457 883 2487 911
rect 2665 883 2695 911
rect 2749 883 2779 911
rect 2853 883 2883 911
rect 2937 883 2967 911
rect 3125 892 3155 918
rect 3209 892 3239 918
rect 3293 892 3323 918
rect 3377 892 3407 918
rect 3529 911 3750 941
rect 2175 873 2497 883
rect 1568 859 1702 869
rect 1568 825 1584 859
rect 1618 825 1652 859
rect 1686 825 1702 859
rect 2175 839 2235 873
rect 2269 839 2303 873
rect 2337 839 2371 873
rect 2405 839 2439 873
rect 2473 839 2497 873
rect 2175 829 2497 839
rect 2655 873 2977 883
rect 2655 839 2679 873
rect 2713 839 2747 873
rect 2781 839 2815 873
rect 2849 839 2883 873
rect 2917 839 2977 873
rect 2655 829 2977 839
rect 3450 859 3584 869
rect 1568 823 1702 825
rect 1568 815 2017 823
rect 1651 793 2017 815
rect 1052 763 1088 778
rect 1146 763 1182 778
rect 1394 763 1430 778
rect 1488 763 1524 778
rect 1697 777 1733 793
rect 1791 777 1827 793
rect 1885 777 1921 793
rect 1979 777 2015 793
rect 2177 791 2213 829
rect 2271 791 2307 829
rect 2365 791 2401 829
rect 2459 791 2495 829
rect 2657 791 2693 829
rect 2751 791 2787 829
rect 2845 791 2881 829
rect 2939 791 2975 829
rect 3450 825 3466 859
rect 3500 825 3534 859
rect 3568 825 3584 859
rect 3450 823 3584 825
rect 3135 815 3584 823
rect 3135 793 3501 815
rect 81 565 117 591
rect 175 565 211 591
rect 269 565 305 591
rect 363 565 399 591
rect 561 565 597 613
rect 655 565 691 613
rect 749 565 785 613
rect 843 565 879 613
rect 1052 565 1088 599
rect 1146 565 1182 599
rect 1394 565 1430 599
rect 1488 565 1524 599
rect 1697 565 1733 613
rect 1791 565 1827 613
rect 1885 565 1921 613
rect 1979 565 2015 613
rect 3137 777 3173 793
rect 3231 777 3267 793
rect 3325 777 3361 793
rect 3419 777 3455 793
rect 3626 778 3666 911
rect 3720 889 3750 911
rect 3978 941 4008 957
rect 4062 941 4092 957
rect 4169 941 4199 1037
rect 4321 1022 4351 1037
rect 4405 1022 4435 1037
rect 4489 1022 4519 1037
rect 4573 1022 4603 1037
rect 3978 911 4199 941
rect 3978 889 4008 911
rect 3720 873 3843 889
rect 3720 839 3731 873
rect 3765 839 3799 873
rect 3833 839 3843 873
rect 3720 823 3843 839
rect 3885 873 4008 889
rect 3885 839 3895 873
rect 3929 839 3963 873
rect 3997 839 4008 873
rect 3885 823 4008 839
rect 3720 778 3760 823
rect 3968 778 4008 823
rect 4062 778 4102 911
rect 4321 892 4351 918
rect 4405 892 4435 918
rect 4489 892 4519 918
rect 4573 892 4603 918
rect 5793 1037 6227 1067
rect 6304 1041 6334 1067
rect 6388 1041 6418 1067
rect 6646 1041 6676 1067
rect 6730 1041 6760 1067
rect 5793 1022 5823 1037
rect 5877 1022 5907 1037
rect 5961 1022 5991 1037
rect 6045 1022 6075 1037
rect 6197 941 6227 1037
rect 6837 1037 7271 1067
rect 7429 1041 7459 1067
rect 7513 1041 7543 1069
rect 7617 1041 7647 1067
rect 7701 1041 7731 1069
rect 7909 1041 7939 1069
rect 7993 1041 8023 1067
rect 8097 1041 8127 1069
rect 8181 1041 8211 1067
rect 6304 941 6334 957
rect 6388 941 6418 957
rect 4761 883 4791 911
rect 4845 883 4875 911
rect 4949 883 4979 911
rect 5033 883 5063 911
rect 5333 883 5363 911
rect 5417 883 5447 911
rect 5521 883 5551 911
rect 5605 883 5635 911
rect 5793 892 5823 918
rect 5877 892 5907 918
rect 5961 892 5991 918
rect 6045 892 6075 918
rect 6197 911 6418 941
rect 4751 873 5073 883
rect 4144 859 4278 869
rect 4144 825 4160 859
rect 4194 825 4228 859
rect 4262 825 4278 859
rect 4751 839 4811 873
rect 4845 839 4879 873
rect 4913 839 4947 873
rect 4981 839 5015 873
rect 5049 839 5073 873
rect 4751 829 5073 839
rect 5323 873 5645 883
rect 5323 839 5347 873
rect 5381 839 5415 873
rect 5449 839 5483 873
rect 5517 839 5551 873
rect 5585 839 5645 873
rect 5323 829 5645 839
rect 6118 859 6252 869
rect 4144 823 4278 825
rect 4144 815 4593 823
rect 4227 793 4593 815
rect 3628 763 3664 778
rect 3722 763 3758 778
rect 3970 763 4006 778
rect 4064 763 4100 778
rect 4273 777 4309 793
rect 4367 777 4403 793
rect 4461 777 4497 793
rect 4555 777 4591 793
rect 4753 791 4789 829
rect 4847 791 4883 829
rect 4941 791 4977 829
rect 5035 791 5071 829
rect 5325 791 5361 829
rect 5419 791 5455 829
rect 5513 791 5549 829
rect 5607 791 5643 829
rect 6118 825 6134 859
rect 6168 825 6202 859
rect 6236 825 6252 859
rect 6118 823 6252 825
rect 5803 815 6252 823
rect 5803 793 6169 815
rect 2177 565 2213 591
rect 2271 565 2307 591
rect 2365 565 2401 591
rect 2459 565 2495 591
rect 2657 565 2693 591
rect 2751 565 2787 591
rect 2845 565 2881 591
rect 2939 565 2975 591
rect 3137 565 3173 613
rect 3231 565 3267 613
rect 3325 565 3361 613
rect 3419 565 3455 613
rect 3628 565 3664 599
rect 3722 565 3758 599
rect 3970 565 4006 599
rect 4064 565 4100 599
rect 4273 565 4309 613
rect 4367 565 4403 613
rect 4461 565 4497 613
rect 4555 565 4591 613
rect 5805 777 5841 793
rect 5899 777 5935 793
rect 5993 777 6029 793
rect 6087 777 6123 793
rect 6294 778 6334 911
rect 6388 889 6418 911
rect 6646 941 6676 957
rect 6730 941 6760 957
rect 6837 941 6867 1037
rect 6989 1022 7019 1037
rect 7073 1022 7103 1037
rect 7157 1022 7187 1037
rect 7241 1022 7271 1037
rect 6646 911 6867 941
rect 6646 889 6676 911
rect 6388 873 6511 889
rect 6388 839 6399 873
rect 6433 839 6467 873
rect 6501 839 6511 873
rect 6388 823 6511 839
rect 6553 873 6676 889
rect 6553 839 6563 873
rect 6597 839 6631 873
rect 6665 839 6676 873
rect 6553 823 6676 839
rect 6388 778 6428 823
rect 6636 778 6676 823
rect 6730 778 6770 911
rect 6989 892 7019 918
rect 7073 892 7103 918
rect 7157 892 7187 918
rect 7241 892 7271 918
rect 8369 1037 8803 1067
rect 8880 1041 8910 1067
rect 8964 1041 8994 1067
rect 9222 1041 9252 1067
rect 9306 1041 9336 1067
rect 8369 1022 8399 1037
rect 8453 1022 8483 1037
rect 8537 1022 8567 1037
rect 8621 1022 8651 1037
rect 8773 941 8803 1037
rect 9413 1037 9847 1067
rect 10005 1041 10035 1067
rect 10089 1041 10119 1069
rect 10193 1041 10223 1067
rect 10277 1041 10307 1069
rect 8880 941 8910 957
rect 8964 941 8994 957
rect 7429 883 7459 911
rect 7513 883 7543 911
rect 7617 883 7647 911
rect 7701 883 7731 911
rect 7909 883 7939 911
rect 7993 883 8023 911
rect 8097 883 8127 911
rect 8181 883 8211 911
rect 8369 892 8399 918
rect 8453 892 8483 918
rect 8537 892 8567 918
rect 8621 892 8651 918
rect 8773 911 8994 941
rect 7419 873 7741 883
rect 6812 859 6946 869
rect 6812 825 6828 859
rect 6862 825 6896 859
rect 6930 825 6946 859
rect 7419 839 7479 873
rect 7513 839 7547 873
rect 7581 839 7615 873
rect 7649 839 7683 873
rect 7717 839 7741 873
rect 7419 829 7741 839
rect 7899 873 8221 883
rect 7899 839 7923 873
rect 7957 839 7991 873
rect 8025 839 8059 873
rect 8093 839 8127 873
rect 8161 839 8221 873
rect 7899 829 8221 839
rect 8694 859 8828 869
rect 6812 823 6946 825
rect 6812 815 7261 823
rect 6895 793 7261 815
rect 6296 763 6332 778
rect 6390 763 6426 778
rect 6638 763 6674 778
rect 6732 763 6768 778
rect 6941 777 6977 793
rect 7035 777 7071 793
rect 7129 777 7165 793
rect 7223 777 7259 793
rect 7421 791 7457 829
rect 7515 791 7551 829
rect 7609 791 7645 829
rect 7703 791 7739 829
rect 7901 791 7937 829
rect 7995 791 8031 829
rect 8089 791 8125 829
rect 8183 791 8219 829
rect 8694 825 8710 859
rect 8744 825 8778 859
rect 8812 825 8828 859
rect 8694 823 8828 825
rect 8379 815 8828 823
rect 8379 793 8745 815
rect 4753 565 4789 591
rect 4847 565 4883 591
rect 4941 565 4977 591
rect 5035 565 5071 591
rect 5325 565 5361 591
rect 5419 565 5455 591
rect 5513 565 5549 591
rect 5607 565 5643 591
rect 5805 565 5841 613
rect 5899 565 5935 613
rect 5993 565 6029 613
rect 6087 565 6123 613
rect 6296 565 6332 599
rect 6390 565 6426 599
rect 6638 565 6674 599
rect 6732 565 6768 599
rect 6941 565 6977 613
rect 7035 565 7071 613
rect 7129 565 7165 613
rect 7223 565 7259 613
rect 8381 777 8417 793
rect 8475 777 8511 793
rect 8569 777 8605 793
rect 8663 777 8699 793
rect 8870 778 8910 911
rect 8964 889 8994 911
rect 9222 941 9252 957
rect 9306 941 9336 957
rect 9413 941 9443 1037
rect 9565 1022 9595 1037
rect 9649 1022 9679 1037
rect 9733 1022 9763 1037
rect 9817 1022 9847 1037
rect 9222 911 9443 941
rect 9222 889 9252 911
rect 8964 873 9087 889
rect 8964 839 8975 873
rect 9009 839 9043 873
rect 9077 839 9087 873
rect 8964 823 9087 839
rect 9129 873 9252 889
rect 9129 839 9139 873
rect 9173 839 9207 873
rect 9241 839 9252 873
rect 9129 823 9252 839
rect 8964 778 9004 823
rect 9212 778 9252 823
rect 9306 778 9346 911
rect 9565 892 9595 918
rect 9649 892 9679 918
rect 9733 892 9763 918
rect 9817 892 9847 918
rect 10005 883 10035 911
rect 10089 883 10119 911
rect 10193 883 10223 911
rect 10277 883 10307 911
rect 9995 873 10317 883
rect 9388 859 9522 869
rect 9388 825 9404 859
rect 9438 825 9472 859
rect 9506 825 9522 859
rect 9995 839 10055 873
rect 10089 839 10123 873
rect 10157 839 10191 873
rect 10225 839 10259 873
rect 10293 839 10317 873
rect 9995 829 10317 839
rect 9388 823 9522 825
rect 9388 815 9837 823
rect 9471 793 9837 815
rect 8872 763 8908 778
rect 8966 763 9002 778
rect 9214 763 9250 778
rect 9308 763 9344 778
rect 9517 777 9553 793
rect 9611 777 9647 793
rect 9705 777 9741 793
rect 9799 777 9835 793
rect 9997 791 10033 829
rect 10091 791 10127 829
rect 10185 791 10221 829
rect 10279 791 10315 829
rect 7421 565 7457 591
rect 7515 565 7551 591
rect 7609 565 7645 591
rect 7703 565 7739 591
rect 7901 565 7937 591
rect 7995 565 8031 591
rect 8089 565 8125 591
rect 8183 565 8219 591
rect 8381 565 8417 613
rect 8475 565 8511 613
rect 8569 565 8605 613
rect 8663 565 8699 613
rect 8872 565 8908 599
rect 8966 565 9002 599
rect 9214 565 9250 599
rect 9308 565 9344 599
rect 9517 565 9553 613
rect 9611 565 9647 613
rect 9705 565 9741 613
rect 9799 565 9835 613
rect 9997 565 10033 591
rect 10091 565 10127 591
rect 10185 565 10221 591
rect 10279 565 10315 591
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 561 475 597 523
rect 655 475 691 523
rect 749 475 785 523
rect 843 475 879 523
rect 1052 489 1088 523
rect 1146 489 1182 523
rect 1394 489 1430 523
rect 1488 489 1524 523
rect 1697 475 1733 523
rect 1791 475 1827 523
rect 1885 475 1921 523
rect 1979 475 2015 523
rect 2177 497 2213 523
rect 2271 497 2307 523
rect 2365 497 2401 523
rect 2459 497 2495 523
rect 2657 497 2693 523
rect 2751 497 2787 523
rect 2845 497 2881 523
rect 2939 497 2975 523
rect 81 259 117 297
rect 175 259 211 297
rect 269 259 305 297
rect 363 259 399 297
rect 561 295 597 311
rect 655 295 691 311
rect 749 295 785 311
rect 843 295 879 311
rect 1052 310 1088 325
rect 1146 310 1182 325
rect 1394 310 1430 325
rect 1488 310 1524 325
rect 559 273 925 295
rect 559 265 1008 273
rect 874 263 1008 265
rect 79 249 401 259
rect 79 215 103 249
rect 137 215 171 249
rect 205 215 239 249
rect 273 215 307 249
rect 341 215 401 249
rect 874 229 890 263
rect 924 229 958 263
rect 992 229 1008 263
rect 874 219 1008 229
rect 79 205 401 215
rect 89 177 119 205
rect 173 177 203 205
rect 277 177 307 205
rect 361 177 391 205
rect 549 170 579 196
rect 633 170 663 196
rect 717 170 747 196
rect 801 170 831 196
rect 1050 177 1090 310
rect 1144 265 1184 310
rect 1392 265 1432 310
rect 1144 249 1267 265
rect 1144 215 1155 249
rect 1189 215 1223 249
rect 1257 215 1267 249
rect 1144 199 1267 215
rect 1309 249 1432 265
rect 1309 215 1319 249
rect 1353 215 1387 249
rect 1421 215 1432 249
rect 1309 199 1432 215
rect 1144 177 1174 199
rect 953 147 1174 177
rect 549 51 579 66
rect 633 51 663 66
rect 717 51 747 66
rect 801 51 831 66
rect 953 51 983 147
rect 1060 131 1090 147
rect 1144 131 1174 147
rect 1402 177 1432 199
rect 1486 177 1526 310
rect 1697 295 1733 311
rect 1791 295 1827 311
rect 1885 295 1921 311
rect 1979 295 2015 311
rect 3137 475 3173 523
rect 3231 475 3267 523
rect 3325 475 3361 523
rect 3419 475 3455 523
rect 3628 489 3664 523
rect 3722 489 3758 523
rect 3970 489 4006 523
rect 4064 489 4100 523
rect 4273 475 4309 523
rect 4367 475 4403 523
rect 4461 475 4497 523
rect 4555 475 4591 523
rect 4753 497 4789 523
rect 4847 497 4883 523
rect 4941 497 4977 523
rect 5035 497 5071 523
rect 5325 497 5361 523
rect 5419 497 5455 523
rect 5513 497 5549 523
rect 5607 497 5643 523
rect 1651 273 2017 295
rect 1568 265 2017 273
rect 1568 263 1702 265
rect 1568 229 1584 263
rect 1618 229 1652 263
rect 1686 229 1702 263
rect 2177 259 2213 297
rect 2271 259 2307 297
rect 2365 259 2401 297
rect 2459 259 2495 297
rect 2657 259 2693 297
rect 2751 259 2787 297
rect 2845 259 2881 297
rect 2939 259 2975 297
rect 3137 295 3173 311
rect 3231 295 3267 311
rect 3325 295 3361 311
rect 3419 295 3455 311
rect 3628 310 3664 325
rect 3722 310 3758 325
rect 3970 310 4006 325
rect 4064 310 4100 325
rect 3135 273 3501 295
rect 3135 265 3584 273
rect 3450 263 3584 265
rect 1568 219 1702 229
rect 2175 249 2497 259
rect 2175 215 2235 249
rect 2269 215 2303 249
rect 2337 215 2371 249
rect 2405 215 2439 249
rect 2473 215 2497 249
rect 2175 205 2497 215
rect 2655 249 2977 259
rect 2655 215 2679 249
rect 2713 215 2747 249
rect 2781 215 2815 249
rect 2849 215 2883 249
rect 2917 215 2977 249
rect 3450 229 3466 263
rect 3500 229 3534 263
rect 3568 229 3584 263
rect 3450 219 3584 229
rect 2655 205 2977 215
rect 1402 147 1623 177
rect 1745 170 1775 196
rect 1829 170 1859 196
rect 1913 170 1943 196
rect 1997 170 2027 196
rect 2185 177 2215 205
rect 2269 177 2299 205
rect 2373 177 2403 205
rect 2457 177 2487 205
rect 2665 177 2695 205
rect 2749 177 2779 205
rect 2853 177 2883 205
rect 2937 177 2967 205
rect 1402 131 1432 147
rect 1486 131 1516 147
rect 89 19 119 47
rect 173 21 203 47
rect 277 19 307 47
rect 361 21 391 47
rect 549 21 983 51
rect 1593 51 1623 147
rect 1745 51 1775 66
rect 1829 51 1859 66
rect 1913 51 1943 66
rect 1997 51 2027 66
rect 1060 21 1090 47
rect 1144 21 1174 47
rect 1402 21 1432 47
rect 1486 21 1516 47
rect 1593 21 2027 51
rect 3125 170 3155 196
rect 3209 170 3239 196
rect 3293 170 3323 196
rect 3377 170 3407 196
rect 3626 177 3666 310
rect 3720 265 3760 310
rect 3968 265 4008 310
rect 3720 249 3843 265
rect 3720 215 3731 249
rect 3765 215 3799 249
rect 3833 215 3843 249
rect 3720 199 3843 215
rect 3885 249 4008 265
rect 3885 215 3895 249
rect 3929 215 3963 249
rect 3997 215 4008 249
rect 3885 199 4008 215
rect 3720 177 3750 199
rect 3529 147 3750 177
rect 3125 51 3155 66
rect 3209 51 3239 66
rect 3293 51 3323 66
rect 3377 51 3407 66
rect 3529 51 3559 147
rect 3636 131 3666 147
rect 3720 131 3750 147
rect 3978 177 4008 199
rect 4062 177 4102 310
rect 4273 295 4309 311
rect 4367 295 4403 311
rect 4461 295 4497 311
rect 4555 295 4591 311
rect 5805 475 5841 523
rect 5899 475 5935 523
rect 5993 475 6029 523
rect 6087 475 6123 523
rect 6296 489 6332 523
rect 6390 489 6426 523
rect 6638 489 6674 523
rect 6732 489 6768 523
rect 6941 475 6977 523
rect 7035 475 7071 523
rect 7129 475 7165 523
rect 7223 475 7259 523
rect 7421 497 7457 523
rect 7515 497 7551 523
rect 7609 497 7645 523
rect 7703 497 7739 523
rect 7901 497 7937 523
rect 7995 497 8031 523
rect 8089 497 8125 523
rect 8183 497 8219 523
rect 4227 273 4593 295
rect 4144 265 4593 273
rect 4144 263 4278 265
rect 4144 229 4160 263
rect 4194 229 4228 263
rect 4262 229 4278 263
rect 4753 259 4789 297
rect 4847 259 4883 297
rect 4941 259 4977 297
rect 5035 259 5071 297
rect 5325 259 5361 297
rect 5419 259 5455 297
rect 5513 259 5549 297
rect 5607 259 5643 297
rect 5805 295 5841 311
rect 5899 295 5935 311
rect 5993 295 6029 311
rect 6087 295 6123 311
rect 6296 310 6332 325
rect 6390 310 6426 325
rect 6638 310 6674 325
rect 6732 310 6768 325
rect 5803 273 6169 295
rect 5803 265 6252 273
rect 6118 263 6252 265
rect 4144 219 4278 229
rect 4751 249 5073 259
rect 4751 215 4811 249
rect 4845 215 4879 249
rect 4913 215 4947 249
rect 4981 215 5015 249
rect 5049 215 5073 249
rect 4751 205 5073 215
rect 5323 249 5645 259
rect 5323 215 5347 249
rect 5381 215 5415 249
rect 5449 215 5483 249
rect 5517 215 5551 249
rect 5585 215 5645 249
rect 6118 229 6134 263
rect 6168 229 6202 263
rect 6236 229 6252 263
rect 6118 219 6252 229
rect 5323 205 5645 215
rect 3978 147 4199 177
rect 4321 170 4351 196
rect 4405 170 4435 196
rect 4489 170 4519 196
rect 4573 170 4603 196
rect 4761 177 4791 205
rect 4845 177 4875 205
rect 4949 177 4979 205
rect 5033 177 5063 205
rect 5333 177 5363 205
rect 5417 177 5447 205
rect 5521 177 5551 205
rect 5605 177 5635 205
rect 3978 131 4008 147
rect 4062 131 4092 147
rect 2185 21 2215 47
rect 2269 19 2299 47
rect 2373 21 2403 47
rect 2457 19 2487 47
rect 2665 19 2695 47
rect 2749 21 2779 47
rect 2853 19 2883 47
rect 2937 21 2967 47
rect 3125 21 3559 51
rect 4169 51 4199 147
rect 4321 51 4351 66
rect 4405 51 4435 66
rect 4489 51 4519 66
rect 4573 51 4603 66
rect 3636 21 3666 47
rect 3720 21 3750 47
rect 3978 21 4008 47
rect 4062 21 4092 47
rect 4169 21 4603 51
rect 5793 170 5823 196
rect 5877 170 5907 196
rect 5961 170 5991 196
rect 6045 170 6075 196
rect 6294 177 6334 310
rect 6388 265 6428 310
rect 6636 265 6676 310
rect 6388 249 6511 265
rect 6388 215 6399 249
rect 6433 215 6467 249
rect 6501 215 6511 249
rect 6388 199 6511 215
rect 6553 249 6676 265
rect 6553 215 6563 249
rect 6597 215 6631 249
rect 6665 215 6676 249
rect 6553 199 6676 215
rect 6388 177 6418 199
rect 6197 147 6418 177
rect 5793 51 5823 66
rect 5877 51 5907 66
rect 5961 51 5991 66
rect 6045 51 6075 66
rect 6197 51 6227 147
rect 6304 131 6334 147
rect 6388 131 6418 147
rect 6646 177 6676 199
rect 6730 177 6770 310
rect 6941 295 6977 311
rect 7035 295 7071 311
rect 7129 295 7165 311
rect 7223 295 7259 311
rect 8381 475 8417 523
rect 8475 475 8511 523
rect 8569 475 8605 523
rect 8663 475 8699 523
rect 8872 489 8908 523
rect 8966 489 9002 523
rect 9214 489 9250 523
rect 9308 489 9344 523
rect 9517 475 9553 523
rect 9611 475 9647 523
rect 9705 475 9741 523
rect 9799 475 9835 523
rect 9997 497 10033 523
rect 10091 497 10127 523
rect 10185 497 10221 523
rect 10279 497 10315 523
rect 6895 273 7261 295
rect 6812 265 7261 273
rect 6812 263 6946 265
rect 6812 229 6828 263
rect 6862 229 6896 263
rect 6930 229 6946 263
rect 7421 259 7457 297
rect 7515 259 7551 297
rect 7609 259 7645 297
rect 7703 259 7739 297
rect 7901 259 7937 297
rect 7995 259 8031 297
rect 8089 259 8125 297
rect 8183 259 8219 297
rect 8381 295 8417 311
rect 8475 295 8511 311
rect 8569 295 8605 311
rect 8663 295 8699 311
rect 8872 310 8908 325
rect 8966 310 9002 325
rect 9214 310 9250 325
rect 9308 310 9344 325
rect 8379 273 8745 295
rect 8379 265 8828 273
rect 8694 263 8828 265
rect 6812 219 6946 229
rect 7419 249 7741 259
rect 7419 215 7479 249
rect 7513 215 7547 249
rect 7581 215 7615 249
rect 7649 215 7683 249
rect 7717 215 7741 249
rect 7419 205 7741 215
rect 7899 249 8221 259
rect 7899 215 7923 249
rect 7957 215 7991 249
rect 8025 215 8059 249
rect 8093 215 8127 249
rect 8161 215 8221 249
rect 8694 229 8710 263
rect 8744 229 8778 263
rect 8812 229 8828 263
rect 8694 219 8828 229
rect 7899 205 8221 215
rect 6646 147 6867 177
rect 6989 170 7019 196
rect 7073 170 7103 196
rect 7157 170 7187 196
rect 7241 170 7271 196
rect 7429 177 7459 205
rect 7513 177 7543 205
rect 7617 177 7647 205
rect 7701 177 7731 205
rect 7909 177 7939 205
rect 7993 177 8023 205
rect 8097 177 8127 205
rect 8181 177 8211 205
rect 6646 131 6676 147
rect 6730 131 6760 147
rect 4761 21 4791 47
rect 4845 19 4875 47
rect 4949 21 4979 47
rect 5033 19 5063 47
rect 5333 19 5363 47
rect 5417 21 5447 47
rect 5521 19 5551 47
rect 5605 21 5635 47
rect 5793 21 6227 51
rect 6837 51 6867 147
rect 6989 51 7019 66
rect 7073 51 7103 66
rect 7157 51 7187 66
rect 7241 51 7271 66
rect 6304 21 6334 47
rect 6388 21 6418 47
rect 6646 21 6676 47
rect 6730 21 6760 47
rect 6837 21 7271 51
rect 8369 170 8399 196
rect 8453 170 8483 196
rect 8537 170 8567 196
rect 8621 170 8651 196
rect 8870 177 8910 310
rect 8964 265 9004 310
rect 9212 265 9252 310
rect 8964 249 9087 265
rect 8964 215 8975 249
rect 9009 215 9043 249
rect 9077 215 9087 249
rect 8964 199 9087 215
rect 9129 249 9252 265
rect 9129 215 9139 249
rect 9173 215 9207 249
rect 9241 215 9252 249
rect 9129 199 9252 215
rect 8964 177 8994 199
rect 8773 147 8994 177
rect 8369 51 8399 66
rect 8453 51 8483 66
rect 8537 51 8567 66
rect 8621 51 8651 66
rect 8773 51 8803 147
rect 8880 131 8910 147
rect 8964 131 8994 147
rect 9222 177 9252 199
rect 9306 177 9346 310
rect 9517 295 9553 311
rect 9611 295 9647 311
rect 9705 295 9741 311
rect 9799 295 9835 311
rect 9471 273 9837 295
rect 9388 265 9837 273
rect 9388 263 9522 265
rect 9388 229 9404 263
rect 9438 229 9472 263
rect 9506 229 9522 263
rect 9997 259 10033 297
rect 10091 259 10127 297
rect 10185 259 10221 297
rect 10279 259 10315 297
rect 9388 219 9522 229
rect 9995 249 10317 259
rect 9995 215 10055 249
rect 10089 215 10123 249
rect 10157 215 10191 249
rect 10225 215 10259 249
rect 10293 215 10317 249
rect 9995 205 10317 215
rect 9222 147 9443 177
rect 9565 170 9595 196
rect 9649 170 9679 196
rect 9733 170 9763 196
rect 9817 170 9847 196
rect 10005 177 10035 205
rect 10089 177 10119 205
rect 10193 177 10223 205
rect 10277 177 10307 205
rect 9222 131 9252 147
rect 9306 131 9336 147
rect 7429 21 7459 47
rect 7513 19 7543 47
rect 7617 21 7647 47
rect 7701 19 7731 47
rect 7909 19 7939 47
rect 7993 21 8023 47
rect 8097 19 8127 47
rect 8181 21 8211 47
rect 8369 21 8803 51
rect 9413 51 9443 147
rect 9565 51 9595 66
rect 9649 51 9679 66
rect 9733 51 9763 66
rect 9817 51 9847 66
rect 8880 21 8910 47
rect 8964 21 8994 47
rect 9222 21 9252 47
rect 9306 21 9336 47
rect 9413 21 9847 51
rect 10005 21 10035 47
rect 10089 19 10119 47
rect 10193 21 10223 47
rect 10277 19 10307 47
<< polycont >>
rect 103 839 137 873
rect 171 839 205 873
rect 239 839 273 873
rect 307 839 341 873
rect 890 825 924 859
rect 958 825 992 859
rect 1155 839 1189 873
rect 1223 839 1257 873
rect 1319 839 1353 873
rect 1387 839 1421 873
rect 1584 825 1618 859
rect 1652 825 1686 859
rect 2235 839 2269 873
rect 2303 839 2337 873
rect 2371 839 2405 873
rect 2439 839 2473 873
rect 2679 839 2713 873
rect 2747 839 2781 873
rect 2815 839 2849 873
rect 2883 839 2917 873
rect 3466 825 3500 859
rect 3534 825 3568 859
rect 3731 839 3765 873
rect 3799 839 3833 873
rect 3895 839 3929 873
rect 3963 839 3997 873
rect 4160 825 4194 859
rect 4228 825 4262 859
rect 4811 839 4845 873
rect 4879 839 4913 873
rect 4947 839 4981 873
rect 5015 839 5049 873
rect 5347 839 5381 873
rect 5415 839 5449 873
rect 5483 839 5517 873
rect 5551 839 5585 873
rect 6134 825 6168 859
rect 6202 825 6236 859
rect 6399 839 6433 873
rect 6467 839 6501 873
rect 6563 839 6597 873
rect 6631 839 6665 873
rect 6828 825 6862 859
rect 6896 825 6930 859
rect 7479 839 7513 873
rect 7547 839 7581 873
rect 7615 839 7649 873
rect 7683 839 7717 873
rect 7923 839 7957 873
rect 7991 839 8025 873
rect 8059 839 8093 873
rect 8127 839 8161 873
rect 8710 825 8744 859
rect 8778 825 8812 859
rect 8975 839 9009 873
rect 9043 839 9077 873
rect 9139 839 9173 873
rect 9207 839 9241 873
rect 9404 825 9438 859
rect 9472 825 9506 859
rect 10055 839 10089 873
rect 10123 839 10157 873
rect 10191 839 10225 873
rect 10259 839 10293 873
rect 103 215 137 249
rect 171 215 205 249
rect 239 215 273 249
rect 307 215 341 249
rect 890 229 924 263
rect 958 229 992 263
rect 1155 215 1189 249
rect 1223 215 1257 249
rect 1319 215 1353 249
rect 1387 215 1421 249
rect 1584 229 1618 263
rect 1652 229 1686 263
rect 2235 215 2269 249
rect 2303 215 2337 249
rect 2371 215 2405 249
rect 2439 215 2473 249
rect 2679 215 2713 249
rect 2747 215 2781 249
rect 2815 215 2849 249
rect 2883 215 2917 249
rect 3466 229 3500 263
rect 3534 229 3568 263
rect 3731 215 3765 249
rect 3799 215 3833 249
rect 3895 215 3929 249
rect 3963 215 3997 249
rect 4160 229 4194 263
rect 4228 229 4262 263
rect 4811 215 4845 249
rect 4879 215 4913 249
rect 4947 215 4981 249
rect 5015 215 5049 249
rect 5347 215 5381 249
rect 5415 215 5449 249
rect 5483 215 5517 249
rect 5551 215 5585 249
rect 6134 229 6168 263
rect 6202 229 6236 263
rect 6399 215 6433 249
rect 6467 215 6501 249
rect 6563 215 6597 249
rect 6631 215 6665 249
rect 6828 229 6862 263
rect 6896 229 6930 263
rect 7479 215 7513 249
rect 7547 215 7581 249
rect 7615 215 7649 249
rect 7683 215 7717 249
rect 7923 215 7957 249
rect 7991 215 8025 249
rect 8059 215 8093 249
rect 8127 215 8161 249
rect 8710 229 8744 263
rect 8778 229 8812 263
rect 8975 215 9009 249
rect 9043 215 9077 249
rect 9139 215 9173 249
rect 9207 215 9241 249
rect 9404 229 9438 263
rect 9472 229 9506 263
rect 10055 215 10089 249
rect 10123 215 10157 249
rect 10191 215 10225 249
rect 10259 215 10293 249
<< locali >>
rect 0 1071 29 1105
rect 63 1071 121 1105
rect 155 1071 213 1105
rect 247 1071 305 1105
rect 339 1071 397 1105
rect 431 1071 489 1105
rect 523 1071 581 1105
rect 615 1071 673 1105
rect 707 1071 765 1105
rect 799 1071 857 1105
rect 891 1071 949 1105
rect 983 1071 1041 1105
rect 1075 1071 1133 1105
rect 1167 1071 1225 1105
rect 1259 1071 1317 1105
rect 1351 1071 1409 1105
rect 1443 1071 1501 1105
rect 1535 1071 1593 1105
rect 1627 1071 1685 1105
rect 1719 1071 1777 1105
rect 1811 1071 1869 1105
rect 1903 1071 1961 1105
rect 1995 1071 2053 1105
rect 2087 1071 2145 1105
rect 2179 1071 2237 1105
rect 2271 1071 2329 1105
rect 2363 1071 2421 1105
rect 2455 1071 2513 1105
rect 2547 1071 2605 1105
rect 2639 1071 2697 1105
rect 2731 1071 2789 1105
rect 2823 1071 2881 1105
rect 2915 1071 2973 1105
rect 3007 1071 3065 1105
rect 3099 1071 3157 1105
rect 3191 1071 3249 1105
rect 3283 1071 3341 1105
rect 3375 1071 3433 1105
rect 3467 1071 3525 1105
rect 3559 1071 3617 1105
rect 3651 1071 3709 1105
rect 3743 1071 3801 1105
rect 3835 1071 3893 1105
rect 3927 1071 3985 1105
rect 4019 1071 4077 1105
rect 4111 1071 4169 1105
rect 4203 1071 4261 1105
rect 4295 1071 4353 1105
rect 4387 1071 4445 1105
rect 4479 1071 4537 1105
rect 4571 1071 4629 1105
rect 4663 1071 4721 1105
rect 4755 1071 4813 1105
rect 4847 1071 4905 1105
rect 4939 1071 4997 1105
rect 5031 1071 5089 1105
rect 5123 1071 5181 1105
rect 5215 1071 5273 1105
rect 5307 1071 5365 1105
rect 5399 1071 5457 1105
rect 5491 1071 5549 1105
rect 5583 1071 5641 1105
rect 5675 1071 5733 1105
rect 5767 1071 5825 1105
rect 5859 1071 5917 1105
rect 5951 1071 6009 1105
rect 6043 1071 6101 1105
rect 6135 1071 6193 1105
rect 6227 1071 6285 1105
rect 6319 1071 6377 1105
rect 6411 1071 6469 1105
rect 6503 1071 6561 1105
rect 6595 1071 6653 1105
rect 6687 1071 6745 1105
rect 6779 1071 6837 1105
rect 6871 1071 6929 1105
rect 6963 1071 7021 1105
rect 7055 1071 7113 1105
rect 7147 1071 7205 1105
rect 7239 1071 7297 1105
rect 7331 1071 7389 1105
rect 7423 1071 7481 1105
rect 7515 1071 7573 1105
rect 7607 1071 7665 1105
rect 7699 1071 7757 1105
rect 7791 1071 7849 1105
rect 7883 1071 7941 1105
rect 7975 1071 8033 1105
rect 8067 1071 8125 1105
rect 8159 1071 8217 1105
rect 8251 1071 8309 1105
rect 8343 1071 8401 1105
rect 8435 1071 8493 1105
rect 8527 1071 8585 1105
rect 8619 1071 8677 1105
rect 8711 1071 8769 1105
rect 8803 1071 8861 1105
rect 8895 1071 8953 1105
rect 8987 1071 9045 1105
rect 9079 1071 9137 1105
rect 9171 1071 9229 1105
rect 9263 1071 9321 1105
rect 9355 1071 9413 1105
rect 9447 1071 9505 1105
rect 9539 1071 9597 1105
rect 9631 1071 9689 1105
rect 9723 1071 9781 1105
rect 9815 1071 9873 1105
rect 9907 1071 9965 1105
rect 9999 1071 10057 1105
rect 10091 1071 10149 1105
rect 10183 1071 10241 1105
rect 10275 1071 10333 1105
rect 10367 1071 10396 1105
rect 29 1029 79 1071
rect 29 995 45 1029
rect 29 961 79 995
rect 29 927 45 961
rect 29 911 79 927
rect 113 1029 179 1037
rect 113 995 129 1029
rect 163 995 179 1029
rect 113 961 179 995
rect 213 1029 267 1071
rect 213 995 223 1029
rect 257 995 267 1029
rect 213 979 267 995
rect 301 1029 367 1037
rect 301 995 317 1029
rect 351 995 367 1029
rect 113 927 129 961
rect 163 945 179 961
rect 301 961 367 995
rect 401 1029 451 1071
rect 435 995 451 1029
rect 401 979 451 995
rect 485 1003 891 1037
rect 485 987 539 1003
rect 301 945 317 961
rect 163 927 317 945
rect 351 945 367 961
rect 485 953 505 987
rect 673 987 707 1003
rect 485 945 539 953
rect 351 927 539 945
rect 113 911 539 927
rect 573 935 589 969
rect 623 935 639 969
rect 573 911 639 935
rect 841 987 891 1003
rect 673 934 707 953
rect 741 935 757 969
rect 791 935 807 969
rect 79 873 357 877
rect 79 839 103 873
rect 137 839 171 873
rect 205 839 239 873
rect 273 839 307 873
rect 341 839 357 873
rect 79 823 357 839
rect 593 875 639 911
rect 741 875 807 935
rect 875 953 891 987
rect 992 1016 1050 1071
rect 992 982 1016 1016
rect 992 966 1050 982
rect 1084 1016 1134 1032
rect 1084 982 1100 1016
rect 841 934 891 953
rect 1084 923 1134 982
rect 1176 1016 1234 1071
rect 1176 982 1184 1016
rect 1218 982 1234 1016
rect 1176 966 1234 982
rect 1342 1016 1400 1071
rect 1342 982 1358 1016
rect 1392 982 1400 1016
rect 1342 966 1400 982
rect 1442 1016 1492 1032
rect 1476 982 1492 1016
rect 1442 923 1492 982
rect 1526 1016 1584 1071
rect 1560 982 1584 1016
rect 1526 966 1584 982
rect 1685 1003 2091 1037
rect 1685 987 1735 1003
rect 1685 953 1701 987
rect 1869 987 1903 1003
rect 1685 934 1735 953
rect 1769 935 1785 969
rect 1819 935 1835 969
rect 1084 875 1118 923
rect 593 815 847 875
rect 25 773 79 789
rect 25 739 35 773
rect 69 739 79 773
rect 25 705 79 739
rect 25 671 35 705
rect 69 671 79 705
rect 25 637 79 671
rect 25 603 35 637
rect 69 603 79 637
rect 25 561 79 603
rect 113 773 559 789
rect 113 739 129 773
rect 163 755 317 773
rect 163 739 179 755
rect 113 705 179 739
rect 301 739 317 755
rect 351 765 559 773
rect 351 755 515 765
rect 351 739 367 755
rect 113 671 129 705
rect 163 671 179 705
rect 113 660 179 671
rect 113 603 129 660
rect 163 603 179 660
rect 113 595 179 603
rect 213 705 267 721
rect 213 671 223 705
rect 257 671 267 705
rect 213 637 267 671
rect 213 603 223 637
rect 257 603 267 637
rect 213 561 267 603
rect 301 705 367 739
rect 499 731 515 755
rect 549 731 559 765
rect 301 671 317 705
rect 351 671 367 705
rect 301 660 367 671
rect 301 603 317 660
rect 351 603 367 660
rect 301 595 367 603
rect 401 705 455 721
rect 401 671 411 705
rect 445 671 455 705
rect 401 637 455 671
rect 401 603 411 637
rect 445 603 455 637
rect 401 561 455 603
rect 499 660 559 731
rect 499 626 513 660
rect 547 659 559 660
rect 499 625 515 626
rect 549 625 559 659
rect 499 595 559 625
rect 593 765 659 815
rect 593 697 609 765
rect 643 697 659 765
rect 593 659 659 697
rect 593 625 609 659
rect 643 625 659 659
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 559 561
rect 25 485 79 527
rect 25 451 35 485
rect 69 451 79 485
rect 25 417 79 451
rect 25 383 35 417
rect 69 383 79 417
rect 25 349 79 383
rect 25 315 35 349
rect 69 315 79 349
rect 25 299 79 315
rect 113 485 179 493
rect 113 428 129 485
rect 163 428 179 485
rect 113 417 179 428
rect 113 383 129 417
rect 163 383 179 417
rect 113 349 179 383
rect 213 485 267 527
rect 213 451 223 485
rect 257 451 267 485
rect 213 417 267 451
rect 213 383 223 417
rect 257 383 267 417
rect 213 367 267 383
rect 301 485 367 493
rect 301 428 317 485
rect 351 428 367 485
rect 301 417 367 428
rect 301 383 317 417
rect 351 383 367 417
rect 113 315 129 349
rect 163 333 179 349
rect 301 349 367 383
rect 401 485 455 527
rect 401 451 411 485
rect 445 451 455 485
rect 401 417 455 451
rect 401 383 411 417
rect 445 383 455 417
rect 401 367 455 383
rect 499 463 559 493
rect 499 462 515 463
rect 499 428 513 462
rect 549 429 559 463
rect 547 428 559 429
rect 301 333 317 349
rect 163 315 317 333
rect 351 333 367 349
rect 499 357 559 428
rect 499 333 515 357
rect 351 323 515 333
rect 549 323 559 357
rect 351 315 559 323
rect 113 299 559 315
rect 593 463 659 625
rect 693 765 747 781
rect 693 731 703 765
rect 737 731 747 765
rect 693 660 747 731
rect 693 625 703 660
rect 737 625 747 660
rect 693 595 747 625
rect 781 765 847 815
rect 881 859 1118 875
rect 881 825 890 859
rect 924 825 958 859
rect 992 825 1118 859
rect 881 809 1118 825
rect 1152 873 1271 889
rect 1152 839 1155 873
rect 1189 839 1223 873
rect 1257 839 1271 873
rect 1152 823 1271 839
rect 1305 873 1424 889
rect 1305 839 1319 873
rect 1353 839 1387 873
rect 1421 839 1424 873
rect 1305 823 1424 839
rect 1458 875 1492 923
rect 1769 875 1835 935
rect 2037 987 2091 1003
rect 1869 934 1903 953
rect 1937 935 1953 969
rect 1987 935 2003 969
rect 1937 911 2003 935
rect 2071 953 2091 987
rect 2125 1029 2175 1071
rect 2125 995 2141 1029
rect 2125 979 2175 995
rect 2209 1029 2275 1037
rect 2209 995 2225 1029
rect 2259 995 2275 1029
rect 2037 945 2091 953
rect 2209 961 2275 995
rect 2309 1029 2363 1071
rect 2309 995 2319 1029
rect 2353 995 2363 1029
rect 2309 979 2363 995
rect 2397 1029 2463 1037
rect 2397 995 2413 1029
rect 2447 995 2463 1029
rect 2209 945 2225 961
rect 2037 927 2225 945
rect 2259 945 2275 961
rect 2397 961 2463 995
rect 2397 945 2413 961
rect 2259 927 2413 945
rect 2447 927 2463 961
rect 2037 911 2463 927
rect 2497 1029 2547 1071
rect 2531 995 2547 1029
rect 2497 961 2547 995
rect 2531 927 2547 961
rect 2497 911 2547 927
rect 2605 1029 2655 1071
rect 2605 995 2621 1029
rect 2605 961 2655 995
rect 2605 927 2621 961
rect 2605 911 2655 927
rect 2689 1029 2755 1037
rect 2689 995 2705 1029
rect 2739 995 2755 1029
rect 2689 961 2755 995
rect 2789 1029 2843 1071
rect 2789 995 2799 1029
rect 2833 995 2843 1029
rect 2789 979 2843 995
rect 2877 1029 2943 1037
rect 2877 995 2893 1029
rect 2927 995 2943 1029
rect 2689 927 2705 961
rect 2739 945 2755 961
rect 2877 961 2943 995
rect 2977 1029 3027 1071
rect 3011 995 3027 1029
rect 2977 979 3027 995
rect 3061 1003 3467 1037
rect 3061 987 3115 1003
rect 2877 945 2893 961
rect 2739 927 2893 945
rect 2927 945 2943 961
rect 3061 953 3081 987
rect 3249 987 3283 1003
rect 3061 945 3115 953
rect 2927 927 3115 945
rect 2689 911 3115 927
rect 3149 935 3165 969
rect 3199 935 3215 969
rect 3149 911 3215 935
rect 3417 987 3467 1003
rect 3249 934 3283 953
rect 3317 935 3333 969
rect 3367 935 3383 969
rect 1937 875 1983 911
rect 1458 859 1695 875
rect 1458 825 1584 859
rect 1618 825 1652 859
rect 1686 825 1695 859
rect 781 697 797 765
rect 831 697 847 765
rect 781 659 847 697
rect 781 625 797 659
rect 831 625 847 659
rect 593 429 609 463
rect 643 429 659 463
rect 593 391 659 429
rect 593 323 609 391
rect 643 323 659 391
rect 593 273 659 323
rect 693 463 747 493
rect 693 428 703 463
rect 737 428 747 463
rect 693 357 747 428
rect 693 323 703 357
rect 737 323 747 357
rect 693 307 747 323
rect 781 463 847 625
rect 881 759 941 775
rect 1084 767 1118 809
rect 1458 809 1695 825
rect 1729 815 1983 875
rect 2219 873 2497 877
rect 2219 839 2235 873
rect 2269 839 2303 873
rect 2337 839 2371 873
rect 2405 839 2439 873
rect 2473 839 2497 873
rect 2219 823 2497 839
rect 2655 873 2933 877
rect 2655 839 2679 873
rect 2713 839 2747 873
rect 2781 839 2815 873
rect 2849 839 2883 873
rect 2917 839 2933 873
rect 2655 823 2933 839
rect 3169 875 3215 911
rect 3317 875 3383 935
rect 3451 953 3467 987
rect 3568 1016 3626 1071
rect 3568 982 3592 1016
rect 3568 966 3626 982
rect 3660 1016 3710 1032
rect 3660 982 3676 1016
rect 3417 934 3467 953
rect 3660 923 3710 982
rect 3752 1016 3810 1071
rect 3752 982 3760 1016
rect 3794 982 3810 1016
rect 3752 966 3810 982
rect 3918 1016 3976 1071
rect 3918 982 3934 1016
rect 3968 982 3976 1016
rect 3918 966 3976 982
rect 4018 1016 4068 1032
rect 4052 982 4068 1016
rect 4018 923 4068 982
rect 4102 1016 4160 1071
rect 4136 982 4160 1016
rect 4102 966 4160 982
rect 4261 1003 4667 1037
rect 4261 987 4311 1003
rect 4261 953 4277 987
rect 4445 987 4479 1003
rect 4261 934 4311 953
rect 4345 935 4361 969
rect 4395 935 4411 969
rect 3660 875 3694 923
rect 1458 767 1492 809
rect 881 725 891 759
rect 925 725 941 759
rect 881 660 941 725
rect 881 659 893 660
rect 881 625 891 659
rect 927 626 941 660
rect 925 625 941 626
rect 881 595 941 625
rect 990 751 1045 767
rect 990 717 1006 751
rect 1040 717 1045 751
rect 990 645 1045 717
rect 990 611 1006 645
rect 1040 611 1045 645
rect 990 561 1045 611
rect 1084 751 1150 767
rect 1084 717 1100 751
rect 1134 717 1150 751
rect 1084 645 1150 717
rect 1084 611 1100 645
rect 1134 611 1150 645
rect 1084 595 1150 611
rect 1184 751 1244 767
rect 1184 717 1194 751
rect 1228 717 1244 751
rect 1184 645 1244 717
rect 1184 611 1194 645
rect 1228 611 1244 645
rect 1184 561 1244 611
rect 1332 751 1392 767
rect 1332 717 1348 751
rect 1382 717 1392 751
rect 1332 645 1392 717
rect 1332 611 1348 645
rect 1382 611 1392 645
rect 1332 561 1392 611
rect 1426 751 1492 767
rect 1426 717 1442 751
rect 1476 717 1492 751
rect 1426 645 1492 717
rect 1426 611 1442 645
rect 1476 611 1492 645
rect 1426 595 1492 611
rect 1531 751 1586 767
rect 1531 717 1536 751
rect 1570 717 1586 751
rect 1531 645 1586 717
rect 1531 611 1536 645
rect 1570 611 1586 645
rect 1531 561 1586 611
rect 1635 759 1695 775
rect 1635 725 1651 759
rect 1685 725 1695 759
rect 1635 660 1695 725
rect 1635 626 1649 660
rect 1683 659 1695 660
rect 1635 625 1651 626
rect 1685 625 1695 659
rect 1635 595 1695 625
rect 1729 765 1795 815
rect 1729 697 1745 765
rect 1779 697 1795 765
rect 1729 659 1795 697
rect 1729 625 1745 659
rect 1779 625 1795 659
rect 881 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1695 561
rect 781 429 797 463
rect 831 429 847 463
rect 781 391 847 429
rect 781 323 797 391
rect 831 323 847 391
rect 781 273 847 323
rect 881 463 941 493
rect 881 429 891 463
rect 925 462 941 463
rect 881 428 893 429
rect 927 428 941 462
rect 881 363 941 428
rect 881 329 891 363
rect 925 329 941 363
rect 881 313 941 329
rect 990 477 1045 527
rect 990 443 1006 477
rect 1040 443 1045 477
rect 990 371 1045 443
rect 990 337 1006 371
rect 1040 337 1045 371
rect 990 321 1045 337
rect 1084 477 1150 493
rect 1084 443 1100 477
rect 1134 443 1150 477
rect 1084 371 1150 443
rect 1084 337 1100 371
rect 1134 337 1150 371
rect 1084 321 1150 337
rect 1184 477 1244 527
rect 1184 443 1194 477
rect 1228 443 1244 477
rect 1184 371 1244 443
rect 1184 337 1194 371
rect 1228 337 1244 371
rect 1184 321 1244 337
rect 1332 477 1392 527
rect 1332 443 1348 477
rect 1382 443 1392 477
rect 1332 371 1392 443
rect 1332 337 1348 371
rect 1382 337 1392 371
rect 1332 321 1392 337
rect 1426 477 1492 493
rect 1426 443 1442 477
rect 1476 443 1492 477
rect 1426 371 1492 443
rect 1426 337 1442 371
rect 1476 337 1492 371
rect 1426 321 1492 337
rect 1531 477 1586 527
rect 1531 443 1536 477
rect 1570 443 1586 477
rect 1531 371 1586 443
rect 1531 337 1536 371
rect 1570 337 1586 371
rect 1531 321 1586 337
rect 1635 463 1695 493
rect 1635 462 1651 463
rect 1635 428 1649 462
rect 1685 429 1695 463
rect 1683 428 1695 429
rect 1635 363 1695 428
rect 1635 329 1651 363
rect 1685 329 1695 363
rect 1084 279 1118 321
rect 79 249 357 265
rect 79 215 103 249
rect 137 215 171 249
rect 205 215 239 249
rect 273 215 307 249
rect 341 215 357 249
rect 79 211 357 215
rect 593 213 847 273
rect 881 263 1118 279
rect 1458 279 1492 321
rect 1635 313 1695 329
rect 1729 463 1795 625
rect 1829 765 1883 781
rect 1829 731 1839 765
rect 1873 731 1883 765
rect 1829 660 1883 731
rect 1829 625 1839 660
rect 1873 625 1883 660
rect 1829 595 1883 625
rect 1917 765 1983 815
rect 3169 815 3423 875
rect 1917 697 1933 765
rect 1967 697 1983 765
rect 1917 659 1983 697
rect 1917 625 1933 659
rect 1967 625 1983 659
rect 1729 429 1745 463
rect 1779 429 1795 463
rect 1729 391 1795 429
rect 1729 323 1745 391
rect 1779 323 1795 391
rect 881 229 890 263
rect 924 229 958 263
rect 992 229 1118 263
rect 881 213 1118 229
rect 593 177 639 213
rect 29 161 79 177
rect 29 127 45 161
rect 29 93 79 127
rect 29 59 45 93
rect 29 17 79 59
rect 113 161 539 177
rect 113 127 129 161
rect 163 143 317 161
rect 163 127 179 143
rect 113 93 179 127
rect 301 127 317 143
rect 351 143 539 161
rect 351 127 367 143
rect 113 59 129 93
rect 163 59 179 93
rect 113 51 179 59
rect 213 93 267 109
rect 213 59 223 93
rect 257 59 267 93
rect 213 17 267 59
rect 301 93 367 127
rect 485 135 539 143
rect 301 59 317 93
rect 351 59 367 93
rect 301 51 367 59
rect 401 93 451 109
rect 435 59 451 93
rect 401 17 451 59
rect 485 101 505 135
rect 573 153 639 177
rect 573 119 589 153
rect 623 119 639 153
rect 673 135 707 154
rect 485 85 539 101
rect 741 153 807 213
rect 1084 165 1118 213
rect 1152 249 1271 265
rect 1152 215 1155 249
rect 1189 215 1223 249
rect 1257 215 1271 249
rect 1152 199 1271 215
rect 1305 249 1424 265
rect 1305 215 1319 249
rect 1353 215 1387 249
rect 1421 215 1424 249
rect 1305 199 1424 215
rect 1458 263 1695 279
rect 1458 229 1584 263
rect 1618 229 1652 263
rect 1686 229 1695 263
rect 1458 213 1695 229
rect 1729 273 1795 323
rect 1829 463 1883 493
rect 1829 428 1839 463
rect 1873 428 1883 463
rect 1829 357 1883 428
rect 1829 323 1839 357
rect 1873 323 1883 357
rect 1829 307 1883 323
rect 1917 463 1983 625
rect 2017 773 2463 789
rect 2017 765 2225 773
rect 2017 731 2027 765
rect 2061 755 2225 765
rect 2061 731 2077 755
rect 2017 660 2077 731
rect 2209 739 2225 755
rect 2259 755 2413 773
rect 2259 739 2275 755
rect 2017 659 2029 660
rect 2017 625 2027 659
rect 2063 626 2077 660
rect 2061 625 2077 626
rect 2017 595 2077 625
rect 2121 705 2175 721
rect 2121 671 2131 705
rect 2165 671 2175 705
rect 2121 637 2175 671
rect 2121 603 2131 637
rect 2165 603 2175 637
rect 2121 561 2175 603
rect 2209 705 2275 739
rect 2397 739 2413 755
rect 2447 739 2463 773
rect 2209 671 2225 705
rect 2259 671 2275 705
rect 2209 660 2275 671
rect 2209 603 2225 660
rect 2259 603 2275 660
rect 2209 595 2275 603
rect 2309 705 2363 721
rect 2309 671 2319 705
rect 2353 671 2363 705
rect 2309 637 2363 671
rect 2309 603 2319 637
rect 2353 603 2363 637
rect 2309 561 2363 603
rect 2397 705 2463 739
rect 2397 671 2413 705
rect 2447 671 2463 705
rect 2397 660 2463 671
rect 2397 603 2413 660
rect 2447 603 2463 660
rect 2397 595 2463 603
rect 2497 773 2551 789
rect 2497 739 2507 773
rect 2541 739 2551 773
rect 2497 705 2551 739
rect 2497 671 2507 705
rect 2541 671 2551 705
rect 2497 637 2551 671
rect 2497 603 2507 637
rect 2541 603 2551 637
rect 2497 561 2551 603
rect 2601 773 2655 789
rect 2601 739 2611 773
rect 2645 739 2655 773
rect 2601 705 2655 739
rect 2601 671 2611 705
rect 2645 671 2655 705
rect 2601 637 2655 671
rect 2601 603 2611 637
rect 2645 603 2655 637
rect 2601 561 2655 603
rect 2689 773 3135 789
rect 2689 739 2705 773
rect 2739 755 2893 773
rect 2739 739 2755 755
rect 2689 705 2755 739
rect 2877 739 2893 755
rect 2927 765 3135 773
rect 2927 755 3091 765
rect 2927 739 2943 755
rect 2689 671 2705 705
rect 2739 671 2755 705
rect 2689 660 2755 671
rect 2689 603 2705 660
rect 2739 603 2755 660
rect 2689 595 2755 603
rect 2789 705 2843 721
rect 2789 671 2799 705
rect 2833 671 2843 705
rect 2789 637 2843 671
rect 2789 603 2799 637
rect 2833 603 2843 637
rect 2789 561 2843 603
rect 2877 705 2943 739
rect 3075 731 3091 755
rect 3125 731 3135 765
rect 2877 671 2893 705
rect 2927 671 2943 705
rect 2877 660 2943 671
rect 2877 603 2893 660
rect 2927 603 2943 660
rect 2877 595 2943 603
rect 2977 705 3031 721
rect 2977 671 2987 705
rect 3021 671 3031 705
rect 2977 637 3031 671
rect 2977 603 2987 637
rect 3021 603 3031 637
rect 2977 561 3031 603
rect 3075 660 3135 731
rect 3075 626 3089 660
rect 3123 659 3135 660
rect 3075 625 3091 626
rect 3125 625 3135 659
rect 3075 595 3135 625
rect 3169 765 3235 815
rect 3169 697 3185 765
rect 3219 697 3235 765
rect 3169 659 3235 697
rect 3169 625 3185 659
rect 3219 625 3235 659
rect 2017 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3135 561
rect 1917 429 1933 463
rect 1967 429 1983 463
rect 1917 391 1983 429
rect 1917 323 1933 391
rect 1967 323 1983 391
rect 1917 273 1983 323
rect 2017 463 2077 493
rect 2017 429 2027 463
rect 2061 462 2077 463
rect 2017 428 2029 429
rect 2063 428 2077 462
rect 2017 357 2077 428
rect 2121 485 2175 527
rect 2121 451 2131 485
rect 2165 451 2175 485
rect 2121 417 2175 451
rect 2121 383 2131 417
rect 2165 383 2175 417
rect 2121 367 2175 383
rect 2209 485 2275 493
rect 2209 428 2225 485
rect 2259 428 2275 485
rect 2209 417 2275 428
rect 2209 383 2225 417
rect 2259 383 2275 417
rect 2017 323 2027 357
rect 2061 333 2077 357
rect 2209 349 2275 383
rect 2309 485 2363 527
rect 2309 451 2319 485
rect 2353 451 2363 485
rect 2309 417 2363 451
rect 2309 383 2319 417
rect 2353 383 2363 417
rect 2309 367 2363 383
rect 2397 485 2463 493
rect 2397 428 2413 485
rect 2447 428 2463 485
rect 2397 417 2463 428
rect 2397 383 2413 417
rect 2447 383 2463 417
rect 2209 333 2225 349
rect 2061 323 2225 333
rect 2017 315 2225 323
rect 2259 333 2275 349
rect 2397 349 2463 383
rect 2397 333 2413 349
rect 2259 315 2413 333
rect 2447 315 2463 349
rect 2017 299 2463 315
rect 2497 485 2551 527
rect 2497 451 2507 485
rect 2541 451 2551 485
rect 2497 417 2551 451
rect 2497 383 2507 417
rect 2541 383 2551 417
rect 2497 349 2551 383
rect 2497 315 2507 349
rect 2541 315 2551 349
rect 2497 299 2551 315
rect 2601 485 2655 527
rect 2601 451 2611 485
rect 2645 451 2655 485
rect 2601 417 2655 451
rect 2601 383 2611 417
rect 2645 383 2655 417
rect 2601 349 2655 383
rect 2601 315 2611 349
rect 2645 315 2655 349
rect 2601 299 2655 315
rect 2689 485 2755 493
rect 2689 428 2705 485
rect 2739 428 2755 485
rect 2689 417 2755 428
rect 2689 383 2705 417
rect 2739 383 2755 417
rect 2689 349 2755 383
rect 2789 485 2843 527
rect 2789 451 2799 485
rect 2833 451 2843 485
rect 2789 417 2843 451
rect 2789 383 2799 417
rect 2833 383 2843 417
rect 2789 367 2843 383
rect 2877 485 2943 493
rect 2877 428 2893 485
rect 2927 428 2943 485
rect 2877 417 2943 428
rect 2877 383 2893 417
rect 2927 383 2943 417
rect 2689 315 2705 349
rect 2739 333 2755 349
rect 2877 349 2943 383
rect 2977 485 3031 527
rect 2977 451 2987 485
rect 3021 451 3031 485
rect 2977 417 3031 451
rect 2977 383 2987 417
rect 3021 383 3031 417
rect 2977 367 3031 383
rect 3075 463 3135 493
rect 3075 462 3091 463
rect 3075 428 3089 462
rect 3125 429 3135 463
rect 3123 428 3135 429
rect 2877 333 2893 349
rect 2739 315 2893 333
rect 2927 333 2943 349
rect 3075 357 3135 428
rect 3075 333 3091 357
rect 2927 323 3091 333
rect 3125 323 3135 357
rect 2927 315 3135 323
rect 2689 299 3135 315
rect 3169 463 3235 625
rect 3269 765 3323 781
rect 3269 731 3279 765
rect 3313 731 3323 765
rect 3269 660 3323 731
rect 3269 625 3279 660
rect 3313 625 3323 660
rect 3269 595 3323 625
rect 3357 765 3423 815
rect 3457 859 3694 875
rect 3457 825 3466 859
rect 3500 825 3534 859
rect 3568 825 3694 859
rect 3457 809 3694 825
rect 3728 873 3847 889
rect 3728 839 3731 873
rect 3765 839 3799 873
rect 3833 839 3847 873
rect 3728 823 3847 839
rect 3881 873 4000 889
rect 3881 839 3895 873
rect 3929 839 3963 873
rect 3997 839 4000 873
rect 3881 823 4000 839
rect 4034 875 4068 923
rect 4345 875 4411 935
rect 4613 987 4667 1003
rect 4445 934 4479 953
rect 4513 935 4529 969
rect 4563 935 4579 969
rect 4513 911 4579 935
rect 4647 953 4667 987
rect 4701 1029 4751 1071
rect 4701 995 4717 1029
rect 4701 979 4751 995
rect 4785 1029 4851 1037
rect 4785 995 4801 1029
rect 4835 995 4851 1029
rect 4613 945 4667 953
rect 4785 961 4851 995
rect 4885 1029 4939 1071
rect 4885 995 4895 1029
rect 4929 995 4939 1029
rect 4885 979 4939 995
rect 4973 1029 5039 1037
rect 4973 995 4989 1029
rect 5023 995 5039 1029
rect 4785 945 4801 961
rect 4613 927 4801 945
rect 4835 945 4851 961
rect 4973 961 5039 995
rect 4973 945 4989 961
rect 4835 927 4989 945
rect 5023 927 5039 961
rect 4613 911 5039 927
rect 5073 1029 5123 1071
rect 5107 995 5123 1029
rect 5073 961 5123 995
rect 5107 927 5123 961
rect 5073 911 5123 927
rect 5169 977 5227 1035
rect 5169 943 5181 977
rect 5215 943 5227 977
rect 5169 926 5227 943
rect 5273 1029 5323 1071
rect 5273 995 5289 1029
rect 5273 961 5323 995
rect 5273 927 5289 961
rect 5273 911 5323 927
rect 5357 1029 5423 1037
rect 5357 995 5373 1029
rect 5407 995 5423 1029
rect 5357 961 5423 995
rect 5457 1029 5511 1071
rect 5457 995 5467 1029
rect 5501 995 5511 1029
rect 5457 979 5511 995
rect 5545 1029 5611 1037
rect 5545 995 5561 1029
rect 5595 995 5611 1029
rect 5357 927 5373 961
rect 5407 945 5423 961
rect 5545 961 5611 995
rect 5645 1029 5695 1071
rect 5679 995 5695 1029
rect 5645 979 5695 995
rect 5729 1003 6135 1037
rect 5729 987 5783 1003
rect 5545 945 5561 961
rect 5407 927 5561 945
rect 5595 945 5611 961
rect 5729 953 5749 987
rect 5917 987 5951 1003
rect 5729 945 5783 953
rect 5595 927 5783 945
rect 5357 911 5783 927
rect 5817 935 5833 969
rect 5867 935 5883 969
rect 5817 911 5883 935
rect 6085 987 6135 1003
rect 5917 934 5951 953
rect 5985 935 6001 969
rect 6035 935 6051 969
rect 4513 875 4559 911
rect 4034 859 4271 875
rect 4034 825 4160 859
rect 4194 825 4228 859
rect 4262 825 4271 859
rect 3357 697 3373 765
rect 3407 697 3423 765
rect 3357 659 3423 697
rect 3357 625 3373 659
rect 3407 625 3423 659
rect 3169 429 3185 463
rect 3219 429 3235 463
rect 3169 391 3235 429
rect 3169 323 3185 391
rect 3219 323 3235 391
rect 1729 213 1983 273
rect 3169 273 3235 323
rect 3269 463 3323 493
rect 3269 428 3279 463
rect 3313 428 3323 463
rect 3269 357 3323 428
rect 3269 323 3279 357
rect 3313 323 3323 357
rect 3269 307 3323 323
rect 3357 463 3423 625
rect 3457 759 3517 775
rect 3660 767 3694 809
rect 4034 809 4271 825
rect 4305 815 4559 875
rect 4795 873 5073 877
rect 4795 839 4811 873
rect 4845 839 4879 873
rect 4913 839 4947 873
rect 4981 839 5015 873
rect 5049 839 5073 873
rect 4795 823 5073 839
rect 5323 873 5601 877
rect 5323 839 5347 873
rect 5381 839 5415 873
rect 5449 839 5483 873
rect 5517 839 5551 873
rect 5585 839 5601 873
rect 5323 823 5601 839
rect 5837 875 5883 911
rect 5985 875 6051 935
rect 6119 953 6135 987
rect 6236 1016 6294 1071
rect 6236 982 6260 1016
rect 6236 966 6294 982
rect 6328 1016 6378 1032
rect 6328 982 6344 1016
rect 6085 934 6135 953
rect 6328 923 6378 982
rect 6420 1016 6478 1071
rect 6420 982 6428 1016
rect 6462 982 6478 1016
rect 6420 966 6478 982
rect 6586 1016 6644 1071
rect 6586 982 6602 1016
rect 6636 982 6644 1016
rect 6586 966 6644 982
rect 6686 1016 6736 1032
rect 6720 982 6736 1016
rect 6686 923 6736 982
rect 6770 1016 6828 1071
rect 6804 982 6828 1016
rect 6770 966 6828 982
rect 6929 1003 7335 1037
rect 6929 987 6979 1003
rect 6929 953 6945 987
rect 7113 987 7147 1003
rect 6929 934 6979 953
rect 7013 935 7029 969
rect 7063 935 7079 969
rect 6328 875 6362 923
rect 4034 767 4068 809
rect 3457 725 3467 759
rect 3501 725 3517 759
rect 3457 660 3517 725
rect 3457 659 3469 660
rect 3457 625 3467 659
rect 3503 626 3517 660
rect 3501 625 3517 626
rect 3457 595 3517 625
rect 3566 751 3621 767
rect 3566 717 3582 751
rect 3616 717 3621 751
rect 3566 645 3621 717
rect 3566 611 3582 645
rect 3616 611 3621 645
rect 3566 561 3621 611
rect 3660 751 3726 767
rect 3660 717 3676 751
rect 3710 717 3726 751
rect 3660 645 3726 717
rect 3660 611 3676 645
rect 3710 611 3726 645
rect 3660 595 3726 611
rect 3760 751 3820 767
rect 3760 717 3770 751
rect 3804 717 3820 751
rect 3760 645 3820 717
rect 3760 611 3770 645
rect 3804 611 3820 645
rect 3760 561 3820 611
rect 3908 751 3968 767
rect 3908 717 3924 751
rect 3958 717 3968 751
rect 3908 645 3968 717
rect 3908 611 3924 645
rect 3958 611 3968 645
rect 3908 561 3968 611
rect 4002 751 4068 767
rect 4002 717 4018 751
rect 4052 717 4068 751
rect 4002 645 4068 717
rect 4002 611 4018 645
rect 4052 611 4068 645
rect 4002 595 4068 611
rect 4107 751 4162 767
rect 4107 717 4112 751
rect 4146 717 4162 751
rect 4107 645 4162 717
rect 4107 611 4112 645
rect 4146 611 4162 645
rect 4107 561 4162 611
rect 4211 759 4271 775
rect 4211 725 4227 759
rect 4261 725 4271 759
rect 4211 660 4271 725
rect 4211 626 4225 660
rect 4259 659 4271 660
rect 4211 625 4227 626
rect 4261 625 4271 659
rect 4211 595 4271 625
rect 4305 765 4371 815
rect 4305 697 4321 765
rect 4355 697 4371 765
rect 4305 659 4371 697
rect 4305 625 4321 659
rect 4355 625 4371 659
rect 3457 527 3525 561
rect 3559 527 3617 561
rect 3651 527 3709 561
rect 3743 527 3801 561
rect 3835 527 3893 561
rect 3927 527 3985 561
rect 4019 527 4077 561
rect 4111 527 4169 561
rect 4203 527 4271 561
rect 3357 429 3373 463
rect 3407 429 3423 463
rect 3357 391 3423 429
rect 3357 323 3373 391
rect 3407 323 3423 391
rect 3357 273 3423 323
rect 3457 463 3517 493
rect 3457 429 3467 463
rect 3501 462 3517 463
rect 3457 428 3469 429
rect 3503 428 3517 462
rect 3457 363 3517 428
rect 3457 329 3467 363
rect 3501 329 3517 363
rect 3457 313 3517 329
rect 3566 477 3621 527
rect 3566 443 3582 477
rect 3616 443 3621 477
rect 3566 371 3621 443
rect 3566 337 3582 371
rect 3616 337 3621 371
rect 3566 321 3621 337
rect 3660 477 3726 493
rect 3660 443 3676 477
rect 3710 443 3726 477
rect 3660 371 3726 443
rect 3660 337 3676 371
rect 3710 337 3726 371
rect 3660 321 3726 337
rect 3760 477 3820 527
rect 3760 443 3770 477
rect 3804 443 3820 477
rect 3760 371 3820 443
rect 3760 337 3770 371
rect 3804 337 3820 371
rect 3760 321 3820 337
rect 3908 477 3968 527
rect 3908 443 3924 477
rect 3958 443 3968 477
rect 3908 371 3968 443
rect 3908 337 3924 371
rect 3958 337 3968 371
rect 3908 321 3968 337
rect 4002 477 4068 493
rect 4002 443 4018 477
rect 4052 443 4068 477
rect 4002 371 4068 443
rect 4002 337 4018 371
rect 4052 337 4068 371
rect 4002 321 4068 337
rect 4107 477 4162 527
rect 4107 443 4112 477
rect 4146 443 4162 477
rect 4107 371 4162 443
rect 4107 337 4112 371
rect 4146 337 4162 371
rect 4107 321 4162 337
rect 4211 463 4271 493
rect 4211 462 4227 463
rect 4211 428 4225 462
rect 4261 429 4271 463
rect 4259 428 4271 429
rect 4211 363 4271 428
rect 4211 329 4227 363
rect 4261 329 4271 363
rect 3660 279 3694 321
rect 1458 165 1492 213
rect 741 119 757 153
rect 791 119 807 153
rect 841 135 891 154
rect 673 85 707 101
rect 875 101 891 135
rect 841 85 891 101
rect 485 51 891 85
rect 992 106 1050 122
rect 992 72 1016 106
rect 992 17 1050 72
rect 1084 106 1134 165
rect 1084 72 1100 106
rect 1084 56 1134 72
rect 1176 106 1234 122
rect 1176 72 1184 106
rect 1218 72 1234 106
rect 1176 17 1234 72
rect 1342 106 1400 122
rect 1342 72 1358 106
rect 1392 72 1400 106
rect 1342 17 1400 72
rect 1442 106 1492 165
rect 1685 135 1735 154
rect 1476 72 1492 106
rect 1442 56 1492 72
rect 1526 106 1584 122
rect 1560 72 1584 106
rect 1526 17 1584 72
rect 1685 101 1701 135
rect 1769 153 1835 213
rect 1937 177 1983 213
rect 2219 249 2497 265
rect 2219 215 2235 249
rect 2269 215 2303 249
rect 2337 215 2371 249
rect 2405 215 2439 249
rect 2473 215 2497 249
rect 2219 211 2497 215
rect 2655 249 2933 265
rect 2655 215 2679 249
rect 2713 215 2747 249
rect 2781 215 2815 249
rect 2849 215 2883 249
rect 2917 215 2933 249
rect 2655 211 2933 215
rect 3169 213 3423 273
rect 3457 263 3694 279
rect 4034 279 4068 321
rect 4211 313 4271 329
rect 4305 463 4371 625
rect 4405 765 4459 781
rect 4405 731 4415 765
rect 4449 731 4459 765
rect 4405 660 4459 731
rect 4405 625 4415 660
rect 4449 625 4459 660
rect 4405 595 4459 625
rect 4493 765 4559 815
rect 5837 815 6091 875
rect 4493 697 4509 765
rect 4543 697 4559 765
rect 4493 659 4559 697
rect 4493 625 4509 659
rect 4543 625 4559 659
rect 4305 429 4321 463
rect 4355 429 4371 463
rect 4305 391 4371 429
rect 4305 323 4321 391
rect 4355 323 4371 391
rect 3457 229 3466 263
rect 3500 229 3534 263
rect 3568 229 3694 263
rect 3457 213 3694 229
rect 3169 177 3215 213
rect 1769 119 1785 153
rect 1819 119 1835 153
rect 1869 135 1903 154
rect 1685 85 1735 101
rect 1937 153 2003 177
rect 1937 119 1953 153
rect 1987 119 2003 153
rect 2037 161 2463 177
rect 2037 143 2225 161
rect 2037 135 2091 143
rect 1869 85 1903 101
rect 2071 101 2091 135
rect 2209 127 2225 143
rect 2259 143 2413 161
rect 2259 127 2275 143
rect 2037 85 2091 101
rect 1685 51 2091 85
rect 2125 93 2175 109
rect 2125 59 2141 93
rect 2125 17 2175 59
rect 2209 93 2275 127
rect 2397 127 2413 143
rect 2447 127 2463 161
rect 2209 59 2225 93
rect 2259 59 2275 93
rect 2209 51 2275 59
rect 2309 93 2363 109
rect 2309 59 2319 93
rect 2353 59 2363 93
rect 2309 17 2363 59
rect 2397 93 2463 127
rect 2397 59 2413 93
rect 2447 59 2463 93
rect 2397 51 2463 59
rect 2497 161 2547 177
rect 2531 127 2547 161
rect 2497 93 2547 127
rect 2531 59 2547 93
rect 2497 17 2547 59
rect 2605 161 2655 177
rect 2605 127 2621 161
rect 2605 93 2655 127
rect 2605 59 2621 93
rect 2605 17 2655 59
rect 2689 161 3115 177
rect 2689 127 2705 161
rect 2739 143 2893 161
rect 2739 127 2755 143
rect 2689 93 2755 127
rect 2877 127 2893 143
rect 2927 143 3115 161
rect 2927 127 2943 143
rect 2689 59 2705 93
rect 2739 59 2755 93
rect 2689 51 2755 59
rect 2789 93 2843 109
rect 2789 59 2799 93
rect 2833 59 2843 93
rect 2789 17 2843 59
rect 2877 93 2943 127
rect 3061 135 3115 143
rect 2877 59 2893 93
rect 2927 59 2943 93
rect 2877 51 2943 59
rect 2977 93 3027 109
rect 3011 59 3027 93
rect 2977 17 3027 59
rect 3061 101 3081 135
rect 3149 153 3215 177
rect 3149 119 3165 153
rect 3199 119 3215 153
rect 3249 135 3283 154
rect 3061 85 3115 101
rect 3317 153 3383 213
rect 3660 165 3694 213
rect 3728 249 3847 265
rect 3728 215 3731 249
rect 3765 215 3799 249
rect 3833 215 3847 249
rect 3728 199 3847 215
rect 3881 249 4000 265
rect 3881 215 3895 249
rect 3929 215 3963 249
rect 3997 215 4000 249
rect 3881 199 4000 215
rect 4034 263 4271 279
rect 4034 229 4160 263
rect 4194 229 4228 263
rect 4262 229 4271 263
rect 4034 213 4271 229
rect 4305 273 4371 323
rect 4405 463 4459 493
rect 4405 428 4415 463
rect 4449 428 4459 463
rect 4405 357 4459 428
rect 4405 323 4415 357
rect 4449 323 4459 357
rect 4405 307 4459 323
rect 4493 463 4559 625
rect 4593 773 5039 789
rect 4593 765 4801 773
rect 4593 731 4603 765
rect 4637 755 4801 765
rect 4637 731 4653 755
rect 4593 660 4653 731
rect 4785 739 4801 755
rect 4835 755 4989 773
rect 4835 739 4851 755
rect 4593 659 4605 660
rect 4593 625 4603 659
rect 4639 626 4653 660
rect 4637 625 4653 626
rect 4593 595 4653 625
rect 4697 705 4751 721
rect 4697 671 4707 705
rect 4741 671 4751 705
rect 4697 637 4751 671
rect 4697 603 4707 637
rect 4741 603 4751 637
rect 4697 561 4751 603
rect 4785 705 4851 739
rect 4973 739 4989 755
rect 5023 739 5039 773
rect 4785 671 4801 705
rect 4835 671 4851 705
rect 4785 660 4851 671
rect 4785 603 4801 660
rect 4835 603 4851 660
rect 4785 595 4851 603
rect 4885 705 4939 721
rect 4885 671 4895 705
rect 4929 671 4939 705
rect 4885 637 4939 671
rect 4885 603 4895 637
rect 4929 603 4939 637
rect 4885 561 4939 603
rect 4973 705 5039 739
rect 4973 671 4989 705
rect 5023 671 5039 705
rect 4973 660 5039 671
rect 4973 603 4989 660
rect 5023 603 5039 660
rect 4973 595 5039 603
rect 5073 773 5127 789
rect 5073 739 5083 773
rect 5117 739 5127 773
rect 5073 705 5127 739
rect 5073 671 5083 705
rect 5117 671 5127 705
rect 5073 637 5127 671
rect 5073 603 5083 637
rect 5117 603 5127 637
rect 5073 561 5127 603
rect 5169 759 5227 794
rect 5169 725 5181 759
rect 5215 725 5227 759
rect 5169 675 5227 725
rect 5169 641 5181 675
rect 5215 641 5227 675
rect 5169 597 5227 641
rect 5269 773 5323 789
rect 5269 739 5279 773
rect 5313 739 5323 773
rect 5269 705 5323 739
rect 5269 671 5279 705
rect 5313 671 5323 705
rect 5269 637 5323 671
rect 5269 603 5279 637
rect 5313 603 5323 637
rect 5269 561 5323 603
rect 5357 773 5803 789
rect 5357 739 5373 773
rect 5407 755 5561 773
rect 5407 739 5423 755
rect 5357 705 5423 739
rect 5545 739 5561 755
rect 5595 765 5803 773
rect 5595 755 5759 765
rect 5595 739 5611 755
rect 5357 671 5373 705
rect 5407 671 5423 705
rect 5357 660 5423 671
rect 5357 603 5373 660
rect 5407 603 5423 660
rect 5357 595 5423 603
rect 5457 705 5511 721
rect 5457 671 5467 705
rect 5501 671 5511 705
rect 5457 637 5511 671
rect 5457 603 5467 637
rect 5501 603 5511 637
rect 5457 561 5511 603
rect 5545 705 5611 739
rect 5743 731 5759 755
rect 5793 731 5803 765
rect 5545 671 5561 705
rect 5595 671 5611 705
rect 5545 660 5611 671
rect 5545 603 5561 660
rect 5595 603 5611 660
rect 5545 595 5611 603
rect 5645 705 5699 721
rect 5645 671 5655 705
rect 5689 671 5699 705
rect 5645 637 5699 671
rect 5645 603 5655 637
rect 5689 603 5699 637
rect 5645 561 5699 603
rect 5743 660 5803 731
rect 5743 626 5757 660
rect 5791 659 5803 660
rect 5743 625 5759 626
rect 5793 625 5803 659
rect 5743 595 5803 625
rect 5837 765 5903 815
rect 5837 697 5853 765
rect 5887 697 5903 765
rect 5837 659 5903 697
rect 5837 625 5853 659
rect 5887 625 5903 659
rect 4593 527 4629 561
rect 4663 527 4721 561
rect 4755 527 4813 561
rect 4847 527 4905 561
rect 4939 527 4997 561
rect 5031 527 5089 561
rect 5123 527 5181 561
rect 5215 527 5273 561
rect 5307 527 5365 561
rect 5399 527 5457 561
rect 5491 527 5549 561
rect 5583 527 5641 561
rect 5675 527 5733 561
rect 5767 527 5803 561
rect 4493 429 4509 463
rect 4543 429 4559 463
rect 4493 391 4559 429
rect 4493 323 4509 391
rect 4543 323 4559 391
rect 4493 273 4559 323
rect 4593 463 4653 493
rect 4593 429 4603 463
rect 4637 462 4653 463
rect 4593 428 4605 429
rect 4639 428 4653 462
rect 4593 357 4653 428
rect 4697 485 4751 527
rect 4697 451 4707 485
rect 4741 451 4751 485
rect 4697 417 4751 451
rect 4697 383 4707 417
rect 4741 383 4751 417
rect 4697 367 4751 383
rect 4785 485 4851 493
rect 4785 428 4801 485
rect 4835 428 4851 485
rect 4785 417 4851 428
rect 4785 383 4801 417
rect 4835 383 4851 417
rect 4593 323 4603 357
rect 4637 333 4653 357
rect 4785 349 4851 383
rect 4885 485 4939 527
rect 4885 451 4895 485
rect 4929 451 4939 485
rect 4885 417 4939 451
rect 4885 383 4895 417
rect 4929 383 4939 417
rect 4885 367 4939 383
rect 4973 485 5039 493
rect 4973 428 4989 485
rect 5023 428 5039 485
rect 4973 417 5039 428
rect 4973 383 4989 417
rect 5023 383 5039 417
rect 4785 333 4801 349
rect 4637 323 4801 333
rect 4593 315 4801 323
rect 4835 333 4851 349
rect 4973 349 5039 383
rect 4973 333 4989 349
rect 4835 315 4989 333
rect 5023 315 5039 349
rect 4593 299 5039 315
rect 5073 485 5127 527
rect 5073 451 5083 485
rect 5117 451 5127 485
rect 5073 417 5127 451
rect 5073 383 5083 417
rect 5117 383 5127 417
rect 5073 349 5127 383
rect 5073 315 5083 349
rect 5117 315 5127 349
rect 5073 299 5127 315
rect 5169 447 5227 491
rect 5169 413 5181 447
rect 5215 413 5227 447
rect 5169 363 5227 413
rect 5169 329 5181 363
rect 5215 329 5227 363
rect 5169 294 5227 329
rect 5269 485 5323 527
rect 5269 451 5279 485
rect 5313 451 5323 485
rect 5269 417 5323 451
rect 5269 383 5279 417
rect 5313 383 5323 417
rect 5269 349 5323 383
rect 5269 315 5279 349
rect 5313 315 5323 349
rect 5269 299 5323 315
rect 5357 485 5423 493
rect 5357 428 5373 485
rect 5407 428 5423 485
rect 5357 417 5423 428
rect 5357 383 5373 417
rect 5407 383 5423 417
rect 5357 349 5423 383
rect 5457 485 5511 527
rect 5457 451 5467 485
rect 5501 451 5511 485
rect 5457 417 5511 451
rect 5457 383 5467 417
rect 5501 383 5511 417
rect 5457 367 5511 383
rect 5545 485 5611 493
rect 5545 428 5561 485
rect 5595 428 5611 485
rect 5545 417 5611 428
rect 5545 383 5561 417
rect 5595 383 5611 417
rect 5357 315 5373 349
rect 5407 333 5423 349
rect 5545 349 5611 383
rect 5645 485 5699 527
rect 5645 451 5655 485
rect 5689 451 5699 485
rect 5645 417 5699 451
rect 5645 383 5655 417
rect 5689 383 5699 417
rect 5645 367 5699 383
rect 5743 463 5803 493
rect 5743 462 5759 463
rect 5743 428 5757 462
rect 5793 429 5803 463
rect 5791 428 5803 429
rect 5545 333 5561 349
rect 5407 315 5561 333
rect 5595 333 5611 349
rect 5743 357 5803 428
rect 5743 333 5759 357
rect 5595 323 5759 333
rect 5793 323 5803 357
rect 5595 315 5803 323
rect 5357 299 5803 315
rect 5837 463 5903 625
rect 5937 765 5991 781
rect 5937 731 5947 765
rect 5981 731 5991 765
rect 5937 660 5991 731
rect 5937 625 5947 660
rect 5981 625 5991 660
rect 5937 595 5991 625
rect 6025 765 6091 815
rect 6125 859 6362 875
rect 6125 825 6134 859
rect 6168 825 6202 859
rect 6236 825 6362 859
rect 6125 809 6362 825
rect 6396 873 6515 889
rect 6396 839 6399 873
rect 6433 839 6467 873
rect 6501 839 6515 873
rect 6396 823 6515 839
rect 6549 873 6668 889
rect 6549 839 6563 873
rect 6597 839 6631 873
rect 6665 839 6668 873
rect 6549 823 6668 839
rect 6702 875 6736 923
rect 7013 875 7079 935
rect 7281 987 7335 1003
rect 7113 934 7147 953
rect 7181 935 7197 969
rect 7231 935 7247 969
rect 7181 911 7247 935
rect 7315 953 7335 987
rect 7369 1029 7419 1071
rect 7369 995 7385 1029
rect 7369 979 7419 995
rect 7453 1029 7519 1037
rect 7453 995 7469 1029
rect 7503 995 7519 1029
rect 7281 945 7335 953
rect 7453 961 7519 995
rect 7553 1029 7607 1071
rect 7553 995 7563 1029
rect 7597 995 7607 1029
rect 7553 979 7607 995
rect 7641 1029 7707 1037
rect 7641 995 7657 1029
rect 7691 995 7707 1029
rect 7453 945 7469 961
rect 7281 927 7469 945
rect 7503 945 7519 961
rect 7641 961 7707 995
rect 7641 945 7657 961
rect 7503 927 7657 945
rect 7691 927 7707 961
rect 7281 911 7707 927
rect 7741 1029 7791 1071
rect 7775 995 7791 1029
rect 7741 961 7791 995
rect 7775 927 7791 961
rect 7741 911 7791 927
rect 7849 1029 7899 1071
rect 7849 995 7865 1029
rect 7849 961 7899 995
rect 7849 927 7865 961
rect 7849 911 7899 927
rect 7933 1029 7999 1037
rect 7933 995 7949 1029
rect 7983 995 7999 1029
rect 7933 961 7999 995
rect 8033 1029 8087 1071
rect 8033 995 8043 1029
rect 8077 995 8087 1029
rect 8033 979 8087 995
rect 8121 1029 8187 1037
rect 8121 995 8137 1029
rect 8171 995 8187 1029
rect 7933 927 7949 961
rect 7983 945 7999 961
rect 8121 961 8187 995
rect 8221 1029 8271 1071
rect 8255 995 8271 1029
rect 8221 979 8271 995
rect 8305 1003 8711 1037
rect 8305 987 8359 1003
rect 8121 945 8137 961
rect 7983 927 8137 945
rect 8171 945 8187 961
rect 8305 953 8325 987
rect 8493 987 8527 1003
rect 8305 945 8359 953
rect 8171 927 8359 945
rect 7933 911 8359 927
rect 8393 935 8409 969
rect 8443 935 8459 969
rect 8393 911 8459 935
rect 8661 987 8711 1003
rect 8493 934 8527 953
rect 8561 935 8577 969
rect 8611 935 8627 969
rect 7181 875 7227 911
rect 6702 859 6939 875
rect 6702 825 6828 859
rect 6862 825 6896 859
rect 6930 825 6939 859
rect 6025 697 6041 765
rect 6075 697 6091 765
rect 6025 659 6091 697
rect 6025 625 6041 659
rect 6075 625 6091 659
rect 5837 429 5853 463
rect 5887 429 5903 463
rect 5837 391 5903 429
rect 5837 323 5853 391
rect 5887 323 5903 391
rect 4305 213 4559 273
rect 5837 273 5903 323
rect 5937 463 5991 493
rect 5937 428 5947 463
rect 5981 428 5991 463
rect 5937 357 5991 428
rect 5937 323 5947 357
rect 5981 323 5991 357
rect 5937 307 5991 323
rect 6025 463 6091 625
rect 6125 759 6185 775
rect 6328 767 6362 809
rect 6702 809 6939 825
rect 6973 815 7227 875
rect 7463 873 7741 877
rect 7463 839 7479 873
rect 7513 839 7547 873
rect 7581 839 7615 873
rect 7649 839 7683 873
rect 7717 839 7741 873
rect 7463 823 7741 839
rect 7899 873 8177 877
rect 7899 839 7923 873
rect 7957 839 7991 873
rect 8025 839 8059 873
rect 8093 839 8127 873
rect 8161 839 8177 873
rect 7899 823 8177 839
rect 8413 875 8459 911
rect 8561 875 8627 935
rect 8695 953 8711 987
rect 8812 1016 8870 1071
rect 8812 982 8836 1016
rect 8812 966 8870 982
rect 8904 1016 8954 1032
rect 8904 982 8920 1016
rect 8661 934 8711 953
rect 8904 923 8954 982
rect 8996 1016 9054 1071
rect 8996 982 9004 1016
rect 9038 982 9054 1016
rect 8996 966 9054 982
rect 9162 1016 9220 1071
rect 9162 982 9178 1016
rect 9212 982 9220 1016
rect 9162 966 9220 982
rect 9262 1016 9312 1032
rect 9296 982 9312 1016
rect 9262 923 9312 982
rect 9346 1016 9404 1071
rect 9380 982 9404 1016
rect 9346 966 9404 982
rect 9505 1003 9911 1037
rect 9505 987 9555 1003
rect 9505 953 9521 987
rect 9689 987 9723 1003
rect 9505 934 9555 953
rect 9589 935 9605 969
rect 9639 935 9655 969
rect 8904 875 8938 923
rect 6702 767 6736 809
rect 6125 725 6135 759
rect 6169 725 6185 759
rect 6125 660 6185 725
rect 6125 659 6137 660
rect 6125 625 6135 659
rect 6171 626 6185 660
rect 6169 625 6185 626
rect 6125 595 6185 625
rect 6234 751 6289 767
rect 6234 717 6250 751
rect 6284 717 6289 751
rect 6234 645 6289 717
rect 6234 611 6250 645
rect 6284 611 6289 645
rect 6234 561 6289 611
rect 6328 751 6394 767
rect 6328 717 6344 751
rect 6378 717 6394 751
rect 6328 645 6394 717
rect 6328 611 6344 645
rect 6378 611 6394 645
rect 6328 595 6394 611
rect 6428 751 6488 767
rect 6428 717 6438 751
rect 6472 717 6488 751
rect 6428 645 6488 717
rect 6428 611 6438 645
rect 6472 611 6488 645
rect 6428 561 6488 611
rect 6576 751 6636 767
rect 6576 717 6592 751
rect 6626 717 6636 751
rect 6576 645 6636 717
rect 6576 611 6592 645
rect 6626 611 6636 645
rect 6576 561 6636 611
rect 6670 751 6736 767
rect 6670 717 6686 751
rect 6720 717 6736 751
rect 6670 645 6736 717
rect 6670 611 6686 645
rect 6720 611 6736 645
rect 6670 595 6736 611
rect 6775 751 6830 767
rect 6775 717 6780 751
rect 6814 717 6830 751
rect 6775 645 6830 717
rect 6775 611 6780 645
rect 6814 611 6830 645
rect 6775 561 6830 611
rect 6879 759 6939 775
rect 6879 725 6895 759
rect 6929 725 6939 759
rect 6879 660 6939 725
rect 6879 626 6893 660
rect 6927 659 6939 660
rect 6879 625 6895 626
rect 6929 625 6939 659
rect 6879 595 6939 625
rect 6973 765 7039 815
rect 6973 697 6989 765
rect 7023 697 7039 765
rect 6973 659 7039 697
rect 6973 625 6989 659
rect 7023 625 7039 659
rect 6125 527 6193 561
rect 6227 527 6285 561
rect 6319 527 6377 561
rect 6411 527 6469 561
rect 6503 527 6561 561
rect 6595 527 6653 561
rect 6687 527 6745 561
rect 6779 527 6837 561
rect 6871 527 6939 561
rect 6025 429 6041 463
rect 6075 429 6091 463
rect 6025 391 6091 429
rect 6025 323 6041 391
rect 6075 323 6091 391
rect 6025 273 6091 323
rect 6125 463 6185 493
rect 6125 429 6135 463
rect 6169 462 6185 463
rect 6125 428 6137 429
rect 6171 428 6185 462
rect 6125 363 6185 428
rect 6125 329 6135 363
rect 6169 329 6185 363
rect 6125 313 6185 329
rect 6234 477 6289 527
rect 6234 443 6250 477
rect 6284 443 6289 477
rect 6234 371 6289 443
rect 6234 337 6250 371
rect 6284 337 6289 371
rect 6234 321 6289 337
rect 6328 477 6394 493
rect 6328 443 6344 477
rect 6378 443 6394 477
rect 6328 371 6394 443
rect 6328 337 6344 371
rect 6378 337 6394 371
rect 6328 321 6394 337
rect 6428 477 6488 527
rect 6428 443 6438 477
rect 6472 443 6488 477
rect 6428 371 6488 443
rect 6428 337 6438 371
rect 6472 337 6488 371
rect 6428 321 6488 337
rect 6576 477 6636 527
rect 6576 443 6592 477
rect 6626 443 6636 477
rect 6576 371 6636 443
rect 6576 337 6592 371
rect 6626 337 6636 371
rect 6576 321 6636 337
rect 6670 477 6736 493
rect 6670 443 6686 477
rect 6720 443 6736 477
rect 6670 371 6736 443
rect 6670 337 6686 371
rect 6720 337 6736 371
rect 6670 321 6736 337
rect 6775 477 6830 527
rect 6775 443 6780 477
rect 6814 443 6830 477
rect 6775 371 6830 443
rect 6775 337 6780 371
rect 6814 337 6830 371
rect 6775 321 6830 337
rect 6879 463 6939 493
rect 6879 462 6895 463
rect 6879 428 6893 462
rect 6929 429 6939 463
rect 6927 428 6939 429
rect 6879 363 6939 428
rect 6879 329 6895 363
rect 6929 329 6939 363
rect 6328 279 6362 321
rect 4034 165 4068 213
rect 3317 119 3333 153
rect 3367 119 3383 153
rect 3417 135 3467 154
rect 3249 85 3283 101
rect 3451 101 3467 135
rect 3417 85 3467 101
rect 3061 51 3467 85
rect 3568 106 3626 122
rect 3568 72 3592 106
rect 3568 17 3626 72
rect 3660 106 3710 165
rect 3660 72 3676 106
rect 3660 56 3710 72
rect 3752 106 3810 122
rect 3752 72 3760 106
rect 3794 72 3810 106
rect 3752 17 3810 72
rect 3918 106 3976 122
rect 3918 72 3934 106
rect 3968 72 3976 106
rect 3918 17 3976 72
rect 4018 106 4068 165
rect 4261 135 4311 154
rect 4052 72 4068 106
rect 4018 56 4068 72
rect 4102 106 4160 122
rect 4136 72 4160 106
rect 4102 17 4160 72
rect 4261 101 4277 135
rect 4345 153 4411 213
rect 4513 177 4559 213
rect 4795 249 5073 265
rect 4795 215 4811 249
rect 4845 215 4879 249
rect 4913 215 4947 249
rect 4981 215 5015 249
rect 5049 215 5073 249
rect 4795 211 5073 215
rect 5323 249 5601 265
rect 5323 215 5347 249
rect 5381 215 5415 249
rect 5449 215 5483 249
rect 5517 215 5551 249
rect 5585 215 5601 249
rect 5323 211 5601 215
rect 5837 213 6091 273
rect 6125 263 6362 279
rect 6702 279 6736 321
rect 6879 313 6939 329
rect 6973 463 7039 625
rect 7073 765 7127 781
rect 7073 731 7083 765
rect 7117 731 7127 765
rect 7073 660 7127 731
rect 7073 625 7083 660
rect 7117 625 7127 660
rect 7073 595 7127 625
rect 7161 765 7227 815
rect 8413 815 8667 875
rect 7161 697 7177 765
rect 7211 697 7227 765
rect 7161 659 7227 697
rect 7161 625 7177 659
rect 7211 625 7227 659
rect 6973 429 6989 463
rect 7023 429 7039 463
rect 6973 391 7039 429
rect 6973 323 6989 391
rect 7023 323 7039 391
rect 6125 229 6134 263
rect 6168 229 6202 263
rect 6236 229 6362 263
rect 6125 213 6362 229
rect 5837 177 5883 213
rect 4345 119 4361 153
rect 4395 119 4411 153
rect 4445 135 4479 154
rect 4261 85 4311 101
rect 4513 153 4579 177
rect 4513 119 4529 153
rect 4563 119 4579 153
rect 4613 161 5039 177
rect 4613 143 4801 161
rect 4613 135 4667 143
rect 4445 85 4479 101
rect 4647 101 4667 135
rect 4785 127 4801 143
rect 4835 143 4989 161
rect 4835 127 4851 143
rect 4613 85 4667 101
rect 4261 51 4667 85
rect 4701 93 4751 109
rect 4701 59 4717 93
rect 4701 17 4751 59
rect 4785 93 4851 127
rect 4973 127 4989 143
rect 5023 127 5039 161
rect 4785 59 4801 93
rect 4835 59 4851 93
rect 4785 51 4851 59
rect 4885 93 4939 109
rect 4885 59 4895 93
rect 4929 59 4939 93
rect 4885 17 4939 59
rect 4973 93 5039 127
rect 4973 59 4989 93
rect 5023 59 5039 93
rect 4973 51 5039 59
rect 5073 161 5123 177
rect 5107 127 5123 161
rect 5073 93 5123 127
rect 5107 59 5123 93
rect 5073 17 5123 59
rect 5169 145 5227 162
rect 5169 111 5181 145
rect 5215 111 5227 145
rect 5169 53 5227 111
rect 5273 161 5323 177
rect 5273 127 5289 161
rect 5273 93 5323 127
rect 5273 59 5289 93
rect 5273 17 5323 59
rect 5357 161 5783 177
rect 5357 127 5373 161
rect 5407 143 5561 161
rect 5407 127 5423 143
rect 5357 93 5423 127
rect 5545 127 5561 143
rect 5595 143 5783 161
rect 5595 127 5611 143
rect 5357 59 5373 93
rect 5407 59 5423 93
rect 5357 51 5423 59
rect 5457 93 5511 109
rect 5457 59 5467 93
rect 5501 59 5511 93
rect 5457 17 5511 59
rect 5545 93 5611 127
rect 5729 135 5783 143
rect 5545 59 5561 93
rect 5595 59 5611 93
rect 5545 51 5611 59
rect 5645 93 5695 109
rect 5679 59 5695 93
rect 5645 17 5695 59
rect 5729 101 5749 135
rect 5817 153 5883 177
rect 5817 119 5833 153
rect 5867 119 5883 153
rect 5917 135 5951 154
rect 5729 85 5783 101
rect 5985 153 6051 213
rect 6328 165 6362 213
rect 6396 249 6515 265
rect 6396 215 6399 249
rect 6433 215 6467 249
rect 6501 215 6515 249
rect 6396 199 6515 215
rect 6549 249 6668 265
rect 6549 215 6563 249
rect 6597 215 6631 249
rect 6665 215 6668 249
rect 6549 199 6668 215
rect 6702 263 6939 279
rect 6702 229 6828 263
rect 6862 229 6896 263
rect 6930 229 6939 263
rect 6702 213 6939 229
rect 6973 273 7039 323
rect 7073 463 7127 493
rect 7073 428 7083 463
rect 7117 428 7127 463
rect 7073 357 7127 428
rect 7073 323 7083 357
rect 7117 323 7127 357
rect 7073 307 7127 323
rect 7161 463 7227 625
rect 7261 773 7707 789
rect 7261 765 7469 773
rect 7261 731 7271 765
rect 7305 755 7469 765
rect 7305 731 7321 755
rect 7261 660 7321 731
rect 7453 739 7469 755
rect 7503 755 7657 773
rect 7503 739 7519 755
rect 7261 659 7273 660
rect 7261 625 7271 659
rect 7307 626 7321 660
rect 7305 625 7321 626
rect 7261 595 7321 625
rect 7365 705 7419 721
rect 7365 671 7375 705
rect 7409 671 7419 705
rect 7365 637 7419 671
rect 7365 603 7375 637
rect 7409 603 7419 637
rect 7365 561 7419 603
rect 7453 705 7519 739
rect 7641 739 7657 755
rect 7691 739 7707 773
rect 7453 671 7469 705
rect 7503 671 7519 705
rect 7453 660 7519 671
rect 7453 603 7469 660
rect 7503 603 7519 660
rect 7453 595 7519 603
rect 7553 705 7607 721
rect 7553 671 7563 705
rect 7597 671 7607 705
rect 7553 637 7607 671
rect 7553 603 7563 637
rect 7597 603 7607 637
rect 7553 561 7607 603
rect 7641 705 7707 739
rect 7641 671 7657 705
rect 7691 671 7707 705
rect 7641 660 7707 671
rect 7641 603 7657 660
rect 7691 603 7707 660
rect 7641 595 7707 603
rect 7741 773 7795 789
rect 7741 739 7751 773
rect 7785 739 7795 773
rect 7741 705 7795 739
rect 7741 671 7751 705
rect 7785 671 7795 705
rect 7741 637 7795 671
rect 7741 603 7751 637
rect 7785 603 7795 637
rect 7741 561 7795 603
rect 7845 773 7899 789
rect 7845 739 7855 773
rect 7889 739 7899 773
rect 7845 705 7899 739
rect 7845 671 7855 705
rect 7889 671 7899 705
rect 7845 637 7899 671
rect 7845 603 7855 637
rect 7889 603 7899 637
rect 7845 561 7899 603
rect 7933 773 8379 789
rect 7933 739 7949 773
rect 7983 755 8137 773
rect 7983 739 7999 755
rect 7933 705 7999 739
rect 8121 739 8137 755
rect 8171 765 8379 773
rect 8171 755 8335 765
rect 8171 739 8187 755
rect 7933 671 7949 705
rect 7983 671 7999 705
rect 7933 660 7999 671
rect 7933 603 7949 660
rect 7983 603 7999 660
rect 7933 595 7999 603
rect 8033 705 8087 721
rect 8033 671 8043 705
rect 8077 671 8087 705
rect 8033 637 8087 671
rect 8033 603 8043 637
rect 8077 603 8087 637
rect 8033 561 8087 603
rect 8121 705 8187 739
rect 8319 731 8335 755
rect 8369 731 8379 765
rect 8121 671 8137 705
rect 8171 671 8187 705
rect 8121 660 8187 671
rect 8121 603 8137 660
rect 8171 603 8187 660
rect 8121 595 8187 603
rect 8221 705 8275 721
rect 8221 671 8231 705
rect 8265 671 8275 705
rect 8221 637 8275 671
rect 8221 603 8231 637
rect 8265 603 8275 637
rect 8221 561 8275 603
rect 8319 660 8379 731
rect 8319 626 8333 660
rect 8367 659 8379 660
rect 8319 625 8335 626
rect 8369 625 8379 659
rect 8319 595 8379 625
rect 8413 765 8479 815
rect 8413 697 8429 765
rect 8463 697 8479 765
rect 8413 659 8479 697
rect 8413 625 8429 659
rect 8463 625 8479 659
rect 7261 527 7297 561
rect 7331 527 7389 561
rect 7423 527 7481 561
rect 7515 527 7573 561
rect 7607 527 7665 561
rect 7699 527 7757 561
rect 7791 527 7849 561
rect 7883 527 7941 561
rect 7975 527 8033 561
rect 8067 527 8125 561
rect 8159 527 8217 561
rect 8251 527 8309 561
rect 8343 527 8379 561
rect 7161 429 7177 463
rect 7211 429 7227 463
rect 7161 391 7227 429
rect 7161 323 7177 391
rect 7211 323 7227 391
rect 7161 273 7227 323
rect 7261 463 7321 493
rect 7261 429 7271 463
rect 7305 462 7321 463
rect 7261 428 7273 429
rect 7307 428 7321 462
rect 7261 357 7321 428
rect 7365 485 7419 527
rect 7365 451 7375 485
rect 7409 451 7419 485
rect 7365 417 7419 451
rect 7365 383 7375 417
rect 7409 383 7419 417
rect 7365 367 7419 383
rect 7453 485 7519 493
rect 7453 428 7469 485
rect 7503 428 7519 485
rect 7453 417 7519 428
rect 7453 383 7469 417
rect 7503 383 7519 417
rect 7261 323 7271 357
rect 7305 333 7321 357
rect 7453 349 7519 383
rect 7553 485 7607 527
rect 7553 451 7563 485
rect 7597 451 7607 485
rect 7553 417 7607 451
rect 7553 383 7563 417
rect 7597 383 7607 417
rect 7553 367 7607 383
rect 7641 485 7707 493
rect 7641 428 7657 485
rect 7691 428 7707 485
rect 7641 417 7707 428
rect 7641 383 7657 417
rect 7691 383 7707 417
rect 7453 333 7469 349
rect 7305 323 7469 333
rect 7261 315 7469 323
rect 7503 333 7519 349
rect 7641 349 7707 383
rect 7641 333 7657 349
rect 7503 315 7657 333
rect 7691 315 7707 349
rect 7261 299 7707 315
rect 7741 485 7795 527
rect 7741 451 7751 485
rect 7785 451 7795 485
rect 7741 417 7795 451
rect 7741 383 7751 417
rect 7785 383 7795 417
rect 7741 349 7795 383
rect 7741 315 7751 349
rect 7785 315 7795 349
rect 7741 299 7795 315
rect 7845 485 7899 527
rect 7845 451 7855 485
rect 7889 451 7899 485
rect 7845 417 7899 451
rect 7845 383 7855 417
rect 7889 383 7899 417
rect 7845 349 7899 383
rect 7845 315 7855 349
rect 7889 315 7899 349
rect 7845 299 7899 315
rect 7933 485 7999 493
rect 7933 428 7949 485
rect 7983 428 7999 485
rect 7933 417 7999 428
rect 7933 383 7949 417
rect 7983 383 7999 417
rect 7933 349 7999 383
rect 8033 485 8087 527
rect 8033 451 8043 485
rect 8077 451 8087 485
rect 8033 417 8087 451
rect 8033 383 8043 417
rect 8077 383 8087 417
rect 8033 367 8087 383
rect 8121 485 8187 493
rect 8121 428 8137 485
rect 8171 428 8187 485
rect 8121 417 8187 428
rect 8121 383 8137 417
rect 8171 383 8187 417
rect 7933 315 7949 349
rect 7983 333 7999 349
rect 8121 349 8187 383
rect 8221 485 8275 527
rect 8221 451 8231 485
rect 8265 451 8275 485
rect 8221 417 8275 451
rect 8221 383 8231 417
rect 8265 383 8275 417
rect 8221 367 8275 383
rect 8319 463 8379 493
rect 8319 462 8335 463
rect 8319 428 8333 462
rect 8369 429 8379 463
rect 8367 428 8379 429
rect 8121 333 8137 349
rect 7983 315 8137 333
rect 8171 333 8187 349
rect 8319 357 8379 428
rect 8319 333 8335 357
rect 8171 323 8335 333
rect 8369 323 8379 357
rect 8171 315 8379 323
rect 7933 299 8379 315
rect 8413 463 8479 625
rect 8513 765 8567 781
rect 8513 731 8523 765
rect 8557 731 8567 765
rect 8513 660 8567 731
rect 8513 625 8523 660
rect 8557 625 8567 660
rect 8513 595 8567 625
rect 8601 765 8667 815
rect 8701 859 8938 875
rect 8701 825 8710 859
rect 8744 825 8778 859
rect 8812 825 8938 859
rect 8701 809 8938 825
rect 8972 873 9091 889
rect 8972 839 8975 873
rect 9009 839 9043 873
rect 9077 839 9091 873
rect 8972 823 9091 839
rect 9125 873 9244 889
rect 9125 839 9139 873
rect 9173 839 9207 873
rect 9241 839 9244 873
rect 9125 823 9244 839
rect 9278 875 9312 923
rect 9589 875 9655 935
rect 9857 987 9911 1003
rect 9689 934 9723 953
rect 9757 935 9773 969
rect 9807 935 9823 969
rect 9757 911 9823 935
rect 9891 953 9911 987
rect 9945 1029 9995 1071
rect 9945 995 9961 1029
rect 9945 979 9995 995
rect 10029 1029 10095 1037
rect 10029 995 10045 1029
rect 10079 995 10095 1029
rect 9857 945 9911 953
rect 10029 961 10095 995
rect 10129 1029 10183 1071
rect 10129 995 10139 1029
rect 10173 995 10183 1029
rect 10129 979 10183 995
rect 10217 1029 10283 1037
rect 10217 995 10233 1029
rect 10267 995 10283 1029
rect 10029 945 10045 961
rect 9857 927 10045 945
rect 10079 945 10095 961
rect 10217 961 10283 995
rect 10217 945 10233 961
rect 10079 927 10233 945
rect 10267 927 10283 961
rect 9857 911 10283 927
rect 10317 1029 10367 1071
rect 10351 995 10367 1029
rect 10317 961 10367 995
rect 10351 927 10367 961
rect 10317 911 10367 927
rect 9757 875 9803 911
rect 9278 859 9515 875
rect 9278 825 9404 859
rect 9438 825 9472 859
rect 9506 825 9515 859
rect 8601 697 8617 765
rect 8651 697 8667 765
rect 8601 659 8667 697
rect 8601 625 8617 659
rect 8651 625 8667 659
rect 8413 429 8429 463
rect 8463 429 8479 463
rect 8413 391 8479 429
rect 8413 323 8429 391
rect 8463 323 8479 391
rect 6973 213 7227 273
rect 8413 273 8479 323
rect 8513 463 8567 493
rect 8513 428 8523 463
rect 8557 428 8567 463
rect 8513 357 8567 428
rect 8513 323 8523 357
rect 8557 323 8567 357
rect 8513 307 8567 323
rect 8601 463 8667 625
rect 8701 759 8761 775
rect 8904 767 8938 809
rect 9278 809 9515 825
rect 9549 815 9803 875
rect 10039 873 10317 877
rect 10039 839 10055 873
rect 10089 839 10123 873
rect 10157 839 10191 873
rect 10225 839 10259 873
rect 10293 839 10317 873
rect 10039 823 10317 839
rect 9278 767 9312 809
rect 8701 725 8711 759
rect 8745 725 8761 759
rect 8701 660 8761 725
rect 8701 659 8713 660
rect 8701 625 8711 659
rect 8747 626 8761 660
rect 8745 625 8761 626
rect 8701 595 8761 625
rect 8810 751 8865 767
rect 8810 717 8826 751
rect 8860 717 8865 751
rect 8810 645 8865 717
rect 8810 611 8826 645
rect 8860 611 8865 645
rect 8810 561 8865 611
rect 8904 751 8970 767
rect 8904 717 8920 751
rect 8954 717 8970 751
rect 8904 645 8970 717
rect 8904 611 8920 645
rect 8954 611 8970 645
rect 8904 595 8970 611
rect 9004 751 9064 767
rect 9004 717 9014 751
rect 9048 717 9064 751
rect 9004 645 9064 717
rect 9004 611 9014 645
rect 9048 611 9064 645
rect 9004 561 9064 611
rect 9152 751 9212 767
rect 9152 717 9168 751
rect 9202 717 9212 751
rect 9152 645 9212 717
rect 9152 611 9168 645
rect 9202 611 9212 645
rect 9152 561 9212 611
rect 9246 751 9312 767
rect 9246 717 9262 751
rect 9296 717 9312 751
rect 9246 645 9312 717
rect 9246 611 9262 645
rect 9296 611 9312 645
rect 9246 595 9312 611
rect 9351 751 9406 767
rect 9351 717 9356 751
rect 9390 717 9406 751
rect 9351 645 9406 717
rect 9351 611 9356 645
rect 9390 611 9406 645
rect 9351 561 9406 611
rect 9455 759 9515 775
rect 9455 725 9471 759
rect 9505 725 9515 759
rect 9455 660 9515 725
rect 9455 626 9469 660
rect 9503 659 9515 660
rect 9455 625 9471 626
rect 9505 625 9515 659
rect 9455 595 9515 625
rect 9549 765 9615 815
rect 9549 697 9565 765
rect 9599 697 9615 765
rect 9549 659 9615 697
rect 9549 625 9565 659
rect 9599 625 9615 659
rect 8701 527 8769 561
rect 8803 527 8861 561
rect 8895 527 8953 561
rect 8987 527 9045 561
rect 9079 527 9137 561
rect 9171 527 9229 561
rect 9263 527 9321 561
rect 9355 527 9413 561
rect 9447 527 9515 561
rect 8601 429 8617 463
rect 8651 429 8667 463
rect 8601 391 8667 429
rect 8601 323 8617 391
rect 8651 323 8667 391
rect 8601 273 8667 323
rect 8701 463 8761 493
rect 8701 429 8711 463
rect 8745 462 8761 463
rect 8701 428 8713 429
rect 8747 428 8761 462
rect 8701 363 8761 428
rect 8701 329 8711 363
rect 8745 329 8761 363
rect 8701 313 8761 329
rect 8810 477 8865 527
rect 8810 443 8826 477
rect 8860 443 8865 477
rect 8810 371 8865 443
rect 8810 337 8826 371
rect 8860 337 8865 371
rect 8810 321 8865 337
rect 8904 477 8970 493
rect 8904 443 8920 477
rect 8954 443 8970 477
rect 8904 371 8970 443
rect 8904 337 8920 371
rect 8954 337 8970 371
rect 8904 321 8970 337
rect 9004 477 9064 527
rect 9004 443 9014 477
rect 9048 443 9064 477
rect 9004 371 9064 443
rect 9004 337 9014 371
rect 9048 337 9064 371
rect 9004 321 9064 337
rect 9152 477 9212 527
rect 9152 443 9168 477
rect 9202 443 9212 477
rect 9152 371 9212 443
rect 9152 337 9168 371
rect 9202 337 9212 371
rect 9152 321 9212 337
rect 9246 477 9312 493
rect 9246 443 9262 477
rect 9296 443 9312 477
rect 9246 371 9312 443
rect 9246 337 9262 371
rect 9296 337 9312 371
rect 9246 321 9312 337
rect 9351 477 9406 527
rect 9351 443 9356 477
rect 9390 443 9406 477
rect 9351 371 9406 443
rect 9351 337 9356 371
rect 9390 337 9406 371
rect 9351 321 9406 337
rect 9455 463 9515 493
rect 9455 462 9471 463
rect 9455 428 9469 462
rect 9505 429 9515 463
rect 9503 428 9515 429
rect 9455 363 9515 428
rect 9455 329 9471 363
rect 9505 329 9515 363
rect 8904 279 8938 321
rect 6702 165 6736 213
rect 5985 119 6001 153
rect 6035 119 6051 153
rect 6085 135 6135 154
rect 5917 85 5951 101
rect 6119 101 6135 135
rect 6085 85 6135 101
rect 5729 51 6135 85
rect 6236 106 6294 122
rect 6236 72 6260 106
rect 6236 17 6294 72
rect 6328 106 6378 165
rect 6328 72 6344 106
rect 6328 56 6378 72
rect 6420 106 6478 122
rect 6420 72 6428 106
rect 6462 72 6478 106
rect 6420 17 6478 72
rect 6586 106 6644 122
rect 6586 72 6602 106
rect 6636 72 6644 106
rect 6586 17 6644 72
rect 6686 106 6736 165
rect 6929 135 6979 154
rect 6720 72 6736 106
rect 6686 56 6736 72
rect 6770 106 6828 122
rect 6804 72 6828 106
rect 6770 17 6828 72
rect 6929 101 6945 135
rect 7013 153 7079 213
rect 7181 177 7227 213
rect 7463 249 7741 265
rect 7463 215 7479 249
rect 7513 215 7547 249
rect 7581 215 7615 249
rect 7649 215 7683 249
rect 7717 215 7741 249
rect 7463 211 7741 215
rect 7899 249 8177 265
rect 7899 215 7923 249
rect 7957 215 7991 249
rect 8025 215 8059 249
rect 8093 215 8127 249
rect 8161 215 8177 249
rect 7899 211 8177 215
rect 8413 213 8667 273
rect 8701 263 8938 279
rect 9278 279 9312 321
rect 9455 313 9515 329
rect 9549 463 9615 625
rect 9649 765 9703 781
rect 9649 731 9659 765
rect 9693 731 9703 765
rect 9649 660 9703 731
rect 9649 625 9659 660
rect 9693 625 9703 660
rect 9649 595 9703 625
rect 9737 765 9803 815
rect 9737 697 9753 765
rect 9787 697 9803 765
rect 9737 659 9803 697
rect 9737 625 9753 659
rect 9787 625 9803 659
rect 9549 429 9565 463
rect 9599 429 9615 463
rect 9549 391 9615 429
rect 9549 323 9565 391
rect 9599 323 9615 391
rect 8701 229 8710 263
rect 8744 229 8778 263
rect 8812 229 8938 263
rect 8701 213 8938 229
rect 8413 177 8459 213
rect 7013 119 7029 153
rect 7063 119 7079 153
rect 7113 135 7147 154
rect 6929 85 6979 101
rect 7181 153 7247 177
rect 7181 119 7197 153
rect 7231 119 7247 153
rect 7281 161 7707 177
rect 7281 143 7469 161
rect 7281 135 7335 143
rect 7113 85 7147 101
rect 7315 101 7335 135
rect 7453 127 7469 143
rect 7503 143 7657 161
rect 7503 127 7519 143
rect 7281 85 7335 101
rect 6929 51 7335 85
rect 7369 93 7419 109
rect 7369 59 7385 93
rect 7369 17 7419 59
rect 7453 93 7519 127
rect 7641 127 7657 143
rect 7691 127 7707 161
rect 7453 59 7469 93
rect 7503 59 7519 93
rect 7453 51 7519 59
rect 7553 93 7607 109
rect 7553 59 7563 93
rect 7597 59 7607 93
rect 7553 17 7607 59
rect 7641 93 7707 127
rect 7641 59 7657 93
rect 7691 59 7707 93
rect 7641 51 7707 59
rect 7741 161 7791 177
rect 7775 127 7791 161
rect 7741 93 7791 127
rect 7775 59 7791 93
rect 7741 17 7791 59
rect 7849 161 7899 177
rect 7849 127 7865 161
rect 7849 93 7899 127
rect 7849 59 7865 93
rect 7849 17 7899 59
rect 7933 161 8359 177
rect 7933 127 7949 161
rect 7983 143 8137 161
rect 7983 127 7999 143
rect 7933 93 7999 127
rect 8121 127 8137 143
rect 8171 143 8359 161
rect 8171 127 8187 143
rect 7933 59 7949 93
rect 7983 59 7999 93
rect 7933 51 7999 59
rect 8033 93 8087 109
rect 8033 59 8043 93
rect 8077 59 8087 93
rect 8033 17 8087 59
rect 8121 93 8187 127
rect 8305 135 8359 143
rect 8121 59 8137 93
rect 8171 59 8187 93
rect 8121 51 8187 59
rect 8221 93 8271 109
rect 8255 59 8271 93
rect 8221 17 8271 59
rect 8305 101 8325 135
rect 8393 153 8459 177
rect 8393 119 8409 153
rect 8443 119 8459 153
rect 8493 135 8527 154
rect 8305 85 8359 101
rect 8561 153 8627 213
rect 8904 165 8938 213
rect 8972 249 9091 265
rect 8972 215 8975 249
rect 9009 215 9043 249
rect 9077 215 9091 249
rect 8972 199 9091 215
rect 9125 249 9244 265
rect 9125 215 9139 249
rect 9173 215 9207 249
rect 9241 215 9244 249
rect 9125 199 9244 215
rect 9278 263 9515 279
rect 9278 229 9404 263
rect 9438 229 9472 263
rect 9506 229 9515 263
rect 9278 213 9515 229
rect 9549 273 9615 323
rect 9649 463 9703 493
rect 9649 428 9659 463
rect 9693 428 9703 463
rect 9649 357 9703 428
rect 9649 323 9659 357
rect 9693 323 9703 357
rect 9649 307 9703 323
rect 9737 463 9803 625
rect 9837 773 10283 789
rect 9837 765 10045 773
rect 9837 731 9847 765
rect 9881 755 10045 765
rect 9881 731 9897 755
rect 9837 660 9897 731
rect 10029 739 10045 755
rect 10079 755 10233 773
rect 10079 739 10095 755
rect 9837 659 9849 660
rect 9837 625 9847 659
rect 9883 626 9897 660
rect 9881 625 9897 626
rect 9837 595 9897 625
rect 9941 705 9995 721
rect 9941 671 9951 705
rect 9985 671 9995 705
rect 9941 637 9995 671
rect 9941 603 9951 637
rect 9985 603 9995 637
rect 9941 561 9995 603
rect 10029 705 10095 739
rect 10217 739 10233 755
rect 10267 739 10283 773
rect 10029 671 10045 705
rect 10079 671 10095 705
rect 10029 660 10095 671
rect 10029 603 10045 660
rect 10079 603 10095 660
rect 10029 595 10095 603
rect 10129 705 10183 721
rect 10129 671 10139 705
rect 10173 671 10183 705
rect 10129 637 10183 671
rect 10129 603 10139 637
rect 10173 603 10183 637
rect 10129 561 10183 603
rect 10217 705 10283 739
rect 10217 671 10233 705
rect 10267 671 10283 705
rect 10217 660 10283 671
rect 10217 603 10233 660
rect 10267 603 10283 660
rect 10217 595 10283 603
rect 10317 773 10371 789
rect 10317 739 10327 773
rect 10361 739 10371 773
rect 10317 705 10371 739
rect 10317 671 10327 705
rect 10361 671 10371 705
rect 10317 637 10371 671
rect 10317 603 10327 637
rect 10361 603 10371 637
rect 10317 561 10371 603
rect 9837 527 9873 561
rect 9907 527 9965 561
rect 9999 527 10057 561
rect 10091 527 10149 561
rect 10183 527 10241 561
rect 10275 527 10333 561
rect 10367 527 10396 561
rect 9737 429 9753 463
rect 9787 429 9803 463
rect 9737 391 9803 429
rect 9737 323 9753 391
rect 9787 323 9803 391
rect 9737 273 9803 323
rect 9837 463 9897 493
rect 9837 429 9847 463
rect 9881 462 9897 463
rect 9837 428 9849 429
rect 9883 428 9897 462
rect 9837 357 9897 428
rect 9941 485 9995 527
rect 9941 451 9951 485
rect 9985 451 9995 485
rect 9941 417 9995 451
rect 9941 383 9951 417
rect 9985 383 9995 417
rect 9941 367 9995 383
rect 10029 485 10095 493
rect 10029 428 10045 485
rect 10079 428 10095 485
rect 10029 417 10095 428
rect 10029 383 10045 417
rect 10079 383 10095 417
rect 9837 323 9847 357
rect 9881 333 9897 357
rect 10029 349 10095 383
rect 10129 485 10183 527
rect 10129 451 10139 485
rect 10173 451 10183 485
rect 10129 417 10183 451
rect 10129 383 10139 417
rect 10173 383 10183 417
rect 10129 367 10183 383
rect 10217 485 10283 493
rect 10217 428 10233 485
rect 10267 428 10283 485
rect 10217 417 10283 428
rect 10217 383 10233 417
rect 10267 383 10283 417
rect 10029 333 10045 349
rect 9881 323 10045 333
rect 9837 315 10045 323
rect 10079 333 10095 349
rect 10217 349 10283 383
rect 10217 333 10233 349
rect 10079 315 10233 333
rect 10267 315 10283 349
rect 9837 299 10283 315
rect 10317 485 10371 527
rect 10317 451 10327 485
rect 10361 451 10371 485
rect 10317 417 10371 451
rect 10317 383 10327 417
rect 10361 383 10371 417
rect 10317 349 10371 383
rect 10317 315 10327 349
rect 10361 315 10371 349
rect 10317 299 10371 315
rect 9549 213 9803 273
rect 9278 165 9312 213
rect 8561 119 8577 153
rect 8611 119 8627 153
rect 8661 135 8711 154
rect 8493 85 8527 101
rect 8695 101 8711 135
rect 8661 85 8711 101
rect 8305 51 8711 85
rect 8812 106 8870 122
rect 8812 72 8836 106
rect 8812 17 8870 72
rect 8904 106 8954 165
rect 8904 72 8920 106
rect 8904 56 8954 72
rect 8996 106 9054 122
rect 8996 72 9004 106
rect 9038 72 9054 106
rect 8996 17 9054 72
rect 9162 106 9220 122
rect 9162 72 9178 106
rect 9212 72 9220 106
rect 9162 17 9220 72
rect 9262 106 9312 165
rect 9505 135 9555 154
rect 9296 72 9312 106
rect 9262 56 9312 72
rect 9346 106 9404 122
rect 9380 72 9404 106
rect 9346 17 9404 72
rect 9505 101 9521 135
rect 9589 153 9655 213
rect 9757 177 9803 213
rect 10039 249 10317 265
rect 10039 215 10055 249
rect 10089 215 10123 249
rect 10157 215 10191 249
rect 10225 215 10259 249
rect 10293 215 10317 249
rect 10039 211 10317 215
rect 9589 119 9605 153
rect 9639 119 9655 153
rect 9689 135 9723 154
rect 9505 85 9555 101
rect 9757 153 9823 177
rect 9757 119 9773 153
rect 9807 119 9823 153
rect 9857 161 10283 177
rect 9857 143 10045 161
rect 9857 135 9911 143
rect 9689 85 9723 101
rect 9891 101 9911 135
rect 10029 127 10045 143
rect 10079 143 10233 161
rect 10079 127 10095 143
rect 9857 85 9911 101
rect 9505 51 9911 85
rect 9945 93 9995 109
rect 9945 59 9961 93
rect 9945 17 9995 59
rect 10029 93 10095 127
rect 10217 127 10233 143
rect 10267 127 10283 161
rect 10029 59 10045 93
rect 10079 59 10095 93
rect 10029 51 10095 59
rect 10129 93 10183 109
rect 10129 59 10139 93
rect 10173 59 10183 93
rect 10129 17 10183 59
rect 10217 93 10283 127
rect 10217 59 10233 93
rect 10267 59 10283 93
rect 10217 51 10283 59
rect 10317 161 10367 177
rect 10351 127 10367 161
rect 10317 93 10367 127
rect 10351 59 10367 93
rect 10317 17 10367 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3341 17
rect 3375 -17 3433 17
rect 3467 -17 3525 17
rect 3559 -17 3617 17
rect 3651 -17 3709 17
rect 3743 -17 3801 17
rect 3835 -17 3893 17
rect 3927 -17 3985 17
rect 4019 -17 4077 17
rect 4111 -17 4169 17
rect 4203 -17 4261 17
rect 4295 -17 4353 17
rect 4387 -17 4445 17
rect 4479 -17 4537 17
rect 4571 -17 4629 17
rect 4663 -17 4721 17
rect 4755 -17 4813 17
rect 4847 -17 4905 17
rect 4939 -17 4997 17
rect 5031 -17 5089 17
rect 5123 -17 5181 17
rect 5215 -17 5273 17
rect 5307 -17 5365 17
rect 5399 -17 5457 17
rect 5491 -17 5549 17
rect 5583 -17 5641 17
rect 5675 -17 5733 17
rect 5767 -17 5825 17
rect 5859 -17 5917 17
rect 5951 -17 6009 17
rect 6043 -17 6101 17
rect 6135 -17 6193 17
rect 6227 -17 6285 17
rect 6319 -17 6377 17
rect 6411 -17 6469 17
rect 6503 -17 6561 17
rect 6595 -17 6653 17
rect 6687 -17 6745 17
rect 6779 -17 6837 17
rect 6871 -17 6929 17
rect 6963 -17 7021 17
rect 7055 -17 7113 17
rect 7147 -17 7205 17
rect 7239 -17 7297 17
rect 7331 -17 7389 17
rect 7423 -17 7481 17
rect 7515 -17 7573 17
rect 7607 -17 7665 17
rect 7699 -17 7757 17
rect 7791 -17 7849 17
rect 7883 -17 7941 17
rect 7975 -17 8033 17
rect 8067 -17 8125 17
rect 8159 -17 8217 17
rect 8251 -17 8309 17
rect 8343 -17 8401 17
rect 8435 -17 8493 17
rect 8527 -17 8585 17
rect 8619 -17 8677 17
rect 8711 -17 8769 17
rect 8803 -17 8861 17
rect 8895 -17 8953 17
rect 8987 -17 9045 17
rect 9079 -17 9137 17
rect 9171 -17 9229 17
rect 9263 -17 9321 17
rect 9355 -17 9413 17
rect 9447 -17 9505 17
rect 9539 -17 9597 17
rect 9631 -17 9689 17
rect 9723 -17 9781 17
rect 9815 -17 9873 17
rect 9907 -17 9965 17
rect 9999 -17 10057 17
rect 10091 -17 10149 17
rect 10183 -17 10241 17
rect 10275 -17 10333 17
rect 10367 -17 10396 17
<< viali >>
rect 29 1071 63 1105
rect 121 1071 155 1105
rect 213 1071 247 1105
rect 305 1071 339 1105
rect 397 1071 431 1105
rect 489 1071 523 1105
rect 581 1071 615 1105
rect 673 1071 707 1105
rect 765 1071 799 1105
rect 857 1071 891 1105
rect 949 1071 983 1105
rect 1041 1071 1075 1105
rect 1133 1071 1167 1105
rect 1225 1071 1259 1105
rect 1317 1071 1351 1105
rect 1409 1071 1443 1105
rect 1501 1071 1535 1105
rect 1593 1071 1627 1105
rect 1685 1071 1719 1105
rect 1777 1071 1811 1105
rect 1869 1071 1903 1105
rect 1961 1071 1995 1105
rect 2053 1071 2087 1105
rect 2145 1071 2179 1105
rect 2237 1071 2271 1105
rect 2329 1071 2363 1105
rect 2421 1071 2455 1105
rect 2513 1071 2547 1105
rect 2605 1071 2639 1105
rect 2697 1071 2731 1105
rect 2789 1071 2823 1105
rect 2881 1071 2915 1105
rect 2973 1071 3007 1105
rect 3065 1071 3099 1105
rect 3157 1071 3191 1105
rect 3249 1071 3283 1105
rect 3341 1071 3375 1105
rect 3433 1071 3467 1105
rect 3525 1071 3559 1105
rect 3617 1071 3651 1105
rect 3709 1071 3743 1105
rect 3801 1071 3835 1105
rect 3893 1071 3927 1105
rect 3985 1071 4019 1105
rect 4077 1071 4111 1105
rect 4169 1071 4203 1105
rect 4261 1071 4295 1105
rect 4353 1071 4387 1105
rect 4445 1071 4479 1105
rect 4537 1071 4571 1105
rect 4629 1071 4663 1105
rect 4721 1071 4755 1105
rect 4813 1071 4847 1105
rect 4905 1071 4939 1105
rect 4997 1071 5031 1105
rect 5089 1071 5123 1105
rect 5181 1071 5215 1105
rect 5273 1071 5307 1105
rect 5365 1071 5399 1105
rect 5457 1071 5491 1105
rect 5549 1071 5583 1105
rect 5641 1071 5675 1105
rect 5733 1071 5767 1105
rect 5825 1071 5859 1105
rect 5917 1071 5951 1105
rect 6009 1071 6043 1105
rect 6101 1071 6135 1105
rect 6193 1071 6227 1105
rect 6285 1071 6319 1105
rect 6377 1071 6411 1105
rect 6469 1071 6503 1105
rect 6561 1071 6595 1105
rect 6653 1071 6687 1105
rect 6745 1071 6779 1105
rect 6837 1071 6871 1105
rect 6929 1071 6963 1105
rect 7021 1071 7055 1105
rect 7113 1071 7147 1105
rect 7205 1071 7239 1105
rect 7297 1071 7331 1105
rect 7389 1071 7423 1105
rect 7481 1071 7515 1105
rect 7573 1071 7607 1105
rect 7665 1071 7699 1105
rect 7757 1071 7791 1105
rect 7849 1071 7883 1105
rect 7941 1071 7975 1105
rect 8033 1071 8067 1105
rect 8125 1071 8159 1105
rect 8217 1071 8251 1105
rect 8309 1071 8343 1105
rect 8401 1071 8435 1105
rect 8493 1071 8527 1105
rect 8585 1071 8619 1105
rect 8677 1071 8711 1105
rect 8769 1071 8803 1105
rect 8861 1071 8895 1105
rect 8953 1071 8987 1105
rect 9045 1071 9079 1105
rect 9137 1071 9171 1105
rect 9229 1071 9263 1105
rect 9321 1071 9355 1105
rect 9413 1071 9447 1105
rect 9505 1071 9539 1105
rect 9597 1071 9631 1105
rect 9689 1071 9723 1105
rect 9781 1071 9815 1105
rect 9873 1071 9907 1105
rect 9965 1071 9999 1105
rect 10057 1071 10091 1105
rect 10149 1071 10183 1105
rect 10241 1071 10275 1105
rect 10333 1071 10367 1105
rect 129 637 163 660
rect 129 626 163 637
rect 317 637 351 660
rect 317 626 351 637
rect 513 659 547 660
rect 513 626 515 659
rect 515 626 547 659
rect 609 697 643 731
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 129 451 163 462
rect 129 428 163 451
rect 317 451 351 462
rect 317 428 351 451
rect 513 429 515 462
rect 515 429 547 462
rect 513 428 547 429
rect 703 659 737 660
rect 703 626 737 659
rect 797 697 831 731
rect 609 357 643 391
rect 703 429 737 462
rect 703 428 737 429
rect 893 659 927 660
rect 893 626 925 659
rect 925 626 927 659
rect 1649 659 1683 660
rect 1649 626 1651 659
rect 1651 626 1683 659
rect 1745 697 1779 731
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 797 357 831 391
rect 893 429 925 462
rect 925 429 927 462
rect 893 428 927 429
rect 1649 429 1651 462
rect 1651 429 1683 462
rect 1649 428 1683 429
rect 1839 659 1873 660
rect 1839 626 1873 659
rect 1933 697 1967 731
rect 1745 357 1779 391
rect 1839 429 1873 462
rect 1839 428 1873 429
rect 2029 659 2063 660
rect 2029 626 2061 659
rect 2061 626 2063 659
rect 2225 637 2259 660
rect 2225 626 2259 637
rect 2413 637 2447 660
rect 2413 626 2447 637
rect 2705 637 2739 660
rect 2705 626 2739 637
rect 2893 637 2927 660
rect 2893 626 2927 637
rect 3089 659 3123 660
rect 3089 626 3091 659
rect 3091 626 3123 659
rect 3185 697 3219 731
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 2881 527 2915 561
rect 2973 527 3007 561
rect 3065 527 3099 561
rect 1933 357 1967 391
rect 2029 429 2061 462
rect 2061 429 2063 462
rect 2029 428 2063 429
rect 2225 451 2259 462
rect 2225 428 2259 451
rect 2413 451 2447 462
rect 2413 428 2447 451
rect 2705 451 2739 462
rect 2705 428 2739 451
rect 2893 451 2927 462
rect 2893 428 2927 451
rect 3089 429 3091 462
rect 3091 429 3123 462
rect 3089 428 3123 429
rect 3279 659 3313 660
rect 3279 626 3313 659
rect 3373 697 3407 731
rect 3185 357 3219 391
rect 3279 429 3313 462
rect 3279 428 3313 429
rect 3469 659 3503 660
rect 3469 626 3501 659
rect 3501 626 3503 659
rect 4225 659 4259 660
rect 4225 626 4227 659
rect 4227 626 4259 659
rect 4321 697 4355 731
rect 3525 527 3559 561
rect 3617 527 3651 561
rect 3709 527 3743 561
rect 3801 527 3835 561
rect 3893 527 3927 561
rect 3985 527 4019 561
rect 4077 527 4111 561
rect 4169 527 4203 561
rect 3373 357 3407 391
rect 3469 429 3501 462
rect 3501 429 3503 462
rect 3469 428 3503 429
rect 4225 429 4227 462
rect 4227 429 4259 462
rect 4225 428 4259 429
rect 4415 659 4449 660
rect 4415 626 4449 659
rect 4509 697 4543 731
rect 4321 357 4355 391
rect 4415 429 4449 462
rect 4415 428 4449 429
rect 4605 659 4639 660
rect 4605 626 4637 659
rect 4637 626 4639 659
rect 4801 637 4835 660
rect 4801 626 4835 637
rect 4989 637 5023 660
rect 4989 626 5023 637
rect 5373 637 5407 660
rect 5373 626 5407 637
rect 5561 637 5595 660
rect 5561 626 5595 637
rect 5757 659 5791 660
rect 5757 626 5759 659
rect 5759 626 5791 659
rect 5853 697 5887 731
rect 4629 527 4663 561
rect 4721 527 4755 561
rect 4813 527 4847 561
rect 4905 527 4939 561
rect 4997 527 5031 561
rect 5089 527 5123 561
rect 5181 527 5215 561
rect 5273 527 5307 561
rect 5365 527 5399 561
rect 5457 527 5491 561
rect 5549 527 5583 561
rect 5641 527 5675 561
rect 5733 527 5767 561
rect 4509 357 4543 391
rect 4605 429 4637 462
rect 4637 429 4639 462
rect 4605 428 4639 429
rect 4801 451 4835 462
rect 4801 428 4835 451
rect 4989 451 5023 462
rect 4989 428 5023 451
rect 5373 451 5407 462
rect 5373 428 5407 451
rect 5561 451 5595 462
rect 5561 428 5595 451
rect 5757 429 5759 462
rect 5759 429 5791 462
rect 5757 428 5791 429
rect 5947 659 5981 660
rect 5947 626 5981 659
rect 6041 697 6075 731
rect 5853 357 5887 391
rect 5947 429 5981 462
rect 5947 428 5981 429
rect 6137 659 6171 660
rect 6137 626 6169 659
rect 6169 626 6171 659
rect 6893 659 6927 660
rect 6893 626 6895 659
rect 6895 626 6927 659
rect 6989 697 7023 731
rect 6193 527 6227 561
rect 6285 527 6319 561
rect 6377 527 6411 561
rect 6469 527 6503 561
rect 6561 527 6595 561
rect 6653 527 6687 561
rect 6745 527 6779 561
rect 6837 527 6871 561
rect 6041 357 6075 391
rect 6137 429 6169 462
rect 6169 429 6171 462
rect 6137 428 6171 429
rect 6893 429 6895 462
rect 6895 429 6927 462
rect 6893 428 6927 429
rect 7083 659 7117 660
rect 7083 626 7117 659
rect 7177 697 7211 731
rect 6989 357 7023 391
rect 7083 429 7117 462
rect 7083 428 7117 429
rect 7273 659 7307 660
rect 7273 626 7305 659
rect 7305 626 7307 659
rect 7469 637 7503 660
rect 7469 626 7503 637
rect 7657 637 7691 660
rect 7657 626 7691 637
rect 7949 637 7983 660
rect 7949 626 7983 637
rect 8137 637 8171 660
rect 8137 626 8171 637
rect 8333 659 8367 660
rect 8333 626 8335 659
rect 8335 626 8367 659
rect 8429 697 8463 731
rect 7297 527 7331 561
rect 7389 527 7423 561
rect 7481 527 7515 561
rect 7573 527 7607 561
rect 7665 527 7699 561
rect 7757 527 7791 561
rect 7849 527 7883 561
rect 7941 527 7975 561
rect 8033 527 8067 561
rect 8125 527 8159 561
rect 8217 527 8251 561
rect 8309 527 8343 561
rect 7177 357 7211 391
rect 7273 429 7305 462
rect 7305 429 7307 462
rect 7273 428 7307 429
rect 7469 451 7503 462
rect 7469 428 7503 451
rect 7657 451 7691 462
rect 7657 428 7691 451
rect 7949 451 7983 462
rect 7949 428 7983 451
rect 8137 451 8171 462
rect 8137 428 8171 451
rect 8333 429 8335 462
rect 8335 429 8367 462
rect 8333 428 8367 429
rect 8523 659 8557 660
rect 8523 626 8557 659
rect 8617 697 8651 731
rect 8429 357 8463 391
rect 8523 429 8557 462
rect 8523 428 8557 429
rect 8713 659 8747 660
rect 8713 626 8745 659
rect 8745 626 8747 659
rect 9469 659 9503 660
rect 9469 626 9471 659
rect 9471 626 9503 659
rect 9565 697 9599 731
rect 8769 527 8803 561
rect 8861 527 8895 561
rect 8953 527 8987 561
rect 9045 527 9079 561
rect 9137 527 9171 561
rect 9229 527 9263 561
rect 9321 527 9355 561
rect 9413 527 9447 561
rect 8617 357 8651 391
rect 8713 429 8745 462
rect 8745 429 8747 462
rect 8713 428 8747 429
rect 9469 429 9471 462
rect 9471 429 9503 462
rect 9469 428 9503 429
rect 9659 659 9693 660
rect 9659 626 9693 659
rect 9753 697 9787 731
rect 9565 357 9599 391
rect 9659 429 9693 462
rect 9659 428 9693 429
rect 9849 659 9883 660
rect 9849 626 9881 659
rect 9881 626 9883 659
rect 10045 637 10079 660
rect 10045 626 10079 637
rect 10233 637 10267 660
rect 10233 626 10267 637
rect 9873 527 9907 561
rect 9965 527 9999 561
rect 10057 527 10091 561
rect 10149 527 10183 561
rect 10241 527 10275 561
rect 10333 527 10367 561
rect 9753 357 9787 391
rect 9849 429 9881 462
rect 9881 429 9883 462
rect 9849 428 9883 429
rect 10045 451 10079 462
rect 10045 428 10079 451
rect 10233 451 10267 462
rect 10233 428 10267 451
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
rect 2881 -17 2915 17
rect 2973 -17 3007 17
rect 3065 -17 3099 17
rect 3157 -17 3191 17
rect 3249 -17 3283 17
rect 3341 -17 3375 17
rect 3433 -17 3467 17
rect 3525 -17 3559 17
rect 3617 -17 3651 17
rect 3709 -17 3743 17
rect 3801 -17 3835 17
rect 3893 -17 3927 17
rect 3985 -17 4019 17
rect 4077 -17 4111 17
rect 4169 -17 4203 17
rect 4261 -17 4295 17
rect 4353 -17 4387 17
rect 4445 -17 4479 17
rect 4537 -17 4571 17
rect 4629 -17 4663 17
rect 4721 -17 4755 17
rect 4813 -17 4847 17
rect 4905 -17 4939 17
rect 4997 -17 5031 17
rect 5089 -17 5123 17
rect 5181 -17 5215 17
rect 5273 -17 5307 17
rect 5365 -17 5399 17
rect 5457 -17 5491 17
rect 5549 -17 5583 17
rect 5641 -17 5675 17
rect 5733 -17 5767 17
rect 5825 -17 5859 17
rect 5917 -17 5951 17
rect 6009 -17 6043 17
rect 6101 -17 6135 17
rect 6193 -17 6227 17
rect 6285 -17 6319 17
rect 6377 -17 6411 17
rect 6469 -17 6503 17
rect 6561 -17 6595 17
rect 6653 -17 6687 17
rect 6745 -17 6779 17
rect 6837 -17 6871 17
rect 6929 -17 6963 17
rect 7021 -17 7055 17
rect 7113 -17 7147 17
rect 7205 -17 7239 17
rect 7297 -17 7331 17
rect 7389 -17 7423 17
rect 7481 -17 7515 17
rect 7573 -17 7607 17
rect 7665 -17 7699 17
rect 7757 -17 7791 17
rect 7849 -17 7883 17
rect 7941 -17 7975 17
rect 8033 -17 8067 17
rect 8125 -17 8159 17
rect 8217 -17 8251 17
rect 8309 -17 8343 17
rect 8401 -17 8435 17
rect 8493 -17 8527 17
rect 8585 -17 8619 17
rect 8677 -17 8711 17
rect 8769 -17 8803 17
rect 8861 -17 8895 17
rect 8953 -17 8987 17
rect 9045 -17 9079 17
rect 9137 -17 9171 17
rect 9229 -17 9263 17
rect 9321 -17 9355 17
rect 9413 -17 9447 17
rect 9505 -17 9539 17
rect 9597 -17 9631 17
rect 9689 -17 9723 17
rect 9781 -17 9815 17
rect 9873 -17 9907 17
rect 9965 -17 9999 17
rect 10057 -17 10091 17
rect 10149 -17 10183 17
rect 10241 -17 10275 17
rect 10333 -17 10367 17
<< metal1 >>
rect 0 1105 10396 1136
rect 0 1071 29 1105
rect 63 1071 121 1105
rect 155 1071 213 1105
rect 247 1071 305 1105
rect 339 1071 397 1105
rect 431 1071 489 1105
rect 523 1071 581 1105
rect 615 1071 673 1105
rect 707 1071 765 1105
rect 799 1071 857 1105
rect 891 1071 949 1105
rect 983 1071 1041 1105
rect 1075 1071 1133 1105
rect 1167 1071 1225 1105
rect 1259 1071 1317 1105
rect 1351 1071 1409 1105
rect 1443 1071 1501 1105
rect 1535 1071 1593 1105
rect 1627 1071 1685 1105
rect 1719 1071 1777 1105
rect 1811 1071 1869 1105
rect 1903 1071 1961 1105
rect 1995 1071 2053 1105
rect 2087 1071 2145 1105
rect 2179 1071 2237 1105
rect 2271 1071 2329 1105
rect 2363 1071 2421 1105
rect 2455 1071 2513 1105
rect 2547 1071 2605 1105
rect 2639 1071 2697 1105
rect 2731 1071 2789 1105
rect 2823 1071 2881 1105
rect 2915 1071 2973 1105
rect 3007 1071 3065 1105
rect 3099 1071 3157 1105
rect 3191 1071 3249 1105
rect 3283 1071 3341 1105
rect 3375 1071 3433 1105
rect 3467 1071 3525 1105
rect 3559 1071 3617 1105
rect 3651 1071 3709 1105
rect 3743 1071 3801 1105
rect 3835 1071 3893 1105
rect 3927 1071 3985 1105
rect 4019 1071 4077 1105
rect 4111 1071 4169 1105
rect 4203 1071 4261 1105
rect 4295 1071 4353 1105
rect 4387 1071 4445 1105
rect 4479 1071 4537 1105
rect 4571 1071 4629 1105
rect 4663 1071 4721 1105
rect 4755 1071 4813 1105
rect 4847 1071 4905 1105
rect 4939 1071 4997 1105
rect 5031 1071 5089 1105
rect 5123 1071 5181 1105
rect 5215 1071 5273 1105
rect 5307 1071 5365 1105
rect 5399 1071 5457 1105
rect 5491 1071 5549 1105
rect 5583 1071 5641 1105
rect 5675 1071 5733 1105
rect 5767 1071 5825 1105
rect 5859 1071 5917 1105
rect 5951 1071 6009 1105
rect 6043 1071 6101 1105
rect 6135 1071 6193 1105
rect 6227 1071 6285 1105
rect 6319 1071 6377 1105
rect 6411 1071 6469 1105
rect 6503 1071 6561 1105
rect 6595 1071 6653 1105
rect 6687 1071 6745 1105
rect 6779 1071 6837 1105
rect 6871 1071 6929 1105
rect 6963 1071 7021 1105
rect 7055 1071 7113 1105
rect 7147 1071 7205 1105
rect 7239 1071 7297 1105
rect 7331 1071 7389 1105
rect 7423 1071 7481 1105
rect 7515 1071 7573 1105
rect 7607 1071 7665 1105
rect 7699 1071 7757 1105
rect 7791 1071 7849 1105
rect 7883 1071 7941 1105
rect 7975 1071 8033 1105
rect 8067 1071 8125 1105
rect 8159 1071 8217 1105
rect 8251 1071 8309 1105
rect 8343 1071 8401 1105
rect 8435 1071 8493 1105
rect 8527 1071 8585 1105
rect 8619 1071 8677 1105
rect 8711 1071 8769 1105
rect 8803 1071 8861 1105
rect 8895 1071 8953 1105
rect 8987 1071 9045 1105
rect 9079 1071 9137 1105
rect 9171 1071 9229 1105
rect 9263 1071 9321 1105
rect 9355 1071 9413 1105
rect 9447 1071 9505 1105
rect 9539 1071 9597 1105
rect 9631 1071 9689 1105
rect 9723 1071 9781 1105
rect 9815 1071 9873 1105
rect 9907 1071 9965 1105
rect 9999 1071 10057 1105
rect 10091 1071 10149 1105
rect 10183 1071 10241 1105
rect 10275 1071 10333 1105
rect 10367 1071 10396 1105
rect 0 1040 10396 1071
rect 597 731 655 737
rect 597 697 609 731
rect 643 728 655 731
rect 785 731 843 737
rect 785 728 797 731
rect 643 700 797 728
rect 643 697 655 700
rect 597 691 655 697
rect 785 697 797 700
rect 831 728 843 731
rect 1733 731 1791 737
rect 1733 728 1745 731
rect 831 700 1745 728
rect 831 697 843 700
rect 785 691 843 697
rect 1733 697 1745 700
rect 1779 728 1791 731
rect 1921 731 1979 737
rect 1921 728 1933 731
rect 1779 700 1933 728
rect 1779 697 1791 700
rect 1733 691 1791 697
rect 1921 697 1933 700
rect 1967 728 1979 731
rect 3173 731 3231 737
rect 3173 728 3185 731
rect 1967 700 3185 728
rect 1967 697 1979 700
rect 1921 691 1979 697
rect 3173 697 3185 700
rect 3219 728 3231 731
rect 3361 731 3419 737
rect 3361 728 3373 731
rect 3219 700 3373 728
rect 3219 697 3231 700
rect 3173 691 3231 697
rect 3361 697 3373 700
rect 3407 728 3419 731
rect 4309 731 4367 737
rect 4309 728 4321 731
rect 3407 700 4321 728
rect 3407 697 3419 700
rect 3361 691 3419 697
rect 4309 697 4321 700
rect 4355 728 4367 731
rect 4497 731 4555 737
rect 4497 728 4509 731
rect 4355 700 4509 728
rect 4355 697 4367 700
rect 4309 691 4367 697
rect 4497 697 4509 700
rect 4543 728 4555 731
rect 5841 731 5899 737
rect 5841 728 5853 731
rect 4543 700 5853 728
rect 4543 697 4555 700
rect 4497 691 4555 697
rect 5841 697 5853 700
rect 5887 728 5899 731
rect 6029 731 6087 737
rect 6029 728 6041 731
rect 5887 700 6041 728
rect 5887 697 5899 700
rect 5841 691 5899 697
rect 6029 697 6041 700
rect 6075 728 6087 731
rect 6977 731 7035 737
rect 6977 728 6989 731
rect 6075 700 6989 728
rect 6075 697 6087 700
rect 6029 691 6087 697
rect 6977 697 6989 700
rect 7023 728 7035 731
rect 7165 731 7223 737
rect 7165 728 7177 731
rect 7023 700 7177 728
rect 7023 697 7035 700
rect 6977 691 7035 697
rect 7165 697 7177 700
rect 7211 728 7223 731
rect 8417 731 8475 737
rect 8417 728 8429 731
rect 7211 700 8429 728
rect 7211 697 7223 700
rect 7165 691 7223 697
rect 8417 697 8429 700
rect 8463 728 8475 731
rect 8605 731 8663 737
rect 8605 728 8617 731
rect 8463 700 8617 728
rect 8463 697 8475 700
rect 8417 691 8475 697
rect 8605 697 8617 700
rect 8651 728 8663 731
rect 9553 731 9611 737
rect 9553 728 9565 731
rect 8651 700 9565 728
rect 8651 697 8663 700
rect 8605 691 8663 697
rect 9553 697 9565 700
rect 9599 728 9611 731
rect 9741 731 9799 737
rect 9741 728 9753 731
rect 9599 700 9753 728
rect 9599 697 9611 700
rect 9553 691 9611 697
rect 9741 697 9753 700
rect 9787 697 9799 731
rect 9741 691 9799 697
rect 117 660 175 666
rect 117 626 129 660
rect 163 657 175 660
rect 305 660 363 666
rect 305 657 317 660
rect 163 629 317 657
rect 163 626 175 629
rect 117 620 175 626
rect 305 626 317 629
rect 351 657 363 660
rect 501 660 559 666
rect 501 657 513 660
rect 351 629 513 657
rect 351 626 363 629
rect 305 620 363 626
rect 501 626 513 629
rect 547 657 559 660
rect 691 660 749 666
rect 691 657 703 660
rect 547 629 703 657
rect 547 626 559 629
rect 501 620 559 626
rect 691 626 703 629
rect 737 657 749 660
rect 881 660 939 666
rect 881 657 893 660
rect 737 629 893 657
rect 737 626 749 629
rect 691 620 749 626
rect 881 626 893 629
rect 927 626 939 660
rect 881 620 939 626
rect 1637 660 1695 666
rect 1637 626 1649 660
rect 1683 657 1695 660
rect 1827 660 1885 666
rect 1827 657 1839 660
rect 1683 629 1839 657
rect 1683 626 1695 629
rect 1637 620 1695 626
rect 1827 626 1839 629
rect 1873 657 1885 660
rect 2017 660 2075 666
rect 2017 657 2029 660
rect 1873 629 2029 657
rect 1873 626 1885 629
rect 1827 620 1885 626
rect 2017 626 2029 629
rect 2063 657 2075 660
rect 2213 660 2271 666
rect 2213 657 2225 660
rect 2063 629 2225 657
rect 2063 626 2075 629
rect 2017 620 2075 626
rect 2213 626 2225 629
rect 2259 657 2271 660
rect 2401 660 2459 666
rect 2401 657 2413 660
rect 2259 629 2413 657
rect 2259 626 2271 629
rect 2213 620 2271 626
rect 2401 626 2413 629
rect 2447 626 2459 660
rect 2401 620 2459 626
rect 2693 660 2751 666
rect 2693 626 2705 660
rect 2739 657 2751 660
rect 2881 660 2939 666
rect 2881 657 2893 660
rect 2739 629 2893 657
rect 2739 626 2751 629
rect 2693 620 2751 626
rect 2881 626 2893 629
rect 2927 657 2939 660
rect 3077 660 3135 666
rect 3077 657 3089 660
rect 2927 629 3089 657
rect 2927 626 2939 629
rect 2881 620 2939 626
rect 3077 626 3089 629
rect 3123 657 3135 660
rect 3267 660 3325 666
rect 3267 657 3279 660
rect 3123 629 3279 657
rect 3123 626 3135 629
rect 3077 620 3135 626
rect 3267 626 3279 629
rect 3313 657 3325 660
rect 3457 660 3515 666
rect 3457 657 3469 660
rect 3313 629 3469 657
rect 3313 626 3325 629
rect 3267 620 3325 626
rect 3457 626 3469 629
rect 3503 626 3515 660
rect 3457 620 3515 626
rect 4213 660 4271 666
rect 4213 626 4225 660
rect 4259 657 4271 660
rect 4403 660 4461 666
rect 4403 657 4415 660
rect 4259 629 4415 657
rect 4259 626 4271 629
rect 4213 620 4271 626
rect 4403 626 4415 629
rect 4449 657 4461 660
rect 4593 660 4651 666
rect 4593 657 4605 660
rect 4449 629 4605 657
rect 4449 626 4461 629
rect 4403 620 4461 626
rect 4593 626 4605 629
rect 4639 657 4651 660
rect 4789 660 4847 666
rect 4789 657 4801 660
rect 4639 629 4801 657
rect 4639 626 4651 629
rect 4593 620 4651 626
rect 4789 626 4801 629
rect 4835 657 4847 660
rect 4977 660 5035 666
rect 4977 657 4989 660
rect 4835 629 4989 657
rect 4835 626 4847 629
rect 4789 620 4847 626
rect 4977 626 4989 629
rect 5023 626 5035 660
rect 4977 620 5035 626
rect 5361 660 5419 666
rect 5361 626 5373 660
rect 5407 657 5419 660
rect 5549 660 5607 666
rect 5549 657 5561 660
rect 5407 629 5561 657
rect 5407 626 5419 629
rect 5361 620 5419 626
rect 5549 626 5561 629
rect 5595 657 5607 660
rect 5745 660 5803 666
rect 5745 657 5757 660
rect 5595 629 5757 657
rect 5595 626 5607 629
rect 5549 620 5607 626
rect 5745 626 5757 629
rect 5791 657 5803 660
rect 5935 660 5993 666
rect 5935 657 5947 660
rect 5791 629 5947 657
rect 5791 626 5803 629
rect 5745 620 5803 626
rect 5935 626 5947 629
rect 5981 657 5993 660
rect 6125 660 6183 666
rect 6125 657 6137 660
rect 5981 629 6137 657
rect 5981 626 5993 629
rect 5935 620 5993 626
rect 6125 626 6137 629
rect 6171 626 6183 660
rect 6125 620 6183 626
rect 6881 660 6939 666
rect 6881 626 6893 660
rect 6927 657 6939 660
rect 7071 660 7129 666
rect 7071 657 7083 660
rect 6927 629 7083 657
rect 6927 626 6939 629
rect 6881 620 6939 626
rect 7071 626 7083 629
rect 7117 657 7129 660
rect 7261 660 7319 666
rect 7261 657 7273 660
rect 7117 629 7273 657
rect 7117 626 7129 629
rect 7071 620 7129 626
rect 7261 626 7273 629
rect 7307 657 7319 660
rect 7457 660 7515 666
rect 7457 657 7469 660
rect 7307 629 7469 657
rect 7307 626 7319 629
rect 7261 620 7319 626
rect 7457 626 7469 629
rect 7503 657 7515 660
rect 7645 660 7703 666
rect 7645 657 7657 660
rect 7503 629 7657 657
rect 7503 626 7515 629
rect 7457 620 7515 626
rect 7645 626 7657 629
rect 7691 626 7703 660
rect 7645 620 7703 626
rect 7937 660 7995 666
rect 7937 626 7949 660
rect 7983 657 7995 660
rect 8125 660 8183 666
rect 8125 657 8137 660
rect 7983 629 8137 657
rect 7983 626 7995 629
rect 7937 620 7995 626
rect 8125 626 8137 629
rect 8171 657 8183 660
rect 8321 660 8379 666
rect 8321 657 8333 660
rect 8171 629 8333 657
rect 8171 626 8183 629
rect 8125 620 8183 626
rect 8321 626 8333 629
rect 8367 657 8379 660
rect 8511 660 8569 666
rect 8511 657 8523 660
rect 8367 629 8523 657
rect 8367 626 8379 629
rect 8321 620 8379 626
rect 8511 626 8523 629
rect 8557 657 8569 660
rect 8701 660 8759 666
rect 8701 657 8713 660
rect 8557 629 8713 657
rect 8557 626 8569 629
rect 8511 620 8569 626
rect 8701 626 8713 629
rect 8747 626 8759 660
rect 8701 620 8759 626
rect 9457 660 9515 666
rect 9457 626 9469 660
rect 9503 657 9515 660
rect 9647 660 9705 666
rect 9647 657 9659 660
rect 9503 629 9659 657
rect 9503 626 9515 629
rect 9457 620 9515 626
rect 9647 626 9659 629
rect 9693 657 9705 660
rect 9837 660 9895 666
rect 9837 657 9849 660
rect 9693 629 9849 657
rect 9693 626 9705 629
rect 9647 620 9705 626
rect 9837 626 9849 629
rect 9883 657 9895 660
rect 10033 660 10091 666
rect 10033 657 10045 660
rect 9883 629 10045 657
rect 9883 626 9895 629
rect 9837 620 9895 626
rect 10033 626 10045 629
rect 10079 657 10091 660
rect 10221 660 10279 666
rect 10221 657 10233 660
rect 10079 629 10233 657
rect 10079 626 10091 629
rect 10033 620 10091 626
rect 10221 626 10233 629
rect 10267 626 10279 660
rect 10221 620 10279 626
rect 0 561 10396 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3525 561
rect 3559 527 3617 561
rect 3651 527 3709 561
rect 3743 527 3801 561
rect 3835 527 3893 561
rect 3927 527 3985 561
rect 4019 527 4077 561
rect 4111 527 4169 561
rect 4203 527 4629 561
rect 4663 527 4721 561
rect 4755 527 4813 561
rect 4847 527 4905 561
rect 4939 527 4997 561
rect 5031 527 5089 561
rect 5123 527 5181 561
rect 5215 527 5273 561
rect 5307 527 5365 561
rect 5399 527 5457 561
rect 5491 527 5549 561
rect 5583 527 5641 561
rect 5675 527 5733 561
rect 5767 527 6193 561
rect 6227 527 6285 561
rect 6319 527 6377 561
rect 6411 527 6469 561
rect 6503 527 6561 561
rect 6595 527 6653 561
rect 6687 527 6745 561
rect 6779 527 6837 561
rect 6871 527 7297 561
rect 7331 527 7389 561
rect 7423 527 7481 561
rect 7515 527 7573 561
rect 7607 527 7665 561
rect 7699 527 7757 561
rect 7791 527 7849 561
rect 7883 527 7941 561
rect 7975 527 8033 561
rect 8067 527 8125 561
rect 8159 527 8217 561
rect 8251 527 8309 561
rect 8343 527 8769 561
rect 8803 527 8861 561
rect 8895 527 8953 561
rect 8987 527 9045 561
rect 9079 527 9137 561
rect 9171 527 9229 561
rect 9263 527 9321 561
rect 9355 527 9413 561
rect 9447 527 9873 561
rect 9907 527 9965 561
rect 9999 527 10057 561
rect 10091 527 10149 561
rect 10183 527 10241 561
rect 10275 527 10333 561
rect 10367 527 10396 561
rect 0 496 10396 527
rect 117 462 175 468
rect 117 428 129 462
rect 163 459 175 462
rect 305 462 363 468
rect 305 459 317 462
rect 163 431 317 459
rect 163 428 175 431
rect 117 422 175 428
rect 305 428 317 431
rect 351 459 363 462
rect 501 462 559 468
rect 501 459 513 462
rect 351 431 513 459
rect 351 428 363 431
rect 305 422 363 428
rect 501 428 513 431
rect 547 459 559 462
rect 691 462 749 468
rect 691 459 703 462
rect 547 431 703 459
rect 547 428 559 431
rect 501 422 559 428
rect 691 428 703 431
rect 737 459 749 462
rect 881 462 939 468
rect 881 459 893 462
rect 737 431 893 459
rect 737 428 749 431
rect 691 422 749 428
rect 881 428 893 431
rect 927 428 939 462
rect 881 422 939 428
rect 1637 462 1695 468
rect 1637 428 1649 462
rect 1683 459 1695 462
rect 1827 462 1885 468
rect 1827 459 1839 462
rect 1683 431 1839 459
rect 1683 428 1695 431
rect 1637 422 1695 428
rect 1827 428 1839 431
rect 1873 459 1885 462
rect 2017 462 2075 468
rect 2017 459 2029 462
rect 1873 431 2029 459
rect 1873 428 1885 431
rect 1827 422 1885 428
rect 2017 428 2029 431
rect 2063 459 2075 462
rect 2213 462 2271 468
rect 2213 459 2225 462
rect 2063 431 2225 459
rect 2063 428 2075 431
rect 2017 422 2075 428
rect 2213 428 2225 431
rect 2259 459 2271 462
rect 2401 462 2459 468
rect 2401 459 2413 462
rect 2259 431 2413 459
rect 2259 428 2271 431
rect 2213 422 2271 428
rect 2401 428 2413 431
rect 2447 428 2459 462
rect 2401 422 2459 428
rect 2693 462 2751 468
rect 2693 428 2705 462
rect 2739 459 2751 462
rect 2881 462 2939 468
rect 2881 459 2893 462
rect 2739 431 2893 459
rect 2739 428 2751 431
rect 2693 422 2751 428
rect 2881 428 2893 431
rect 2927 459 2939 462
rect 3077 462 3135 468
rect 3077 459 3089 462
rect 2927 431 3089 459
rect 2927 428 2939 431
rect 2881 422 2939 428
rect 3077 428 3089 431
rect 3123 459 3135 462
rect 3267 462 3325 468
rect 3267 459 3279 462
rect 3123 431 3279 459
rect 3123 428 3135 431
rect 3077 422 3135 428
rect 3267 428 3279 431
rect 3313 459 3325 462
rect 3457 462 3515 468
rect 3457 459 3469 462
rect 3313 431 3469 459
rect 3313 428 3325 431
rect 3267 422 3325 428
rect 3457 428 3469 431
rect 3503 428 3515 462
rect 3457 422 3515 428
rect 4213 462 4271 468
rect 4213 428 4225 462
rect 4259 459 4271 462
rect 4403 462 4461 468
rect 4403 459 4415 462
rect 4259 431 4415 459
rect 4259 428 4271 431
rect 4213 422 4271 428
rect 4403 428 4415 431
rect 4449 459 4461 462
rect 4593 462 4651 468
rect 4593 459 4605 462
rect 4449 431 4605 459
rect 4449 428 4461 431
rect 4403 422 4461 428
rect 4593 428 4605 431
rect 4639 459 4651 462
rect 4789 462 4847 468
rect 4789 459 4801 462
rect 4639 431 4801 459
rect 4639 428 4651 431
rect 4593 422 4651 428
rect 4789 428 4801 431
rect 4835 459 4847 462
rect 4977 462 5035 468
rect 4977 459 4989 462
rect 4835 431 4989 459
rect 4835 428 4847 431
rect 4789 422 4847 428
rect 4977 428 4989 431
rect 5023 428 5035 462
rect 4977 422 5035 428
rect 5361 462 5419 468
rect 5361 428 5373 462
rect 5407 459 5419 462
rect 5549 462 5607 468
rect 5549 459 5561 462
rect 5407 431 5561 459
rect 5407 428 5419 431
rect 5361 422 5419 428
rect 5549 428 5561 431
rect 5595 459 5607 462
rect 5745 462 5803 468
rect 5745 459 5757 462
rect 5595 431 5757 459
rect 5595 428 5607 431
rect 5549 422 5607 428
rect 5745 428 5757 431
rect 5791 459 5803 462
rect 5935 462 5993 468
rect 5935 459 5947 462
rect 5791 431 5947 459
rect 5791 428 5803 431
rect 5745 422 5803 428
rect 5935 428 5947 431
rect 5981 459 5993 462
rect 6125 462 6183 468
rect 6125 459 6137 462
rect 5981 431 6137 459
rect 5981 428 5993 431
rect 5935 422 5993 428
rect 6125 428 6137 431
rect 6171 428 6183 462
rect 6125 422 6183 428
rect 6881 462 6939 468
rect 6881 428 6893 462
rect 6927 459 6939 462
rect 7071 462 7129 468
rect 7071 459 7083 462
rect 6927 431 7083 459
rect 6927 428 6939 431
rect 6881 422 6939 428
rect 7071 428 7083 431
rect 7117 459 7129 462
rect 7261 462 7319 468
rect 7261 459 7273 462
rect 7117 431 7273 459
rect 7117 428 7129 431
rect 7071 422 7129 428
rect 7261 428 7273 431
rect 7307 459 7319 462
rect 7457 462 7515 468
rect 7457 459 7469 462
rect 7307 431 7469 459
rect 7307 428 7319 431
rect 7261 422 7319 428
rect 7457 428 7469 431
rect 7503 459 7515 462
rect 7645 462 7703 468
rect 7645 459 7657 462
rect 7503 431 7657 459
rect 7503 428 7515 431
rect 7457 422 7515 428
rect 7645 428 7657 431
rect 7691 428 7703 462
rect 7645 422 7703 428
rect 7937 462 7995 468
rect 7937 428 7949 462
rect 7983 459 7995 462
rect 8125 462 8183 468
rect 8125 459 8137 462
rect 7983 431 8137 459
rect 7983 428 7995 431
rect 7937 422 7995 428
rect 8125 428 8137 431
rect 8171 459 8183 462
rect 8321 462 8379 468
rect 8321 459 8333 462
rect 8171 431 8333 459
rect 8171 428 8183 431
rect 8125 422 8183 428
rect 8321 428 8333 431
rect 8367 459 8379 462
rect 8511 462 8569 468
rect 8511 459 8523 462
rect 8367 431 8523 459
rect 8367 428 8379 431
rect 8321 422 8379 428
rect 8511 428 8523 431
rect 8557 459 8569 462
rect 8701 462 8759 468
rect 8701 459 8713 462
rect 8557 431 8713 459
rect 8557 428 8569 431
rect 8511 422 8569 428
rect 8701 428 8713 431
rect 8747 428 8759 462
rect 8701 422 8759 428
rect 9457 462 9515 468
rect 9457 428 9469 462
rect 9503 459 9515 462
rect 9647 462 9705 468
rect 9647 459 9659 462
rect 9503 431 9659 459
rect 9503 428 9515 431
rect 9457 422 9515 428
rect 9647 428 9659 431
rect 9693 459 9705 462
rect 9837 462 9895 468
rect 9837 459 9849 462
rect 9693 431 9849 459
rect 9693 428 9705 431
rect 9647 422 9705 428
rect 9837 428 9849 431
rect 9883 459 9895 462
rect 10033 462 10091 468
rect 10033 459 10045 462
rect 9883 431 10045 459
rect 9883 428 9895 431
rect 9837 422 9895 428
rect 10033 428 10045 431
rect 10079 459 10091 462
rect 10221 462 10279 468
rect 10221 459 10233 462
rect 10079 431 10233 459
rect 10079 428 10091 431
rect 10033 422 10091 428
rect 10221 428 10233 431
rect 10267 428 10279 462
rect 10221 422 10279 428
rect 597 391 655 397
rect 597 357 609 391
rect 643 388 655 391
rect 785 391 843 397
rect 785 388 797 391
rect 643 360 797 388
rect 643 357 655 360
rect 597 351 655 357
rect 785 357 797 360
rect 831 388 843 391
rect 1733 391 1791 397
rect 1733 388 1745 391
rect 831 360 1745 388
rect 831 357 843 360
rect 785 351 843 357
rect 1733 357 1745 360
rect 1779 388 1791 391
rect 1921 391 1979 397
rect 1921 388 1933 391
rect 1779 360 1933 388
rect 1779 357 1791 360
rect 1733 351 1791 357
rect 1921 357 1933 360
rect 1967 388 1979 391
rect 3173 391 3231 397
rect 3173 388 3185 391
rect 1967 360 3185 388
rect 1967 357 1979 360
rect 1921 351 1979 357
rect 3173 357 3185 360
rect 3219 388 3231 391
rect 3361 391 3419 397
rect 3361 388 3373 391
rect 3219 360 3373 388
rect 3219 357 3231 360
rect 3173 351 3231 357
rect 3361 357 3373 360
rect 3407 388 3419 391
rect 4309 391 4367 397
rect 4309 388 4321 391
rect 3407 360 4321 388
rect 3407 357 3419 360
rect 3361 351 3419 357
rect 4309 357 4321 360
rect 4355 388 4367 391
rect 4497 391 4555 397
rect 4497 388 4509 391
rect 4355 360 4509 388
rect 4355 357 4367 360
rect 4309 351 4367 357
rect 4497 357 4509 360
rect 4543 388 4555 391
rect 5841 391 5899 397
rect 5841 388 5853 391
rect 4543 360 5853 388
rect 4543 357 4555 360
rect 4497 351 4555 357
rect 5841 357 5853 360
rect 5887 388 5899 391
rect 6029 391 6087 397
rect 6029 388 6041 391
rect 5887 360 6041 388
rect 5887 357 5899 360
rect 5841 351 5899 357
rect 6029 357 6041 360
rect 6075 388 6087 391
rect 6977 391 7035 397
rect 6977 388 6989 391
rect 6075 360 6989 388
rect 6075 357 6087 360
rect 6029 351 6087 357
rect 6977 357 6989 360
rect 7023 388 7035 391
rect 7165 391 7223 397
rect 7165 388 7177 391
rect 7023 360 7177 388
rect 7023 357 7035 360
rect 6977 351 7035 357
rect 7165 357 7177 360
rect 7211 388 7223 391
rect 8417 391 8475 397
rect 8417 388 8429 391
rect 7211 360 8429 388
rect 7211 357 7223 360
rect 7165 351 7223 357
rect 8417 357 8429 360
rect 8463 388 8475 391
rect 8605 391 8663 397
rect 8605 388 8617 391
rect 8463 360 8617 388
rect 8463 357 8475 360
rect 8417 351 8475 357
rect 8605 357 8617 360
rect 8651 388 8663 391
rect 9553 391 9611 397
rect 9553 388 9565 391
rect 8651 360 9565 388
rect 8651 357 8663 360
rect 8605 351 8663 357
rect 9553 357 9565 360
rect 9599 388 9611 391
rect 9741 391 9799 397
rect 9741 388 9753 391
rect 9599 360 9753 388
rect 9599 357 9611 360
rect 9553 351 9611 357
rect 9741 357 9753 360
rect 9787 357 9799 391
rect 9741 351 9799 357
rect 0 17 10396 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3341 17
rect 3375 -17 3433 17
rect 3467 -17 3525 17
rect 3559 -17 3617 17
rect 3651 -17 3709 17
rect 3743 -17 3801 17
rect 3835 -17 3893 17
rect 3927 -17 3985 17
rect 4019 -17 4077 17
rect 4111 -17 4169 17
rect 4203 -17 4261 17
rect 4295 -17 4353 17
rect 4387 -17 4445 17
rect 4479 -17 4537 17
rect 4571 -17 4629 17
rect 4663 -17 4721 17
rect 4755 -17 4813 17
rect 4847 -17 4905 17
rect 4939 -17 4997 17
rect 5031 -17 5089 17
rect 5123 -17 5181 17
rect 5215 -17 5273 17
rect 5307 -17 5365 17
rect 5399 -17 5457 17
rect 5491 -17 5549 17
rect 5583 -17 5641 17
rect 5675 -17 5733 17
rect 5767 -17 5825 17
rect 5859 -17 5917 17
rect 5951 -17 6009 17
rect 6043 -17 6101 17
rect 6135 -17 6193 17
rect 6227 -17 6285 17
rect 6319 -17 6377 17
rect 6411 -17 6469 17
rect 6503 -17 6561 17
rect 6595 -17 6653 17
rect 6687 -17 6745 17
rect 6779 -17 6837 17
rect 6871 -17 6929 17
rect 6963 -17 7021 17
rect 7055 -17 7113 17
rect 7147 -17 7205 17
rect 7239 -17 7297 17
rect 7331 -17 7389 17
rect 7423 -17 7481 17
rect 7515 -17 7573 17
rect 7607 -17 7665 17
rect 7699 -17 7757 17
rect 7791 -17 7849 17
rect 7883 -17 7941 17
rect 7975 -17 8033 17
rect 8067 -17 8125 17
rect 8159 -17 8217 17
rect 8251 -17 8309 17
rect 8343 -17 8401 17
rect 8435 -17 8493 17
rect 8527 -17 8585 17
rect 8619 -17 8677 17
rect 8711 -17 8769 17
rect 8803 -17 8861 17
rect 8895 -17 8953 17
rect 8987 -17 9045 17
rect 9079 -17 9137 17
rect 9171 -17 9229 17
rect 9263 -17 9321 17
rect 9355 -17 9413 17
rect 9447 -17 9505 17
rect 9539 -17 9597 17
rect 9631 -17 9689 17
rect 9723 -17 9781 17
rect 9815 -17 9873 17
rect 9907 -17 9965 17
rect 9999 -17 10057 17
rect 10091 -17 10149 17
rect 10183 -17 10241 17
rect 10275 -17 10333 17
rect 10367 -17 10396 17
rect 0 -48 10396 -17
<< labels >>
rlabel comment s 7820 0 7820 0 4 muxb4to1_1
rlabel comment s 7820 1088 7820 1088 4 muxb4to1_1
rlabel comment s 5244 1088 5244 1088 4 muxb4to1_1
rlabel comment s 5152 0 5152 0 4 tap_1
rlabel comment s 5244 0 5244 0 4 muxb4to1_1
rlabel comment s 5152 0 5152 0 4 muxb4to1_1
rlabel comment s 5152 1088 5152 1088 4 muxb4to1_1
rlabel comment s 5152 1088 5152 1088 4 tap_1
rlabel comment s 2576 0 2576 0 4 muxb4to1_1
rlabel comment s 2576 1088 2576 1088 4 muxb4to1_1
rlabel comment s 2576 1088 2576 1088 4 muxb4to1_1
rlabel comment s 2576 0 2576 0 4 muxb4to1_1
rlabel comment s 0 1088 0 1088 4 muxb4to1_1
rlabel comment s 0 0 0 0 4 muxb4to1_1
rlabel comment s 7820 1088 7820 1088 4 muxb4to1_1
rlabel comment s 7820 0 7820 0 4 muxb4to1_1
rlabel comment s 10396 1088 10396 1088 4 muxb4to1_1
rlabel comment s 10396 0 10396 0 4 muxb4to1_1
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 33 nsew
flabel metal1 s 609 697 643 731 0 FreeSans 200 0 0 0 Z
port 37 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 36 nsew
flabel metal1 s 609 357 643 391 0 FreeSans 200 0 0 0 Z
port 37 nsew
flabel metal1 s 29 1071 63 1105 0 FreeSans 200 0 0 0 VGND
port 33 nsew
flabel metal1 s 7757 527 7791 561 0 FreeSans 200 180 0 0 VPWR
port 36 nsew
flabel metal1 s 7757 -17 7791 17 0 FreeSans 200 180 0 0 VGND
port 33 nsew
flabel metal1 s 7774 544 7774 544 0 FreeSans 200 180 0 0 VPWR
port 36 nsew
flabel metal1 s 7757 1071 7791 1105 0 FreeSans 200 180 0 0 VGND
port 33 nsew
flabel metal1 s 5178 533 5221 555 0 FreeSans 200 0 0 0 VPWR
port 36 nsew
flabel metal1 s 5180 -10 5220 14 0 FreeSans 200 0 0 0 VGND
port 33 nsew
flabel metal1 s 5273 527 5307 561 0 FreeSans 200 0 0 0 VPWR
port 36 nsew
flabel metal1 s 5273 -17 5307 17 0 FreeSans 200 0 0 0 VGND
port 33 nsew
flabel metal1 s 5290 544 5290 544 0 FreeSans 200 0 0 0 VPWR
port 36 nsew
flabel metal1 s 5273 1071 5307 1105 0 FreeSans 200 0 0 0 VGND
port 33 nsew
flabel metal1 s 5089 527 5123 561 0 FreeSans 200 180 0 0 VPWR
port 36 nsew
flabel metal1 s 5089 -17 5123 17 0 FreeSans 200 180 0 0 VGND
port 33 nsew
flabel metal1 s 5106 544 5106 544 0 FreeSans 200 180 0 0 VPWR
port 36 nsew
flabel metal1 s 5089 1071 5123 1105 0 FreeSans 200 180 0 0 VGND
port 33 nsew
flabel metal1 s 5198 544 5198 544 0 FreeSans 200 0 0 0 VPWR
port 36 nsew
flabel metal1 s 5180 1074 5220 1098 0 FreeSans 200 0 0 0 VGND
port 33 nsew
flabel metal1 s 2513 527 2547 561 0 FreeSans 200 180 0 0 VPWR
port 36 nsew
flabel metal1 s 2513 -17 2547 17 0 FreeSans 200 180 0 0 VGND
port 33 nsew
flabel metal1 s 2530 544 2530 544 0 FreeSans 200 180 0 0 VPWR
port 36 nsew
flabel metal1 s 2513 1071 2547 1105 0 FreeSans 200 180 0 0 VGND
port 33 nsew
flabel metal1 s 2605 527 2639 561 0 FreeSans 200 0 0 0 VPWR
port 36 nsew
flabel metal1 s 2605 1071 2639 1105 0 FreeSans 200 0 0 0 VGND
port 33 nsew
flabel metal1 s 2622 544 2622 544 0 FreeSans 200 0 0 0 VPWR
port 36 nsew
flabel metal1 s 2605 -17 2639 17 0 FreeSans 200 0 0 0 VGND
port 33 nsew
flabel metal1 s 46 544 46 544 0 FreeSans 200 0 0 0 VPWR
port 36 nsew
flabel metal1 s 46 1088 46 1088 0 FreeSans 200 0 0 0 VGND
port 33 nsew
flabel metal1 s 46 544 46 544 0 FreeSans 200 0 0 0 VPWR
port 36 nsew
flabel metal1 s 46 0 46 0 0 FreeSans 200 0 0 0 VGND
port 33 nsew
flabel metal1 s 7849 527 7883 561 0 FreeSans 200 0 0 0 VPWR
port 36 nsew
flabel metal1 s 7849 1071 7883 1105 0 FreeSans 200 0 0 0 VGND
port 33 nsew
flabel metal1 s 7866 544 7866 544 0 FreeSans 200 0 0 0 VPWR
port 36 nsew
flabel metal1 s 7849 -17 7883 17 0 FreeSans 200 0 0 0 VGND
port 33 nsew
flabel metal1 s 10333 527 10367 561 0 FreeSans 200 180 0 0 VPWR
port 36 nsew
flabel metal1 s 10333 1071 10367 1105 0 FreeSans 200 180 0 0 VGND
port 33 nsew
flabel metal1 s 10350 544 10350 544 0 FreeSans 200 180 0 0 VPWR
port 36 nsew
flabel metal1 s 10333 -17 10367 17 0 FreeSans 200 180 0 0 VGND
port 33 nsew
flabel pwell s 7757 -17 7791 17 0 FreeSans 200 180 0 0 VNB
port 34 nsew
flabel pwell s 7757 1071 7791 1105 0 FreeSans 200 180 0 0 VNB
port 34 nsew
flabel pwell s 5273 -17 5307 17 0 FreeSans 200 0 0 0 VNB
port 34 nsew
flabel pwell s 5273 1071 5307 1105 0 FreeSans 200 0 0 0 VNB
port 34 nsew
flabel pwell s 5089 -17 5123 17 0 FreeSans 200 180 0 0 VNB
port 34 nsew
flabel pwell s 5089 1071 5123 1105 0 FreeSans 200 180 0 0 VNB
port 34 nsew
flabel pwell s 2513 -17 2547 17 0 FreeSans 200 180 0 0 VNB
port 34 nsew
flabel pwell s 2513 1071 2547 1105 0 FreeSans 200 180 0 0 VNB
port 34 nsew
flabel pwell s 2605 1071 2639 1105 0 FreeSans 200 0 0 0 VNB
port 34 nsew
flabel pwell s 2605 -17 2639 17 0 FreeSans 200 0 0 0 VNB
port 34 nsew
flabel pwell s 29 1071 63 1105 0 FreeSans 200 0 0 0 VNB
port 34 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 34 nsew
flabel pwell s 7849 1071 7883 1105 0 FreeSans 200 0 0 0 VNB
port 34 nsew
flabel pwell s 7849 -17 7883 17 0 FreeSans 200 0 0 0 VNB
port 34 nsew
flabel pwell s 10333 1071 10367 1105 0 FreeSans 200 180 0 0 VNB
port 34 nsew
flabel pwell s 10333 -17 10367 17 0 FreeSans 200 180 0 0 VNB
port 34 nsew
flabel nbase s 7757 527 7791 561 0 FreeSans 200 180 0 0 VPB
port 35 nsew
flabel nbase s 7774 544 7774 544 0 FreeSans 200 180 0 0 VPB
port 35 nsew
flabel nbase s 5273 527 5307 561 0 FreeSans 200 0 0 0 VPB
port 35 nsew
flabel nbase s 5290 544 5290 544 0 FreeSans 200 0 0 0 VPB
port 35 nsew
flabel nbase s 5089 527 5123 561 0 FreeSans 200 180 0 0 VPB
port 35 nsew
flabel nbase s 5106 544 5106 544 0 FreeSans 200 180 0 0 VPB
port 35 nsew
flabel nbase s 2513 527 2547 561 0 FreeSans 200 180 0 0 VPB
port 35 nsew
flabel nbase s 2530 544 2530 544 0 FreeSans 200 180 0 0 VPB
port 35 nsew
flabel nbase s 2605 527 2639 561 0 FreeSans 200 0 0 0 VPB
port 35 nsew
flabel nbase s 2622 544 2622 544 0 FreeSans 200 0 0 0 VPB
port 35 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 35 nsew
flabel nbase s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
port 35 nsew
flabel nbase s 7849 527 7883 561 0 FreeSans 200 0 0 0 VPB
port 35 nsew
flabel nbase s 7866 544 7866 544 0 FreeSans 200 0 0 0 VPB
port 35 nsew
flabel nbase s 10333 527 10367 561 0 FreeSans 200 180 0 0 VPB
port 35 nsew
flabel nbase s 10350 544 10350 544 0 FreeSans 200 180 0 0 VPB
port 35 nsew
flabel corelocali s 5181 969 5215 1003 0 FreeSans 200 0 0 0 VNB
port 34 nsew
flabel corelocali s 5181 425 5215 459 0 FreeSans 200 0 0 0 VPB
port 35 nsew
flabel corelocali s 9045 221 9079 255 0 FreeSans 200 0 0 0 S[6]
port 26 nsew
flabel corelocali s 3801 833 3835 867 0 FreeSans 200 0 0 0 S[10]
port 22 nsew
flabel corelocali s 5365 833 5399 867 0 FreeSans 200 0 0 0 D[12]
port 4 nsew
flabel corelocali s 7665 833 7699 867 0 FreeSans 200 0 0 0 D[13]
port 3 nsew
flabel corelocali s 121 833 155 867 0 FreeSans 200 0 0 0 D[8]
port 8 nsew
flabel corelocali s 10241 833 10275 867 0 FreeSans 200 0 0 0 D[15]
port 1 nsew
flabel corelocali s 2697 833 2731 867 0 FreeSans 200 0 0 0 D[10]
port 6 nsew
flabel corelocali s 2421 833 2455 867 0 FreeSans 200 0 0 0 D[9]
port 7 nsew
flabel corelocali s 7941 833 7975 867 0 FreeSans 200 0 0 0 D[14]
port 2 nsew
flabel corelocali s 9045 833 9079 867 0 FreeSans 200 0 0 0 S[14]
port 18 nsew
flabel corelocali s 4997 833 5031 867 0 FreeSans 200 0 0 0 D[11]
port 5 nsew
flabel corelocali s 3893 833 3927 867 0 FreeSans 200 0 0 0 S[11]
port 21 nsew
flabel corelocali s 1225 833 1259 867 0 FreeSans 200 0 0 0 S[8]
port 24 nsew
flabel corelocali s 9137 833 9171 867 0 FreeSans 200 0 0 0 S[15]
port 17 nsew
flabel corelocali s 6469 833 6503 867 0 FreeSans 200 0 0 0 S[12]
port 20 nsew
flabel corelocali s 1317 833 1351 867 0 FreeSans 200 0 0 0 S[9]
port 23 nsew
flabel corelocali s 6561 833 6595 867 0 FreeSans 200 0 0 0 S[13]
port 19 nsew
flabel corelocali s 4997 221 5031 255 0 FreeSans 200 0 0 0 D[3]
port 13 nsew
flabel corelocali s 121 221 155 255 0 FreeSans 200 0 0 0 D[0]
port 16 nsew
flabel corelocali s 5365 221 5399 255 0 FreeSans 200 0 0 0 D[4]
port 12 nsew
flabel corelocali s 7665 221 7699 255 0 FreeSans 200 0 0 0 D[5]
port 11 nsew
flabel corelocali s 2697 221 2731 255 0 FreeSans 200 0 0 0 D[2]
port 14 nsew
flabel corelocali s 2421 221 2455 255 0 FreeSans 200 0 0 0 D[1]
port 15 nsew
flabel corelocali s 7941 221 7975 255 0 FreeSans 200 0 0 0 D[6]
port 10 nsew
flabel corelocali s 3801 221 3835 255 0 FreeSans 200 0 0 0 S[2]
port 30 nsew
flabel corelocali s 3893 221 3927 255 0 FreeSans 200 0 0 0 S[3]
port 29 nsew
flabel corelocali s 9137 221 9171 255 0 FreeSans 200 0 0 0 S[7]
port 25 nsew
flabel corelocali s 1225 221 1259 255 0 FreeSans 200 0 0 0 S[0]
port 32 nsew
flabel corelocali s 1317 221 1351 255 0 FreeSans 200 0 0 0 S[1]
port 31 nsew
flabel corelocali s 6469 221 6503 255 0 FreeSans 200 0 0 0 S[4]
port 28 nsew
flabel corelocali s 6561 221 6595 255 0 FreeSans 200 0 0 0 S[5]
port 27 nsew
flabel corelocali s 10241 221 10275 255 0 FreeSans 200 0 0 0 D[7]
port 9 nsew
flabel corelocali s 5181 629 5215 663 0 FreeSans 200 0 0 0 VPB
port 35 nsew
flabel corelocali s 5181 85 5215 119 0 FreeSans 200 0 0 0 VNB
port 34 nsew
flabel corelocali s 5181 362 5209 386 0 FreeSans 250 0 0 0 VPB
port 35 nsew
flabel corelocali s 5198 102 5198 102 0 FreeSans 250 0 0 0 VNB
port 34 nsew
flabel corelocali s 5181 702 5209 726 0 FreeSans 250 0 0 0 VPB
port 35 nsew
flabel corelocali s 5190 975 5206 994 0 FreeSans 250 0 0 0 VNB
port 34 nsew
<< properties >>
string FIXED_BBOX 0 0 10396 1088
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3268980
string GDS_START 3118284
string path 128.800 13.600 131.100 13.600 
<< end >>
