magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 2208 561
rect 28 299 81 527
rect 115 333 166 493
rect 200 367 252 527
rect 287 333 338 490
rect 373 367 424 527
rect 465 333 510 493
rect 544 367 596 527
rect 631 333 682 490
rect 717 367 768 527
rect 803 333 851 490
rect 893 367 944 527
rect 981 333 1056 490
rect 1098 424 1150 527
rect 1098 367 1149 424
rect 1185 333 1235 490
rect 1271 367 1322 527
rect 1357 333 1407 490
rect 1443 367 1494 527
rect 1529 333 1579 490
rect 1615 367 1666 527
rect 1701 333 1751 490
rect 1787 367 1838 527
rect 1873 333 1921 490
rect 1959 367 2010 527
rect 2045 333 2096 490
rect 2130 367 2182 527
rect 115 291 2096 333
rect 465 283 1751 291
rect 69 179 431 255
rect 371 17 425 122
rect 465 56 510 283
rect 544 17 597 122
rect 631 56 682 283
rect 716 17 769 122
rect 803 56 851 283
rect 893 17 946 122
rect 981 56 1051 283
rect 1098 17 1151 122
rect 1185 56 1235 283
rect 1270 17 1315 122
rect 1357 56 1407 283
rect 1442 17 1495 122
rect 1529 56 1579 283
rect 1614 17 1667 122
rect 1701 56 1751 283
rect 1786 179 2142 255
rect 1786 17 1839 122
rect 0 -17 2208 17
<< metal1 >>
rect 0 496 2208 592
rect 293 252 443 261
rect 1857 252 2007 261
rect 293 224 2007 252
rect 293 215 443 224
rect 1857 215 2007 224
rect 0 -48 2208 48
<< labels >>
rlabel locali s 69 179 431 255 6 A
port 1 nsew signal input
rlabel locali s 1786 179 2142 255 6 A
port 1 nsew signal input
rlabel metal1 s 1857 252 2007 261 6 A
port 1 nsew signal input
rlabel metal1 s 1857 215 2007 224 6 A
port 1 nsew signal input
rlabel metal1 s 293 252 443 261 6 A
port 1 nsew signal input
rlabel metal1 s 293 224 2007 252 6 A
port 1 nsew signal input
rlabel metal1 s 293 215 443 224 6 A
port 1 nsew signal input
rlabel locali s 2045 333 2096 490 6 Y
port 2 nsew signal output
rlabel locali s 1873 333 1921 490 6 Y
port 2 nsew signal output
rlabel locali s 1701 333 1751 490 6 Y
port 2 nsew signal output
rlabel locali s 1701 56 1751 283 6 Y
port 2 nsew signal output
rlabel locali s 1529 333 1579 490 6 Y
port 2 nsew signal output
rlabel locali s 1529 56 1579 283 6 Y
port 2 nsew signal output
rlabel locali s 1357 333 1407 490 6 Y
port 2 nsew signal output
rlabel locali s 1357 56 1407 283 6 Y
port 2 nsew signal output
rlabel locali s 1185 333 1235 490 6 Y
port 2 nsew signal output
rlabel locali s 1185 56 1235 283 6 Y
port 2 nsew signal output
rlabel locali s 981 333 1056 490 6 Y
port 2 nsew signal output
rlabel locali s 981 56 1051 283 6 Y
port 2 nsew signal output
rlabel locali s 803 333 851 490 6 Y
port 2 nsew signal output
rlabel locali s 803 56 851 283 6 Y
port 2 nsew signal output
rlabel locali s 631 333 682 490 6 Y
port 2 nsew signal output
rlabel locali s 631 56 682 283 6 Y
port 2 nsew signal output
rlabel locali s 465 333 510 493 6 Y
port 2 nsew signal output
rlabel locali s 465 283 1751 291 6 Y
port 2 nsew signal output
rlabel locali s 465 56 510 283 6 Y
port 2 nsew signal output
rlabel locali s 287 333 338 490 6 Y
port 2 nsew signal output
rlabel locali s 115 333 166 493 6 Y
port 2 nsew signal output
rlabel locali s 115 291 2096 333 6 Y
port 2 nsew signal output
rlabel locali s 1786 17 1839 122 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1614 17 1667 122 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1442 17 1495 122 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1270 17 1315 122 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1098 17 1151 122 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 893 17 946 122 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 716 17 769 122 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 544 17 597 122 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 371 17 425 122 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 0 -17 2208 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 2208 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 2130 367 2182 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1959 367 2010 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1787 367 1838 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1615 367 1666 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1443 367 1494 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1271 367 1322 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1098 424 1150 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1098 367 1149 424 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 893 367 944 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 717 367 768 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 544 367 596 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 373 367 424 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 200 367 252 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 28 299 81 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 0 527 2208 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 496 2208 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2208 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3215186
string GDS_START 3202198
<< end >>
