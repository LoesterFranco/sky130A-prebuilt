magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 89 47 119 131
rect 287 47 317 177
rect 381 47 411 177
rect 465 47 495 177
rect 559 47 589 177
rect 767 47 797 177
rect 861 47 891 177
rect 973 47 1003 177
rect 1067 47 1097 177
<< pmoshvt >>
rect 81 413 117 497
rect 279 297 315 497
rect 373 297 409 497
rect 467 297 503 497
rect 561 297 597 497
rect 749 297 785 497
rect 843 297 879 497
rect 955 297 991 497
rect 1049 297 1085 497
<< ndiff >>
rect 225 161 287 177
rect 27 103 89 131
rect 27 69 35 103
rect 69 69 89 103
rect 27 47 89 69
rect 119 93 171 131
rect 119 59 129 93
rect 163 59 171 93
rect 119 47 171 59
rect 225 127 233 161
rect 267 127 287 161
rect 225 93 287 127
rect 225 59 233 93
rect 267 59 287 93
rect 225 47 287 59
rect 317 161 381 177
rect 317 127 327 161
rect 361 127 381 161
rect 317 47 381 127
rect 411 127 465 177
rect 411 93 421 127
rect 455 93 465 127
rect 411 47 465 93
rect 495 93 559 177
rect 495 59 515 93
rect 549 59 559 93
rect 495 47 559 59
rect 589 161 651 177
rect 589 127 609 161
rect 643 127 651 161
rect 589 47 651 127
rect 705 161 767 177
rect 705 127 713 161
rect 747 127 767 161
rect 705 47 767 127
rect 797 93 861 177
rect 797 59 807 93
rect 841 59 861 93
rect 797 47 861 59
rect 891 169 973 177
rect 891 135 910 169
rect 944 135 973 169
rect 891 101 973 135
rect 891 67 910 101
rect 944 67 973 101
rect 891 47 973 67
rect 1003 93 1067 177
rect 1003 59 1013 93
rect 1047 59 1067 93
rect 1003 47 1067 59
rect 1097 161 1149 177
rect 1097 127 1107 161
rect 1141 127 1149 161
rect 1097 93 1149 127
rect 1097 59 1107 93
rect 1141 59 1149 93
rect 1097 47 1149 59
<< pdiff >>
rect 27 475 81 497
rect 27 441 35 475
rect 69 441 81 475
rect 27 413 81 441
rect 117 485 171 497
rect 117 451 129 485
rect 163 451 171 485
rect 117 413 171 451
rect 225 485 279 497
rect 225 451 233 485
rect 267 451 279 485
rect 225 417 279 451
rect 225 383 233 417
rect 267 383 279 417
rect 225 349 279 383
rect 225 315 233 349
rect 267 315 279 349
rect 225 297 279 315
rect 315 485 373 497
rect 315 451 327 485
rect 361 451 373 485
rect 315 417 373 451
rect 315 383 327 417
rect 361 383 373 417
rect 315 349 373 383
rect 315 315 327 349
rect 361 315 373 349
rect 315 297 373 315
rect 409 485 467 497
rect 409 451 421 485
rect 455 451 467 485
rect 409 417 467 451
rect 409 383 421 417
rect 455 383 467 417
rect 409 297 467 383
rect 503 485 561 497
rect 503 451 515 485
rect 549 451 561 485
rect 503 417 561 451
rect 503 383 515 417
rect 549 383 561 417
rect 503 349 561 383
rect 503 315 515 349
rect 549 315 561 349
rect 503 297 561 315
rect 597 485 749 497
rect 597 451 609 485
rect 643 451 687 485
rect 721 451 749 485
rect 597 417 749 451
rect 597 383 609 417
rect 643 383 687 417
rect 721 383 749 417
rect 597 297 749 383
rect 785 485 843 497
rect 785 451 797 485
rect 831 451 843 485
rect 785 417 843 451
rect 785 383 797 417
rect 831 383 843 417
rect 785 349 843 383
rect 785 315 797 349
rect 831 315 843 349
rect 785 297 843 315
rect 879 485 955 497
rect 879 451 898 485
rect 932 451 955 485
rect 879 417 955 451
rect 879 383 898 417
rect 932 383 955 417
rect 879 297 955 383
rect 991 485 1049 497
rect 991 451 1003 485
rect 1037 451 1049 485
rect 991 417 1049 451
rect 991 383 1003 417
rect 1037 383 1049 417
rect 991 297 1049 383
rect 1085 485 1167 497
rect 1085 451 1113 485
rect 1147 451 1167 485
rect 1085 417 1167 451
rect 1085 383 1113 417
rect 1147 383 1167 417
rect 1085 349 1167 383
rect 1085 315 1113 349
rect 1147 315 1167 349
rect 1085 297 1167 315
<< ndiffc >>
rect 35 69 69 103
rect 129 59 163 93
rect 233 127 267 161
rect 233 59 267 93
rect 327 127 361 161
rect 421 93 455 127
rect 515 59 549 93
rect 609 127 643 161
rect 713 127 747 161
rect 807 59 841 93
rect 910 135 944 169
rect 910 67 944 101
rect 1013 59 1047 93
rect 1107 127 1141 161
rect 1107 59 1141 93
<< pdiffc >>
rect 35 441 69 475
rect 129 451 163 485
rect 233 451 267 485
rect 233 383 267 417
rect 233 315 267 349
rect 327 451 361 485
rect 327 383 361 417
rect 327 315 361 349
rect 421 451 455 485
rect 421 383 455 417
rect 515 451 549 485
rect 515 383 549 417
rect 515 315 549 349
rect 609 451 643 485
rect 687 451 721 485
rect 609 383 643 417
rect 687 383 721 417
rect 797 451 831 485
rect 797 383 831 417
rect 797 315 831 349
rect 898 451 932 485
rect 898 383 932 417
rect 1003 451 1037 485
rect 1003 383 1037 417
rect 1113 451 1147 485
rect 1113 383 1147 417
rect 1113 315 1147 349
<< poly >>
rect 81 497 117 523
rect 279 497 315 523
rect 373 497 409 523
rect 467 497 503 523
rect 561 497 597 523
rect 749 497 785 523
rect 843 497 879 523
rect 955 497 991 523
rect 1049 497 1085 523
rect 81 398 117 413
rect 79 265 119 398
rect 279 282 315 297
rect 373 282 409 297
rect 467 282 503 297
rect 561 282 597 297
rect 749 282 785 297
rect 843 282 879 297
rect 955 282 991 297
rect 1049 282 1085 297
rect 277 265 317 282
rect 371 265 411 282
rect 22 249 119 265
rect 22 215 32 249
rect 66 215 119 249
rect 22 199 119 215
rect 201 249 411 265
rect 201 215 217 249
rect 251 215 411 249
rect 201 199 411 215
rect 89 131 119 199
rect 287 177 317 199
rect 381 177 411 199
rect 465 265 505 282
rect 559 265 599 282
rect 747 265 787 282
rect 841 265 881 282
rect 953 265 993 282
rect 1047 265 1087 282
rect 465 249 656 265
rect 465 215 485 249
rect 519 215 606 249
rect 640 215 656 249
rect 465 199 656 215
rect 747 249 911 265
rect 747 215 763 249
rect 797 215 847 249
rect 881 215 911 249
rect 747 199 911 215
rect 953 249 1172 265
rect 953 215 1020 249
rect 1054 215 1122 249
rect 1156 215 1172 249
rect 953 199 1172 215
rect 465 177 495 199
rect 559 177 589 199
rect 767 177 797 199
rect 861 177 891 199
rect 973 177 1003 199
rect 1067 177 1097 199
rect 89 21 119 47
rect 287 21 317 47
rect 381 21 411 47
rect 465 21 495 47
rect 559 21 589 47
rect 767 21 797 47
rect 861 21 891 47
rect 973 21 1003 47
rect 1067 21 1097 47
<< polycont >>
rect 32 215 66 249
rect 217 215 251 249
rect 485 215 519 249
rect 606 215 640 249
rect 763 215 797 249
rect 847 215 881 249
rect 1020 215 1054 249
rect 1122 215 1156 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 18 475 69 493
rect 18 441 35 475
rect 103 485 267 527
rect 103 451 129 485
rect 163 451 233 485
rect 18 417 69 441
rect 217 417 267 451
rect 18 383 144 417
rect 18 249 66 323
rect 18 215 32 249
rect 18 199 66 215
rect 100 249 144 383
rect 217 383 233 417
rect 217 349 267 383
rect 217 315 233 349
rect 217 289 267 315
rect 301 485 377 493
rect 301 451 327 485
rect 361 451 377 485
rect 301 417 377 451
rect 301 383 327 417
rect 361 383 377 417
rect 301 349 377 383
rect 421 485 455 527
rect 421 417 455 451
rect 421 367 455 383
rect 489 485 565 493
rect 489 451 515 485
rect 549 451 565 485
rect 489 417 565 451
rect 489 383 515 417
rect 549 383 565 417
rect 301 315 327 349
rect 361 333 377 349
rect 489 349 565 383
rect 609 485 737 527
rect 643 451 687 485
rect 721 451 737 485
rect 609 417 737 451
rect 643 383 687 417
rect 721 383 737 417
rect 609 367 737 383
rect 771 485 847 493
rect 771 451 797 485
rect 831 451 847 485
rect 771 417 847 451
rect 771 383 797 417
rect 831 383 847 417
rect 489 333 515 349
rect 361 315 515 333
rect 549 333 565 349
rect 771 349 847 383
rect 891 485 943 527
rect 891 451 898 485
rect 932 451 943 485
rect 891 417 943 451
rect 891 383 898 417
rect 932 383 943 417
rect 891 367 943 383
rect 977 485 1053 493
rect 977 451 1003 485
rect 1037 451 1053 485
rect 977 417 1053 451
rect 977 383 1003 417
rect 1037 383 1053 417
rect 771 333 797 349
rect 549 315 797 333
rect 831 333 847 349
rect 977 333 1053 383
rect 831 315 1053 333
rect 301 289 1053 315
rect 1097 485 1176 527
rect 1097 451 1113 485
rect 1147 451 1176 485
rect 1097 417 1176 451
rect 1097 383 1113 417
rect 1147 383 1176 417
rect 1097 349 1176 383
rect 1097 315 1113 349
rect 1147 315 1176 349
rect 1097 299 1176 315
rect 100 215 217 249
rect 251 215 267 249
rect 100 161 144 215
rect 18 127 144 161
rect 217 161 267 181
rect 217 127 233 161
rect 301 161 377 289
rect 432 249 670 255
rect 432 215 485 249
rect 519 215 606 249
rect 640 215 670 249
rect 722 249 937 255
rect 722 215 763 249
rect 797 215 847 249
rect 881 215 937 249
rect 1004 249 1177 255
rect 1004 215 1020 249
rect 1054 215 1122 249
rect 1156 215 1177 249
rect 301 127 327 161
rect 361 127 377 161
rect 421 161 659 181
rect 421 127 609 161
rect 643 127 659 161
rect 697 169 1158 181
rect 697 161 910 169
rect 697 127 713 161
rect 747 135 910 161
rect 944 161 1158 169
rect 944 143 1107 161
rect 944 135 961 143
rect 747 127 961 135
rect 18 103 69 127
rect 18 69 35 103
rect 217 93 267 127
rect 901 123 961 127
rect 1091 127 1107 143
rect 1141 127 1158 161
rect 901 101 953 123
rect 18 51 69 69
rect 103 59 129 93
rect 163 59 179 93
rect 103 17 179 59
rect 217 59 233 93
rect 267 59 455 93
rect 217 51 455 59
rect 489 59 515 93
rect 549 59 807 93
rect 841 59 857 93
rect 489 51 857 59
rect 901 67 910 101
rect 944 67 953 101
rect 901 51 953 67
rect 1013 93 1047 109
rect 1013 17 1047 59
rect 1091 93 1158 127
rect 1091 59 1107 93
rect 1141 59 1158 93
rect 1091 51 1158 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
flabel corelocali s 1036 221 1070 255 0 FreeSans 250 0 0 0 D
port 4 nsew
flabel corelocali s 1130 221 1164 255 0 FreeSans 250 0 0 0 D
port 4 nsew
flabel corelocali s 855 221 889 255 0 FreeSans 250 0 0 0 C
port 3 nsew
flabel corelocali s 763 221 797 255 0 FreeSans 250 0 0 0 C
port 3 nsew
flabel corelocali s 587 221 621 255 0 FreeSans 250 0 0 0 B
port 2 nsew
flabel corelocali s 491 221 525 255 0 FreeSans 250 0 0 0 B
port 2 nsew
flabel corelocali s 309 153 343 187 0 FreeSans 250 0 0 0 Y
port 9 nsew
flabel corelocali s 310 221 344 255 0 FreeSans 250 0 0 0 Y
port 9 nsew
flabel corelocali s 310 289 344 323 0 FreeSans 250 0 0 0 Y
port 9 nsew
flabel corelocali s 30 289 64 323 0 FreeSans 250 0 0 0 A_N
port 1 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 250 0 0 0 A_N
port 1 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
rlabel comment s 0 0 0 0 4 nand4b_2
<< properties >>
string FIXED_BBOX 0 0 1196 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2331924
string GDS_START 2321864
<< end >>
