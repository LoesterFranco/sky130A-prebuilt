magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 373 518 439 602
rect 133 484 439 518
rect 133 366 167 484
rect 373 468 439 484
rect 85 300 167 366
rect 201 300 359 366
rect 647 364 751 596
rect 717 226 751 364
rect 642 70 751 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 17 400 89 576
rect 130 552 196 649
rect 17 264 51 400
rect 237 434 339 450
rect 237 400 427 434
rect 473 410 539 649
rect 393 376 427 400
rect 393 342 613 376
rect 492 330 613 342
rect 374 264 440 268
rect 17 230 440 264
rect 492 264 683 330
rect 17 91 106 230
rect 492 196 532 264
rect 140 17 197 170
rect 231 162 532 196
rect 231 91 290 162
rect 478 17 544 128
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel locali s 201 300 359 366 6 A
port 1 nsew signal input
rlabel locali s 373 518 439 602 6 TE_B
port 2 nsew signal input
rlabel locali s 373 468 439 484 6 TE_B
port 2 nsew signal input
rlabel locali s 133 484 439 518 6 TE_B
port 2 nsew signal input
rlabel locali s 133 366 167 484 6 TE_B
port 2 nsew signal input
rlabel locali s 85 300 167 366 6 TE_B
port 2 nsew signal input
rlabel locali s 717 226 751 364 6 Z
port 3 nsew signal output
rlabel locali s 647 364 751 596 6 Z
port 3 nsew signal output
rlabel locali s 642 70 751 226 6 Z
port 3 nsew signal output
rlabel metal1 s 0 -49 768 49 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 617 768 715 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2043556
string GDS_START 2037166
<< end >>
