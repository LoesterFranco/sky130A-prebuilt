magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 1694 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 83 47 113 177
rect 177 47 207 177
rect 271 47 301 177
rect 365 47 395 177
rect 459 47 489 177
rect 553 47 583 177
rect 647 47 677 177
rect 751 47 781 177
rect 835 47 865 177
rect 929 47 959 177
rect 1023 47 1053 177
rect 1117 47 1147 177
rect 1211 47 1241 177
rect 1305 47 1335 177
rect 1399 47 1429 177
rect 1503 47 1533 177
<< pmoshvt >>
rect 85 297 121 497
rect 179 297 215 497
rect 273 297 309 497
rect 367 297 403 497
rect 461 297 497 497
rect 555 297 591 497
rect 649 297 685 497
rect 743 297 779 497
rect 837 297 873 497
rect 931 297 967 497
rect 1025 297 1061 497
rect 1119 297 1155 497
rect 1213 297 1249 497
rect 1307 297 1343 497
rect 1401 297 1437 497
rect 1495 297 1531 497
<< ndiff >>
rect 27 163 83 177
rect 27 129 39 163
rect 73 129 83 163
rect 27 95 83 129
rect 27 61 39 95
rect 73 61 83 95
rect 27 47 83 61
rect 113 163 177 177
rect 113 129 133 163
rect 167 129 177 163
rect 113 95 177 129
rect 113 61 133 95
rect 167 61 177 95
rect 113 47 177 61
rect 207 95 271 177
rect 207 61 227 95
rect 261 61 271 95
rect 207 47 271 61
rect 301 163 365 177
rect 301 129 321 163
rect 355 129 365 163
rect 301 95 365 129
rect 301 61 321 95
rect 355 61 365 95
rect 301 47 365 61
rect 395 95 459 177
rect 395 61 415 95
rect 449 61 459 95
rect 395 47 459 61
rect 489 163 553 177
rect 489 129 509 163
rect 543 129 553 163
rect 489 95 553 129
rect 489 61 509 95
rect 543 61 553 95
rect 489 47 553 61
rect 583 95 647 177
rect 583 61 603 95
rect 637 61 647 95
rect 583 47 647 61
rect 677 163 751 177
rect 677 129 697 163
rect 731 129 751 163
rect 677 95 751 129
rect 677 61 697 95
rect 731 61 751 95
rect 677 47 751 61
rect 781 95 835 177
rect 781 61 791 95
rect 825 61 835 95
rect 781 47 835 61
rect 865 163 929 177
rect 865 129 885 163
rect 919 129 929 163
rect 865 95 929 129
rect 865 61 885 95
rect 919 61 929 95
rect 865 47 929 61
rect 959 95 1023 177
rect 959 61 979 95
rect 1013 61 1023 95
rect 959 47 1023 61
rect 1053 163 1117 177
rect 1053 129 1073 163
rect 1107 129 1117 163
rect 1053 95 1117 129
rect 1053 61 1073 95
rect 1107 61 1117 95
rect 1053 47 1117 61
rect 1147 95 1211 177
rect 1147 61 1167 95
rect 1201 61 1211 95
rect 1147 47 1211 61
rect 1241 163 1305 177
rect 1241 129 1261 163
rect 1295 129 1305 163
rect 1241 95 1305 129
rect 1241 61 1261 95
rect 1295 61 1305 95
rect 1241 47 1305 61
rect 1335 95 1399 177
rect 1335 61 1355 95
rect 1389 61 1399 95
rect 1335 47 1399 61
rect 1429 163 1503 177
rect 1429 129 1449 163
rect 1483 129 1503 163
rect 1429 95 1503 129
rect 1429 61 1449 95
rect 1483 61 1503 95
rect 1429 47 1503 61
rect 1533 95 1585 177
rect 1533 61 1543 95
rect 1577 61 1585 95
rect 1533 47 1585 61
<< pdiff >>
rect 27 477 85 497
rect 27 443 39 477
rect 73 443 85 477
rect 27 409 85 443
rect 27 375 39 409
rect 73 375 85 409
rect 27 341 85 375
rect 27 307 39 341
rect 73 307 85 341
rect 27 297 85 307
rect 121 485 179 497
rect 121 451 133 485
rect 167 451 179 485
rect 121 417 179 451
rect 121 383 133 417
rect 167 383 179 417
rect 121 297 179 383
rect 215 477 273 497
rect 215 443 227 477
rect 261 443 273 477
rect 215 409 273 443
rect 215 375 227 409
rect 261 375 273 409
rect 215 341 273 375
rect 215 307 227 341
rect 261 307 273 341
rect 215 297 273 307
rect 309 485 367 497
rect 309 451 321 485
rect 355 451 367 485
rect 309 417 367 451
rect 309 383 321 417
rect 355 383 367 417
rect 309 297 367 383
rect 403 477 461 497
rect 403 443 415 477
rect 449 443 461 477
rect 403 409 461 443
rect 403 375 415 409
rect 449 375 461 409
rect 403 341 461 375
rect 403 307 415 341
rect 449 307 461 341
rect 403 297 461 307
rect 497 485 555 497
rect 497 451 509 485
rect 543 451 555 485
rect 497 417 555 451
rect 497 383 509 417
rect 543 383 555 417
rect 497 297 555 383
rect 591 477 649 497
rect 591 443 603 477
rect 637 443 649 477
rect 591 409 649 443
rect 591 375 603 409
rect 637 375 649 409
rect 591 341 649 375
rect 591 307 603 341
rect 637 307 649 341
rect 591 297 649 307
rect 685 485 743 497
rect 685 451 697 485
rect 731 451 743 485
rect 685 417 743 451
rect 685 383 697 417
rect 731 383 743 417
rect 685 297 743 383
rect 779 477 837 497
rect 779 443 791 477
rect 825 443 837 477
rect 779 409 837 443
rect 779 375 791 409
rect 825 375 837 409
rect 779 341 837 375
rect 779 307 791 341
rect 825 307 837 341
rect 779 297 837 307
rect 873 409 931 497
rect 873 375 885 409
rect 919 375 931 409
rect 873 341 931 375
rect 873 307 885 341
rect 919 307 931 341
rect 873 297 931 307
rect 967 477 1025 497
rect 967 443 979 477
rect 1013 443 1025 477
rect 967 409 1025 443
rect 967 375 979 409
rect 1013 375 1025 409
rect 967 297 1025 375
rect 1061 409 1119 497
rect 1061 375 1073 409
rect 1107 375 1119 409
rect 1061 341 1119 375
rect 1061 307 1073 341
rect 1107 307 1119 341
rect 1061 297 1119 307
rect 1155 477 1213 497
rect 1155 443 1167 477
rect 1201 443 1213 477
rect 1155 409 1213 443
rect 1155 375 1167 409
rect 1201 375 1213 409
rect 1155 297 1213 375
rect 1249 409 1307 497
rect 1249 375 1261 409
rect 1295 375 1307 409
rect 1249 341 1307 375
rect 1249 307 1261 341
rect 1295 307 1307 341
rect 1249 297 1307 307
rect 1343 477 1401 497
rect 1343 443 1355 477
rect 1389 443 1401 477
rect 1343 409 1401 443
rect 1343 375 1355 409
rect 1389 375 1401 409
rect 1343 297 1401 375
rect 1437 409 1495 497
rect 1437 375 1449 409
rect 1483 375 1495 409
rect 1437 341 1495 375
rect 1437 307 1449 341
rect 1483 307 1495 341
rect 1437 297 1495 307
rect 1531 477 1587 497
rect 1531 443 1543 477
rect 1577 443 1587 477
rect 1531 409 1587 443
rect 1531 375 1543 409
rect 1577 375 1587 409
rect 1531 297 1587 375
<< ndiffc >>
rect 39 129 73 163
rect 39 61 73 95
rect 133 129 167 163
rect 133 61 167 95
rect 227 61 261 95
rect 321 129 355 163
rect 321 61 355 95
rect 415 61 449 95
rect 509 129 543 163
rect 509 61 543 95
rect 603 61 637 95
rect 697 129 731 163
rect 697 61 731 95
rect 791 61 825 95
rect 885 129 919 163
rect 885 61 919 95
rect 979 61 1013 95
rect 1073 129 1107 163
rect 1073 61 1107 95
rect 1167 61 1201 95
rect 1261 129 1295 163
rect 1261 61 1295 95
rect 1355 61 1389 95
rect 1449 129 1483 163
rect 1449 61 1483 95
rect 1543 61 1577 95
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 133 451 167 485
rect 133 383 167 417
rect 227 443 261 477
rect 227 375 261 409
rect 227 307 261 341
rect 321 451 355 485
rect 321 383 355 417
rect 415 443 449 477
rect 415 375 449 409
rect 415 307 449 341
rect 509 451 543 485
rect 509 383 543 417
rect 603 443 637 477
rect 603 375 637 409
rect 603 307 637 341
rect 697 451 731 485
rect 697 383 731 417
rect 791 443 825 477
rect 791 375 825 409
rect 791 307 825 341
rect 885 375 919 409
rect 885 307 919 341
rect 979 443 1013 477
rect 979 375 1013 409
rect 1073 375 1107 409
rect 1073 307 1107 341
rect 1167 443 1201 477
rect 1167 375 1201 409
rect 1261 375 1295 409
rect 1261 307 1295 341
rect 1355 443 1389 477
rect 1355 375 1389 409
rect 1449 375 1483 409
rect 1449 307 1483 341
rect 1543 443 1577 477
rect 1543 375 1577 409
<< poly >>
rect 85 497 121 523
rect 179 497 215 523
rect 273 497 309 523
rect 367 497 403 523
rect 461 497 497 523
rect 555 497 591 523
rect 649 497 685 523
rect 743 497 779 523
rect 837 497 873 523
rect 931 497 967 523
rect 1025 497 1061 523
rect 1119 497 1155 523
rect 1213 497 1249 523
rect 1307 497 1343 523
rect 1401 497 1437 523
rect 1495 497 1531 523
rect 85 282 121 297
rect 179 282 215 297
rect 273 282 309 297
rect 367 282 403 297
rect 461 282 497 297
rect 555 282 591 297
rect 649 282 685 297
rect 743 282 779 297
rect 837 282 873 297
rect 931 282 967 297
rect 1025 282 1061 297
rect 1119 282 1155 297
rect 1213 282 1249 297
rect 1307 282 1343 297
rect 1401 282 1437 297
rect 1495 282 1531 297
rect 83 265 123 282
rect 177 265 217 282
rect 271 265 311 282
rect 365 265 405 282
rect 459 265 499 282
rect 553 265 593 282
rect 647 265 687 282
rect 741 265 781 282
rect 83 249 781 265
rect 83 215 103 249
rect 137 215 181 249
rect 215 215 259 249
rect 293 215 337 249
rect 371 215 415 249
rect 449 215 483 249
rect 517 215 561 249
rect 595 215 639 249
rect 673 215 717 249
rect 751 215 781 249
rect 83 199 781 215
rect 83 177 113 199
rect 177 177 207 199
rect 271 177 301 199
rect 365 177 395 199
rect 459 177 489 199
rect 553 177 583 199
rect 647 177 677 199
rect 751 177 781 199
rect 835 265 875 282
rect 929 265 969 282
rect 1023 265 1063 282
rect 1117 265 1157 282
rect 1211 265 1251 282
rect 1305 265 1345 282
rect 1399 265 1439 282
rect 1493 265 1533 282
rect 835 249 1533 265
rect 835 215 858 249
rect 892 215 936 249
rect 970 215 1014 249
rect 1048 215 1092 249
rect 1126 215 1170 249
rect 1204 215 1238 249
rect 1272 215 1316 249
rect 1350 215 1394 249
rect 1428 215 1533 249
rect 835 199 1533 215
rect 835 177 865 199
rect 929 177 959 199
rect 1023 177 1053 199
rect 1117 177 1147 199
rect 1211 177 1241 199
rect 1305 177 1335 199
rect 1399 177 1429 199
rect 1503 177 1533 199
rect 83 21 113 47
rect 177 21 207 47
rect 271 21 301 47
rect 365 21 395 47
rect 459 21 489 47
rect 553 21 583 47
rect 647 21 677 47
rect 751 21 781 47
rect 835 21 865 47
rect 929 21 959 47
rect 1023 21 1053 47
rect 1117 21 1147 47
rect 1211 21 1241 47
rect 1305 21 1335 47
rect 1399 21 1429 47
rect 1503 21 1533 47
<< polycont >>
rect 103 215 137 249
rect 181 215 215 249
rect 259 215 293 249
rect 337 215 371 249
rect 415 215 449 249
rect 483 215 517 249
rect 561 215 595 249
rect 639 215 673 249
rect 717 215 751 249
rect 858 215 892 249
rect 936 215 970 249
rect 1014 215 1048 249
rect 1092 215 1126 249
rect 1170 215 1204 249
rect 1238 215 1272 249
rect 1316 215 1350 249
rect 1394 215 1428 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 18 477 81 493
rect 18 443 39 477
rect 73 443 81 477
rect 18 409 81 443
rect 18 375 39 409
rect 73 375 81 409
rect 18 341 81 375
rect 125 485 175 527
rect 125 451 133 485
rect 167 451 175 485
rect 125 417 175 451
rect 125 383 133 417
rect 167 383 175 417
rect 125 367 175 383
rect 219 477 269 493
rect 219 443 227 477
rect 261 443 269 477
rect 219 409 269 443
rect 219 375 227 409
rect 261 375 269 409
rect 18 307 39 341
rect 73 333 81 341
rect 219 341 269 375
rect 313 485 363 527
rect 313 451 321 485
rect 355 451 363 485
rect 313 417 363 451
rect 313 383 321 417
rect 355 383 363 417
rect 313 367 363 383
rect 407 477 457 493
rect 407 443 415 477
rect 449 443 457 477
rect 407 409 457 443
rect 407 375 415 409
rect 449 375 457 409
rect 219 333 227 341
rect 73 307 227 333
rect 261 333 269 341
rect 407 341 457 375
rect 501 485 551 527
rect 501 451 509 485
rect 543 451 551 485
rect 501 417 551 451
rect 501 383 509 417
rect 543 383 551 417
rect 501 367 551 383
rect 595 477 645 493
rect 595 443 603 477
rect 637 443 645 477
rect 595 409 645 443
rect 595 375 603 409
rect 637 375 645 409
rect 407 333 415 341
rect 261 307 415 333
rect 449 333 457 341
rect 595 341 645 375
rect 689 485 739 527
rect 689 451 697 485
rect 731 451 739 485
rect 689 417 739 451
rect 689 383 697 417
rect 731 383 739 417
rect 689 367 739 383
rect 783 477 1585 493
rect 783 443 791 477
rect 825 459 979 477
rect 825 443 833 459
rect 783 409 833 443
rect 971 443 979 459
rect 1013 459 1167 477
rect 1013 443 1021 459
rect 783 375 791 409
rect 825 375 833 409
rect 595 333 603 341
rect 449 307 603 333
rect 637 333 645 341
rect 783 341 833 375
rect 783 333 791 341
rect 637 307 791 333
rect 825 307 833 341
rect 18 291 833 307
rect 877 409 927 425
rect 877 375 885 409
rect 919 375 927 409
rect 877 341 927 375
rect 971 409 1021 443
rect 1159 443 1167 459
rect 1201 459 1355 477
rect 1201 443 1209 459
rect 971 375 979 409
rect 1013 375 1021 409
rect 971 357 1021 375
rect 1065 409 1115 425
rect 1065 375 1073 409
rect 1107 375 1115 409
rect 877 307 885 341
rect 919 323 927 341
rect 1065 341 1115 375
rect 1159 409 1209 443
rect 1347 443 1355 459
rect 1389 459 1543 477
rect 1389 443 1397 459
rect 1159 375 1167 409
rect 1201 375 1209 409
rect 1159 357 1209 375
rect 1253 409 1303 425
rect 1253 375 1261 409
rect 1295 375 1303 409
rect 1065 323 1073 341
rect 919 307 1073 323
rect 1107 323 1115 341
rect 1253 341 1303 375
rect 1347 409 1397 443
rect 1535 443 1543 459
rect 1577 443 1585 477
rect 1347 375 1355 409
rect 1389 375 1397 409
rect 1347 357 1397 375
rect 1441 409 1491 425
rect 1441 375 1449 409
rect 1483 375 1491 409
rect 1253 323 1261 341
rect 1107 307 1261 323
rect 1295 323 1303 341
rect 1441 341 1491 375
rect 1535 409 1585 443
rect 1535 375 1543 409
rect 1577 375 1585 409
rect 1535 357 1585 375
rect 1441 323 1449 341
rect 1295 307 1449 323
rect 1483 323 1491 341
rect 1483 307 1605 323
rect 877 289 1605 307
rect 72 249 786 255
rect 72 215 103 249
rect 137 215 181 249
rect 215 215 259 249
rect 293 215 337 249
rect 371 215 415 249
rect 449 215 483 249
rect 517 215 561 249
rect 595 215 639 249
rect 673 215 717 249
rect 751 215 786 249
rect 840 249 1458 255
rect 840 215 858 249
rect 892 215 936 249
rect 970 215 1014 249
rect 1048 215 1092 249
rect 1126 215 1170 249
rect 1204 215 1238 249
rect 1272 215 1316 249
rect 1350 215 1394 249
rect 1428 215 1458 249
rect 1492 181 1605 289
rect 18 163 73 181
rect 18 129 39 163
rect 18 95 73 129
rect 18 61 39 95
rect 18 17 73 61
rect 107 163 1605 181
rect 107 129 133 163
rect 167 145 321 163
rect 167 129 183 145
rect 107 95 183 129
rect 295 129 321 145
rect 355 145 509 163
rect 355 129 371 145
rect 107 61 133 95
rect 167 61 183 95
rect 107 51 183 61
rect 227 95 261 111
rect 227 17 261 61
rect 295 95 371 129
rect 483 129 509 145
rect 543 145 697 163
rect 543 129 559 145
rect 295 61 321 95
rect 355 61 371 95
rect 295 51 371 61
rect 415 95 449 111
rect 415 17 449 61
rect 483 95 559 129
rect 671 129 697 145
rect 731 145 885 163
rect 731 129 747 145
rect 483 61 509 95
rect 543 61 559 95
rect 483 51 559 61
rect 603 95 637 111
rect 603 17 637 61
rect 671 95 747 129
rect 859 129 885 145
rect 919 145 1073 163
rect 919 129 935 145
rect 671 61 697 95
rect 731 61 747 95
rect 671 51 747 61
rect 791 95 825 111
rect 791 17 825 61
rect 859 95 935 129
rect 1047 129 1073 145
rect 1107 145 1261 163
rect 1107 129 1123 145
rect 859 61 885 95
rect 919 61 935 95
rect 859 51 935 61
rect 979 95 1013 111
rect 979 17 1013 61
rect 1047 95 1123 129
rect 1235 129 1261 145
rect 1295 145 1449 163
rect 1295 129 1311 145
rect 1047 61 1073 95
rect 1107 61 1123 95
rect 1047 51 1123 61
rect 1167 95 1201 111
rect 1167 17 1201 61
rect 1235 95 1311 129
rect 1423 129 1449 145
rect 1483 145 1605 163
rect 1483 129 1499 145
rect 1235 61 1261 95
rect 1295 61 1311 95
rect 1235 51 1311 61
rect 1355 95 1389 111
rect 1355 17 1389 61
rect 1423 95 1499 129
rect 1423 61 1449 95
rect 1483 61 1499 95
rect 1423 51 1499 61
rect 1543 95 1601 111
rect 1577 61 1601 95
rect 1543 17 1601 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
<< metal1 >>
rect 0 561 1656 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 0 496 1656 527
rect 0 17 1656 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
rect 0 -48 1656 -17
<< labels >>
flabel corelocali s 1500 289 1534 323 0 FreeSans 400 0 0 0 Y
port 7 nsew
flabel corelocali s 131 221 165 255 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 1049 221 1083 255 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew
rlabel comment s 0 0 0 0 4 nor2_8
<< properties >>
string FIXED_BBOX 0 0 1656 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2410014
string GDS_START 2397816
<< end >>
