magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 308 401 384 493
rect 308 367 483 401
rect 25 153 69 265
rect 183 153 275 265
rect 387 165 483 367
rect 334 131 483 165
rect 334 77 368 131
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 31 333 103 368
rect 240 367 274 527
rect 428 435 462 527
rect 31 299 353 333
rect 103 119 149 299
rect 309 199 353 299
rect 21 17 69 119
rect 103 51 171 119
rect 227 17 290 119
rect 402 17 478 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
rlabel locali s 183 153 275 265 6 A
port 1 nsew signal input
rlabel locali s 25 153 69 265 6 B
port 2 nsew signal input
rlabel locali s 387 165 483 367 6 X
port 3 nsew signal output
rlabel locali s 334 131 483 165 6 X
port 3 nsew signal output
rlabel locali s 334 77 368 131 6 X
port 3 nsew signal output
rlabel locali s 308 401 384 493 6 X
port 3 nsew signal output
rlabel locali s 308 367 483 401 6 X
port 3 nsew signal output
rlabel metal1 s 0 -48 552 48 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 496 552 592 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 552 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 617370
string GDS_START 612600
<< end >>
