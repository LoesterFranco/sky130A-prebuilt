magic
tech sky130A
magscale 1 2
timestamp 1599588232
<< locali >>
rect 85 222 161 356
rect 303 264 369 356
rect 880 236 946 302
rect 985 236 1056 349
rect 1266 236 1332 310
rect 2895 70 2963 596
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3072 683
rect 17 492 87 596
rect 189 526 239 649
rect 273 581 443 615
rect 273 492 307 581
rect 17 458 307 492
rect 17 162 51 458
rect 341 424 375 547
rect 409 492 443 581
rect 477 526 527 649
rect 629 492 679 595
rect 409 458 679 492
rect 195 390 477 424
rect 195 230 261 390
rect 411 304 477 390
rect 511 350 611 367
rect 545 316 611 350
rect 511 301 611 316
rect 645 267 679 458
rect 578 233 679 267
rect 713 581 942 615
rect 713 459 769 581
rect 195 199 362 230
rect 195 196 378 199
rect 17 96 118 162
rect 216 17 282 162
rect 328 107 378 196
rect 414 17 480 199
rect 578 107 644 233
rect 713 199 747 459
rect 803 451 874 547
rect 908 485 942 581
rect 976 519 1026 649
rect 1128 500 1198 587
rect 1232 534 1298 649
rect 1502 534 1568 649
rect 1602 546 1763 596
rect 1602 500 1636 546
rect 1797 512 1863 596
rect 1973 546 2039 649
rect 2181 546 2247 649
rect 1128 485 1636 500
rect 908 466 1636 485
rect 1767 478 1863 512
rect 1897 478 2440 512
rect 908 451 1232 466
rect 803 417 837 451
rect 678 107 747 199
rect 781 383 1164 417
rect 781 202 837 383
rect 1098 283 1164 383
rect 1198 249 1232 451
rect 1322 366 1478 432
rect 1322 352 1400 366
rect 1093 215 1232 249
rect 781 121 915 202
rect 781 51 837 121
rect 951 17 1001 202
rect 1093 121 1159 215
rect 1366 202 1400 352
rect 1524 330 1558 466
rect 1681 432 1733 467
rect 1592 398 1733 432
rect 1592 364 1715 398
rect 1524 296 1647 330
rect 1204 17 1256 181
rect 1290 168 1400 202
rect 1290 70 1356 168
rect 1401 17 1467 134
rect 1503 85 1553 226
rect 1597 119 1647 296
rect 1681 85 1715 364
rect 1767 358 1801 478
rect 1897 444 1931 478
rect 1835 392 1931 444
rect 2077 394 2161 444
rect 2027 358 2093 359
rect 1749 324 2093 358
rect 1749 119 1783 324
rect 2027 307 2093 324
rect 2127 305 2161 394
rect 1913 273 1979 290
rect 2127 273 2277 305
rect 1817 204 1868 269
rect 1913 239 2277 273
rect 2312 256 2372 360
rect 2406 347 2440 478
rect 2474 388 2561 596
rect 2666 530 2757 649
rect 2791 476 2857 596
rect 2613 415 2857 476
rect 2527 381 2561 388
rect 2527 347 2757 381
rect 2406 290 2493 347
rect 2535 256 2601 311
rect 1913 238 1979 239
rect 1817 170 2068 204
rect 1817 85 1851 170
rect 1503 51 1851 85
rect 1950 17 2000 136
rect 2034 85 2068 170
rect 2102 119 2136 239
rect 2312 222 2601 256
rect 2312 205 2346 222
rect 2170 171 2346 205
rect 2635 188 2669 347
rect 2723 276 2757 347
rect 2809 350 2857 415
rect 2809 316 2815 350
rect 2849 316 2857 350
rect 2809 310 2857 316
rect 2723 210 2789 276
rect 2170 85 2204 171
rect 2380 154 2669 188
rect 2823 162 2857 310
rect 2034 51 2204 85
rect 2238 17 2288 137
rect 2380 70 2446 154
rect 2560 17 2751 120
rect 2785 70 2857 162
rect 3001 364 3051 649
rect 2999 17 3049 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3072 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 511 316 545 350
rect 2815 316 2849 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
<< metal1 >>
rect 0 683 3072 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3072 683
rect 0 617 3072 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 3072 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3072 17
rect 0 -49 3072 -17
<< obsm1 >>
rect 499 350 557 356
rect 499 316 511 350
rect 545 347 557 350
rect 2803 350 2861 356
rect 2803 347 2815 350
rect 545 319 2815 347
rect 545 316 557 319
rect 499 310 557 316
rect 2803 316 2815 319
rect 2849 316 2861 350
rect 2803 310 2861 316
<< labels >>
rlabel locali s 85 222 161 356 6 D
port 1 nsew signal input
rlabel locali s 303 264 369 356 6 DE
port 2 nsew signal input
rlabel locali s 2895 70 2963 596 6 Q
port 3 nsew signal output
rlabel locali s 985 236 1056 349 6 SCD
port 4 nsew signal input
rlabel locali s 880 236 946 302 6 SCE
port 5 nsew signal input
rlabel locali s 1266 236 1332 310 6 CLK
port 6 nsew clock input
rlabel metal1 s 0 -49 3072 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 8 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 9 nsew power bidirectional
rlabel metal1 s 0 617 3072 715 6 VPWR
port 10 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 3072 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 414626
string GDS_START 392362
<< end >>
