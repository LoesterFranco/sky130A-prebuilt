magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 1602 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 89 47 119 177
rect 183 47 213 177
rect 277 47 307 177
rect 361 47 391 177
rect 465 47 495 177
rect 559 47 589 177
rect 757 47 787 177
rect 841 47 871 177
rect 945 47 975 177
rect 1039 47 1069 177
rect 1123 47 1153 177
rect 1217 47 1247 177
rect 1311 47 1341 177
rect 1415 47 1445 177
<< pmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 457 297 493 497
rect 551 297 587 497
rect 749 297 785 497
rect 843 297 879 497
rect 937 297 973 497
rect 1031 297 1067 497
rect 1125 297 1161 497
rect 1219 297 1255 497
rect 1313 297 1349 497
rect 1407 297 1443 497
<< ndiff >>
rect 27 163 89 177
rect 27 129 35 163
rect 69 129 89 163
rect 27 95 89 129
rect 27 61 35 95
rect 69 61 89 95
rect 27 47 89 61
rect 119 163 183 177
rect 119 129 129 163
rect 163 129 183 163
rect 119 47 183 129
rect 213 163 277 177
rect 213 129 223 163
rect 257 129 277 163
rect 213 95 277 129
rect 213 61 223 95
rect 257 61 277 95
rect 213 47 277 61
rect 307 163 361 177
rect 307 129 317 163
rect 351 129 361 163
rect 307 47 361 129
rect 391 95 465 177
rect 391 61 411 95
rect 445 61 465 95
rect 391 47 465 61
rect 495 163 559 177
rect 495 129 505 163
rect 539 129 559 163
rect 495 47 559 129
rect 589 93 641 177
rect 589 59 599 93
rect 633 59 641 93
rect 589 47 641 59
rect 695 93 757 177
rect 695 59 703 93
rect 737 59 757 93
rect 695 47 757 59
rect 787 169 841 177
rect 787 135 797 169
rect 831 135 841 169
rect 787 101 841 135
rect 787 67 797 101
rect 831 67 841 101
rect 787 47 841 67
rect 871 95 945 177
rect 871 61 891 95
rect 925 61 945 95
rect 871 47 945 61
rect 975 163 1039 177
rect 975 129 985 163
rect 1019 129 1039 163
rect 975 95 1039 129
rect 975 61 985 95
rect 1019 61 1039 95
rect 975 47 1039 61
rect 1069 163 1123 177
rect 1069 129 1079 163
rect 1113 129 1123 163
rect 1069 95 1123 129
rect 1069 61 1079 95
rect 1113 61 1123 95
rect 1069 47 1123 61
rect 1153 163 1217 177
rect 1153 129 1173 163
rect 1207 129 1217 163
rect 1153 95 1217 129
rect 1153 61 1173 95
rect 1207 61 1217 95
rect 1153 47 1217 61
rect 1247 95 1311 177
rect 1247 61 1267 95
rect 1301 61 1311 95
rect 1247 47 1311 61
rect 1341 163 1415 177
rect 1341 129 1361 163
rect 1395 129 1415 163
rect 1341 95 1415 129
rect 1341 61 1361 95
rect 1395 61 1415 95
rect 1341 47 1415 61
rect 1445 95 1497 177
rect 1445 61 1455 95
rect 1489 61 1497 95
rect 1445 47 1497 61
<< pdiff >>
rect 27 483 81 497
rect 27 449 35 483
rect 69 449 81 483
rect 27 415 81 449
rect 27 381 35 415
rect 69 381 81 415
rect 27 347 81 381
rect 27 313 35 347
rect 69 313 81 347
rect 27 297 81 313
rect 117 477 175 497
rect 117 443 129 477
rect 163 443 175 477
rect 117 409 175 443
rect 117 375 129 409
rect 163 375 175 409
rect 117 341 175 375
rect 117 307 129 341
rect 163 307 175 341
rect 117 297 175 307
rect 211 477 269 497
rect 211 443 223 477
rect 257 443 269 477
rect 211 297 269 443
rect 305 477 363 497
rect 305 443 317 477
rect 351 443 363 477
rect 305 297 363 443
rect 399 391 457 497
rect 399 357 411 391
rect 445 357 457 391
rect 399 297 457 357
rect 493 477 551 497
rect 493 443 505 477
rect 539 443 551 477
rect 493 297 551 443
rect 587 477 749 497
rect 587 443 601 477
rect 635 443 703 477
rect 737 443 749 477
rect 587 297 749 443
rect 785 477 843 497
rect 785 443 797 477
rect 831 443 843 477
rect 785 297 843 443
rect 879 391 937 497
rect 879 357 891 391
rect 925 357 937 391
rect 879 297 937 357
rect 973 477 1031 497
rect 973 443 985 477
rect 1019 443 1031 477
rect 973 297 1031 443
rect 1067 477 1125 497
rect 1067 443 1079 477
rect 1113 443 1125 477
rect 1067 297 1125 443
rect 1161 477 1219 497
rect 1161 443 1173 477
rect 1207 443 1219 477
rect 1161 409 1219 443
rect 1161 375 1173 409
rect 1207 375 1219 409
rect 1161 297 1219 375
rect 1255 477 1313 497
rect 1255 443 1267 477
rect 1301 443 1313 477
rect 1255 297 1313 443
rect 1349 477 1407 497
rect 1349 443 1361 477
rect 1395 443 1407 477
rect 1349 409 1407 443
rect 1349 375 1361 409
rect 1395 375 1407 409
rect 1349 341 1407 375
rect 1349 307 1361 341
rect 1395 307 1407 341
rect 1349 297 1407 307
rect 1443 477 1497 497
rect 1443 443 1455 477
rect 1489 443 1497 477
rect 1443 409 1497 443
rect 1443 375 1455 409
rect 1489 375 1497 409
rect 1443 297 1497 375
<< ndiffc >>
rect 35 129 69 163
rect 35 61 69 95
rect 129 129 163 163
rect 223 129 257 163
rect 223 61 257 95
rect 317 129 351 163
rect 411 61 445 95
rect 505 129 539 163
rect 599 59 633 93
rect 703 59 737 93
rect 797 135 831 169
rect 797 67 831 101
rect 891 61 925 95
rect 985 129 1019 163
rect 985 61 1019 95
rect 1079 129 1113 163
rect 1079 61 1113 95
rect 1173 129 1207 163
rect 1173 61 1207 95
rect 1267 61 1301 95
rect 1361 129 1395 163
rect 1361 61 1395 95
rect 1455 61 1489 95
<< pdiffc >>
rect 35 449 69 483
rect 35 381 69 415
rect 35 313 69 347
rect 129 443 163 477
rect 129 375 163 409
rect 129 307 163 341
rect 223 443 257 477
rect 317 443 351 477
rect 411 357 445 391
rect 505 443 539 477
rect 601 443 635 477
rect 703 443 737 477
rect 797 443 831 477
rect 891 357 925 391
rect 985 443 1019 477
rect 1079 443 1113 477
rect 1173 443 1207 477
rect 1173 375 1207 409
rect 1267 443 1301 477
rect 1361 443 1395 477
rect 1361 375 1395 409
rect 1361 307 1395 341
rect 1455 443 1489 477
rect 1455 375 1489 409
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 457 497 493 523
rect 551 497 587 523
rect 749 497 785 523
rect 843 497 879 523
rect 937 497 973 523
rect 1031 497 1067 523
rect 1125 497 1161 523
rect 1219 497 1255 523
rect 1313 497 1349 523
rect 1407 497 1443 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 457 282 493 297
rect 551 282 587 297
rect 749 282 785 297
rect 843 282 879 297
rect 937 282 973 297
rect 1031 282 1067 297
rect 1125 282 1161 297
rect 1219 282 1255 297
rect 1313 282 1349 297
rect 1407 282 1443 297
rect 79 265 119 282
rect 173 265 213 282
rect 267 265 307 282
rect 361 265 401 282
rect 455 265 495 282
rect 549 265 589 282
rect 747 265 787 282
rect 22 249 213 265
rect 22 215 38 249
rect 72 215 213 249
rect 22 199 213 215
rect 255 249 319 265
rect 255 215 265 249
rect 299 215 319 249
rect 255 199 319 215
rect 361 249 495 265
rect 361 215 411 249
rect 445 215 495 249
rect 361 199 495 215
rect 539 249 603 265
rect 539 215 549 249
rect 583 215 603 249
rect 539 199 603 215
rect 721 249 787 265
rect 721 215 731 249
rect 765 215 787 249
rect 721 199 787 215
rect 89 177 119 199
rect 183 177 213 199
rect 277 177 307 199
rect 361 177 391 199
rect 465 177 495 199
rect 559 177 589 199
rect 757 177 787 199
rect 841 265 881 282
rect 935 265 975 282
rect 1029 265 1069 282
rect 1123 265 1163 282
rect 1217 265 1257 282
rect 1311 265 1351 282
rect 1405 265 1445 282
rect 841 249 975 265
rect 841 215 891 249
rect 925 215 975 249
rect 841 199 975 215
rect 1017 249 1081 265
rect 1017 215 1027 249
rect 1061 215 1081 249
rect 1017 199 1081 215
rect 1123 249 1445 265
rect 1123 215 1173 249
rect 1207 215 1261 249
rect 1295 215 1361 249
rect 1395 215 1445 249
rect 1123 199 1445 215
rect 841 177 871 199
rect 945 177 975 199
rect 1039 177 1069 199
rect 1123 177 1153 199
rect 1217 177 1247 199
rect 1311 177 1341 199
rect 1415 177 1445 199
rect 89 21 119 47
rect 183 21 213 47
rect 277 21 307 47
rect 361 21 391 47
rect 465 21 495 47
rect 559 21 589 47
rect 757 21 787 47
rect 841 21 871 47
rect 945 21 975 47
rect 1039 21 1069 47
rect 1123 21 1153 47
rect 1217 21 1247 47
rect 1311 21 1341 47
rect 1415 21 1445 47
<< polycont >>
rect 38 215 72 249
rect 265 215 299 249
rect 411 215 445 249
rect 549 215 583 249
rect 731 215 765 249
rect 891 215 925 249
rect 1027 215 1061 249
rect 1173 215 1207 249
rect 1261 215 1295 249
rect 1361 215 1395 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 29 483 79 527
rect 29 449 35 483
rect 69 449 79 483
rect 29 415 79 449
rect 29 381 35 415
rect 69 381 79 415
rect 29 347 79 381
rect 29 313 35 347
rect 69 313 79 347
rect 29 291 79 313
rect 123 477 173 493
rect 123 443 129 477
rect 163 443 173 477
rect 123 409 173 443
rect 217 477 267 527
rect 217 443 223 477
rect 257 443 267 477
rect 217 425 267 443
rect 311 477 549 493
rect 311 443 317 477
rect 351 459 505 477
rect 351 443 361 459
rect 311 425 361 443
rect 499 443 505 459
rect 539 443 549 477
rect 499 425 549 443
rect 593 477 745 527
rect 593 443 601 477
rect 635 443 703 477
rect 737 443 745 477
rect 593 425 745 443
rect 789 477 1027 493
rect 789 443 797 477
rect 831 459 985 477
rect 831 443 839 459
rect 789 425 839 443
rect 977 443 985 459
rect 1019 443 1027 477
rect 977 425 1027 443
rect 1071 477 1121 527
rect 1071 443 1079 477
rect 1113 443 1121 477
rect 1071 425 1121 443
rect 1173 477 1215 493
rect 1207 443 1215 477
rect 123 375 129 409
rect 163 391 173 409
rect 1173 409 1215 443
rect 1259 477 1309 527
rect 1259 443 1267 477
rect 1301 443 1309 477
rect 1259 425 1309 443
rect 1353 477 1403 493
rect 1353 443 1361 477
rect 1395 443 1403 477
rect 163 375 411 391
rect 123 357 411 375
rect 445 357 891 391
rect 925 357 1129 391
rect 1207 391 1215 409
rect 1353 409 1403 443
rect 1207 375 1300 391
rect 1173 357 1300 375
rect 123 341 179 357
rect 123 307 129 341
rect 163 307 179 341
rect 1095 323 1129 357
rect 1266 323 1300 357
rect 1353 375 1361 409
rect 1395 375 1403 409
rect 1353 341 1403 375
rect 1447 477 1497 527
rect 1447 443 1455 477
rect 1489 443 1497 477
rect 1447 409 1497 443
rect 1447 375 1455 409
rect 1489 375 1497 409
rect 1447 359 1497 375
rect 1353 323 1361 341
rect 18 249 88 255
rect 18 215 38 249
rect 72 215 88 249
rect 17 163 69 179
rect 123 173 179 307
rect 213 289 609 323
rect 213 249 346 289
rect 213 215 265 249
rect 299 215 346 249
rect 390 249 499 255
rect 390 215 411 249
rect 445 215 499 249
rect 533 249 609 289
rect 533 215 549 249
rect 583 215 609 249
rect 661 289 1045 323
rect 1095 289 1185 323
rect 1266 307 1361 323
rect 1395 323 1403 341
rect 1395 307 1542 323
rect 1266 289 1542 307
rect 661 249 791 289
rect 995 255 1045 289
rect 1141 255 1185 289
rect 661 215 731 249
rect 765 215 791 249
rect 825 249 951 255
rect 825 215 891 249
rect 925 215 951 249
rect 995 249 1107 255
rect 995 215 1027 249
rect 1061 215 1107 249
rect 1141 249 1411 255
rect 1141 215 1173 249
rect 1207 215 1261 249
rect 1295 215 1361 249
rect 1395 215 1411 249
rect 1473 181 1542 289
rect 17 129 35 163
rect 103 163 179 173
rect 103 129 129 163
rect 163 129 179 163
rect 223 163 257 181
rect 291 169 1035 181
rect 291 163 797 169
rect 291 129 317 163
rect 351 129 505 163
rect 539 135 797 163
rect 831 163 1035 169
rect 831 145 985 163
rect 831 135 847 145
rect 539 129 847 135
rect 17 95 69 129
rect 223 95 257 129
rect 797 101 847 129
rect 959 129 985 145
rect 1019 129 1035 163
rect 17 61 35 95
rect 69 61 223 95
rect 257 61 411 95
rect 445 93 651 95
rect 445 61 599 93
rect 17 59 599 61
rect 633 59 651 93
rect 17 51 651 59
rect 687 59 703 93
rect 737 59 753 93
rect 687 17 753 59
rect 831 67 847 101
rect 797 51 847 67
rect 891 95 925 111
rect 891 17 925 61
rect 959 95 1035 129
rect 959 61 985 95
rect 1019 61 1035 95
rect 959 51 1035 61
rect 1079 163 1113 181
rect 1079 95 1113 129
rect 1079 17 1113 61
rect 1147 163 1542 181
rect 1147 129 1173 163
rect 1207 145 1361 163
rect 1207 129 1223 145
rect 1147 95 1223 129
rect 1335 129 1361 145
rect 1395 147 1542 163
rect 1395 129 1411 147
rect 1147 61 1173 95
rect 1207 61 1223 95
rect 1147 51 1223 61
rect 1267 95 1301 111
rect 1267 17 1301 61
rect 1335 95 1411 129
rect 1335 61 1361 95
rect 1395 61 1411 95
rect 1335 51 1411 61
rect 1455 95 1506 113
rect 1489 61 1506 95
rect 1455 17 1506 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
<< metal1 >>
rect 0 561 1564 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 0 496 1564 527
rect 0 17 1564 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
rect 0 -48 1564 -17
<< labels >>
flabel corelocali s 30 221 64 255 0 FreeSans 400 0 0 0 C1
port 5 nsew
flabel corelocali s 1042 221 1076 255 0 FreeSans 400 180 0 0 A1
port 1 nsew
flabel corelocali s 848 221 882 255 0 FreeSans 400 180 0 0 A2
port 2 nsew
flabel corelocali s 292 238 292 238 0 FreeSans 400 0 0 0 B1
port 3 nsew
flabel corelocali s 415 238 415 238 0 FreeSans 400 0 0 0 B2
port 4 nsew
flabel corelocali s 1478 289 1512 323 0 FreeSans 400 0 0 0 X
port 10 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew
rlabel comment s 0 0 0 0 4 o221a_4
<< properties >>
string FIXED_BBOX 0 0 1564 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 847230
string GDS_START 835908
<< end >>
