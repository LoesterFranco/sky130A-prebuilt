magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1196 561
rect 108 439 153 527
rect 17 214 66 323
rect 122 268 178 323
rect 112 234 178 268
rect 122 214 178 234
rect 349 299 383 527
rect 417 333 467 493
rect 501 367 551 527
rect 585 333 651 493
rect 685 367 823 527
rect 857 333 923 493
rect 957 367 991 527
rect 1025 333 1091 493
rect 417 289 1091 333
rect 1125 289 1179 527
rect 417 131 483 289
rect 649 215 710 289
rect 744 215 923 255
rect 989 215 1175 255
rect 103 17 153 109
rect 1041 17 1075 113
rect 0 -17 1196 17
<< obsli1 >>
rect 17 396 74 488
rect 187 430 315 493
rect 17 357 246 396
rect 212 255 246 357
rect 212 180 246 221
rect 17 146 246 180
rect 280 282 315 430
rect 17 51 69 146
rect 280 143 316 282
rect 280 112 315 143
rect 549 221 581 255
rect 549 215 615 221
rect 585 131 923 181
rect 957 147 1179 181
rect 187 51 315 112
rect 349 97 383 117
rect 957 97 1007 147
rect 349 51 735 97
rect 773 51 1007 97
rect 1109 51 1179 147
<< obsli1c >>
rect 212 221 246 255
rect 581 221 615 255
<< metal1 >>
rect 0 496 1196 592
rect 0 -48 1196 48
<< obsm1 >>
rect 200 255 627 261
rect 200 221 212 255
rect 246 221 581 255
rect 615 221 627 255
rect 200 215 627 221
<< labels >>
rlabel locali s 122 268 178 323 6 A_N
port 1 nsew signal input
rlabel locali s 122 214 178 234 6 A_N
port 1 nsew signal input
rlabel locali s 112 234 178 268 6 A_N
port 1 nsew signal input
rlabel locali s 17 214 66 323 6 B_N
port 2 nsew signal input
rlabel locali s 744 215 923 255 6 C
port 3 nsew signal input
rlabel locali s 989 215 1175 255 6 D
port 4 nsew signal input
rlabel locali s 1025 333 1091 493 6 Y
port 5 nsew signal output
rlabel locali s 857 333 923 493 6 Y
port 5 nsew signal output
rlabel locali s 649 215 710 289 6 Y
port 5 nsew signal output
rlabel locali s 585 333 651 493 6 Y
port 5 nsew signal output
rlabel locali s 417 333 467 493 6 Y
port 5 nsew signal output
rlabel locali s 417 289 1091 333 6 Y
port 5 nsew signal output
rlabel locali s 417 131 483 289 6 Y
port 5 nsew signal output
rlabel locali s 1041 17 1075 113 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 103 17 153 109 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 1196 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1196 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1125 289 1179 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 957 367 991 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 685 367 823 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 501 367 551 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 349 299 383 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 108 439 153 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 1196 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 1196 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1912254
string GDS_START 1901866
<< end >>
