magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 920 561
rect 103 441 169 527
rect 86 199 156 339
rect 190 199 248 265
rect 501 425 629 491
rect 663 367 719 527
rect 761 299 816 493
rect 528 199 659 265
rect 132 17 166 165
rect 782 152 816 299
rect 850 288 884 527
rect 299 17 370 97
rect 479 17 545 97
rect 647 17 723 97
rect 761 83 816 152
rect 850 17 884 205
rect 0 -17 920 17
<< obsli1 >>
rect 17 407 69 491
rect 307 441 456 475
rect 17 373 388 407
rect 17 165 52 373
rect 199 305 320 339
rect 282 249 320 305
rect 354 317 388 373
rect 422 391 456 441
rect 422 357 629 391
rect 595 333 629 357
rect 354 283 484 317
rect 595 299 727 333
rect 282 215 371 249
rect 282 165 320 215
rect 450 199 484 283
rect 693 265 727 299
rect 693 199 748 265
rect 693 165 727 199
rect 17 90 81 165
rect 216 131 320 165
rect 405 131 727 165
rect 216 90 250 131
rect 405 61 439 131
rect 579 61 613 131
<< metal1 >>
rect 0 496 920 592
rect 0 -48 920 48
<< labels >>
rlabel locali s 528 199 659 265 6 A
port 1 nsew signal input
rlabel locali s 501 425 629 491 6 B
port 2 nsew signal input
rlabel locali s 86 199 156 339 6 C_N
port 3 nsew signal input
rlabel locali s 190 199 248 265 6 D_N
port 4 nsew signal input
rlabel locali s 782 152 816 299 6 X
port 5 nsew signal output
rlabel locali s 761 299 816 493 6 X
port 5 nsew signal output
rlabel locali s 761 83 816 152 6 X
port 5 nsew signal output
rlabel locali s 850 17 884 205 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 647 17 723 97 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 479 17 545 97 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 299 17 370 97 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 132 17 166 165 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 920 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 920 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 850 288 884 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 663 367 719 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 103 441 169 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 920 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 920 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 920 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1120050
string GDS_START 1112442
<< end >>
