magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 89 53 119 137
rect 279 47 309 177
rect 363 47 393 177
rect 471 47 501 177
rect 565 47 595 177
rect 659 47 689 177
rect 763 47 793 177
<< pmoshvt >>
rect 81 413 117 497
rect 283 297 319 497
rect 365 297 401 497
rect 473 297 509 497
rect 567 297 603 497
rect 661 297 697 497
rect 755 297 791 497
<< ndiff >>
rect 192 137 279 177
rect 27 106 89 137
rect 27 72 35 106
rect 69 72 89 106
rect 27 53 89 72
rect 119 97 279 137
rect 119 63 129 97
rect 163 63 225 97
rect 259 63 279 97
rect 119 53 279 63
rect 192 47 279 53
rect 309 165 363 177
rect 309 131 319 165
rect 353 131 363 165
rect 309 97 363 131
rect 309 63 319 97
rect 353 63 363 97
rect 309 47 363 63
rect 393 165 471 177
rect 393 131 427 165
rect 461 131 471 165
rect 393 97 471 131
rect 393 63 427 97
rect 461 63 471 97
rect 393 47 471 63
rect 501 165 565 177
rect 501 131 521 165
rect 555 131 565 165
rect 501 97 565 131
rect 501 63 521 97
rect 555 63 565 97
rect 501 47 565 63
rect 595 94 659 177
rect 595 60 615 94
rect 649 60 659 94
rect 595 47 659 60
rect 689 165 763 177
rect 689 131 709 165
rect 743 131 763 165
rect 689 97 763 131
rect 689 63 709 97
rect 743 63 763 97
rect 689 47 763 63
rect 793 94 859 177
rect 793 60 803 94
rect 837 60 859 94
rect 793 47 859 60
<< pdiff >>
rect 27 475 81 497
rect 27 441 35 475
rect 69 441 81 475
rect 27 413 81 441
rect 117 457 175 497
rect 117 423 129 457
rect 163 423 175 457
rect 117 413 175 423
rect 229 479 283 497
rect 229 445 237 479
rect 271 445 283 479
rect 229 411 283 445
rect 229 377 237 411
rect 271 377 283 411
rect 229 343 283 377
rect 229 309 237 343
rect 271 309 283 343
rect 229 297 283 309
rect 319 297 365 497
rect 401 485 473 497
rect 401 451 426 485
rect 460 451 473 485
rect 401 417 473 451
rect 401 383 426 417
rect 460 383 473 417
rect 401 297 473 383
rect 509 477 567 497
rect 509 443 521 477
rect 555 443 567 477
rect 509 409 567 443
rect 509 375 521 409
rect 555 375 567 409
rect 509 297 567 375
rect 603 477 661 497
rect 603 443 615 477
rect 649 443 661 477
rect 603 297 661 443
rect 697 477 755 497
rect 697 443 709 477
rect 743 443 755 477
rect 697 409 755 443
rect 697 375 709 409
rect 743 375 755 409
rect 697 341 755 375
rect 697 307 709 341
rect 743 307 755 341
rect 697 297 755 307
rect 791 477 852 497
rect 791 443 803 477
rect 837 443 852 477
rect 791 409 852 443
rect 791 375 803 409
rect 837 375 852 409
rect 791 297 852 375
<< ndiffc >>
rect 35 72 69 106
rect 129 63 163 97
rect 225 63 259 97
rect 319 131 353 165
rect 319 63 353 97
rect 427 131 461 165
rect 427 63 461 97
rect 521 131 555 165
rect 521 63 555 97
rect 615 60 649 94
rect 709 131 743 165
rect 709 63 743 97
rect 803 60 837 94
<< pdiffc >>
rect 35 441 69 475
rect 129 423 163 457
rect 237 445 271 479
rect 237 377 271 411
rect 237 309 271 343
rect 426 451 460 485
rect 426 383 460 417
rect 521 443 555 477
rect 521 375 555 409
rect 615 443 649 477
rect 709 443 743 477
rect 709 375 743 409
rect 709 307 743 341
rect 803 443 837 477
rect 803 375 837 409
<< poly >>
rect 81 497 117 523
rect 283 497 319 523
rect 365 497 401 523
rect 473 497 509 523
rect 567 497 603 523
rect 661 497 697 523
rect 755 497 791 523
rect 81 398 117 413
rect 79 265 119 398
rect 283 282 319 297
rect 365 282 401 297
rect 473 282 509 297
rect 567 282 603 297
rect 661 282 697 297
rect 755 282 791 297
rect 281 265 321 282
rect 22 249 119 265
rect 22 215 35 249
rect 69 215 119 249
rect 22 199 119 215
rect 184 249 321 265
rect 184 215 194 249
rect 228 215 321 249
rect 184 199 321 215
rect 363 265 403 282
rect 471 265 511 282
rect 565 265 605 282
rect 659 265 699 282
rect 753 265 793 282
rect 363 249 427 265
rect 363 215 373 249
rect 407 215 427 249
rect 363 199 427 215
rect 471 249 793 265
rect 471 215 554 249
rect 588 215 632 249
rect 666 215 710 249
rect 744 215 793 249
rect 471 199 793 215
rect 89 137 119 199
rect 279 177 309 199
rect 363 177 393 199
rect 471 177 501 199
rect 565 177 595 199
rect 659 177 689 199
rect 763 177 793 199
rect 89 27 119 53
rect 279 21 309 47
rect 363 21 393 47
rect 471 21 501 47
rect 565 21 595 47
rect 659 21 689 47
rect 763 21 793 47
<< polycont >>
rect 35 215 69 249
rect 194 215 228 249
rect 373 215 407 249
rect 554 215 588 249
rect 632 215 666 249
rect 710 215 744 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 18 475 69 527
rect 18 441 35 475
rect 18 425 69 441
rect 129 457 163 493
rect 18 249 85 391
rect 18 215 35 249
rect 69 215 85 249
rect 129 265 163 423
rect 208 479 312 493
rect 208 445 237 479
rect 271 445 312 479
rect 208 411 312 445
rect 208 377 237 411
rect 271 377 312 411
rect 208 343 312 377
rect 413 485 469 527
rect 413 451 426 485
rect 460 451 469 485
rect 413 417 469 451
rect 413 383 426 417
rect 460 383 469 417
rect 413 367 469 383
rect 513 477 563 493
rect 513 443 521 477
rect 555 443 563 477
rect 513 409 563 443
rect 607 477 657 527
rect 607 443 615 477
rect 649 443 657 477
rect 607 427 657 443
rect 701 477 751 493
rect 701 443 709 477
rect 743 443 751 477
rect 513 375 521 409
rect 555 391 563 409
rect 701 409 751 443
rect 701 391 709 409
rect 555 375 709 391
rect 743 375 751 409
rect 513 357 751 375
rect 795 477 845 527
rect 795 443 803 477
rect 837 443 845 477
rect 795 409 845 443
rect 795 375 803 409
rect 837 375 845 409
rect 795 359 845 375
rect 208 309 237 343
rect 271 323 312 343
rect 616 341 751 357
rect 271 309 572 323
rect 208 299 572 309
rect 268 289 572 299
rect 616 307 709 341
rect 743 323 751 341
rect 743 307 898 323
rect 616 289 898 307
rect 129 249 234 265
rect 129 215 194 249
rect 228 215 234 249
rect 129 199 234 215
rect 129 181 179 199
rect 22 147 179 181
rect 268 181 312 289
rect 346 249 494 255
rect 346 215 373 249
rect 407 215 494 249
rect 538 249 572 289
rect 538 215 554 249
rect 588 215 632 249
rect 666 215 710 249
rect 744 215 760 249
rect 821 181 898 289
rect 268 165 369 181
rect 268 147 319 165
rect 22 106 84 147
rect 293 131 319 147
rect 353 131 369 165
rect 22 72 35 106
rect 69 72 84 106
rect 22 53 84 72
rect 128 97 259 113
rect 128 63 129 97
rect 163 63 225 97
rect 128 17 259 63
rect 293 97 369 131
rect 293 63 319 97
rect 353 63 369 97
rect 293 61 369 63
rect 426 165 461 181
rect 426 131 427 165
rect 426 97 461 131
rect 426 63 427 97
rect 426 17 461 63
rect 495 165 898 181
rect 495 131 521 165
rect 555 147 709 165
rect 555 131 571 147
rect 495 97 571 131
rect 683 131 709 147
rect 743 147 898 165
rect 743 131 759 147
rect 495 63 521 97
rect 555 63 571 97
rect 495 58 571 63
rect 615 94 649 110
rect 615 17 649 60
rect 683 97 759 131
rect 683 63 709 97
rect 743 63 759 97
rect 683 58 759 63
rect 803 94 837 110
rect 803 17 837 60
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel corelocali s 414 238 414 238 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 29 221 63 255 0 FreeSans 400 0 0 0 B_N
port 2 nsew
flabel corelocali s 852 223 886 257 0 FreeSans 400 0 0 0 X
port 7 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew
rlabel comment s 0 0 0 0 4 or2b_4
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 661866
string GDS_START 654706
<< end >>
