magic
tech sky130A
magscale 1 2
timestamp 1599588238
<< locali >>
rect 217 291 331 357
rect 487 310 553 430
rect 85 191 439 257
rect 313 162 439 191
rect 655 236 737 310
rect 2137 394 2203 596
rect 2333 403 2371 596
rect 2333 394 2471 403
rect 2137 360 2471 394
rect 2352 226 2471 360
rect 2149 176 2471 226
rect 2149 70 2199 176
rect 2335 70 2373 176
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2496 683
rect 17 425 111 596
rect 145 460 211 649
rect 319 512 385 596
rect 517 546 641 649
rect 777 546 895 649
rect 1031 542 1081 594
rect 929 512 1081 542
rect 319 508 1081 512
rect 319 478 963 508
rect 1115 502 1187 594
rect 1336 571 1402 649
rect 1221 503 1620 537
rect 319 462 385 478
rect 373 425 439 428
rect 17 391 439 425
rect 17 305 183 391
rect 17 157 51 305
rect 373 294 439 391
rect 587 270 621 478
rect 665 398 731 444
rect 665 364 833 398
rect 473 236 621 270
rect 771 260 833 364
rect 867 330 901 478
rect 1015 444 1081 474
rect 935 408 1081 444
rect 935 364 985 408
rect 867 296 985 330
rect 17 70 98 157
rect 132 17 198 157
rect 473 128 507 236
rect 771 202 805 260
rect 625 168 805 202
rect 296 78 507 128
rect 541 17 591 162
rect 625 70 691 168
rect 737 17 803 134
rect 839 85 889 226
rect 935 119 985 296
rect 1019 85 1053 408
rect 1115 356 1149 502
rect 1221 456 1255 503
rect 1183 390 1255 456
rect 1443 435 1552 469
rect 1367 356 1432 388
rect 1087 322 1432 356
rect 1087 119 1121 322
rect 1466 288 1500 435
rect 1586 391 1620 503
rect 1654 438 1720 564
rect 1845 472 1911 649
rect 1654 404 1837 438
rect 1554 325 1620 391
rect 1803 360 1837 404
rect 1946 394 2027 564
rect 1155 188 1215 272
rect 1259 222 1500 288
rect 1707 282 1769 343
rect 1155 154 1432 188
rect 1155 85 1189 154
rect 839 51 1189 85
rect 1298 17 1364 120
rect 1398 93 1432 154
rect 1466 177 1500 222
rect 1534 248 1769 282
rect 1803 294 1959 360
rect 1993 326 2027 394
rect 2061 388 2095 649
rect 2243 428 2293 649
rect 2407 437 2473 649
rect 1534 211 1625 248
rect 1803 214 1837 294
rect 1993 260 2309 326
rect 1466 127 1557 177
rect 1591 93 1625 211
rect 1398 59 1625 93
rect 1659 180 1837 214
rect 1871 226 2027 260
rect 1871 180 1933 226
rect 1659 70 1725 180
rect 1839 17 1905 146
rect 1967 70 2001 226
rect 2037 17 2103 192
rect 2235 17 2301 142
rect 2407 17 2473 142
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2496 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
<< metal1 >>
rect 0 683 2496 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2496 683
rect 0 617 2496 649
rect 0 17 2496 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2496 17
rect 0 -49 2496 -17
<< labels >>
rlabel locali s 217 291 331 357 6 D
port 1 nsew signal input
rlabel locali s 2352 226 2471 360 6 Q
port 2 nsew signal output
rlabel locali s 2335 70 2373 176 6 Q
port 2 nsew signal output
rlabel locali s 2333 403 2371 596 6 Q
port 2 nsew signal output
rlabel locali s 2333 394 2471 403 6 Q
port 2 nsew signal output
rlabel locali s 2149 176 2471 226 6 Q
port 2 nsew signal output
rlabel locali s 2149 70 2199 176 6 Q
port 2 nsew signal output
rlabel locali s 2137 394 2203 596 6 Q
port 2 nsew signal output
rlabel locali s 2137 360 2471 394 6 Q
port 2 nsew signal output
rlabel locali s 487 310 553 430 6 SCD
port 3 nsew signal input
rlabel locali s 313 162 439 191 6 SCE
port 4 nsew signal input
rlabel locali s 85 191 439 257 6 SCE
port 4 nsew signal input
rlabel locali s 655 236 737 310 6 CLK
port 5 nsew clock input
rlabel metal1 s 0 -49 2496 49 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 617 2496 715 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2496 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 224356
string GDS_START 206894
<< end >>
