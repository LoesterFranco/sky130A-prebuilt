magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 644 561
rect 19 333 77 527
rect 111 165 157 493
rect 191 444 257 527
rect 471 425 537 527
rect 293 199 358 282
rect 111 127 191 165
rect 53 17 119 93
rect 153 51 191 127
rect 225 17 291 89
rect 448 73 524 265
rect 562 150 625 265
rect 561 17 627 113
rect 0 -17 644 17
<< obsli1 >>
rect 295 384 358 493
rect 191 338 358 384
rect 392 387 437 493
rect 571 387 615 493
rect 191 199 259 338
rect 392 334 615 387
rect 225 165 259 199
rect 225 131 373 165
rect 335 51 373 131
<< metal1 >>
rect 0 496 644 592
rect 0 -48 644 48
<< labels >>
rlabel locali s 448 73 524 265 6 A1
port 1 nsew signal input
rlabel locali s 562 150 625 265 6 A2
port 2 nsew signal input
rlabel locali s 293 199 358 282 6 B1
port 3 nsew signal input
rlabel locali s 153 51 191 127 6 X
port 4 nsew signal output
rlabel locali s 111 165 157 493 6 X
port 4 nsew signal output
rlabel locali s 111 127 191 165 6 X
port 4 nsew signal output
rlabel locali s 561 17 627 113 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 225 17 291 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 53 17 119 93 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 644 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 644 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 471 425 537 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 191 444 257 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 19 333 77 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 644 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 644 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 4034592
string GDS_START 4029038
<< end >>
