magic
tech sky130A
magscale 1 2
timestamp 1601050082
<< locali >>
rect 95 202 161 404
rect 263 236 359 310
rect 2024 236 2087 596
rect 2311 364 2377 596
rect 2024 226 2063 236
rect 1997 70 2063 226
rect 2343 210 2377 364
rect 2311 70 2377 210
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2400 683
rect 23 472 73 596
rect 113 518 179 649
rect 315 506 381 649
rect 421 581 775 615
rect 421 480 471 581
rect 23 446 359 472
rect 505 459 601 547
rect 635 459 707 547
rect 505 446 539 459
rect 23 438 539 446
rect 23 168 57 438
rect 325 412 539 438
rect 195 378 291 404
rect 195 344 471 378
rect 195 202 229 344
rect 405 260 471 344
rect 23 76 73 168
rect 109 17 159 168
rect 195 70 287 202
rect 321 17 373 202
rect 409 85 459 226
rect 505 169 539 412
rect 573 287 639 421
rect 505 119 571 169
rect 605 85 639 287
rect 409 51 639 85
rect 673 211 707 459
rect 741 467 775 581
rect 809 501 888 649
rect 922 581 1108 615
rect 922 467 956 581
rect 741 433 956 467
rect 741 272 789 433
rect 990 399 1040 547
rect 1074 459 1108 581
rect 1142 493 1210 649
rect 1352 530 1490 581
rect 1614 530 1648 649
rect 1352 496 1580 530
rect 1688 496 1754 596
rect 1074 425 1207 459
rect 846 355 1040 399
rect 1081 350 1139 391
rect 823 287 1047 321
rect 1081 316 1087 350
rect 1121 316 1139 350
rect 1173 358 1207 425
rect 1352 392 1402 496
rect 1446 404 1512 462
rect 1546 444 1754 496
rect 1800 512 1866 596
rect 1912 546 1982 649
rect 1800 478 1947 512
rect 1546 410 1879 444
rect 1368 370 1402 392
rect 1173 324 1321 358
rect 1368 336 1444 370
rect 1081 310 1139 316
rect 1287 290 1321 324
rect 823 211 857 287
rect 990 258 1047 287
rect 1187 258 1253 290
rect 673 177 857 211
rect 891 177 955 253
rect 990 224 1253 258
rect 1287 224 1376 290
rect 990 211 1047 224
rect 673 77 723 177
rect 821 17 887 143
rect 921 87 1036 177
rect 1171 17 1237 190
rect 1287 85 1321 224
rect 1410 185 1444 336
rect 1355 119 1444 185
rect 1478 85 1512 404
rect 1554 202 1620 376
rect 1657 350 1734 356
rect 1657 316 1663 350
rect 1697 316 1734 350
rect 1657 236 1734 316
rect 1813 242 1879 410
rect 1913 202 1947 478
rect 2136 310 2170 575
rect 2210 399 2276 649
rect 2136 244 2308 310
rect 1554 168 1947 202
rect 1287 51 1512 85
rect 1613 17 1751 134
rect 1785 83 1851 168
rect 1897 17 1963 134
rect 2136 188 2175 244
rect 2109 70 2175 188
rect 2211 17 2277 188
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2400 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 1087 316 1121 350
rect 1663 316 1697 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
<< metal1 >>
rect 0 683 2400 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2400 683
rect 0 617 2400 649
rect 1075 350 1133 356
rect 1075 316 1087 350
rect 1121 347 1133 350
rect 1651 350 1709 356
rect 1651 347 1663 350
rect 1121 319 1663 347
rect 1121 316 1133 319
rect 1075 310 1133 316
rect 1651 316 1663 319
rect 1697 316 1709 350
rect 1651 310 1709 316
rect 0 17 2400 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2400 17
rect 0 -49 2400 -17
<< labels >>
rlabel locali s 95 202 161 404 6 D
port 1 nsew signal input
rlabel locali s 2343 210 2377 364 6 Q
port 2 nsew signal output
rlabel locali s 2311 364 2377 596 6 Q
port 2 nsew signal output
rlabel locali s 2311 70 2377 210 6 Q
port 2 nsew signal output
rlabel locali s 2024 236 2087 596 6 Q_N
port 3 nsew signal output
rlabel locali s 2024 226 2063 236 6 Q_N
port 3 nsew signal output
rlabel locali s 1997 70 2063 226 6 Q_N
port 3 nsew signal output
rlabel metal1 s 1651 347 1709 356 6 SET_B
port 4 nsew signal input
rlabel metal1 s 1651 310 1709 319 6 SET_B
port 4 nsew signal input
rlabel metal1 s 1075 347 1133 356 6 SET_B
port 4 nsew signal input
rlabel metal1 s 1075 319 1709 347 6 SET_B
port 4 nsew signal input
rlabel metal1 s 1075 310 1133 319 6 SET_B
port 4 nsew signal input
rlabel locali s 263 236 359 310 6 CLK
port 5 nsew clock input
rlabel metal1 s 0 -49 2400 49 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 617 2400 715 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2400 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2787538
string GDS_START 2769364
<< end >>
