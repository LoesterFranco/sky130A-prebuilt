magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 644 561
rect 17 299 69 527
rect 117 425 440 491
rect 474 367 530 527
rect 305 265 354 323
rect 572 299 627 493
rect 18 215 85 265
rect 305 199 470 265
rect 17 17 69 181
rect 593 152 627 299
rect 291 17 357 97
rect 459 17 534 97
rect 572 83 627 152
rect 0 -17 644 17
<< obsli1 >>
rect 119 265 153 377
rect 205 357 440 391
rect 205 299 271 357
rect 406 333 440 357
rect 406 299 538 333
rect 504 265 538 299
rect 119 199 262 265
rect 504 199 559 265
rect 119 181 169 199
rect 103 97 169 181
rect 504 165 538 199
rect 205 131 538 165
rect 205 51 257 131
rect 391 61 425 131
<< metal1 >>
rect 0 496 644 592
rect 0 -48 644 48
<< labels >>
rlabel locali s 305 265 354 323 6 A
port 1 nsew signal input
rlabel locali s 305 199 470 265 6 A
port 1 nsew signal input
rlabel locali s 117 425 440 491 6 B
port 2 nsew signal input
rlabel locali s 18 215 85 265 6 C_N
port 3 nsew signal input
rlabel locali s 593 152 627 299 6 X
port 4 nsew signal output
rlabel locali s 572 299 627 493 6 X
port 4 nsew signal output
rlabel locali s 572 83 627 152 6 X
port 4 nsew signal output
rlabel locali s 459 17 534 97 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 291 17 357 97 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 17 17 69 181 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 644 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 644 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 474 367 530 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 17 299 69 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 644 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 644 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1050648
string GDS_START 1044442
<< end >>
