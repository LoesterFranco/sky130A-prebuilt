magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 19 211 183 265
rect 558 205 625 259
rect 663 205 730 259
rect 1105 211 1269 265
rect 1307 211 1471 265
rect 1846 205 1913 259
rect 1951 205 2018 259
rect 2393 211 2557 265
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2576 561
rect 19 442 85 493
rect 19 333 79 442
rect 119 421 179 527
rect 113 367 179 421
rect 223 459 456 493
rect 223 333 257 459
rect 293 391 379 425
rect 293 357 305 391
rect 339 357 379 391
rect 293 351 379 357
rect 19 299 257 333
rect 206 177 267 185
rect 317 177 351 351
rect 422 329 456 459
rect 510 327 576 493
rect 490 295 576 327
rect 420 293 576 295
rect 611 293 677 527
rect 712 327 778 493
rect 832 459 1065 493
rect 832 329 866 459
rect 909 391 995 425
rect 909 357 949 391
rect 983 357 995 391
rect 909 351 995 357
rect 712 295 798 327
rect 712 293 868 295
rect 420 261 524 293
rect 764 261 868 293
rect 420 241 503 261
rect 29 143 267 177
rect 29 51 95 143
rect 129 17 172 109
rect 206 85 267 143
rect 301 119 367 177
rect 401 85 435 154
rect 469 151 503 241
rect 785 241 868 261
rect 785 151 819 241
rect 937 177 971 351
rect 1031 333 1065 459
rect 1109 421 1169 527
rect 1203 442 1269 493
rect 1109 367 1175 421
rect 1209 333 1269 442
rect 1031 299 1269 333
rect 1307 442 1373 493
rect 1307 333 1367 442
rect 1407 421 1467 527
rect 1401 367 1467 421
rect 1511 459 1744 493
rect 1511 333 1545 459
rect 1581 391 1667 425
rect 1581 357 1593 391
rect 1627 357 1667 391
rect 1581 351 1667 357
rect 1307 299 1545 333
rect 1021 177 1082 185
rect 1494 177 1555 185
rect 1605 177 1639 351
rect 1710 329 1744 459
rect 1798 327 1864 493
rect 1778 295 1864 327
rect 1708 293 1864 295
rect 1899 293 1965 527
rect 2000 327 2066 493
rect 2120 459 2353 493
rect 2120 329 2154 459
rect 2197 391 2283 425
rect 2197 357 2237 391
rect 2271 357 2283 391
rect 2197 351 2283 357
rect 2000 295 2086 327
rect 2000 293 2156 295
rect 1708 261 1812 293
rect 2052 261 2156 293
rect 1708 241 1791 261
rect 469 117 585 151
rect 206 51 435 85
rect 535 66 585 117
rect 619 17 669 132
rect 703 117 819 151
rect 703 66 753 117
rect 853 85 887 154
rect 921 119 987 177
rect 1021 143 1259 177
rect 1021 85 1082 143
rect 853 51 1082 85
rect 1116 17 1159 109
rect 1193 51 1259 143
rect 1317 143 1555 177
rect 1317 51 1383 143
rect 1417 17 1460 109
rect 1494 85 1555 143
rect 1589 119 1655 177
rect 1689 85 1723 154
rect 1757 151 1791 241
rect 2073 241 2156 261
rect 2073 151 2107 241
rect 2225 177 2259 351
rect 2319 333 2353 459
rect 2397 421 2457 527
rect 2491 442 2557 493
rect 2397 367 2463 421
rect 2497 333 2557 442
rect 2319 299 2557 333
rect 2309 177 2370 185
rect 1757 117 1873 151
rect 1494 51 1723 85
rect 1823 66 1873 117
rect 1907 17 1957 132
rect 1991 117 2107 151
rect 1991 66 2041 117
rect 2141 85 2175 154
rect 2209 119 2275 177
rect 2309 143 2547 177
rect 2309 85 2370 143
rect 2141 51 2370 85
rect 2404 17 2447 109
rect 2481 51 2547 143
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2576 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 305 357 339 391
rect 949 357 983 391
rect 1593 357 1627 391
rect 2237 357 2271 391
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
<< metal1 >>
rect 0 561 2576 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2576 561
rect 0 496 2576 527
rect 293 391 351 397
rect 293 357 305 391
rect 339 388 351 391
rect 937 391 995 397
rect 937 388 949 391
rect 339 360 949 388
rect 339 357 351 360
rect 293 351 351 357
rect 937 357 949 360
rect 983 388 995 391
rect 1581 391 1639 397
rect 1581 388 1593 391
rect 983 360 1593 388
rect 983 357 995 360
rect 937 351 995 357
rect 1581 357 1593 360
rect 1627 388 1639 391
rect 2225 391 2283 397
rect 2225 388 2237 391
rect 1627 360 2237 388
rect 1627 357 1639 360
rect 1581 351 1639 357
rect 2225 357 2237 360
rect 2271 357 2283 391
rect 2225 351 2283 357
rect 0 17 2576 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2576 17
rect 0 -48 2576 -17
<< labels >>
rlabel locali s 19 211 183 265 6 D[0]
port 1 nsew signal input
rlabel locali s 1105 211 1269 265 6 D[1]
port 2 nsew signal input
rlabel locali s 1307 211 1471 265 6 D[2]
port 3 nsew signal input
rlabel locali s 2393 211 2557 265 6 D[3]
port 4 nsew signal input
rlabel locali s 558 205 625 259 6 S[0]
port 5 nsew signal input
rlabel locali s 663 205 730 259 6 S[1]
port 6 nsew signal input
rlabel locali s 1846 205 1913 259 6 S[2]
port 7 nsew signal input
rlabel locali s 1951 205 2018 259 6 S[3]
port 8 nsew signal input
rlabel metal1 s 2225 388 2283 397 6 Z
port 9 nsew signal output
rlabel metal1 s 2225 351 2283 360 6 Z
port 9 nsew signal output
rlabel metal1 s 1581 388 1639 397 6 Z
port 9 nsew signal output
rlabel metal1 s 1581 351 1639 360 6 Z
port 9 nsew signal output
rlabel metal1 s 937 388 995 397 6 Z
port 9 nsew signal output
rlabel metal1 s 937 351 995 360 6 Z
port 9 nsew signal output
rlabel metal1 s 293 388 351 397 6 Z
port 9 nsew signal output
rlabel metal1 s 293 360 2283 388 6 Z
port 9 nsew signal output
rlabel metal1 s 293 351 351 360 6 Z
port 9 nsew signal output
rlabel metal1 s 0 -48 2576 48 8 VGND
port 10 nsew ground bidirectional
rlabel metal1 s 0 496 2576 592 6 VPWR
port 11 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2576 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2741656
string GDS_START 2711914
<< end >>
