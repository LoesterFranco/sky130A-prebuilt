magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 232 406 269 487
rect 232 371 375 406
rect 85 149 167 265
rect 297 165 375 371
rect 228 131 375 165
rect 228 51 269 131
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 17 333 71 487
rect 105 371 181 527
rect 303 442 380 527
rect 17 299 263 333
rect 17 117 51 299
rect 203 199 263 299
rect 17 51 69 117
rect 121 17 176 113
rect 303 17 380 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
rlabel locali s 85 149 167 265 6 A
port 1 nsew signal input
rlabel locali s 297 165 375 371 6 X
port 2 nsew signal output
rlabel locali s 232 406 269 487 6 X
port 2 nsew signal output
rlabel locali s 232 371 375 406 6 X
port 2 nsew signal output
rlabel locali s 228 131 375 165 6 X
port 2 nsew signal output
rlabel locali s 228 51 269 131 6 X
port 2 nsew signal output
rlabel metal1 s 0 -48 460 48 8 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 496 460 592 6 VPWR
port 4 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 460 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1765424
string GDS_START 1760910
<< end >>
