magic
tech sky130A
magscale 1 2
timestamp 1604502729
<< locali >>
rect 123 424 332 596
rect 466 424 741 596
rect 123 390 839 424
rect 217 336 455 356
rect 102 270 455 336
rect 489 270 759 356
rect 793 236 839 390
rect 467 202 839 236
rect 467 122 533 202
rect 667 122 741 202
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 23 370 89 649
rect 366 458 432 649
rect 775 458 841 649
rect 23 202 433 236
rect 23 70 73 202
rect 109 17 175 161
rect 211 70 245 202
rect 281 17 347 161
rect 383 85 433 202
rect 567 85 633 161
rect 775 85 841 161
rect 383 51 841 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel locali s 489 270 759 356 6 A
port 1 nsew signal input
rlabel locali s 217 336 455 356 6 B
port 2 nsew signal input
rlabel locali s 102 270 455 336 6 B
port 2 nsew signal input
rlabel locali s 793 236 839 390 6 Y
port 3 nsew signal output
rlabel locali s 667 122 741 202 6 Y
port 3 nsew signal output
rlabel locali s 467 202 839 236 6 Y
port 3 nsew signal output
rlabel locali s 467 122 533 202 6 Y
port 3 nsew signal output
rlabel locali s 466 424 741 596 6 Y
port 3 nsew signal output
rlabel locali s 123 424 332 596 6 Y
port 3 nsew signal output
rlabel locali s 123 390 839 424 6 Y
port 3 nsew signal output
rlabel metal1 s 0 -49 864 49 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 617 864 715 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1926168
string GDS_START 1918250
<< end >>
