magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 113 333 179 493
rect 301 333 367 493
rect 489 333 555 493
rect 677 333 743 493
rect 865 333 931 493
rect 1053 333 1119 493
rect 113 299 1119 333
rect 79 211 553 265
rect 667 177 727 299
rect 1065 265 1119 299
rect 761 211 1031 265
rect 1065 211 1183 265
rect 1065 177 1119 211
rect 667 127 1119 177
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 25 299 79 527
rect 213 367 267 527
rect 401 367 455 527
rect 589 367 643 527
rect 777 367 831 527
rect 965 367 1019 527
rect 1153 299 1207 527
rect 18 143 633 177
rect 18 51 85 143
rect 119 17 173 109
rect 207 51 273 143
rect 307 17 361 109
rect 395 51 461 143
rect 495 17 549 109
rect 583 93 633 143
rect 1153 93 1213 177
rect 583 51 1213 93
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
rlabel locali s 761 211 1031 265 6 A
port 1 nsew signal input
rlabel locali s 79 211 553 265 6 B
port 2 nsew signal input
rlabel locali s 1065 265 1119 299 6 Y
port 3 nsew signal output
rlabel locali s 1065 211 1183 265 6 Y
port 3 nsew signal output
rlabel locali s 1065 177 1119 211 6 Y
port 3 nsew signal output
rlabel locali s 1053 333 1119 493 6 Y
port 3 nsew signal output
rlabel locali s 865 333 931 493 6 Y
port 3 nsew signal output
rlabel locali s 677 333 743 493 6 Y
port 3 nsew signal output
rlabel locali s 667 177 727 299 6 Y
port 3 nsew signal output
rlabel locali s 667 127 1119 177 6 Y
port 3 nsew signal output
rlabel locali s 489 333 555 493 6 Y
port 3 nsew signal output
rlabel locali s 301 333 367 493 6 Y
port 3 nsew signal output
rlabel locali s 113 333 179 493 6 Y
port 3 nsew signal output
rlabel locali s 113 299 1119 333 6 Y
port 3 nsew signal output
rlabel metal1 s 0 -48 1288 48 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 496 1288 592 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1288 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3440178
string GDS_START 3430442
<< end >>
