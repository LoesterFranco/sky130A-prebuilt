magic
tech sky130A
magscale 1 2
timestamp 1604502701
<< nwell >>
rect -38 332 710 704
<< pwell >>
rect 0 0 672 49
<< scpmos >>
rect 113 368 143 536
rect 230 368 260 592
rect 320 368 350 592
rect 434 368 464 592
rect 524 368 554 592
<< nmoslvt >>
rect 125 112 155 222
rect 233 74 263 222
rect 311 74 341 222
rect 413 74 443 222
rect 521 74 551 222
<< ndiff >>
rect 27 186 125 222
rect 27 152 80 186
rect 114 152 125 186
rect 27 112 125 152
rect 155 127 233 222
rect 155 112 187 127
rect 175 93 187 112
rect 221 93 233 127
rect 175 74 233 93
rect 263 74 311 222
rect 341 74 413 222
rect 443 74 521 222
rect 551 194 643 222
rect 551 160 581 194
rect 615 160 643 194
rect 551 120 643 160
rect 551 86 581 120
rect 615 86 643 120
rect 551 74 643 86
<< pdiff >>
rect 161 580 230 592
rect 161 546 173 580
rect 207 546 230 580
rect 161 536 230 546
rect 54 524 113 536
rect 54 490 66 524
rect 100 490 113 524
rect 54 414 113 490
rect 54 380 66 414
rect 100 380 113 414
rect 54 368 113 380
rect 143 497 230 536
rect 143 463 173 497
rect 207 463 230 497
rect 143 414 230 463
rect 143 380 173 414
rect 207 380 230 414
rect 143 368 230 380
rect 260 580 320 592
rect 260 546 273 580
rect 307 546 320 580
rect 260 497 320 546
rect 260 463 273 497
rect 307 463 320 497
rect 260 414 320 463
rect 260 380 273 414
rect 307 380 320 414
rect 260 368 320 380
rect 350 580 434 592
rect 350 546 373 580
rect 407 546 434 580
rect 350 498 434 546
rect 350 464 373 498
rect 407 464 434 498
rect 350 368 434 464
rect 464 580 524 592
rect 464 546 477 580
rect 511 546 524 580
rect 464 497 524 546
rect 464 463 477 497
rect 511 463 524 497
rect 464 414 524 463
rect 464 380 477 414
rect 511 380 524 414
rect 464 368 524 380
rect 554 582 623 592
rect 554 548 577 582
rect 611 548 623 582
rect 554 514 623 548
rect 554 480 577 514
rect 611 480 623 514
rect 554 446 623 480
rect 554 412 577 446
rect 611 412 623 446
rect 554 368 623 412
<< ndiffc >>
rect 80 152 114 186
rect 187 93 221 127
rect 581 160 615 194
rect 581 86 615 120
<< pdiffc >>
rect 173 546 207 580
rect 66 490 100 524
rect 66 380 100 414
rect 173 463 207 497
rect 173 380 207 414
rect 273 546 307 580
rect 273 463 307 497
rect 273 380 307 414
rect 373 546 407 580
rect 373 464 407 498
rect 477 546 511 580
rect 477 463 511 497
rect 477 380 511 414
rect 577 548 611 582
rect 577 480 611 514
rect 577 412 611 446
<< poly >>
rect 230 592 260 618
rect 320 592 350 618
rect 434 592 464 618
rect 524 592 554 618
rect 113 536 143 562
rect 113 353 143 368
rect 230 353 260 368
rect 320 353 350 368
rect 434 353 464 368
rect 524 353 554 368
rect 110 310 146 353
rect 227 310 263 353
rect 317 310 353 353
rect 431 310 467 353
rect 521 310 557 353
rect 89 294 155 310
rect 89 260 105 294
rect 139 260 155 294
rect 89 244 155 260
rect 197 294 263 310
rect 197 260 213 294
rect 247 260 263 294
rect 197 244 263 260
rect 305 294 371 310
rect 305 260 321 294
rect 355 260 371 294
rect 305 244 371 260
rect 413 294 479 310
rect 413 260 429 294
rect 463 260 479 294
rect 413 244 479 260
rect 521 294 587 310
rect 521 260 537 294
rect 571 260 587 294
rect 521 244 587 260
rect 125 222 155 244
rect 233 222 263 244
rect 311 222 341 244
rect 413 222 443 244
rect 521 222 551 244
rect 125 86 155 112
rect 233 48 263 74
rect 311 48 341 74
rect 413 48 443 74
rect 521 48 551 74
<< polycont >>
rect 105 260 139 294
rect 213 260 247 294
rect 321 260 355 294
rect 429 260 463 294
rect 537 260 571 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 157 580 223 649
rect 157 546 173 580
rect 207 546 223 580
rect 21 524 116 540
rect 21 490 66 524
rect 100 490 116 524
rect 21 414 116 490
rect 21 380 66 414
rect 100 380 116 414
rect 21 364 116 380
rect 157 497 223 546
rect 157 463 173 497
rect 207 463 223 497
rect 157 414 223 463
rect 157 380 173 414
rect 207 380 223 414
rect 157 364 223 380
rect 257 580 323 596
rect 257 546 273 580
rect 307 546 323 580
rect 257 497 323 546
rect 257 463 273 497
rect 307 463 323 497
rect 357 580 423 649
rect 357 546 373 580
rect 407 546 423 580
rect 357 498 423 546
rect 357 464 373 498
rect 407 464 423 498
rect 457 580 527 596
rect 457 546 477 580
rect 511 546 527 580
rect 457 497 527 546
rect 257 430 323 463
rect 457 463 477 497
rect 511 463 527 497
rect 457 430 527 463
rect 257 414 527 430
rect 257 380 273 414
rect 307 380 477 414
rect 511 380 527 414
rect 561 582 627 649
rect 561 548 577 582
rect 611 548 627 582
rect 561 514 627 548
rect 561 480 577 514
rect 611 480 627 514
rect 561 446 627 480
rect 561 412 577 446
rect 611 412 627 446
rect 257 378 527 380
rect 257 364 655 378
rect 21 202 55 364
rect 323 344 655 364
rect 89 294 163 310
rect 89 260 105 294
rect 139 260 163 294
rect 89 236 163 260
rect 197 294 263 310
rect 197 260 213 294
rect 247 260 263 294
rect 197 236 263 260
rect 305 294 371 310
rect 305 260 321 294
rect 355 260 371 294
rect 305 236 371 260
rect 409 294 479 310
rect 409 260 429 294
rect 463 260 479 294
rect 409 236 479 260
rect 513 294 587 310
rect 513 260 537 294
rect 571 260 587 294
rect 513 244 587 260
rect 513 202 547 244
rect 621 210 655 344
rect 21 186 547 202
rect 21 152 80 186
rect 114 168 547 186
rect 581 194 655 210
rect 114 152 130 168
rect 21 136 130 152
rect 615 160 655 194
rect 171 127 237 134
rect 171 93 187 127
rect 221 93 237 127
rect 171 17 237 93
rect 581 120 655 160
rect 615 86 655 120
rect 581 70 655 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel comment s 0 0 0 0 4 nand4b_1
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 127 242 161 276 0 FreeSans 340 0 0 0 A_N
port 1 nsew
flabel corelocali s 223 242 257 276 0 FreeSans 340 0 0 0 D
port 4 nsew
flabel corelocali s 415 390 449 424 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 319 242 353 276 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 415 242 449 276 0 FreeSans 340 0 0 0 B
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 672 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1452656
string GDS_START 1446650
<< end >>
