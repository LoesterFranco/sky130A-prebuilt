magic
tech sky130A
magscale 1 2
timestamp 1604502701
<< nwell >>
rect -38 332 614 704
<< pwell >>
rect 0 0 576 49
<< scpmos >>
rect 90 424 120 592
rect 275 368 305 592
rect 365 368 395 592
rect 461 368 491 592
<< nmoslvt >>
rect 83 74 113 184
rect 278 74 308 222
rect 374 74 404 222
rect 462 74 492 222
<< ndiff >>
rect 222 210 278 222
rect 27 146 83 184
rect 27 112 38 146
rect 72 112 83 146
rect 27 74 83 112
rect 113 146 168 184
rect 113 112 124 146
rect 158 112 168 146
rect 113 74 168 112
rect 222 176 233 210
rect 267 176 278 210
rect 222 120 278 176
rect 222 86 233 120
rect 267 86 278 120
rect 222 74 278 86
rect 308 210 374 222
rect 308 176 329 210
rect 363 176 374 210
rect 308 120 374 176
rect 308 86 329 120
rect 363 86 374 120
rect 308 74 374 86
rect 404 120 462 222
rect 404 86 416 120
rect 450 86 462 120
rect 404 74 462 86
rect 492 210 549 222
rect 492 176 503 210
rect 537 176 549 210
rect 492 120 549 176
rect 492 86 503 120
rect 537 86 549 120
rect 492 74 549 86
<< pdiff >>
rect 31 580 90 592
rect 31 546 43 580
rect 77 546 90 580
rect 31 470 90 546
rect 31 436 43 470
rect 77 436 90 470
rect 31 424 90 436
rect 120 580 275 592
rect 120 546 143 580
rect 177 546 211 580
rect 245 546 275 580
rect 120 508 275 546
rect 120 474 143 508
rect 177 474 211 508
rect 245 474 275 508
rect 120 424 275 474
rect 222 368 275 424
rect 305 580 365 592
rect 305 546 318 580
rect 352 546 365 580
rect 305 497 365 546
rect 305 463 318 497
rect 352 463 365 497
rect 305 414 365 463
rect 305 380 318 414
rect 352 380 365 414
rect 305 368 365 380
rect 395 368 461 592
rect 491 580 549 592
rect 491 546 504 580
rect 538 546 549 580
rect 491 510 549 546
rect 491 476 504 510
rect 538 476 549 510
rect 491 440 549 476
rect 491 406 504 440
rect 538 406 549 440
rect 491 368 549 406
<< ndiffc >>
rect 38 112 72 146
rect 124 112 158 146
rect 233 176 267 210
rect 233 86 267 120
rect 329 176 363 210
rect 329 86 363 120
rect 416 86 450 120
rect 503 176 537 210
rect 503 86 537 120
<< pdiffc >>
rect 43 546 77 580
rect 43 436 77 470
rect 143 546 177 580
rect 211 546 245 580
rect 143 474 177 508
rect 211 474 245 508
rect 318 546 352 580
rect 318 463 352 497
rect 318 380 352 414
rect 504 546 538 580
rect 504 476 538 510
rect 504 406 538 440
<< poly >>
rect 90 592 120 618
rect 275 592 305 618
rect 365 592 395 618
rect 461 592 491 618
rect 90 409 120 424
rect 87 404 123 409
rect 83 374 123 404
rect 83 356 113 374
rect 47 340 113 356
rect 275 353 305 368
rect 365 353 395 368
rect 461 353 491 368
rect 47 306 63 340
rect 97 306 113 340
rect 47 290 113 306
rect 83 184 113 290
rect 161 310 227 326
rect 161 276 177 310
rect 211 290 227 310
rect 272 290 308 353
rect 362 326 398 353
rect 458 326 494 353
rect 211 276 308 290
rect 161 260 308 276
rect 350 310 416 326
rect 350 276 366 310
rect 400 276 416 310
rect 350 260 416 276
rect 458 310 555 326
rect 458 276 505 310
rect 539 276 555 310
rect 458 260 555 276
rect 278 222 308 260
rect 374 222 404 260
rect 462 222 492 260
rect 83 48 113 74
rect 278 48 308 74
rect 374 48 404 74
rect 462 48 492 74
<< polycont >>
rect 63 306 97 340
rect 177 276 211 310
rect 366 276 400 310
rect 505 276 539 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 27 580 93 596
rect 27 546 43 580
rect 77 546 93 580
rect 27 470 93 546
rect 27 436 43 470
rect 77 436 93 470
rect 127 580 261 649
rect 127 546 143 580
rect 177 546 211 580
rect 245 546 261 580
rect 127 508 261 546
rect 127 474 143 508
rect 177 474 211 508
rect 245 474 261 508
rect 127 458 261 474
rect 295 580 368 596
rect 295 546 318 580
rect 352 546 368 580
rect 504 580 554 649
rect 295 497 368 546
rect 295 463 318 497
rect 352 463 368 497
rect 27 424 93 436
rect 27 390 183 424
rect 295 414 368 463
rect 295 398 318 414
rect 25 340 113 356
rect 25 306 63 340
rect 97 306 113 340
rect 25 290 113 306
rect 149 326 183 390
rect 261 380 318 398
rect 352 380 368 414
rect 261 364 368 380
rect 149 310 227 326
rect 149 276 177 310
rect 211 276 227 310
rect 149 260 227 276
rect 149 256 183 260
rect 22 222 183 256
rect 261 226 295 364
rect 409 326 455 578
rect 538 546 554 580
rect 504 510 554 546
rect 538 476 554 510
rect 504 440 554 476
rect 538 406 554 440
rect 504 390 554 406
rect 350 310 455 326
rect 350 276 366 310
rect 400 276 455 310
rect 350 260 455 276
rect 489 310 555 356
rect 489 276 505 310
rect 539 276 555 310
rect 489 260 555 276
rect 22 146 72 222
rect 217 210 295 226
rect 22 112 38 146
rect 22 70 72 112
rect 108 146 174 188
rect 108 112 124 146
rect 158 112 174 146
rect 108 17 174 112
rect 217 176 233 210
rect 267 176 295 210
rect 217 120 295 176
rect 217 86 233 120
rect 267 86 295 120
rect 217 70 295 86
rect 329 210 553 226
rect 363 192 503 210
rect 329 120 363 176
rect 537 176 553 210
rect 329 70 363 86
rect 399 120 467 136
rect 399 86 416 120
rect 450 86 467 120
rect 399 17 467 86
rect 503 120 553 176
rect 537 86 553 120
rect 503 70 553 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o21bai_1
flabel pwell s 0 0 576 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 576 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 576 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 576 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 B1_N
port 3 nsew
flabel corelocali s 319 390 353 424 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 319 464 353 498 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 319 538 353 572 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 415 390 449 424 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 415 464 449 498 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 415 538 449 572 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 576 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1135606
string GDS_START 1129240
<< end >>
