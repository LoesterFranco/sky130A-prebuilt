magic
tech sky130A
magscale 1 2
timestamp 1604502705
<< nwell >>
rect -38 356 2822 704
rect -38 332 1199 356
rect 1945 332 2822 356
rect 750 311 1199 332
<< pwell >>
rect 0 0 2784 49
<< scnmos >>
rect 84 88 114 172
rect 294 81 324 165
rect 366 81 396 165
rect 508 81 538 165
rect 586 81 616 165
rect 674 81 704 165
rect 824 74 854 222
rect 1044 79 1074 227
rect 1242 123 1272 207
rect 1381 123 1411 207
rect 1459 123 1489 207
rect 1537 123 1567 207
rect 1655 144 1685 272
rect 1797 144 1827 272
rect 2043 74 2073 158
rect 2123 74 2153 158
rect 2235 74 2265 158
rect 2313 74 2343 158
rect 2554 74 2584 184
rect 2670 74 2700 222
<< pmoshvt >>
rect 86 464 116 592
rect 176 464 206 592
rect 254 464 284 592
rect 441 464 471 592
rect 519 464 549 592
rect 643 464 673 592
rect 929 347 959 547
rect 1019 347 1049 547
rect 1221 463 1251 547
rect 1311 463 1341 547
rect 1402 463 1432 547
rect 1492 463 1522 547
rect 1722 392 1752 592
rect 1909 392 1939 592
rect 2012 508 2042 592
rect 2094 508 2124 592
rect 2249 508 2279 592
rect 2339 508 2369 592
rect 2551 424 2581 592
rect 2667 368 2697 592
<< ndiff >>
rect 27 147 84 172
rect 27 113 39 147
rect 73 113 84 147
rect 27 88 84 113
rect 114 147 185 172
rect 774 165 824 222
rect 114 113 139 147
rect 173 113 185 147
rect 114 88 185 113
rect 239 132 294 165
rect 239 98 249 132
rect 283 98 294 132
rect 239 81 294 98
rect 324 81 366 165
rect 396 153 508 165
rect 396 119 435 153
rect 469 119 508 153
rect 396 81 508 119
rect 538 81 586 165
rect 616 140 674 165
rect 616 106 628 140
rect 662 106 674 140
rect 616 81 674 106
rect 704 81 824 165
rect 719 74 824 81
rect 854 208 911 222
rect 854 174 865 208
rect 899 174 911 208
rect 854 74 911 174
rect 965 79 1044 227
rect 1074 215 1131 227
rect 1074 181 1085 215
rect 1119 181 1131 215
rect 1605 207 1655 272
rect 1074 79 1131 181
rect 1185 190 1242 207
rect 1185 156 1197 190
rect 1231 156 1242 190
rect 1185 123 1242 156
rect 1272 195 1381 207
rect 1272 161 1334 195
rect 1368 161 1381 195
rect 1272 123 1381 161
rect 1411 123 1459 207
rect 1489 123 1537 207
rect 1567 144 1655 207
rect 1685 260 1797 272
rect 1685 226 1724 260
rect 1758 226 1797 260
rect 1685 144 1797 226
rect 1827 158 1877 272
rect 2599 210 2670 222
rect 2599 184 2625 210
rect 1827 144 2043 158
rect 1567 124 1640 144
rect 1567 123 1594 124
rect 719 72 809 74
rect 719 38 747 72
rect 781 38 809 72
rect 965 72 1029 79
rect 719 27 809 38
rect 965 38 980 72
rect 1014 38 1029 72
rect 965 27 1029 38
rect 1582 90 1594 123
rect 1628 90 1640 124
rect 1582 78 1640 90
rect 1842 108 2043 144
rect 1842 74 1854 108
rect 1888 74 1982 108
rect 2016 74 2043 108
rect 2073 74 2123 158
rect 2153 120 2235 158
rect 2153 86 2176 120
rect 2210 86 2235 120
rect 2153 74 2235 86
rect 2265 74 2313 158
rect 2343 140 2443 158
rect 2343 106 2375 140
rect 2409 106 2443 140
rect 2343 74 2443 106
rect 2497 146 2554 184
rect 2497 112 2509 146
rect 2543 112 2554 146
rect 2497 74 2554 112
rect 2584 176 2625 184
rect 2659 176 2670 210
rect 2584 128 2670 176
rect 2584 94 2611 128
rect 2645 94 2670 128
rect 2584 74 2670 94
rect 2700 210 2757 222
rect 2700 176 2711 210
rect 2745 176 2757 210
rect 2700 120 2757 176
rect 2700 86 2711 120
rect 2745 86 2757 120
rect 2700 74 2757 86
rect 1842 62 2028 74
<< pdiff >>
rect 567 628 625 639
rect 567 594 579 628
rect 613 594 625 628
rect 567 592 625 594
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 510 86 546
rect 27 476 39 510
rect 73 476 86 510
rect 27 464 86 476
rect 116 578 176 592
rect 116 544 129 578
rect 163 544 176 578
rect 116 464 176 544
rect 206 464 254 592
rect 284 576 441 592
rect 284 542 297 576
rect 331 542 394 576
rect 428 542 441 576
rect 284 464 441 542
rect 471 464 519 592
rect 549 464 643 592
rect 673 580 732 592
rect 673 546 686 580
rect 720 546 732 580
rect 1665 580 1722 592
rect 673 510 732 546
rect 673 476 686 510
rect 720 476 732 510
rect 673 464 732 476
rect 862 398 929 547
rect 862 364 882 398
rect 916 364 929 398
rect 862 347 929 364
rect 959 534 1019 547
rect 959 500 972 534
rect 1006 500 1019 534
rect 959 347 1019 500
rect 1049 433 1108 547
rect 1162 526 1221 547
rect 1162 492 1174 526
rect 1208 492 1221 526
rect 1162 463 1221 492
rect 1251 526 1311 547
rect 1251 492 1264 526
rect 1298 492 1311 526
rect 1251 463 1311 492
rect 1341 463 1402 547
rect 1432 526 1492 547
rect 1432 492 1445 526
rect 1479 492 1492 526
rect 1432 463 1492 492
rect 1522 526 1581 547
rect 1522 492 1535 526
rect 1569 492 1581 526
rect 1522 463 1581 492
rect 1665 546 1675 580
rect 1709 546 1722 580
rect 1665 512 1722 546
rect 1665 478 1675 512
rect 1709 478 1722 512
rect 1049 398 1116 433
rect 1049 364 1062 398
rect 1096 364 1116 398
rect 1049 347 1116 364
rect 1665 392 1722 478
rect 1752 580 1909 592
rect 1752 546 1775 580
rect 1809 546 1862 580
rect 1896 546 1909 580
rect 1752 512 1909 546
rect 1752 478 1775 512
rect 1809 478 1862 512
rect 1896 478 1909 512
rect 1752 444 1909 478
rect 1752 410 1775 444
rect 1809 410 1862 444
rect 1896 410 1909 444
rect 1752 392 1909 410
rect 1939 580 2012 592
rect 1939 546 1963 580
rect 1997 546 2012 580
rect 1939 512 2012 546
rect 1939 478 1952 512
rect 1986 508 2012 512
rect 2042 508 2094 592
rect 2124 580 2249 592
rect 2124 546 2164 580
rect 2198 546 2249 580
rect 2124 508 2249 546
rect 2279 567 2339 592
rect 2279 533 2292 567
rect 2326 533 2339 567
rect 2279 508 2339 533
rect 2369 578 2438 592
rect 2369 544 2392 578
rect 2426 544 2438 578
rect 2369 508 2438 544
rect 2492 580 2551 592
rect 2492 546 2504 580
rect 2538 546 2551 580
rect 1986 478 1994 508
rect 1939 444 1994 478
rect 1939 410 1952 444
rect 1986 410 1994 444
rect 1939 392 1994 410
rect 2492 470 2551 546
rect 2492 436 2504 470
rect 2538 436 2551 470
rect 2492 424 2551 436
rect 2581 580 2667 592
rect 2581 546 2611 580
rect 2645 546 2667 580
rect 2581 497 2667 546
rect 2581 463 2611 497
rect 2645 463 2667 497
rect 2581 424 2667 463
rect 2599 414 2667 424
rect 2599 380 2611 414
rect 2645 380 2667 414
rect 2599 368 2667 380
rect 2697 580 2757 592
rect 2697 546 2711 580
rect 2745 546 2757 580
rect 2697 497 2757 546
rect 2697 463 2711 497
rect 2745 463 2757 497
rect 2697 414 2757 463
rect 2697 380 2711 414
rect 2745 380 2757 414
rect 2697 368 2757 380
<< ndiffc >>
rect 39 113 73 147
rect 139 113 173 147
rect 249 98 283 132
rect 435 119 469 153
rect 628 106 662 140
rect 865 174 899 208
rect 1085 181 1119 215
rect 1197 156 1231 190
rect 1334 161 1368 195
rect 1724 226 1758 260
rect 747 38 781 72
rect 980 38 1014 72
rect 1594 90 1628 124
rect 1854 74 1888 108
rect 1982 74 2016 108
rect 2176 86 2210 120
rect 2375 106 2409 140
rect 2509 112 2543 146
rect 2625 176 2659 210
rect 2611 94 2645 128
rect 2711 176 2745 210
rect 2711 86 2745 120
<< pdiffc >>
rect 579 594 613 628
rect 39 546 73 580
rect 39 476 73 510
rect 129 544 163 578
rect 297 542 331 576
rect 394 542 428 576
rect 686 546 720 580
rect 686 476 720 510
rect 882 364 916 398
rect 972 500 1006 534
rect 1174 492 1208 526
rect 1264 492 1298 526
rect 1445 492 1479 526
rect 1535 492 1569 526
rect 1675 546 1709 580
rect 1675 478 1709 512
rect 1062 364 1096 398
rect 1775 546 1809 580
rect 1862 546 1896 580
rect 1775 478 1809 512
rect 1862 478 1896 512
rect 1775 410 1809 444
rect 1862 410 1896 444
rect 1963 546 1997 580
rect 1952 478 1986 512
rect 2164 546 2198 580
rect 2292 533 2326 567
rect 2392 544 2426 578
rect 2504 546 2538 580
rect 1952 410 1986 444
rect 2504 436 2538 470
rect 2611 546 2645 580
rect 2611 463 2645 497
rect 2611 380 2645 414
rect 2711 546 2745 580
rect 2711 463 2745 497
rect 2711 380 2745 414
<< poly >>
rect 86 592 116 618
rect 176 592 206 618
rect 254 592 284 618
rect 441 592 471 618
rect 519 592 549 618
rect 643 615 1522 645
rect 643 592 673 615
rect 929 547 959 573
rect 1019 547 1049 573
rect 1221 547 1251 573
rect 1311 547 1341 573
rect 1402 547 1432 573
rect 1492 547 1522 615
rect 1722 592 1752 618
rect 1909 592 1939 618
rect 2012 592 2042 618
rect 2094 592 2124 618
rect 2249 592 2279 618
rect 2339 592 2369 618
rect 2551 592 2581 618
rect 2667 592 2697 618
rect 86 449 116 464
rect 176 449 206 464
rect 254 449 284 464
rect 441 449 471 464
rect 519 449 549 464
rect 643 449 673 464
rect 83 416 119 449
rect 173 416 209 449
rect 84 400 209 416
rect 84 366 123 400
rect 157 386 209 400
rect 251 422 287 449
rect 251 406 396 422
rect 251 392 346 406
rect 157 366 173 386
rect 84 332 173 366
rect 330 372 346 392
rect 380 372 396 406
rect 330 356 396 372
rect 84 298 123 332
rect 157 298 173 332
rect 84 282 173 298
rect 84 172 114 282
rect 258 237 324 253
rect 258 203 274 237
rect 308 203 324 237
rect 258 187 324 203
rect 294 165 324 187
rect 366 165 396 356
rect 438 377 474 449
rect 516 419 590 449
rect 640 419 704 449
rect 438 361 509 377
rect 438 327 459 361
rect 493 327 509 361
rect 438 311 509 327
rect 560 371 590 419
rect 674 405 704 419
rect 674 389 747 405
rect 560 355 626 371
rect 560 321 576 355
rect 610 321 626 355
rect 560 305 626 321
rect 674 355 697 389
rect 731 355 747 389
rect 674 321 747 355
rect 444 241 538 257
rect 444 207 460 241
rect 494 207 538 241
rect 444 191 538 207
rect 508 165 538 191
rect 586 165 616 305
rect 674 287 697 321
rect 731 287 747 321
rect 929 310 959 347
rect 1019 315 1049 347
rect 674 271 747 287
rect 824 294 959 310
rect 674 165 704 271
rect 824 260 871 294
rect 905 260 959 294
rect 824 244 959 260
rect 1001 305 1067 315
rect 1221 305 1251 463
rect 1311 413 1341 463
rect 1293 397 1359 413
rect 1293 363 1309 397
rect 1343 363 1359 397
rect 1293 347 1359 363
rect 1402 374 1432 463
rect 1492 448 1522 463
rect 1492 416 1567 448
rect 1402 358 1495 374
rect 1402 324 1445 358
rect 1479 324 1495 358
rect 1402 308 1495 324
rect 1537 360 1567 416
rect 2012 493 2042 508
rect 2094 493 2124 508
rect 2249 493 2279 508
rect 2339 493 2369 508
rect 1722 377 1752 392
rect 1909 377 1939 392
rect 1719 360 1755 377
rect 1537 344 1603 360
rect 1537 310 1553 344
rect 1587 310 1603 344
rect 1001 299 1350 305
rect 1001 265 1017 299
rect 1051 275 1350 299
rect 1051 265 1074 275
rect 1001 249 1074 265
rect 824 222 854 244
rect 1044 227 1074 249
rect 1320 260 1350 275
rect 84 62 114 88
rect 294 55 324 81
rect 366 55 396 81
rect 508 55 538 81
rect 586 55 616 81
rect 674 55 704 81
rect 1242 207 1272 233
rect 1320 230 1411 260
rect 1381 207 1411 230
rect 1459 207 1489 308
rect 1537 294 1603 310
rect 1645 344 1755 360
rect 1645 310 1661 344
rect 1695 310 1755 344
rect 1645 294 1755 310
rect 1797 344 1864 360
rect 1797 310 1814 344
rect 1848 310 1864 344
rect 1797 294 1864 310
rect 1537 207 1567 294
rect 1655 272 1685 294
rect 1797 272 1827 294
rect 1906 246 1942 377
rect 2009 311 2045 493
rect 2091 476 2127 493
rect 2246 487 2282 493
rect 2087 460 2153 476
rect 2087 426 2103 460
rect 2137 426 2153 460
rect 2087 410 2153 426
rect 2009 295 2079 311
rect 2009 261 2029 295
rect 2063 261 2079 295
rect 1899 230 1965 246
rect 2009 245 2079 261
rect 1899 196 1915 230
rect 1949 203 1965 230
rect 1949 196 2073 203
rect 1899 173 2073 196
rect 2043 158 2073 173
rect 2123 158 2153 410
rect 2235 457 2282 487
rect 2235 308 2265 457
rect 2336 409 2372 493
rect 2551 409 2581 424
rect 2336 379 2584 409
rect 2336 314 2366 379
rect 2667 353 2697 368
rect 2664 337 2700 353
rect 2496 321 2700 337
rect 2199 292 2265 308
rect 2199 258 2215 292
rect 2249 258 2265 292
rect 2199 242 2265 258
rect 2235 158 2265 242
rect 2313 298 2379 314
rect 2313 264 2329 298
rect 2363 264 2379 298
rect 2496 287 2512 321
rect 2546 287 2700 321
rect 2496 271 2700 287
rect 2313 230 2379 264
rect 2313 196 2329 230
rect 2363 229 2379 230
rect 2363 199 2584 229
rect 2670 222 2700 271
rect 2363 196 2379 199
rect 2313 180 2379 196
rect 2554 184 2584 199
rect 2313 158 2343 180
rect 1242 101 1272 123
rect 1242 85 1331 101
rect 824 48 854 74
rect 1044 53 1074 79
rect 1242 51 1281 85
rect 1315 51 1331 85
rect 1242 33 1331 51
rect 1381 55 1411 123
rect 1459 97 1489 123
rect 1537 97 1567 123
rect 1655 118 1685 144
rect 1797 55 1827 144
rect 1381 25 1827 55
rect 2043 48 2073 74
rect 2123 48 2153 74
rect 2235 48 2265 74
rect 2313 48 2343 74
rect 2554 48 2584 74
rect 2670 48 2700 74
<< polycont >>
rect 123 366 157 400
rect 346 372 380 406
rect 123 298 157 332
rect 274 203 308 237
rect 459 327 493 361
rect 576 321 610 355
rect 697 355 731 389
rect 460 207 494 241
rect 697 287 731 321
rect 871 260 905 294
rect 1309 363 1343 397
rect 1445 324 1479 358
rect 1553 310 1587 344
rect 1017 265 1051 299
rect 1661 310 1695 344
rect 1814 310 1848 344
rect 2103 426 2137 460
rect 2029 261 2063 295
rect 1915 196 1949 230
rect 2215 258 2249 292
rect 2329 264 2363 298
rect 2512 287 2546 321
rect 2329 196 2363 230
rect 1281 51 1315 85
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 23 580 73 596
rect 23 546 39 580
rect 23 510 73 546
rect 113 578 179 649
rect 563 628 629 649
rect 563 594 579 628
rect 613 594 629 628
rect 113 544 129 578
rect 163 544 179 578
rect 113 526 179 544
rect 281 576 444 592
rect 281 542 297 576
rect 331 542 394 576
rect 428 560 444 576
rect 686 580 736 596
rect 428 546 686 560
rect 720 546 736 580
rect 428 542 736 546
rect 281 526 736 542
rect 23 476 39 510
rect 686 510 736 526
rect 73 476 509 492
rect 23 458 509 476
rect 23 248 73 458
rect 107 400 173 416
rect 107 366 123 400
rect 157 366 173 400
rect 107 332 173 366
rect 217 406 396 424
rect 217 372 346 406
rect 380 372 396 406
rect 217 356 396 372
rect 443 361 509 458
rect 720 479 736 510
rect 956 534 1022 649
rect 956 500 972 534
rect 1006 500 1022 534
rect 1171 526 1223 547
rect 1171 492 1174 526
rect 1208 492 1223 526
rect 720 476 929 479
rect 686 470 929 476
rect 686 468 940 470
rect 686 466 944 468
rect 1171 466 1223 492
rect 686 439 1223 466
rect 1257 526 1314 547
rect 1257 492 1264 526
rect 1298 492 1314 526
rect 1257 489 1314 492
rect 1445 526 1479 649
rect 1659 580 1725 649
rect 1257 447 1411 489
rect 1445 476 1479 492
rect 1515 526 1590 547
rect 1515 492 1535 526
rect 1569 492 1590 526
rect 781 434 1223 439
rect 107 298 123 332
rect 157 316 173 332
rect 443 327 459 361
rect 493 327 509 361
rect 443 316 509 327
rect 560 355 647 430
rect 560 321 576 355
rect 610 321 647 355
rect 157 298 409 316
rect 560 305 647 321
rect 681 389 747 405
rect 681 355 697 389
rect 731 355 747 389
rect 681 350 747 355
rect 681 321 703 350
rect 107 282 409 298
rect 681 287 697 321
rect 737 316 747 350
rect 731 287 747 316
rect 23 237 324 248
rect 23 210 274 237
rect 23 147 89 210
rect 258 203 274 210
rect 308 203 324 237
rect 258 187 324 203
rect 375 241 510 282
rect 681 271 747 287
rect 375 207 460 241
rect 494 207 510 241
rect 781 237 815 434
rect 932 432 1223 434
rect 1377 442 1411 447
rect 1515 442 1590 492
rect 1659 546 1675 580
rect 1709 546 1725 580
rect 1659 512 1725 546
rect 1659 478 1675 512
rect 1709 478 1725 512
rect 1659 462 1725 478
rect 1759 580 1913 596
rect 1759 546 1775 580
rect 1809 546 1862 580
rect 1896 546 1913 580
rect 1759 512 1913 546
rect 1759 478 1775 512
rect 1809 478 1862 512
rect 1896 478 1913 512
rect 1377 428 1590 442
rect 1759 444 1913 478
rect 1759 428 1775 444
rect 851 398 920 400
rect 1299 398 1343 413
rect 851 364 882 398
rect 916 364 1006 398
rect 969 321 1006 364
rect 1046 364 1062 398
rect 1096 397 1343 398
rect 1096 364 1309 397
rect 1046 363 1309 364
rect 1046 355 1343 363
rect 1085 347 1343 355
rect 1377 408 1704 428
rect 855 294 935 310
rect 855 260 871 294
rect 905 260 935 294
rect 855 242 935 260
rect 969 299 1051 321
rect 969 265 1017 299
rect 969 247 1051 265
rect 1085 293 1135 347
rect 1085 253 1299 293
rect 375 191 510 207
rect 544 203 815 237
rect 969 208 1033 247
rect 1085 217 1135 253
rect 23 113 39 147
rect 73 113 89 147
rect 23 84 89 113
rect 123 147 189 176
rect 544 153 578 203
rect 123 113 139 147
rect 173 113 189 147
rect 123 17 189 113
rect 233 132 299 153
rect 233 98 249 132
rect 283 98 299 132
rect 391 119 435 153
rect 469 119 578 153
rect 612 140 678 169
rect 233 85 299 98
rect 612 106 628 140
rect 662 106 678 140
rect 781 140 815 203
rect 849 174 865 208
rect 899 174 1033 208
rect 1069 215 1135 217
rect 1069 181 1085 215
rect 1119 181 1135 215
rect 1069 174 1135 181
rect 1181 190 1231 219
rect 1181 156 1197 190
rect 1181 140 1231 156
rect 781 106 1231 140
rect 1265 109 1299 253
rect 1377 219 1411 408
rect 1529 394 1704 408
rect 1445 358 1495 374
rect 1479 324 1495 358
rect 1445 260 1495 324
rect 1537 350 1607 360
rect 1537 344 1567 350
rect 1537 310 1553 344
rect 1601 316 1607 350
rect 1587 310 1607 316
rect 1537 294 1607 310
rect 1645 344 1704 394
rect 1645 310 1661 344
rect 1695 310 1704 344
rect 1645 294 1704 310
rect 1738 410 1775 428
rect 1809 410 1862 444
rect 1896 410 1913 444
rect 1738 394 1913 410
rect 1947 580 2013 596
rect 1947 546 1963 580
rect 1997 546 2013 580
rect 1947 512 2013 546
rect 2121 580 2242 649
rect 2121 546 2164 580
rect 2198 546 2242 580
rect 2121 530 2242 546
rect 2276 567 2342 596
rect 2276 533 2292 567
rect 2326 533 2342 567
rect 1947 478 1952 512
rect 1986 478 2013 512
rect 2276 492 2342 533
rect 2376 578 2442 649
rect 2376 544 2392 578
rect 2426 544 2442 578
rect 2376 526 2442 544
rect 2488 580 2559 596
rect 2488 546 2504 580
rect 2538 546 2559 580
rect 1947 444 2013 478
rect 1947 410 1952 444
rect 1986 410 2013 444
rect 2087 460 2447 492
rect 2087 426 2103 460
rect 2137 458 2447 460
rect 2087 410 2137 426
rect 1738 260 1772 394
rect 1947 376 2013 410
rect 2171 390 2379 424
rect 2171 376 2205 390
rect 1806 344 1870 360
rect 1806 310 1814 344
rect 1848 310 1870 344
rect 1947 342 2205 376
rect 2239 350 2279 356
rect 1806 308 1870 310
rect 2273 316 2279 350
rect 2239 308 2279 316
rect 1806 295 2079 308
rect 1806 294 2029 295
rect 1836 274 2029 294
rect 2013 261 2029 274
rect 2063 261 2079 295
rect 1445 226 1724 260
rect 1758 226 1802 260
rect 2013 245 2079 261
rect 2199 292 2279 308
rect 2199 258 2215 292
rect 2249 258 2279 292
rect 2199 242 2279 258
rect 2313 298 2379 390
rect 2313 264 2329 298
rect 2363 264 2379 298
rect 1899 230 1965 240
rect 1333 195 1411 219
rect 1333 161 1334 195
rect 1368 161 1411 195
rect 1899 196 1915 230
rect 1949 196 1965 230
rect 2313 230 2379 264
rect 2313 208 2329 230
rect 1899 192 1965 196
rect 1333 145 1411 161
rect 1499 158 1965 192
rect 1999 196 2329 208
rect 2363 196 2379 230
rect 1999 174 2379 196
rect 1499 109 1544 158
rect 1999 124 2033 174
rect 2413 140 2447 458
rect 612 85 678 106
rect 233 51 678 85
rect 1265 85 1544 109
rect 715 38 747 72
rect 781 38 813 72
rect 715 17 813 38
rect 961 38 980 72
rect 1014 38 1033 72
rect 1265 51 1281 85
rect 1315 51 1544 85
rect 1578 90 1594 124
rect 1628 90 1644 124
rect 961 17 1033 38
rect 1578 17 1644 90
rect 1838 108 2033 124
rect 1838 74 1854 108
rect 1888 74 1982 108
rect 2016 74 2033 108
rect 1838 58 2033 74
rect 2146 120 2240 136
rect 2146 86 2176 120
rect 2210 86 2240 120
rect 2338 106 2375 140
rect 2409 106 2447 140
rect 2338 90 2447 106
rect 2488 470 2559 546
rect 2488 436 2504 470
rect 2538 436 2559 470
rect 2488 337 2559 436
rect 2595 580 2661 649
rect 2595 546 2611 580
rect 2645 546 2661 580
rect 2595 497 2661 546
rect 2595 463 2611 497
rect 2645 463 2661 497
rect 2595 414 2661 463
rect 2595 380 2611 414
rect 2645 380 2661 414
rect 2595 364 2661 380
rect 2695 580 2761 596
rect 2695 546 2711 580
rect 2745 546 2761 580
rect 2695 497 2761 546
rect 2695 463 2711 497
rect 2745 463 2761 497
rect 2695 414 2761 463
rect 2695 380 2711 414
rect 2745 380 2761 414
rect 2488 321 2562 337
rect 2488 287 2512 321
rect 2546 287 2562 321
rect 2488 271 2562 287
rect 2488 146 2559 271
rect 2488 112 2509 146
rect 2543 112 2559 146
rect 2146 17 2240 86
rect 2488 70 2559 112
rect 2595 210 2661 226
rect 2595 176 2625 210
rect 2659 176 2661 210
rect 2595 128 2661 176
rect 2595 94 2611 128
rect 2645 94 2661 128
rect 2595 17 2661 94
rect 2695 210 2761 380
rect 2695 176 2711 210
rect 2745 176 2761 210
rect 2695 120 2761 176
rect 2695 86 2711 120
rect 2745 86 2761 120
rect 2695 70 2761 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 703 321 737 350
rect 703 316 731 321
rect 731 316 737 321
rect 1567 344 1601 350
rect 1567 316 1587 344
rect 1587 316 1601 344
rect 2239 316 2273 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
<< metal1 >>
rect 0 683 2784 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 0 617 2784 649
rect 691 350 749 356
rect 691 316 703 350
rect 737 347 749 350
rect 1555 350 1613 356
rect 1555 347 1567 350
rect 737 319 1567 347
rect 737 316 749 319
rect 691 310 749 316
rect 1555 316 1567 319
rect 1601 347 1613 350
rect 2227 350 2285 356
rect 2227 347 2239 350
rect 1601 319 2239 347
rect 1601 316 1613 319
rect 1555 310 1613 316
rect 2227 316 2239 319
rect 2273 316 2285 350
rect 2227 310 2285 316
rect 0 17 2784 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
rect 0 -49 2784 -17
<< labels >>
flabel comment s 1182 290 1182 290 0 FreeSans 300 0 0 0 no_jumper_check
flabel comment s 1114 630 1114 630 0 FreeSans 300 0 0 0 no_jumper_check
rlabel comment s 0 0 0 0 4 sdfrtn_1
flabel pwell s 0 0 2784 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 0 617 2784 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 703 316 737 350 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew
flabel metal1 s 0 617 2784 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 2784 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 2719 94 2753 128 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2719 168 2753 202 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2719 242 2753 276 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2719 316 2753 350 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2719 390 2753 424 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2719 464 2753 498 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2719 538 2753 572 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 895 242 929 276 0 FreeSans 340 0 0 0 CLK_N
port 1 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 SCD
port 4 nsew
flabel corelocali s 607 390 641 424 0 FreeSans 340 0 0 0 SCD
port 4 nsew
flabel corelocali s 415 242 449 276 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 223 390 257 424 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 319 390 353 424 0 FreeSans 340 0 0 0 D
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 2784 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 140548
string GDS_START 119354
<< end >>
