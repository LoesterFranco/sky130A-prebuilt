magic
tech sky130A
magscale 1 2
timestamp 1599588209
<< nwell >>
rect -38 332 710 704
<< pwell >>
rect 0 0 672 49
<< scpmos >>
rect 88 368 118 592
rect 226 368 256 568
rect 310 368 340 568
rect 412 368 442 568
rect 520 368 550 536
<< nmoslvt >>
rect 84 74 114 222
rect 200 94 230 222
rect 301 94 331 222
rect 445 94 475 222
rect 544 94 574 222
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 210 200 222
rect 114 176 139 210
rect 173 176 200 210
rect 114 120 200 176
rect 114 86 139 120
rect 173 94 200 120
rect 230 210 301 222
rect 230 176 241 210
rect 275 176 301 210
rect 230 140 301 176
rect 230 106 241 140
rect 275 106 301 140
rect 230 94 301 106
rect 331 140 445 222
rect 331 106 372 140
rect 406 106 445 140
rect 331 94 445 106
rect 475 210 544 222
rect 475 176 499 210
rect 533 176 544 210
rect 475 140 544 176
rect 475 106 499 140
rect 533 106 544 140
rect 475 94 544 106
rect 574 210 645 222
rect 574 176 599 210
rect 633 176 645 210
rect 574 140 645 176
rect 574 106 599 140
rect 633 106 645 140
rect 574 94 645 106
rect 173 86 185 94
rect 114 74 185 86
<< pdiff >>
rect 29 580 88 592
rect 29 546 41 580
rect 75 546 88 580
rect 29 497 88 546
rect 29 463 41 497
rect 75 463 88 497
rect 29 414 88 463
rect 29 380 41 414
rect 75 380 88 414
rect 29 368 88 380
rect 118 580 187 592
rect 118 546 141 580
rect 175 568 187 580
rect 175 546 226 568
rect 118 499 226 546
rect 118 465 168 499
rect 202 465 226 499
rect 118 368 226 465
rect 256 368 310 568
rect 340 368 412 568
rect 442 560 501 568
rect 442 526 455 560
rect 489 536 501 560
rect 489 526 520 536
rect 442 492 520 526
rect 442 458 455 492
rect 489 458 520 492
rect 442 424 520 458
rect 442 390 455 424
rect 489 390 520 424
rect 442 368 520 390
rect 550 508 645 536
rect 550 474 563 508
rect 597 474 645 508
rect 550 368 645 474
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 139 176 173 210
rect 139 86 173 120
rect 241 176 275 210
rect 241 106 275 140
rect 372 106 406 140
rect 499 176 533 210
rect 499 106 533 140
rect 599 176 633 210
rect 599 106 633 140
<< pdiffc >>
rect 41 546 75 580
rect 41 463 75 497
rect 41 380 75 414
rect 141 546 175 580
rect 168 465 202 499
rect 455 526 489 560
rect 455 458 489 492
rect 455 390 489 424
rect 563 474 597 508
<< poly >>
rect 88 592 118 618
rect 226 568 256 594
rect 310 568 340 594
rect 412 568 442 594
rect 520 536 550 562
rect 88 353 118 368
rect 226 353 256 368
rect 310 353 340 368
rect 412 353 442 368
rect 520 353 550 368
rect 85 330 121 353
rect 223 336 259 353
rect 84 314 151 330
rect 84 280 101 314
rect 135 280 151 314
rect 84 264 151 280
rect 193 320 259 336
rect 307 326 343 353
rect 409 336 445 353
rect 517 336 553 353
rect 193 286 209 320
rect 243 286 259 320
rect 193 270 259 286
rect 301 310 367 326
rect 301 276 317 310
rect 351 276 367 310
rect 84 222 114 264
rect 200 222 230 270
rect 301 260 367 276
rect 409 320 475 336
rect 409 286 425 320
rect 459 286 475 320
rect 409 270 475 286
rect 517 320 583 336
rect 517 286 533 320
rect 567 286 583 320
rect 517 270 583 286
rect 301 222 331 260
rect 445 222 475 270
rect 544 222 574 270
rect 84 48 114 74
rect 200 68 230 94
rect 301 68 331 94
rect 445 68 475 94
rect 544 68 574 94
<< polycont >>
rect 101 280 135 314
rect 209 286 243 320
rect 317 276 351 310
rect 425 286 459 320
rect 533 286 567 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 17 580 91 596
rect 17 546 41 580
rect 75 546 91 580
rect 17 497 91 546
rect 17 463 41 497
rect 75 463 91 497
rect 17 414 91 463
rect 125 580 218 649
rect 125 546 141 580
rect 175 546 218 580
rect 125 499 218 546
rect 125 465 168 499
rect 202 465 218 499
rect 125 458 218 465
rect 439 560 505 576
rect 439 526 455 560
rect 489 526 505 560
rect 439 492 505 526
rect 439 458 455 492
rect 489 458 505 492
rect 547 508 610 649
rect 547 474 563 508
rect 597 474 610 508
rect 547 458 610 474
rect 439 424 505 458
rect 17 380 41 414
rect 75 380 91 414
rect 17 364 91 380
rect 125 390 455 424
rect 489 390 651 424
rect 17 226 51 364
rect 125 330 159 390
rect 85 314 159 330
rect 85 280 101 314
rect 135 280 159 314
rect 85 264 159 280
rect 193 320 263 356
rect 193 286 209 320
rect 243 286 263 320
rect 193 270 263 286
rect 301 310 367 356
rect 301 276 317 310
rect 351 276 367 310
rect 301 260 367 276
rect 409 320 475 356
rect 409 286 425 320
rect 459 286 475 320
rect 409 270 475 286
rect 509 320 583 356
rect 509 286 533 320
rect 567 286 583 320
rect 509 270 583 286
rect 617 226 651 390
rect 17 210 89 226
rect 17 176 39 210
rect 73 176 89 210
rect 17 120 89 176
rect 17 86 39 120
rect 73 86 89 120
rect 17 70 89 86
rect 123 210 189 226
rect 123 176 139 210
rect 173 176 189 210
rect 123 120 189 176
rect 123 86 139 120
rect 173 86 189 120
rect 225 210 549 226
rect 225 176 241 210
rect 275 192 499 210
rect 275 176 292 192
rect 225 140 292 176
rect 483 176 499 192
rect 533 176 549 210
rect 225 106 241 140
rect 275 106 292 140
rect 225 90 292 106
rect 353 140 426 156
rect 353 106 372 140
rect 406 106 426 140
rect 123 17 189 86
rect 353 17 426 106
rect 483 140 549 176
rect 483 106 499 140
rect 533 106 549 140
rect 483 90 549 106
rect 583 210 651 226
rect 583 176 599 210
rect 633 176 651 210
rect 583 140 651 176
rect 583 106 599 140
rect 633 106 651 140
rect 583 90 651 106
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o31a_1
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 B1
port 4 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 672 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1369902
string GDS_START 1363536
<< end >>
