magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 141 330 175 596
rect 305 330 371 596
rect 631 387 839 430
rect 631 353 665 387
rect 805 354 839 387
rect 141 282 371 330
rect 25 236 371 282
rect 605 287 665 353
rect 699 287 765 353
rect 805 288 931 354
rect 1081 290 1223 356
rect 25 228 503 236
rect 281 202 503 228
rect 281 96 331 202
rect 453 96 503 202
rect 991 101 1025 134
rect 991 51 1064 101
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 35 380 101 649
rect 215 364 265 649
rect 411 370 461 649
rect 495 596 703 615
rect 495 581 883 596
rect 495 336 529 581
rect 563 498 597 547
rect 637 532 883 581
rect 923 498 973 596
rect 563 464 973 498
rect 563 388 597 464
rect 923 424 973 464
rect 1007 458 1102 649
rect 1136 424 1186 596
rect 1226 458 1292 649
rect 1332 424 1382 596
rect 923 390 1382 424
rect 923 388 973 390
rect 1332 388 1382 390
rect 405 270 571 336
rect 537 253 571 270
rect 1145 253 1211 255
rect 537 219 1211 253
rect 195 17 245 194
rect 367 17 417 168
rect 726 200 792 219
rect 1145 203 1211 219
rect 539 17 605 185
rect 828 166 871 185
rect 640 116 871 166
rect 907 17 957 185
rect 1247 169 1281 255
rect 1059 135 1281 169
rect 1247 119 1281 135
rect 1317 17 1383 255
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 683 1440 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 0 617 1440 649
rect 0 17 1440 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -49 1440 -17
<< labels >>
rlabel locali s 1081 290 1223 356 6 A1
port 1 nsew signal input
rlabel locali s 991 101 1025 134 6 A2
port 2 nsew signal input
rlabel locali s 991 51 1064 101 6 A2
port 2 nsew signal input
rlabel locali s 699 287 765 353 6 B1
port 3 nsew signal input
rlabel locali s 805 354 839 387 6 B2
port 4 nsew signal input
rlabel locali s 805 288 931 354 6 B2
port 4 nsew signal input
rlabel locali s 631 387 839 430 6 B2
port 4 nsew signal input
rlabel locali s 631 353 665 387 6 B2
port 4 nsew signal input
rlabel locali s 605 287 665 353 6 B2
port 4 nsew signal input
rlabel locali s 453 96 503 202 6 X
port 5 nsew signal output
rlabel locali s 305 330 371 596 6 X
port 5 nsew signal output
rlabel locali s 281 202 503 228 6 X
port 5 nsew signal output
rlabel locali s 281 96 331 202 6 X
port 5 nsew signal output
rlabel locali s 141 330 175 596 6 X
port 5 nsew signal output
rlabel locali s 141 282 371 330 6 X
port 5 nsew signal output
rlabel locali s 25 236 371 282 6 X
port 5 nsew signal output
rlabel locali s 25 228 503 236 6 X
port 5 nsew signal output
rlabel metal1 s 0 -49 1440 49 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1440 715 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1440 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3540226
string GDS_START 3528918
<< end >>
