magic
tech sky130A
magscale 1 2
timestamp 1599588232
<< locali >>
rect 217 364 481 444
rect 85 238 167 310
rect 217 230 263 364
rect 583 270 649 356
rect 793 294 1031 360
rect 1369 294 1436 360
rect 217 196 508 230
rect 217 70 294 196
rect 442 70 508 196
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 17 512 89 572
rect 130 546 205 649
rect 319 546 391 649
rect 527 546 596 649
rect 744 546 810 649
rect 1036 546 1106 649
rect 1220 546 1286 649
rect 1400 546 1513 649
rect 17 478 1504 512
rect 17 364 89 478
rect 515 394 1376 444
rect 515 390 703 394
rect 17 204 51 364
rect 515 330 549 390
rect 1130 388 1216 394
rect 297 264 549 330
rect 1182 260 1216 388
rect 1250 294 1335 360
rect 1301 260 1335 294
rect 1470 260 1504 478
rect 692 236 1095 260
rect 17 90 81 204
rect 117 17 183 204
rect 660 226 1095 236
rect 1182 226 1267 260
rect 1301 226 1504 260
rect 334 17 400 162
rect 542 17 608 226
rect 660 121 726 226
rect 762 158 1025 192
rect 762 126 821 158
rect 857 17 923 124
rect 959 121 1025 158
rect 1061 85 1095 226
rect 1131 153 1181 192
rect 1216 187 1267 226
rect 1325 153 1391 187
rect 1131 119 1391 153
rect 1433 85 1499 192
rect 1061 51 1499 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
rlabel locali s 85 238 167 310 6 A_N
port 1 nsew signal input
rlabel locali s 1369 294 1436 360 6 B
port 2 nsew signal input
rlabel locali s 583 270 649 356 6 C
port 3 nsew signal input
rlabel locali s 793 294 1031 360 6 D
port 4 nsew signal input
rlabel locali s 442 70 508 196 6 X
port 5 nsew signal output
rlabel locali s 217 364 481 444 6 X
port 5 nsew signal output
rlabel locali s 217 230 263 364 6 X
port 5 nsew signal output
rlabel locali s 217 196 508 230 6 X
port 5 nsew signal output
rlabel locali s 217 70 294 196 6 X
port 5 nsew signal output
rlabel metal1 s 0 -49 1536 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 7 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 617 1536 715 6 VPWR
port 9 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1536 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3345956
string GDS_START 3334714
<< end >>
