magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 97 93 127 177
rect 186 93 216 177
rect 394 47 424 177
rect 490 47 520 177
rect 594 47 624 177
rect 678 47 708 177
<< pmoshvt >>
rect 81 410 117 494
rect 188 297 224 381
rect 386 297 422 497
rect 482 297 518 497
rect 586 297 622 497
rect 680 297 716 497
<< ndiff >>
rect 35 149 97 177
rect 35 115 43 149
rect 77 115 97 149
rect 35 93 97 115
rect 127 149 186 177
rect 127 115 141 149
rect 175 115 186 149
rect 127 93 186 115
rect 216 149 277 177
rect 216 115 235 149
rect 269 115 277 149
rect 216 93 277 115
rect 332 93 394 177
rect 332 59 340 93
rect 374 59 394 93
rect 332 47 394 59
rect 424 116 490 177
rect 424 82 434 116
rect 468 82 490 116
rect 424 47 490 82
rect 520 95 594 177
rect 520 61 534 95
rect 568 61 594 95
rect 520 47 594 61
rect 624 116 678 177
rect 624 82 634 116
rect 668 82 678 116
rect 624 47 678 82
rect 708 163 770 177
rect 708 129 728 163
rect 762 129 770 163
rect 708 95 770 129
rect 708 61 728 95
rect 762 61 770 95
rect 708 47 770 61
<< pdiff >>
rect 27 475 81 494
rect 27 441 35 475
rect 69 441 81 475
rect 27 410 81 441
rect 117 482 171 494
rect 117 448 129 482
rect 163 448 171 482
rect 117 410 171 448
rect 134 381 171 410
rect 332 425 386 497
rect 332 391 340 425
rect 374 391 386 425
rect 134 297 188 381
rect 224 343 278 381
rect 224 309 236 343
rect 270 309 278 343
rect 224 297 278 309
rect 332 297 386 391
rect 422 297 482 497
rect 518 297 586 497
rect 622 297 680 497
rect 716 485 770 497
rect 716 451 728 485
rect 762 451 770 485
rect 716 417 770 451
rect 716 383 728 417
rect 762 383 770 417
rect 716 297 770 383
<< ndiffc >>
rect 43 115 77 149
rect 141 115 175 149
rect 235 115 269 149
rect 340 59 374 93
rect 434 82 468 116
rect 534 61 568 95
rect 634 82 668 116
rect 728 129 762 163
rect 728 61 762 95
<< pdiffc >>
rect 35 441 69 475
rect 129 448 163 482
rect 340 391 374 425
rect 236 309 270 343
rect 728 451 762 485
rect 728 383 762 417
<< poly >>
rect 81 494 117 520
rect 386 497 422 523
rect 482 497 518 523
rect 586 497 622 523
rect 680 497 716 523
rect 81 395 117 410
rect 79 265 119 395
rect 188 381 224 407
rect 188 282 224 297
rect 386 282 422 297
rect 482 282 518 297
rect 586 282 622 297
rect 680 282 716 297
rect 186 265 226 282
rect 384 265 424 282
rect 480 265 520 282
rect 584 265 624 282
rect 79 249 133 265
rect 79 215 89 249
rect 123 215 133 249
rect 79 199 133 215
rect 186 249 244 265
rect 186 215 200 249
rect 234 215 244 249
rect 186 199 244 215
rect 314 249 424 265
rect 314 215 324 249
rect 358 215 424 249
rect 314 199 424 215
rect 466 249 520 265
rect 466 215 476 249
rect 510 215 520 249
rect 466 199 520 215
rect 570 249 624 265
rect 570 215 580 249
rect 614 215 624 249
rect 570 199 624 215
rect 97 177 127 199
rect 186 177 216 199
rect 394 177 424 199
rect 490 177 520 199
rect 594 177 624 199
rect 678 265 718 282
rect 678 249 732 265
rect 678 215 688 249
rect 722 215 732 249
rect 678 199 732 215
rect 678 177 708 199
rect 97 67 127 93
rect 186 67 216 93
rect 394 21 424 47
rect 490 21 520 47
rect 594 21 624 47
rect 678 21 708 47
<< polycont >>
rect 89 215 123 249
rect 200 215 234 249
rect 324 215 358 249
rect 476 215 510 249
rect 580 215 614 249
rect 688 215 722 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 17 475 69 491
rect 17 441 35 475
rect 103 482 179 527
rect 103 448 129 482
rect 163 448 179 482
rect 227 459 523 493
rect 702 485 798 527
rect 17 414 69 441
rect 227 414 261 459
rect 17 377 261 414
rect 315 391 340 425
rect 374 391 442 425
rect 17 165 52 377
rect 86 249 166 339
rect 220 309 236 343
rect 270 309 358 343
rect 220 305 358 309
rect 86 215 89 249
rect 123 215 166 249
rect 86 199 166 215
rect 200 249 268 265
rect 234 215 268 249
rect 200 199 268 215
rect 324 249 358 305
rect 324 165 358 215
rect 17 149 81 165
rect 17 115 43 149
rect 77 115 81 149
rect 17 90 81 115
rect 141 149 175 165
rect 141 17 175 115
rect 235 149 358 165
rect 269 131 358 149
rect 392 165 442 391
rect 476 249 523 459
rect 510 215 523 249
rect 476 199 523 215
rect 564 249 626 482
rect 702 451 728 485
rect 762 451 798 485
rect 702 417 798 451
rect 702 383 728 417
rect 762 383 798 417
rect 702 375 798 383
rect 564 215 580 249
rect 614 215 626 249
rect 564 199 626 215
rect 672 249 733 341
rect 672 215 688 249
rect 722 215 733 249
rect 672 199 733 215
rect 392 131 668 165
rect 235 90 269 115
rect 434 116 474 131
rect 324 93 390 96
rect 324 59 340 93
rect 374 59 390 93
rect 468 82 474 116
rect 628 116 668 131
rect 434 60 474 82
rect 518 95 584 97
rect 518 61 534 95
rect 568 61 584 95
rect 628 82 634 116
rect 628 62 668 82
rect 702 163 798 165
rect 702 129 728 163
rect 762 129 798 163
rect 702 95 798 129
rect 324 17 390 59
rect 518 17 584 61
rect 702 61 728 95
rect 762 61 798 95
rect 702 17 798 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel corelocali s 688 221 722 255 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 132 289 166 323 0 FreeSans 400 0 0 0 C_N
port 3 nsew
flabel corelocali s 132 221 166 255 0 FreeSans 400 0 0 0 C_N
port 3 nsew
flabel corelocali s 231 238 231 238 0 FreeSans 400 0 0 0 D_N
port 4 nsew
flabel corelocali s 580 289 614 323 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel corelocali s 632 85 666 119 0 FreeSans 200 0 0 0 Y
port 9 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
rlabel comment s 0 0 0 0 4 nor4bb_1
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2537148
string GDS_START 2530660
<< end >>
