magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1472 561
rect 33 289 83 527
rect 201 425 251 527
rect 713 425 757 527
rect 885 425 933 527
rect 369 391 419 425
rect 537 391 587 425
rect 1387 425 1443 527
rect 369 357 783 391
rect 1051 391 1101 425
rect 1219 391 1269 425
rect 1051 357 1455 391
rect 749 323 783 357
rect 230 289 715 323
rect 749 289 825 323
rect 230 255 283 289
rect 17 215 283 255
rect 337 215 619 255
rect 655 249 715 289
rect 655 215 721 249
rect 125 17 159 111
rect 293 17 327 111
rect 461 17 495 111
rect 629 17 663 111
rect 791 164 825 289
rect 859 289 1387 323
rect 859 199 988 289
rect 1022 215 1292 255
rect 1343 199 1387 289
rect 1421 164 1455 357
rect 791 129 1455 164
rect 0 -17 1472 17
<< obsli1 >>
rect 117 391 167 493
rect 285 459 679 493
rect 285 391 335 459
rect 453 425 503 459
rect 621 425 679 459
rect 791 425 851 493
rect 967 459 1353 493
rect 117 357 335 391
rect 817 391 851 425
rect 967 391 1017 459
rect 1135 425 1185 459
rect 1303 427 1353 459
rect 817 357 1017 391
rect 117 289 167 357
rect 25 147 757 181
rect 25 145 259 147
rect 25 51 91 145
rect 193 51 259 145
rect 361 145 595 147
rect 361 51 427 145
rect 529 51 595 145
rect 697 95 757 147
rect 697 51 1449 95
<< metal1 >>
rect 0 496 1472 592
rect 0 -48 1472 48
<< labels >>
rlabel locali s 655 249 715 289 6 A1
port 1 nsew signal input
rlabel locali s 655 215 721 249 6 A1
port 1 nsew signal input
rlabel locali s 230 289 715 323 6 A1
port 1 nsew signal input
rlabel locali s 230 255 283 289 6 A1
port 1 nsew signal input
rlabel locali s 17 215 283 255 6 A1
port 1 nsew signal input
rlabel locali s 337 215 619 255 6 A2
port 2 nsew signal input
rlabel locali s 1343 199 1387 289 6 B1
port 3 nsew signal input
rlabel locali s 859 289 1387 323 6 B1
port 3 nsew signal input
rlabel locali s 859 199 988 289 6 B1
port 3 nsew signal input
rlabel locali s 1022 215 1292 255 6 B2
port 4 nsew signal input
rlabel locali s 1421 164 1455 357 6 Y
port 5 nsew signal output
rlabel locali s 1219 391 1269 425 6 Y
port 5 nsew signal output
rlabel locali s 1051 391 1101 425 6 Y
port 5 nsew signal output
rlabel locali s 1051 357 1455 391 6 Y
port 5 nsew signal output
rlabel locali s 791 164 825 289 6 Y
port 5 nsew signal output
rlabel locali s 791 129 1455 164 6 Y
port 5 nsew signal output
rlabel locali s 749 323 783 357 6 Y
port 5 nsew signal output
rlabel locali s 749 289 825 323 6 Y
port 5 nsew signal output
rlabel locali s 537 391 587 425 6 Y
port 5 nsew signal output
rlabel locali s 369 391 419 425 6 Y
port 5 nsew signal output
rlabel locali s 369 357 783 391 6 Y
port 5 nsew signal output
rlabel locali s 629 17 663 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 461 17 495 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 293 17 327 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 125 17 159 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 1472 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1472 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1387 425 1443 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 885 425 933 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 713 425 757 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 201 425 251 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 33 289 83 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 1472 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 1472 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1472 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1512612
string GDS_START 1502008
<< end >>
