magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 351 370 441 493
rect 20 145 65 265
rect 202 213 285 265
rect 405 163 441 370
rect 257 129 441 163
rect 257 51 327 129
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 83 336 135 381
rect 185 371 251 527
rect 83 302 371 336
rect 99 109 135 302
rect 327 197 371 302
rect 66 74 135 109
rect 181 17 223 179
rect 361 17 427 95
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
rlabel locali s 20 145 65 265 6 A
port 1 nsew signal input
rlabel locali s 202 213 285 265 6 SLEEP
port 2 nsew signal input
rlabel locali s 405 163 441 370 6 X
port 3 nsew signal output
rlabel locali s 351 370 441 493 6 X
port 3 nsew signal output
rlabel locali s 257 129 441 163 6 X
port 3 nsew signal output
rlabel locali s 257 51 327 129 6 X
port 3 nsew signal output
rlabel metal1 s 0 -48 460 48 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 496 460 592 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 460 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2614556
string GDS_START 2610158
<< end >>
