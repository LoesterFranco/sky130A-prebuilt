magic
tech sky130A
magscale 1 2
timestamp 1604502741
<< locali >>
rect 181 236 263 356
rect 297 286 363 356
rect 475 368 545 596
rect 511 234 545 368
rect 25 51 263 134
rect 436 162 551 234
rect 436 78 502 162
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 37 424 103 556
rect 137 458 203 649
rect 241 424 307 556
rect 375 458 441 649
rect 37 390 441 424
rect 37 268 103 390
rect 37 168 108 268
rect 407 334 441 390
rect 407 268 477 334
rect 579 364 645 649
rect 336 17 402 234
rect 585 128 649 234
rect 536 17 649 128
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel locali s 25 51 263 134 6 A
port 1 nsew signal input
rlabel locali s 181 236 263 356 6 B
port 2 nsew signal input
rlabel locali s 297 286 363 356 6 C
port 3 nsew signal input
rlabel locali s 511 234 545 368 6 X
port 4 nsew signal output
rlabel locali s 475 368 545 596 6 X
port 4 nsew signal output
rlabel locali s 436 162 551 234 6 X
port 4 nsew signal output
rlabel locali s 436 78 502 162 6 X
port 4 nsew signal output
rlabel metal1 s 0 -49 672 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 617 672 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3153546
string GDS_START 3147292
<< end >>
