magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 1050 582
<< pwell >>
rect 25 -17 59 17
<< scnmos >>
rect 100 47 130 177
rect 196 47 226 177
rect 282 47 312 177
rect 388 47 418 177
rect 578 47 608 177
rect 684 47 714 177
rect 770 47 800 177
rect 876 47 906 177
<< pmoshvt >>
rect 92 297 128 497
rect 188 297 224 497
rect 284 297 320 497
rect 380 297 416 497
rect 580 297 616 497
rect 676 297 712 497
rect 772 297 808 497
rect 868 297 904 497
<< ndiff >>
rect 37 135 100 177
rect 37 101 45 135
rect 79 101 100 135
rect 37 47 100 101
rect 130 169 196 177
rect 130 135 141 169
rect 175 135 196 169
rect 130 101 196 135
rect 130 67 141 101
rect 175 67 196 101
rect 130 47 196 67
rect 226 93 282 177
rect 226 59 237 93
rect 271 59 282 93
rect 226 47 282 59
rect 312 168 388 177
rect 312 134 333 168
rect 367 134 388 168
rect 312 47 388 134
rect 418 93 471 177
rect 418 59 429 93
rect 463 59 471 93
rect 418 47 471 59
rect 525 93 578 177
rect 525 59 533 93
rect 567 59 578 93
rect 525 47 578 59
rect 608 168 684 177
rect 608 134 629 168
rect 663 134 684 168
rect 608 47 684 134
rect 714 124 770 177
rect 714 90 725 124
rect 759 90 770 124
rect 714 47 770 90
rect 800 89 876 177
rect 800 55 821 89
rect 855 55 876 89
rect 800 47 876 55
rect 906 127 959 177
rect 906 93 917 127
rect 951 93 959 127
rect 906 47 959 93
<< pdiff >>
rect 37 475 92 497
rect 37 441 45 475
rect 79 441 92 475
rect 37 407 92 441
rect 37 373 45 407
rect 79 373 92 407
rect 37 297 92 373
rect 128 407 188 497
rect 128 373 141 407
rect 175 373 188 407
rect 128 339 188 373
rect 128 305 141 339
rect 175 305 188 339
rect 128 297 188 305
rect 224 475 284 497
rect 224 441 237 475
rect 271 441 284 475
rect 224 407 284 441
rect 224 373 237 407
rect 271 373 284 407
rect 224 297 284 373
rect 320 415 380 497
rect 320 381 333 415
rect 367 381 380 415
rect 320 347 380 381
rect 320 313 333 347
rect 367 313 380 347
rect 320 297 380 313
rect 416 485 471 497
rect 416 451 429 485
rect 463 451 471 485
rect 416 417 471 451
rect 416 383 429 417
rect 463 383 471 417
rect 416 297 471 383
rect 525 485 580 497
rect 525 451 533 485
rect 567 451 580 485
rect 525 417 580 451
rect 525 383 533 417
rect 567 383 580 417
rect 525 297 580 383
rect 616 477 676 497
rect 616 443 629 477
rect 663 443 676 477
rect 616 409 676 443
rect 616 375 629 409
rect 663 375 676 409
rect 616 341 676 375
rect 616 307 629 341
rect 663 307 676 341
rect 616 297 676 307
rect 712 485 772 497
rect 712 451 725 485
rect 759 451 772 485
rect 712 417 772 451
rect 712 383 725 417
rect 759 383 772 417
rect 712 297 772 383
rect 808 477 868 497
rect 808 443 821 477
rect 855 443 868 477
rect 808 409 868 443
rect 808 375 821 409
rect 855 375 868 409
rect 808 341 868 375
rect 808 307 821 341
rect 855 307 868 341
rect 808 297 868 307
rect 904 485 959 497
rect 904 451 917 485
rect 951 451 959 485
rect 904 417 959 451
rect 904 383 917 417
rect 951 383 959 417
rect 904 297 959 383
<< ndiffc >>
rect 45 101 79 135
rect 141 135 175 169
rect 141 67 175 101
rect 237 59 271 93
rect 333 134 367 168
rect 429 59 463 93
rect 533 59 567 93
rect 629 134 663 168
rect 725 90 759 124
rect 821 55 855 89
rect 917 93 951 127
<< pdiffc >>
rect 45 441 79 475
rect 45 373 79 407
rect 141 373 175 407
rect 141 305 175 339
rect 237 441 271 475
rect 237 373 271 407
rect 333 381 367 415
rect 333 313 367 347
rect 429 451 463 485
rect 429 383 463 417
rect 533 451 567 485
rect 533 383 567 417
rect 629 443 663 477
rect 629 375 663 409
rect 629 307 663 341
rect 725 451 759 485
rect 725 383 759 417
rect 821 443 855 477
rect 821 375 855 409
rect 821 307 855 341
rect 917 451 951 485
rect 917 383 951 417
<< poly >>
rect 92 497 128 523
rect 188 497 224 523
rect 284 497 320 523
rect 380 497 416 523
rect 580 497 616 523
rect 676 497 712 523
rect 772 497 808 523
rect 868 497 904 523
rect 92 282 128 297
rect 188 282 224 297
rect 284 282 320 297
rect 380 282 416 297
rect 580 282 616 297
rect 676 282 712 297
rect 772 282 808 297
rect 868 282 904 297
rect 90 265 130 282
rect 186 265 226 282
rect 36 249 226 265
rect 36 215 46 249
rect 80 215 226 249
rect 36 199 226 215
rect 100 177 130 199
rect 196 177 226 199
rect 282 265 322 282
rect 378 265 418 282
rect 282 249 418 265
rect 282 215 333 249
rect 367 215 418 249
rect 282 199 418 215
rect 282 177 312 199
rect 388 177 418 199
rect 578 265 618 282
rect 674 265 714 282
rect 578 249 714 265
rect 578 215 596 249
rect 630 215 664 249
rect 698 215 714 249
rect 578 199 714 215
rect 578 177 608 199
rect 684 177 714 199
rect 770 265 810 282
rect 866 265 906 282
rect 770 249 906 265
rect 770 215 794 249
rect 828 215 862 249
rect 896 215 906 249
rect 770 199 906 215
rect 770 177 800 199
rect 876 177 906 199
rect 100 21 130 47
rect 196 21 226 47
rect 282 21 312 47
rect 388 21 418 47
rect 578 21 608 47
rect 684 21 714 47
rect 770 21 800 47
rect 876 21 906 47
<< polycont >>
rect 46 215 80 249
rect 333 215 367 249
rect 596 215 630 249
rect 664 215 698 249
rect 794 215 828 249
rect 862 215 896 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 29 485 483 491
rect 29 475 429 485
rect 29 441 45 475
rect 79 457 237 475
rect 79 441 81 457
rect 29 407 81 441
rect 235 441 237 457
rect 271 451 429 475
rect 463 451 483 485
rect 271 441 273 451
rect 29 373 45 407
rect 79 373 81 407
rect 29 357 81 373
rect 115 407 179 423
rect 115 373 141 407
rect 175 373 179 407
rect 115 339 179 373
rect 235 407 273 441
rect 427 417 483 451
rect 235 373 237 407
rect 271 373 273 407
rect 235 357 273 373
rect 307 381 333 415
rect 367 381 383 415
rect 20 249 81 323
rect 20 215 46 249
rect 80 215 81 249
rect 20 199 81 215
rect 115 305 141 339
rect 175 305 179 339
rect 307 347 383 381
rect 427 383 429 417
rect 463 383 483 417
rect 427 367 483 383
rect 527 485 573 527
rect 527 451 533 485
rect 567 451 573 485
rect 527 417 573 451
rect 527 383 533 417
rect 567 383 573 417
rect 527 367 573 383
rect 619 477 673 493
rect 619 443 629 477
rect 663 443 673 477
rect 619 409 673 443
rect 619 375 629 409
rect 663 375 673 409
rect 115 171 179 305
rect 213 257 257 323
rect 307 313 333 347
rect 367 331 383 347
rect 619 341 673 375
rect 719 485 765 527
rect 719 451 725 485
rect 759 451 765 485
rect 719 417 765 451
rect 719 383 725 417
rect 759 383 765 417
rect 719 367 765 383
rect 811 477 865 493
rect 811 443 821 477
rect 855 443 865 477
rect 811 409 865 443
rect 811 375 821 409
rect 855 375 865 409
rect 619 331 629 341
rect 367 313 629 331
rect 307 307 629 313
rect 663 331 673 341
rect 811 341 865 375
rect 911 485 957 527
rect 911 451 917 485
rect 951 451 957 485
rect 911 417 957 451
rect 911 383 917 417
rect 951 383 957 417
rect 911 367 957 383
rect 811 331 821 341
rect 663 307 821 331
rect 855 307 865 341
rect 307 291 865 307
rect 937 257 983 331
rect 213 249 387 257
rect 213 215 333 249
rect 367 215 387 249
rect 213 207 387 215
rect 562 249 714 257
rect 562 215 596 249
rect 630 215 664 249
rect 698 215 714 249
rect 562 207 714 215
rect 778 249 983 257
rect 778 215 794 249
rect 828 215 862 249
rect 896 215 983 249
rect 778 207 983 215
rect 115 169 679 171
rect 29 135 79 163
rect 29 101 45 135
rect 29 17 79 101
rect 115 135 141 169
rect 175 168 679 169
rect 175 135 333 168
rect 115 134 333 135
rect 367 134 629 168
rect 663 134 679 168
rect 115 131 679 134
rect 115 101 177 131
rect 115 67 141 101
rect 175 67 177 101
rect 725 127 967 171
rect 725 124 759 127
rect 115 51 177 67
rect 211 93 287 95
rect 211 59 237 93
rect 271 59 287 93
rect 211 17 287 59
rect 403 93 479 95
rect 403 59 429 93
rect 463 59 479 93
rect 403 17 479 59
rect 517 93 725 95
rect 517 59 533 93
rect 567 90 725 93
rect 951 93 967 127
rect 567 59 759 90
rect 517 53 759 59
rect 795 89 871 91
rect 795 55 821 89
rect 855 55 871 89
rect 795 17 871 55
rect 917 53 967 93
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
flabel corelocali s 937 221 971 255 0 FreeSans 200 0 0 0 A2
port 2 nsew
flabel corelocali s 25 221 59 255 0 FreeSans 200 0 0 0 C1
port 4 nsew
flabel corelocali s 25 289 59 323 0 FreeSans 200 0 0 0 C1
port 4 nsew
flabel corelocali s 318 238 318 238 0 FreeSans 200 0 0 0 B1
port 3 nsew
flabel corelocali s 117 289 151 323 0 FreeSans 200 0 0 0 Y
port 9 nsew
flabel corelocali s 117 349 151 391 0 FreeSans 200 0 0 0 Y
port 9 nsew
flabel corelocali s 117 221 151 255 0 FreeSans 200 0 0 0 Y
port 9 nsew
flabel corelocali s 117 153 151 187 0 FreeSans 200 0 0 0 Y
port 9 nsew
flabel corelocali s 117 85 151 119 0 FreeSans 200 0 0 0 Y
port 9 nsew
flabel corelocali s 577 221 611 255 0 FreeSans 200 0 0 0 A1
port 1 nsew
flabel corelocali s 944 289 978 323 0 FreeSans 200 0 0 0 A2
port 2 nsew
flabel corelocali s 646 238 646 238 0 FreeSans 200 0 0 0 A1
port 1 nsew
flabel corelocali s 215 221 249 255 0 FreeSans 200 0 0 0 B1
port 3 nsew
flabel corelocali s 834 238 834 238 0 FreeSans 200 0 0 0 A2
port 2 nsew
flabel corelocali s 215 289 249 323 0 FreeSans 200 0 0 0 B1
port 3 nsew
flabel metal1 s 25 527 59 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
flabel metal1 s 25 -17 59 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel nbase s 25 527 59 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel pwell s 25 -17 59 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
rlabel comment s 0 0 0 0 4 a211oi_2
<< properties >>
string FIXED_BBOX 0 0 1012 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1115742
string GDS_START 1106622
<< end >>
