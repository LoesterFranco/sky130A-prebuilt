magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 460 561
rect 220 367 254 527
rect 288 401 354 493
rect 388 435 422 527
rect 288 367 443 401
rect 30 153 69 265
rect 173 153 255 265
rect 357 165 443 367
rect 304 131 443 165
rect 21 17 69 119
rect 207 17 270 119
rect 304 77 338 131
rect 372 17 438 97
rect 0 -17 460 17
<< obsli1 >>
rect 31 333 103 368
rect 31 299 323 333
rect 103 119 139 299
rect 289 199 323 299
rect 103 51 161 119
<< metal1 >>
rect 0 496 460 592
rect 0 -48 460 48
<< labels >>
rlabel locali s 173 153 255 265 6 A
port 1 nsew signal input
rlabel locali s 30 153 69 265 6 B
port 2 nsew signal input
rlabel locali s 357 165 443 367 6 X
port 3 nsew signal output
rlabel locali s 304 131 443 165 6 X
port 3 nsew signal output
rlabel locali s 304 77 338 131 6 X
port 3 nsew signal output
rlabel locali s 288 401 354 493 6 X
port 3 nsew signal output
rlabel locali s 288 367 443 401 6 X
port 3 nsew signal output
rlabel locali s 372 17 438 97 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 207 17 270 119 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 21 17 69 119 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 460 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 460 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 388 435 422 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 220 367 254 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 460 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 460 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 460 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1003430
string GDS_START 999072
<< end >>
