magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 103 333 179 493
rect 291 333 367 493
rect 511 333 587 493
rect 789 333 865 493
rect 103 289 865 333
rect 22 215 179 255
rect 213 215 370 255
rect 487 215 676 255
rect 744 211 865 289
rect 923 215 989 255
rect 789 127 865 211
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 18 299 69 527
rect 223 367 257 527
rect 411 367 477 527
rect 659 367 735 527
rect 909 289 975 527
rect 18 147 257 181
rect 18 51 85 147
rect 129 17 163 109
rect 197 93 257 147
rect 291 127 677 181
rect 721 93 755 177
rect 909 93 975 181
rect 197 51 465 93
rect 503 51 975 93
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
rlabel locali s 923 215 989 255 6 A
port 1 nsew signal input
rlabel locali s 487 215 676 255 6 B
port 2 nsew signal input
rlabel locali s 213 215 370 255 6 C
port 3 nsew signal input
rlabel locali s 22 215 179 255 6 D
port 4 nsew signal input
rlabel locali s 789 333 865 493 6 Y
port 5 nsew signal output
rlabel locali s 789 127 865 211 6 Y
port 5 nsew signal output
rlabel locali s 744 211 865 289 6 Y
port 5 nsew signal output
rlabel locali s 511 333 587 493 6 Y
port 5 nsew signal output
rlabel locali s 291 333 367 493 6 Y
port 5 nsew signal output
rlabel locali s 103 333 179 493 6 Y
port 5 nsew signal output
rlabel locali s 103 289 865 333 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -48 1012 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 1012 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1012 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2301954
string GDS_START 2293066
<< end >>
