magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1196 561
rect 103 391 169 425
rect 119 325 153 391
rect 287 325 321 425
rect 454 451 588 527
rect 710 451 844 527
rect 953 451 1087 527
rect 29 257 65 325
rect 119 291 436 325
rect 29 215 165 257
rect 209 216 345 257
rect 235 215 301 216
rect 393 165 436 291
rect 483 215 644 325
rect 745 215 896 325
rect 943 215 1172 325
rect 119 17 153 109
rect 271 131 620 165
rect 911 17 978 93
rect 1112 17 1177 177
rect 0 -17 1196 17
<< obsli1 >>
rect 35 459 405 493
rect 35 359 69 459
rect 203 359 237 459
rect 371 417 405 459
rect 636 417 670 493
rect 878 417 912 493
rect 1127 417 1161 493
rect 371 383 1161 417
rect 371 359 405 383
rect 636 359 670 383
rect 878 359 912 383
rect 1127 359 1161 383
rect 35 143 237 177
rect 35 93 69 143
rect 19 59 85 93
rect 203 93 237 143
rect 724 127 1078 161
rect 187 59 423 93
rect 470 59 874 93
rect 1012 55 1078 127
<< metal1 >>
rect 0 496 1196 592
rect 0 -48 1196 48
<< labels >>
rlabel locali s 483 215 644 325 6 A1
port 1 nsew signal input
rlabel locali s 745 215 896 325 6 A2
port 2 nsew signal input
rlabel locali s 943 215 1172 325 6 A3
port 3 nsew signal input
rlabel locali s 235 215 301 216 6 B1
port 4 nsew signal input
rlabel locali s 209 216 345 257 6 B1
port 4 nsew signal input
rlabel locali s 29 257 65 325 6 B2
port 5 nsew signal input
rlabel locali s 29 215 165 257 6 B2
port 5 nsew signal input
rlabel locali s 393 165 436 291 6 Y
port 6 nsew signal output
rlabel locali s 287 325 321 425 6 Y
port 6 nsew signal output
rlabel locali s 271 131 620 165 6 Y
port 6 nsew signal output
rlabel locali s 119 325 153 391 6 Y
port 6 nsew signal output
rlabel locali s 119 291 436 325 6 Y
port 6 nsew signal output
rlabel locali s 103 391 169 425 6 Y
port 6 nsew signal output
rlabel locali s 1112 17 1177 177 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 911 17 978 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 119 17 153 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 1196 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1196 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 953 451 1087 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 710 451 844 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 454 451 588 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 1196 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 1196 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3658642
string GDS_START 3647408
<< end >>
