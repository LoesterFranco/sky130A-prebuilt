magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 815 393 857 425
rect 1099 393 1149 425
rect 815 359 1149 393
rect 1099 325 1149 359
rect 168 289 670 323
rect 168 257 202 289
rect 97 215 202 257
rect 636 257 670 289
rect 271 215 581 255
rect 636 215 861 257
rect 1099 283 1268 325
rect 1190 95 1268 283
rect 997 61 1268 95
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 17 393 80 493
rect 124 427 174 527
rect 218 393 268 493
rect 312 427 362 527
rect 406 393 456 493
rect 518 425 568 493
rect 612 427 662 527
rect 706 459 951 493
rect 706 425 771 459
rect 901 427 951 459
rect 1005 427 1055 527
rect 17 391 456 393
rect 17 357 756 391
rect 1193 359 1268 527
rect 17 179 63 357
rect 722 325 756 357
rect 722 291 1041 325
rect 1007 249 1041 291
rect 1007 215 1149 249
rect 17 129 182 179
rect 226 145 464 181
rect 226 95 276 145
rect 21 51 276 95
rect 320 17 354 111
rect 388 51 464 145
rect 526 17 560 181
rect 594 145 1151 181
rect 594 51 670 145
rect 714 17 748 111
rect 782 51 865 145
rect 1081 129 1151 145
rect 909 17 943 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< obsm1 >>
rect 521 456 579 465
rect 725 456 783 465
rect 521 428 783 456
rect 521 419 579 428
rect 725 419 783 428
<< labels >>
rlabel locali s 271 215 581 255 6 A
port 1 nsew signal input
rlabel locali s 636 257 670 289 6 B
port 2 nsew signal input
rlabel locali s 636 215 861 257 6 B
port 2 nsew signal input
rlabel locali s 168 289 670 323 6 B
port 2 nsew signal input
rlabel locali s 168 257 202 289 6 B
port 2 nsew signal input
rlabel locali s 97 215 202 257 6 B
port 2 nsew signal input
rlabel locali s 1190 95 1268 283 6 Y
port 3 nsew signal output
rlabel locali s 1099 393 1149 425 6 Y
port 3 nsew signal output
rlabel locali s 1099 325 1149 359 6 Y
port 3 nsew signal output
rlabel locali s 1099 283 1268 325 6 Y
port 3 nsew signal output
rlabel locali s 997 61 1268 95 6 Y
port 3 nsew signal output
rlabel locali s 815 393 857 425 6 Y
port 3 nsew signal output
rlabel locali s 815 359 1149 393 6 Y
port 3 nsew signal output
rlabel metal1 s 0 -48 1288 48 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 496 1288 592 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1288 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 695744
string GDS_START 686584
<< end >>
