magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 2246 704
<< pwell >>
rect 0 0 2208 49
<< scnmos >>
rect 84 74 114 222
rect 170 74 200 222
rect 270 74 300 222
rect 359 74 389 222
rect 456 74 486 222
rect 556 74 586 222
rect 656 74 686 222
rect 756 74 786 222
rect 856 74 886 222
rect 974 74 1004 222
rect 1073 74 1103 222
rect 1160 74 1190 222
rect 1329 74 1359 222
rect 1443 74 1473 222
rect 1529 74 1559 222
rect 1643 74 1673 222
rect 1743 74 1773 222
rect 1843 74 1873 222
rect 1929 74 1959 222
rect 2029 74 2059 222
<< pmoshvt >>
rect 86 368 116 592
rect 176 368 206 592
rect 266 368 296 592
rect 356 368 386 592
rect 446 368 476 592
rect 536 368 566 592
rect 626 368 656 592
rect 718 368 748 592
rect 920 368 950 592
rect 1010 368 1040 592
rect 1100 368 1130 592
rect 1190 368 1220 592
rect 1300 368 1330 592
rect 1390 368 1420 592
rect 1490 368 1520 592
rect 1590 368 1620 592
rect 1802 368 1832 592
rect 1892 368 1922 592
rect 2002 368 2032 592
rect 2092 368 2122 592
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 189 170 222
rect 114 155 125 189
rect 159 155 170 189
rect 114 74 170 155
rect 200 144 270 222
rect 200 110 225 144
rect 259 110 270 144
rect 200 74 270 110
rect 300 189 359 222
rect 300 155 311 189
rect 345 155 359 189
rect 300 74 359 155
rect 389 144 456 222
rect 389 110 411 144
rect 445 110 456 144
rect 389 74 456 110
rect 486 189 556 222
rect 486 155 511 189
rect 545 155 556 189
rect 486 74 556 155
rect 586 144 656 222
rect 586 110 611 144
rect 645 110 656 144
rect 586 74 656 110
rect 686 189 756 222
rect 686 155 711 189
rect 745 155 756 189
rect 686 74 756 155
rect 786 144 856 222
rect 786 110 811 144
rect 845 110 856 144
rect 786 74 856 110
rect 886 100 974 222
rect 886 74 913 100
rect 901 66 913 74
rect 947 74 974 100
rect 1004 184 1073 222
rect 1004 150 1015 184
rect 1049 150 1073 184
rect 1004 116 1073 150
rect 1004 82 1015 116
rect 1049 82 1073 116
rect 1004 74 1073 82
rect 1103 116 1160 222
rect 1103 82 1115 116
rect 1149 82 1160 116
rect 1103 74 1160 82
rect 1190 197 1329 222
rect 1190 184 1284 197
rect 1190 150 1215 184
rect 1249 163 1284 184
rect 1318 163 1329 197
rect 1249 150 1329 163
rect 1190 116 1329 150
rect 1190 82 1242 116
rect 1276 82 1329 116
rect 1190 74 1329 82
rect 1359 136 1443 222
rect 1359 102 1384 136
rect 1418 102 1443 136
rect 1359 74 1443 102
rect 1473 210 1529 222
rect 1473 176 1484 210
rect 1518 176 1529 210
rect 1473 120 1529 176
rect 1473 86 1484 120
rect 1518 86 1529 120
rect 1473 74 1529 86
rect 1559 136 1643 222
rect 1559 102 1584 136
rect 1618 102 1643 136
rect 1559 74 1643 102
rect 1673 210 1743 222
rect 1673 176 1684 210
rect 1718 176 1743 210
rect 1673 120 1743 176
rect 1673 86 1684 120
rect 1718 86 1743 120
rect 1673 74 1743 86
rect 1773 136 1843 222
rect 1773 102 1784 136
rect 1818 102 1843 136
rect 1773 74 1843 102
rect 1873 210 1929 222
rect 1873 176 1884 210
rect 1918 176 1929 210
rect 1873 120 1929 176
rect 1873 86 1884 120
rect 1918 86 1929 120
rect 1873 74 1929 86
rect 1959 136 2029 222
rect 1959 102 1984 136
rect 2018 102 2029 136
rect 1959 74 2029 102
rect 2059 210 2130 222
rect 2059 176 2084 210
rect 2118 176 2130 210
rect 2059 120 2130 176
rect 2059 86 2084 120
rect 2118 86 2130 120
rect 2059 74 2130 86
rect 947 66 959 74
rect 901 54 959 66
rect 1205 70 1314 74
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 510 86 546
rect 27 476 39 510
rect 73 476 86 510
rect 27 440 86 476
rect 27 406 39 440
rect 73 406 86 440
rect 27 368 86 406
rect 116 531 176 592
rect 116 497 129 531
rect 163 497 176 531
rect 116 440 176 497
rect 116 406 129 440
rect 163 406 176 440
rect 116 368 176 406
rect 206 580 266 592
rect 206 546 219 580
rect 253 546 266 580
rect 206 508 266 546
rect 206 474 219 508
rect 253 474 266 508
rect 206 368 266 474
rect 296 531 356 592
rect 296 497 309 531
rect 343 497 356 531
rect 296 440 356 497
rect 296 406 309 440
rect 343 406 356 440
rect 296 368 356 406
rect 386 580 446 592
rect 386 546 399 580
rect 433 546 446 580
rect 386 508 446 546
rect 386 474 399 508
rect 433 474 446 508
rect 386 368 446 474
rect 476 578 536 592
rect 476 544 489 578
rect 523 544 536 578
rect 476 368 536 544
rect 566 580 626 592
rect 566 546 579 580
rect 613 546 626 580
rect 566 508 626 546
rect 566 474 579 508
rect 613 474 626 508
rect 566 368 626 474
rect 656 578 718 592
rect 656 544 669 578
rect 703 544 718 578
rect 656 368 718 544
rect 748 580 807 592
rect 748 546 761 580
rect 795 546 807 580
rect 748 508 807 546
rect 748 474 761 508
rect 795 474 807 508
rect 748 368 807 474
rect 861 580 920 592
rect 861 546 873 580
rect 907 546 920 580
rect 861 508 920 546
rect 861 474 873 508
rect 907 474 920 508
rect 861 368 920 474
rect 950 531 1010 592
rect 950 497 963 531
rect 997 497 1010 531
rect 950 440 1010 497
rect 950 406 963 440
rect 997 406 1010 440
rect 950 368 1010 406
rect 1040 580 1100 592
rect 1040 546 1053 580
rect 1087 546 1100 580
rect 1040 508 1100 546
rect 1040 474 1053 508
rect 1087 474 1100 508
rect 1040 368 1100 474
rect 1130 531 1190 592
rect 1130 497 1143 531
rect 1177 497 1190 531
rect 1130 440 1190 497
rect 1130 406 1143 440
rect 1177 406 1190 440
rect 1130 368 1190 406
rect 1220 580 1300 592
rect 1220 546 1243 580
rect 1277 546 1300 580
rect 1220 508 1300 546
rect 1220 474 1243 508
rect 1277 474 1300 508
rect 1220 440 1300 474
rect 1220 406 1243 440
rect 1277 406 1300 440
rect 1220 368 1300 406
rect 1330 531 1390 592
rect 1330 497 1343 531
rect 1377 497 1390 531
rect 1330 440 1390 497
rect 1330 406 1343 440
rect 1377 406 1390 440
rect 1330 368 1390 406
rect 1420 580 1490 592
rect 1420 546 1443 580
rect 1477 546 1490 580
rect 1420 508 1490 546
rect 1420 474 1443 508
rect 1477 474 1490 508
rect 1420 368 1490 474
rect 1520 531 1590 592
rect 1520 497 1543 531
rect 1577 497 1590 531
rect 1520 440 1590 497
rect 1520 406 1543 440
rect 1577 406 1590 440
rect 1520 368 1590 406
rect 1620 580 1689 592
rect 1620 546 1643 580
rect 1677 546 1689 580
rect 1620 508 1689 546
rect 1620 474 1643 508
rect 1677 474 1689 508
rect 1620 368 1689 474
rect 1743 580 1802 592
rect 1743 546 1755 580
rect 1789 546 1802 580
rect 1743 508 1802 546
rect 1743 474 1755 508
rect 1789 474 1802 508
rect 1743 368 1802 474
rect 1832 580 1892 592
rect 1832 546 1845 580
rect 1879 546 1892 580
rect 1832 510 1892 546
rect 1832 476 1845 510
rect 1879 476 1892 510
rect 1832 440 1892 476
rect 1832 406 1845 440
rect 1879 406 1892 440
rect 1832 368 1892 406
rect 1922 580 2002 592
rect 1922 546 1945 580
rect 1979 546 2002 580
rect 1922 508 2002 546
rect 1922 474 1945 508
rect 1979 474 2002 508
rect 1922 368 2002 474
rect 2032 580 2092 592
rect 2032 546 2045 580
rect 2079 546 2092 580
rect 2032 510 2092 546
rect 2032 476 2045 510
rect 2079 476 2092 510
rect 2032 440 2092 476
rect 2032 406 2045 440
rect 2079 406 2092 440
rect 2032 368 2092 406
rect 2122 580 2181 592
rect 2122 546 2135 580
rect 2169 546 2181 580
rect 2122 510 2181 546
rect 2122 476 2135 510
rect 2169 476 2181 510
rect 2122 440 2181 476
rect 2122 406 2135 440
rect 2169 406 2181 440
rect 2122 368 2181 406
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 125 155 159 189
rect 225 110 259 144
rect 311 155 345 189
rect 411 110 445 144
rect 511 155 545 189
rect 611 110 645 144
rect 711 155 745 189
rect 811 110 845 144
rect 913 66 947 100
rect 1015 150 1049 184
rect 1015 82 1049 116
rect 1115 82 1149 116
rect 1215 150 1249 184
rect 1284 163 1318 197
rect 1242 82 1276 116
rect 1384 102 1418 136
rect 1484 176 1518 210
rect 1484 86 1518 120
rect 1584 102 1618 136
rect 1684 176 1718 210
rect 1684 86 1718 120
rect 1784 102 1818 136
rect 1884 176 1918 210
rect 1884 86 1918 120
rect 1984 102 2018 136
rect 2084 176 2118 210
rect 2084 86 2118 120
<< pdiffc >>
rect 39 546 73 580
rect 39 476 73 510
rect 39 406 73 440
rect 129 497 163 531
rect 129 406 163 440
rect 219 546 253 580
rect 219 474 253 508
rect 309 497 343 531
rect 309 406 343 440
rect 399 546 433 580
rect 399 474 433 508
rect 489 544 523 578
rect 579 546 613 580
rect 579 474 613 508
rect 669 544 703 578
rect 761 546 795 580
rect 761 474 795 508
rect 873 546 907 580
rect 873 474 907 508
rect 963 497 997 531
rect 963 406 997 440
rect 1053 546 1087 580
rect 1053 474 1087 508
rect 1143 497 1177 531
rect 1143 406 1177 440
rect 1243 546 1277 580
rect 1243 474 1277 508
rect 1243 406 1277 440
rect 1343 497 1377 531
rect 1343 406 1377 440
rect 1443 546 1477 580
rect 1443 474 1477 508
rect 1543 497 1577 531
rect 1543 406 1577 440
rect 1643 546 1677 580
rect 1643 474 1677 508
rect 1755 546 1789 580
rect 1755 474 1789 508
rect 1845 546 1879 580
rect 1845 476 1879 510
rect 1845 406 1879 440
rect 1945 546 1979 580
rect 1945 474 1979 508
rect 2045 546 2079 580
rect 2045 476 2079 510
rect 2045 406 2079 440
rect 2135 546 2169 580
rect 2135 476 2169 510
rect 2135 406 2169 440
<< poly >>
rect 86 592 116 618
rect 176 592 206 618
rect 266 592 296 618
rect 356 592 386 618
rect 446 592 476 618
rect 536 592 566 618
rect 626 592 656 618
rect 718 592 748 618
rect 920 592 950 618
rect 1010 592 1040 618
rect 1100 592 1130 618
rect 1190 592 1220 618
rect 1300 592 1330 618
rect 1390 592 1420 618
rect 1490 592 1520 618
rect 1590 592 1620 618
rect 1802 592 1832 618
rect 1892 592 1922 618
rect 2002 592 2032 618
rect 2092 592 2122 618
rect 86 353 116 368
rect 176 353 206 368
rect 266 353 296 368
rect 356 353 386 368
rect 446 353 476 368
rect 536 353 566 368
rect 626 353 656 368
rect 718 353 748 368
rect 920 353 950 368
rect 1010 353 1040 368
rect 1100 353 1130 368
rect 1190 353 1220 368
rect 1300 353 1330 368
rect 1390 353 1420 368
rect 1490 353 1520 368
rect 1590 353 1620 368
rect 1802 353 1832 368
rect 1892 353 1922 368
rect 2002 353 2032 368
rect 2092 353 2122 368
rect 83 336 119 353
rect 173 336 209 353
rect 263 336 299 353
rect 353 336 389 353
rect 83 320 389 336
rect 83 286 99 320
rect 133 286 167 320
rect 201 286 235 320
rect 269 286 303 320
rect 337 286 389 320
rect 83 270 389 286
rect 443 336 479 353
rect 533 336 569 353
rect 623 336 659 353
rect 715 336 751 353
rect 917 336 953 353
rect 1007 336 1043 353
rect 1097 336 1133 353
rect 1187 336 1223 353
rect 1300 336 1333 353
rect 1387 336 1423 353
rect 1487 336 1523 353
rect 1587 336 1623 353
rect 1799 336 1835 353
rect 1889 336 1925 353
rect 1999 336 2035 353
rect 2089 336 2125 353
rect 443 320 786 336
rect 443 286 459 320
rect 493 286 527 320
rect 561 286 595 320
rect 629 286 663 320
rect 697 286 731 320
rect 765 286 786 320
rect 917 320 1223 336
rect 917 300 933 320
rect 443 270 786 286
rect 84 222 114 270
rect 170 222 200 270
rect 270 222 300 270
rect 359 222 389 270
rect 456 222 486 270
rect 556 222 586 270
rect 656 222 686 270
rect 756 222 786 270
rect 856 286 933 300
rect 967 286 1001 320
rect 1035 286 1069 320
rect 1103 306 1223 320
rect 1303 320 1673 336
rect 1103 286 1190 306
rect 856 270 1190 286
rect 1303 286 1319 320
rect 1353 286 1387 320
rect 1421 286 1455 320
rect 1489 286 1523 320
rect 1557 286 1591 320
rect 1625 286 1673 320
rect 1303 270 1673 286
rect 856 222 886 270
rect 974 222 1004 270
rect 1073 222 1103 270
rect 1160 222 1190 270
rect 1329 222 1359 270
rect 1443 222 1473 270
rect 1529 222 1559 270
rect 1643 222 1673 270
rect 1743 320 2125 336
rect 1743 286 1769 320
rect 1803 286 1837 320
rect 1871 286 1905 320
rect 1939 286 1973 320
rect 2007 306 2125 320
rect 2007 286 2059 306
rect 1743 270 2059 286
rect 1743 222 1773 270
rect 1843 222 1873 270
rect 1929 222 1959 270
rect 2029 222 2059 270
rect 84 48 114 74
rect 170 48 200 74
rect 270 48 300 74
rect 359 48 389 74
rect 456 48 486 74
rect 556 48 586 74
rect 656 48 686 74
rect 756 48 786 74
rect 856 48 886 74
rect 974 48 1004 74
rect 1073 48 1103 74
rect 1160 48 1190 74
rect 1329 48 1359 74
rect 1443 48 1473 74
rect 1529 48 1559 74
rect 1643 48 1673 74
rect 1743 48 1773 74
rect 1843 48 1873 74
rect 1929 48 1959 74
rect 2029 48 2059 74
<< polycont >>
rect 99 286 133 320
rect 167 286 201 320
rect 235 286 269 320
rect 303 286 337 320
rect 459 286 493 320
rect 527 286 561 320
rect 595 286 629 320
rect 663 286 697 320
rect 731 286 765 320
rect 933 286 967 320
rect 1001 286 1035 320
rect 1069 286 1103 320
rect 1319 286 1353 320
rect 1387 286 1421 320
rect 1455 286 1489 320
rect 1523 286 1557 320
rect 1591 286 1625 320
rect 1769 286 1803 320
rect 1837 286 1871 320
rect 1905 286 1939 320
rect 1973 286 2007 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 23 581 449 615
rect 23 580 89 581
rect 23 546 39 580
rect 73 546 89 580
rect 203 580 253 581
rect 23 510 89 546
rect 23 476 39 510
rect 73 476 89 510
rect 23 440 89 476
rect 23 406 39 440
rect 73 406 89 440
rect 23 390 89 406
rect 129 531 163 547
rect 129 440 163 497
rect 203 546 219 580
rect 399 580 449 581
rect 203 508 253 546
rect 203 474 219 508
rect 203 458 253 474
rect 293 531 359 547
rect 293 497 309 531
rect 343 497 359 531
rect 293 440 359 497
rect 433 546 449 580
rect 399 508 449 546
rect 489 578 523 649
rect 489 526 523 544
rect 563 580 629 596
rect 563 546 579 580
rect 613 546 629 580
rect 433 492 449 508
rect 563 508 629 546
rect 669 578 703 649
rect 669 526 703 544
rect 745 580 811 596
rect 745 546 761 580
rect 795 546 811 580
rect 563 492 579 508
rect 433 474 579 492
rect 613 492 629 508
rect 745 508 811 546
rect 745 492 761 508
rect 613 474 761 492
rect 795 474 811 508
rect 399 458 811 474
rect 857 581 1693 615
rect 857 580 907 581
rect 857 546 873 580
rect 1053 580 1087 581
rect 857 508 907 546
rect 857 474 873 508
rect 857 458 907 474
rect 947 531 1013 547
rect 947 497 963 531
rect 997 497 1013 531
rect 293 424 309 440
rect 163 406 309 424
rect 343 424 359 440
rect 947 440 1013 497
rect 1229 580 1293 581
rect 1053 508 1087 546
rect 1053 458 1087 474
rect 1127 531 1193 547
rect 1127 497 1143 531
rect 1177 497 1193 531
rect 947 424 963 440
rect 343 406 963 424
rect 997 424 1013 440
rect 1127 440 1193 497
rect 1127 424 1143 440
rect 997 406 1143 424
rect 1177 424 1193 440
rect 1229 546 1243 580
rect 1277 546 1293 580
rect 1427 580 1493 581
rect 1229 508 1293 546
rect 1229 474 1243 508
rect 1277 474 1293 508
rect 1229 440 1293 474
rect 1177 406 1195 424
rect 129 390 1195 406
rect 1229 406 1243 440
rect 1277 406 1293 440
rect 1229 390 1293 406
rect 1327 531 1393 547
rect 1327 497 1343 531
rect 1377 497 1393 531
rect 1327 440 1393 497
rect 1427 546 1443 580
rect 1477 546 1493 580
rect 1627 580 1693 581
rect 1427 508 1493 546
rect 1427 474 1443 508
rect 1477 474 1493 508
rect 1427 458 1493 474
rect 1527 531 1593 547
rect 1527 497 1543 531
rect 1577 497 1593 531
rect 1327 406 1343 440
rect 1377 424 1393 440
rect 1527 440 1593 497
rect 1627 546 1643 580
rect 1677 546 1693 580
rect 1627 508 1693 546
rect 1627 474 1643 508
rect 1677 474 1693 508
rect 1627 458 1693 474
rect 1739 580 1789 649
rect 1739 546 1755 580
rect 1739 508 1789 546
rect 1739 474 1755 508
rect 1739 458 1789 474
rect 1829 580 1895 596
rect 1829 546 1845 580
rect 1879 546 1895 580
rect 1829 510 1895 546
rect 1829 476 1845 510
rect 1879 476 1895 510
rect 1527 424 1543 440
rect 1377 406 1543 424
rect 1577 424 1593 440
rect 1829 440 1895 476
rect 1929 580 1995 649
rect 1929 546 1945 580
rect 1979 546 1995 580
rect 1929 508 1995 546
rect 1929 474 1945 508
rect 1979 474 1995 508
rect 1929 458 1995 474
rect 2029 580 2095 596
rect 2029 546 2045 580
rect 2079 546 2095 580
rect 2029 510 2095 546
rect 2029 476 2045 510
rect 2079 476 2095 510
rect 1829 424 1845 440
rect 1577 406 1845 424
rect 1879 424 1895 440
rect 2029 440 2095 476
rect 2029 424 2045 440
rect 1879 406 2045 424
rect 2079 406 2095 440
rect 1327 390 2095 406
rect 2135 580 2185 649
rect 2169 546 2185 580
rect 2135 510 2185 546
rect 2169 476 2185 510
rect 2135 440 2185 476
rect 2169 406 2185 440
rect 2135 390 2185 406
rect 25 320 359 356
rect 25 286 99 320
rect 133 286 167 320
rect 201 286 235 320
rect 269 286 303 320
rect 337 286 359 320
rect 409 320 839 356
rect 409 286 459 320
rect 493 286 527 320
rect 561 286 595 320
rect 629 286 663 320
rect 697 286 731 320
rect 765 286 839 320
rect 889 320 1127 356
rect 889 286 933 320
rect 967 286 1001 320
rect 1035 286 1069 320
rect 1103 286 1127 320
rect 1161 252 1195 390
rect 1273 320 1703 356
rect 1273 286 1319 320
rect 1353 286 1387 320
rect 1421 286 1455 320
rect 1489 286 1523 320
rect 1557 286 1591 320
rect 1625 286 1703 320
rect 1273 270 1703 286
rect 1753 320 2183 356
rect 1753 286 1769 320
rect 1803 286 1837 320
rect 1871 286 1905 320
rect 1939 286 1973 320
rect 2007 286 2183 320
rect 1753 270 2183 286
rect 23 210 73 226
rect 23 176 39 210
rect 23 120 73 176
rect 23 86 39 120
rect 109 218 1195 252
rect 109 189 175 218
rect 109 155 125 189
rect 159 155 175 189
rect 311 189 361 218
rect 109 119 175 155
rect 209 144 275 184
rect 23 85 73 86
rect 209 110 225 144
rect 259 110 275 144
rect 345 155 361 189
rect 495 189 561 218
rect 311 119 361 155
rect 395 144 461 184
rect 209 85 275 110
rect 395 110 411 144
rect 445 110 461 144
rect 495 155 511 189
rect 545 155 561 189
rect 695 189 761 218
rect 495 119 561 155
rect 595 144 661 184
rect 395 85 461 110
rect 595 110 611 144
rect 645 110 661 144
rect 695 155 711 189
rect 745 155 761 189
rect 1266 210 2134 236
rect 1266 202 1484 210
rect 1266 197 1334 202
rect 1266 184 1284 197
rect 695 119 761 155
rect 795 150 1015 184
rect 1049 150 1215 184
rect 1249 163 1284 184
rect 1318 163 1334 197
rect 1468 176 1484 202
rect 1518 202 1684 210
rect 1518 176 1534 202
rect 1249 150 1334 163
rect 795 144 861 150
rect 595 85 661 110
rect 795 110 811 144
rect 845 110 861 144
rect 999 116 1065 150
rect 1199 116 1334 150
rect 795 85 861 110
rect 23 51 861 85
rect 897 100 963 116
rect 897 66 913 100
rect 947 66 963 100
rect 999 82 1015 116
rect 1049 82 1065 116
rect 999 66 1065 82
rect 1099 82 1115 116
rect 1149 82 1165 116
rect 897 17 963 66
rect 1099 17 1165 82
rect 1199 82 1242 116
rect 1276 82 1334 116
rect 1199 66 1334 82
rect 1368 136 1434 168
rect 1368 102 1384 136
rect 1418 102 1434 136
rect 1368 17 1434 102
rect 1468 120 1534 176
rect 1668 176 1684 202
rect 1718 202 1884 210
rect 1718 176 1734 202
rect 1468 86 1484 120
rect 1518 86 1534 120
rect 1468 70 1534 86
rect 1568 136 1634 168
rect 1568 102 1584 136
rect 1618 102 1634 136
rect 1568 17 1634 102
rect 1668 120 1734 176
rect 1868 176 1884 202
rect 1918 202 2084 210
rect 1918 176 1934 202
rect 1668 86 1684 120
rect 1718 86 1734 120
rect 1668 70 1734 86
rect 1768 136 1834 168
rect 1768 102 1784 136
rect 1818 102 1834 136
rect 1768 17 1834 102
rect 1868 120 1934 176
rect 2068 176 2084 202
rect 2118 176 2134 210
rect 1868 86 1884 120
rect 1918 86 1934 120
rect 1868 70 1934 86
rect 1968 136 2034 168
rect 1968 102 1984 136
rect 2018 102 2034 136
rect 1968 17 2034 102
rect 2068 120 2134 176
rect 2068 86 2084 120
rect 2118 86 2134 120
rect 2068 70 2134 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
<< metal1 >>
rect 0 683 2208 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 0 617 2208 649
rect 0 17 2208 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
rect 0 -49 2208 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o32ai_4
flabel pwell s 0 0 2208 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 0 617 2208 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 0 617 2208 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 2208 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 319 464 353 498 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 B2
port 5 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 B2
port 5 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 B2
port 5 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 B2
port 5 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 B1
port 4 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 B1
port 4 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 4 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 B1
port 4 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 B1
port 4 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 1279 316 1313 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 1375 316 1409 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 1471 316 1505 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 1567 316 1601 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 1663 316 1697 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 1759 316 1793 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 1855 316 1889 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 1951 316 1985 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 2047 316 2081 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 2143 316 2177 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 2208 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 958918
string GDS_START 940966
<< end >>
