magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1012 561
rect 103 451 169 527
rect 282 451 348 527
rect 450 451 516 527
rect 695 451 761 527
rect 927 451 993 527
rect 88 153 158 327
rect 196 309 432 343
rect 196 164 252 309
rect 196 130 416 164
rect 114 17 180 94
rect 214 51 248 130
rect 282 17 348 94
rect 382 51 416 130
rect 573 199 617 265
rect 669 151 711 265
rect 763 147 829 265
rect 457 17 523 89
rect 0 -17 1012 17
<< obsli1 >>
rect 17 417 69 493
rect 17 383 980 417
rect 17 117 52 383
rect 476 309 909 343
rect 476 249 510 309
rect 288 215 510 249
rect 17 51 69 117
rect 476 157 510 215
rect 476 123 593 157
rect 946 199 980 383
rect 559 94 593 123
rect 878 94 993 162
rect 559 60 993 94
<< metal1 >>
rect 0 496 1012 592
rect 0 -48 1012 48
<< labels >>
rlabel locali s 88 153 158 327 6 A_N
port 1 nsew signal input
rlabel locali s 763 147 829 265 6 B
port 2 nsew signal input
rlabel locali s 669 151 711 265 6 C
port 3 nsew signal input
rlabel locali s 573 199 617 265 6 D
port 4 nsew signal input
rlabel locali s 382 51 416 130 6 X
port 5 nsew signal output
rlabel locali s 214 51 248 130 6 X
port 5 nsew signal output
rlabel locali s 196 309 432 343 6 X
port 5 nsew signal output
rlabel locali s 196 164 252 309 6 X
port 5 nsew signal output
rlabel locali s 196 130 416 164 6 X
port 5 nsew signal output
rlabel locali s 457 17 523 89 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 282 17 348 94 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 114 17 180 94 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 1012 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1012 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 927 451 993 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 695 451 761 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 450 451 516 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 282 451 348 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 103 451 169 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 1012 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 1012 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1012 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3858944
string GDS_START 3851266
<< end >>
