magic
tech sky130A
magscale 1 2
timestamp 1599588238
<< locali >>
rect 113 492 179 596
rect 303 492 369 596
rect 505 492 559 596
rect 113 458 559 492
rect 113 364 219 458
rect 25 236 147 310
rect 185 252 219 364
rect 285 390 565 424
rect 285 336 359 390
rect 253 310 359 336
rect 253 286 319 310
rect 393 286 459 356
rect 531 330 565 390
rect 531 264 613 330
rect 185 218 455 252
rect 389 187 455 218
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 23 364 73 649
rect 213 526 263 649
rect 403 526 469 649
rect 599 364 649 649
rect 20 184 86 202
rect 20 153 274 184
rect 586 153 652 230
rect 20 150 652 153
rect 20 70 70 150
rect 208 119 652 150
rect 106 17 172 116
rect 208 66 242 119
rect 291 51 553 85
rect 589 81 652 119
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel locali s 393 286 459 356 6 A
port 1 nsew signal input
rlabel locali s 531 330 565 390 6 B
port 2 nsew signal input
rlabel locali s 531 264 613 330 6 B
port 2 nsew signal input
rlabel locali s 285 390 565 424 6 B
port 2 nsew signal input
rlabel locali s 285 336 359 390 6 B
port 2 nsew signal input
rlabel locali s 253 310 359 336 6 B
port 2 nsew signal input
rlabel locali s 253 286 319 310 6 B
port 2 nsew signal input
rlabel locali s 25 236 147 310 6 C
port 3 nsew signal input
rlabel locali s 505 492 559 596 6 Y
port 4 nsew signal output
rlabel locali s 389 187 455 218 6 Y
port 4 nsew signal output
rlabel locali s 303 492 369 596 6 Y
port 4 nsew signal output
rlabel locali s 185 252 219 364 6 Y
port 4 nsew signal output
rlabel locali s 185 218 455 252 6 Y
port 4 nsew signal output
rlabel locali s 113 492 179 596 6 Y
port 4 nsew signal output
rlabel locali s 113 458 559 492 6 Y
port 4 nsew signal output
rlabel locali s 113 364 219 458 6 Y
port 4 nsew signal output
rlabel metal1 s 0 -49 672 49 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 617 672 715 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1748528
string GDS_START 1741932
<< end >>
