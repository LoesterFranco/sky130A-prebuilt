magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 2024 561
rect 104 427 170 527
rect 19 195 89 325
rect 103 17 169 93
rect 376 449 442 527
rect 356 157 390 337
rect 751 433 785 527
rect 492 271 558 337
rect 616 157 650 223
rect 706 207 804 331
rect 356 123 650 157
rect 1186 367 1220 527
rect 395 17 461 89
rect 495 61 530 123
rect 1562 427 1623 527
rect 1781 325 1816 527
rect 752 17 792 105
rect 1144 17 1218 117
rect 1852 301 1921 479
rect 1549 17 1623 123
rect 1887 164 1921 301
rect 1955 281 1989 527
rect 1781 17 1815 139
rect 1852 61 1921 164
rect 1955 17 1989 186
rect 0 -17 2024 17
<< obsli1 >>
rect 36 393 70 493
rect 36 391 169 393
rect 36 359 128 391
rect 123 357 128 359
rect 162 357 169 391
rect 123 194 169 357
rect 123 161 162 194
rect 35 127 162 161
rect 204 187 249 493
rect 204 153 210 187
rect 244 153 249 187
rect 204 143 249 153
rect 35 69 69 127
rect 203 69 249 143
rect 287 415 342 489
rect 538 449 717 483
rect 287 372 649 415
rect 287 89 321 372
rect 424 225 458 372
rect 615 337 649 372
rect 683 399 717 449
rect 842 413 889 488
rect 938 438 1152 472
rect 842 399 876 413
rect 683 365 876 399
rect 996 391 1084 402
rect 615 271 654 337
rect 424 191 492 225
rect 842 173 876 365
rect 684 139 876 173
rect 910 207 958 381
rect 996 357 1041 391
rect 1075 357 1084 391
rect 996 331 1084 357
rect 1118 315 1152 438
rect 1254 427 1304 493
rect 1349 433 1526 467
rect 1118 297 1220 315
rect 1060 263 1220 297
rect 910 187 1026 207
rect 910 153 949 187
rect 983 153 1026 187
rect 910 141 1026 153
rect 287 55 361 89
rect 684 89 718 139
rect 842 107 876 139
rect 1060 107 1094 263
rect 1186 249 1220 263
rect 1128 213 1162 219
rect 1254 213 1288 427
rect 1322 391 1360 393
rect 1322 357 1324 391
rect 1358 357 1360 391
rect 1322 249 1360 357
rect 1394 315 1458 381
rect 1128 153 1288 213
rect 1394 207 1432 315
rect 1492 281 1526 433
rect 1693 381 1747 491
rect 1560 315 1747 381
rect 564 55 718 89
rect 842 73 912 107
rect 946 73 1094 107
rect 1254 107 1288 153
rect 1322 187 1432 207
rect 1322 153 1326 187
rect 1360 153 1432 187
rect 1322 141 1432 153
rect 1466 265 1526 281
rect 1713 265 1747 315
rect 1466 199 1679 265
rect 1713 199 1853 265
rect 1466 107 1500 199
rect 1713 165 1747 199
rect 1254 73 1346 107
rect 1392 73 1500 107
rect 1677 60 1747 165
<< obsli1c >>
rect 128 357 162 391
rect 210 153 244 187
rect 1041 357 1075 391
rect 949 153 983 187
rect 1324 357 1358 391
rect 1326 153 1360 187
<< metal1 >>
rect 0 496 2024 592
rect 0 -48 2024 48
<< obsm1 >>
rect 116 391 174 397
rect 116 357 128 391
rect 162 388 174 391
rect 1029 391 1087 397
rect 1029 388 1041 391
rect 162 360 1041 388
rect 162 357 174 360
rect 116 351 174 357
rect 1029 357 1041 360
rect 1075 388 1087 391
rect 1312 391 1370 397
rect 1312 388 1324 391
rect 1075 360 1324 388
rect 1075 357 1087 360
rect 1029 351 1087 357
rect 1312 357 1324 360
rect 1358 357 1370 391
rect 1312 351 1370 357
rect 198 187 256 193
rect 198 153 210 187
rect 244 184 256 187
rect 937 187 995 193
rect 937 184 949 187
rect 244 156 949 184
rect 244 153 256 156
rect 198 147 256 153
rect 937 153 949 156
rect 983 184 995 187
rect 1314 187 1372 193
rect 1314 184 1326 187
rect 983 156 1326 184
rect 983 153 995 156
rect 937 147 995 153
rect 1314 153 1326 156
rect 1360 153 1372 187
rect 1314 147 1372 153
<< labels >>
rlabel locali s 492 271 558 337 6 D
port 1 nsew signal input
rlabel locali s 1887 164 1921 301 6 Q
port 2 nsew signal output
rlabel locali s 1852 301 1921 479 6 Q
port 2 nsew signal output
rlabel locali s 1852 61 1921 164 6 Q
port 2 nsew signal output
rlabel locali s 706 207 804 331 6 SCD
port 3 nsew signal input
rlabel locali s 616 157 650 223 6 SCE
port 4 nsew signal input
rlabel locali s 495 61 530 123 6 SCE
port 4 nsew signal input
rlabel locali s 356 157 390 337 6 SCE
port 4 nsew signal input
rlabel locali s 356 123 650 157 6 SCE
port 4 nsew signal input
rlabel locali s 19 195 89 325 6 CLK
port 5 nsew clock input
rlabel locali s 1955 17 1989 186 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1781 17 1815 139 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1549 17 1623 123 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1144 17 1218 117 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 752 17 792 105 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 395 17 461 89 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 103 17 169 93 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 2024 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 2024 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1955 281 1989 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1781 325 1816 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1562 427 1623 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1186 367 1220 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 751 433 785 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 376 449 442 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 104 427 170 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 2024 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 2024 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2024 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 392160
string GDS_START 376362
<< end >>
