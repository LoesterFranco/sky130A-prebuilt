magic
tech sky130A
magscale 1 2
timestamp 1601050058
<< locali >>
rect 119 401 170 485
rect 30 367 170 401
rect 30 177 76 367
rect 214 207 305 265
rect 266 199 305 207
rect 30 143 170 177
rect 104 63 170 143
rect 537 199 620 323
rect 654 199 712 323
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 18 451 85 527
rect 208 455 274 527
rect 395 421 445 493
rect 223 379 445 421
rect 223 333 257 379
rect 114 299 257 333
rect 291 311 373 345
rect 114 215 180 299
rect 339 265 373 311
rect 411 335 445 379
rect 479 403 545 493
rect 579 437 613 527
rect 647 403 713 493
rect 479 369 713 403
rect 411 301 503 335
rect 339 199 435 265
rect 18 17 69 109
rect 204 17 244 173
rect 339 165 373 199
rect 291 131 373 165
rect 469 165 503 301
rect 469 127 548 165
rect 395 17 461 93
rect 647 17 713 165
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel locali s 537 199 620 323 6 A1
port 1 nsew signal input
rlabel locali s 654 199 712 323 6 A2
port 2 nsew signal input
rlabel locali s 266 199 305 207 6 B1_N
port 3 nsew signal input
rlabel locali s 214 207 305 265 6 B1_N
port 3 nsew signal input
rlabel locali s 119 401 170 485 6 X
port 4 nsew signal output
rlabel locali s 104 63 170 143 6 X
port 4 nsew signal output
rlabel locali s 30 367 170 401 6 X
port 4 nsew signal output
rlabel locali s 30 177 76 367 6 X
port 4 nsew signal output
rlabel locali s 30 143 170 177 6 X
port 4 nsew signal output
rlabel metal1 s 0 -48 736 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 736 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3989514
string GDS_START 3983218
<< end >>
