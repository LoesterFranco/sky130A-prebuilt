magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 79 47 109 177
rect 287 47 317 177
rect 381 47 411 177
rect 475 47 505 177
rect 569 47 599 177
rect 674 47 704 177
rect 768 47 798 177
rect 862 47 892 177
rect 956 47 986 177
<< pmoshvt >>
rect 81 297 117 497
rect 186 309 222 497
rect 280 309 316 497
rect 374 309 410 497
rect 468 309 504 497
rect 676 297 712 497
rect 770 297 806 497
rect 864 297 900 497
rect 958 297 994 497
<< ndiff >>
rect 27 129 79 177
rect 27 95 35 129
rect 69 95 79 129
rect 27 47 79 95
rect 109 93 171 177
rect 109 59 129 93
rect 163 59 171 93
rect 109 47 171 59
rect 235 129 287 177
rect 235 95 243 129
rect 277 95 287 129
rect 235 47 287 95
rect 317 89 381 177
rect 317 55 337 89
rect 371 55 381 89
rect 317 47 381 55
rect 411 129 475 177
rect 411 95 431 129
rect 465 95 475 129
rect 411 47 475 95
rect 505 89 569 177
rect 505 55 525 89
rect 559 55 569 89
rect 505 47 569 55
rect 599 129 674 177
rect 599 95 625 129
rect 659 95 674 129
rect 599 47 674 95
rect 704 165 768 177
rect 704 131 724 165
rect 758 131 768 165
rect 704 47 768 131
rect 798 90 862 177
rect 798 56 818 90
rect 852 56 862 90
rect 798 47 862 56
rect 892 165 956 177
rect 892 131 912 165
rect 946 131 956 165
rect 892 47 956 131
rect 986 90 1052 177
rect 986 56 1006 90
rect 1040 56 1052 90
rect 986 47 1052 56
<< pdiff >>
rect 27 448 81 497
rect 27 414 35 448
rect 69 414 81 448
rect 27 380 81 414
rect 27 346 35 380
rect 69 346 81 380
rect 27 297 81 346
rect 117 489 186 497
rect 117 455 129 489
rect 163 455 186 489
rect 117 421 186 455
rect 117 387 129 421
rect 163 387 186 421
rect 117 309 186 387
rect 222 448 280 497
rect 222 414 234 448
rect 268 414 280 448
rect 222 380 280 414
rect 222 346 234 380
rect 268 346 280 380
rect 222 309 280 346
rect 316 489 374 497
rect 316 455 328 489
rect 362 455 374 489
rect 316 421 374 455
rect 316 387 328 421
rect 362 387 374 421
rect 316 309 374 387
rect 410 448 468 497
rect 410 414 422 448
rect 456 414 468 448
rect 410 380 468 414
rect 410 346 422 380
rect 456 346 468 380
rect 410 309 468 346
rect 504 485 558 497
rect 504 451 516 485
rect 550 451 558 485
rect 504 417 558 451
rect 504 383 516 417
rect 550 383 558 417
rect 504 309 558 383
rect 622 448 676 497
rect 622 414 630 448
rect 664 414 676 448
rect 622 380 676 414
rect 622 346 630 380
rect 664 346 676 380
rect 117 297 169 309
rect 622 297 676 346
rect 712 407 770 497
rect 712 373 724 407
rect 758 373 770 407
rect 712 339 770 373
rect 712 305 724 339
rect 758 305 770 339
rect 712 297 770 305
rect 806 448 864 497
rect 806 414 818 448
rect 852 414 864 448
rect 806 380 864 414
rect 806 346 818 380
rect 852 346 864 380
rect 806 297 864 346
rect 900 407 958 497
rect 900 373 912 407
rect 946 373 958 407
rect 900 339 958 373
rect 900 305 912 339
rect 946 305 958 339
rect 900 297 958 305
rect 994 448 1048 497
rect 994 414 1006 448
rect 1040 414 1048 448
rect 994 380 1048 414
rect 994 346 1006 380
rect 1040 346 1048 380
rect 994 297 1048 346
<< ndiffc >>
rect 35 95 69 129
rect 129 59 163 93
rect 243 95 277 129
rect 337 55 371 89
rect 431 95 465 129
rect 525 55 559 89
rect 625 95 659 129
rect 724 131 758 165
rect 818 56 852 90
rect 912 131 946 165
rect 1006 56 1040 90
<< pdiffc >>
rect 35 414 69 448
rect 35 346 69 380
rect 129 455 163 489
rect 129 387 163 421
rect 234 414 268 448
rect 234 346 268 380
rect 328 455 362 489
rect 328 387 362 421
rect 422 414 456 448
rect 422 346 456 380
rect 516 451 550 485
rect 516 383 550 417
rect 630 414 664 448
rect 630 346 664 380
rect 724 373 758 407
rect 724 305 758 339
rect 818 414 852 448
rect 818 346 852 380
rect 912 373 946 407
rect 912 305 946 339
rect 1006 414 1040 448
rect 1006 346 1040 380
<< poly >>
rect 81 497 117 523
rect 186 497 222 523
rect 280 497 316 523
rect 374 497 410 523
rect 468 497 504 523
rect 676 497 712 523
rect 770 497 806 523
rect 864 497 900 523
rect 958 497 994 523
rect 81 282 117 297
rect 186 294 222 309
rect 280 294 316 309
rect 374 294 410 309
rect 468 294 504 309
rect 79 265 119 282
rect 184 265 506 294
rect 676 282 712 297
rect 770 282 806 297
rect 864 282 900 297
rect 958 282 994 297
rect 674 265 714 282
rect 768 265 808 282
rect 862 265 902 282
rect 956 265 996 282
rect 22 264 506 265
rect 22 249 224 264
rect 22 215 32 249
rect 66 235 224 249
rect 548 249 612 265
rect 66 215 109 235
rect 548 222 558 249
rect 22 199 109 215
rect 79 177 109 199
rect 287 215 558 222
rect 592 215 612 249
rect 287 199 612 215
rect 674 249 1056 265
rect 674 215 1012 249
rect 1046 215 1056 249
rect 674 199 1056 215
rect 287 192 599 199
rect 287 177 317 192
rect 381 177 411 192
rect 475 177 505 192
rect 569 177 599 192
rect 674 177 704 199
rect 768 177 798 199
rect 862 177 892 199
rect 956 177 986 199
rect 79 21 109 47
rect 287 21 317 47
rect 381 21 411 47
rect 475 21 505 47
rect 569 21 599 47
rect 674 21 704 47
rect 768 21 798 47
rect 862 21 892 47
rect 956 21 986 47
<< polycont >>
rect 32 215 66 249
rect 558 215 592 249
rect 1012 215 1046 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 17 448 69 493
rect 17 414 35 448
rect 17 380 69 414
rect 17 346 35 380
rect 103 489 179 527
rect 103 455 129 489
rect 163 455 179 489
rect 103 421 179 455
rect 103 387 129 421
rect 163 387 179 421
rect 103 367 179 387
rect 213 448 268 493
rect 213 414 234 448
rect 213 380 268 414
rect 17 333 69 346
rect 213 346 234 380
rect 302 489 378 527
rect 302 455 328 489
rect 362 455 378 489
rect 302 421 378 455
rect 302 387 328 421
rect 362 387 378 421
rect 302 367 378 387
rect 422 448 456 493
rect 422 380 456 414
rect 213 333 268 346
rect 490 485 578 527
rect 490 451 516 485
rect 550 451 578 485
rect 490 417 578 451
rect 490 383 516 417
rect 550 383 578 417
rect 490 367 578 383
rect 622 459 1040 493
rect 622 448 664 459
rect 622 414 630 448
rect 818 448 852 459
rect 622 380 664 414
rect 422 333 456 346
rect 622 346 630 380
rect 622 333 664 346
rect 17 299 179 333
rect 213 299 664 333
rect 698 407 774 415
rect 698 373 724 407
rect 758 373 774 407
rect 698 339 774 373
rect 698 305 724 339
rect 758 305 774 339
rect 1006 448 1040 459
rect 818 380 852 414
rect 818 330 852 346
rect 886 407 962 415
rect 886 373 912 407
rect 946 373 962 407
rect 886 339 962 373
rect 103 265 179 299
rect 698 296 774 305
rect 886 305 912 339
rect 946 305 962 339
rect 1006 380 1040 414
rect 1006 330 1040 346
rect 886 296 962 305
rect 17 249 69 265
rect 17 215 32 249
rect 66 215 69 249
rect 17 199 69 215
rect 103 249 664 265
rect 103 215 558 249
rect 592 215 664 249
rect 103 199 664 215
rect 103 165 179 199
rect 698 165 962 296
rect 17 131 179 165
rect 213 131 659 165
rect 17 129 69 131
rect 17 95 35 129
rect 213 129 277 131
rect 17 51 69 95
rect 103 93 179 97
rect 103 59 129 93
rect 163 59 179 93
rect 103 17 179 59
rect 213 95 243 129
rect 431 129 465 131
rect 213 51 277 95
rect 321 89 387 97
rect 321 55 337 89
rect 371 55 387 89
rect 321 17 387 55
rect 625 129 659 131
rect 431 51 465 95
rect 509 89 575 97
rect 509 55 525 89
rect 559 55 575 89
rect 509 17 575 55
rect 698 131 724 165
rect 758 131 912 165
rect 946 131 962 165
rect 698 124 962 131
rect 996 249 1083 265
rect 996 215 1012 249
rect 1046 215 1083 249
rect 996 124 1083 215
rect 625 90 659 95
rect 625 56 818 90
rect 852 56 1006 90
rect 1040 56 1087 90
rect 625 51 1087 56
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
flabel corelocali s 30 221 64 255 0 FreeSans 200 0 0 0 TE_B
port 2 nsew
flabel corelocali s 858 153 892 187 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 858 221 892 255 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 766 221 800 255 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 766 153 800 187 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 1039 153 1073 187 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 1039 221 1073 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew
rlabel comment s 0 0 0 0 4 einvn_4
<< properties >>
string FIXED_BBOX 0 0 1104 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2025302
string GDS_START 2017172
<< end >>
