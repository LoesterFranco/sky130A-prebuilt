magic
tech sky130A
magscale 1 2
timestamp 1599588209
<< nwell >>
rect -38 332 998 704
<< pwell >>
rect 0 0 960 49
<< scpmos >>
rect 122 368 152 568
rect 206 368 236 568
rect 320 368 350 568
rect 448 368 478 568
rect 548 368 578 568
rect 744 368 774 592
rect 834 368 864 592
<< nmoslvt >>
rect 125 74 155 222
rect 239 74 269 222
rect 339 74 369 222
rect 431 74 461 222
rect 545 74 575 222
rect 757 74 787 222
rect 843 74 873 222
<< ndiff >>
rect 54 202 125 222
rect 54 168 80 202
rect 114 168 125 202
rect 54 120 125 168
rect 54 86 80 120
rect 114 86 125 120
rect 54 74 125 86
rect 155 126 239 222
rect 155 92 180 126
rect 214 92 239 126
rect 155 74 239 92
rect 269 202 339 222
rect 269 168 294 202
rect 328 168 339 202
rect 269 120 339 168
rect 269 86 294 120
rect 328 86 339 120
rect 269 74 339 86
rect 369 74 431 222
rect 461 74 545 222
rect 575 210 632 222
rect 575 176 586 210
rect 620 176 632 210
rect 575 120 632 176
rect 575 86 586 120
rect 620 86 632 120
rect 575 74 632 86
rect 686 143 757 222
rect 686 109 712 143
rect 746 109 757 143
rect 686 74 757 109
rect 787 210 843 222
rect 787 176 798 210
rect 832 176 843 210
rect 787 120 843 176
rect 787 86 798 120
rect 832 86 843 120
rect 787 74 843 86
rect 873 210 933 222
rect 873 176 885 210
rect 919 176 933 210
rect 873 120 933 176
rect 873 86 885 120
rect 919 86 933 120
rect 873 74 933 86
<< pdiff >>
rect 691 568 744 592
rect 63 556 122 568
rect 63 522 75 556
rect 109 522 122 556
rect 63 485 122 522
rect 63 451 75 485
rect 109 451 122 485
rect 63 414 122 451
rect 63 380 75 414
rect 109 380 122 414
rect 63 368 122 380
rect 152 368 206 568
rect 236 556 320 568
rect 236 522 273 556
rect 307 522 320 556
rect 236 485 320 522
rect 236 451 273 485
rect 307 451 320 485
rect 236 414 320 451
rect 236 380 273 414
rect 307 380 320 414
rect 236 368 320 380
rect 350 560 448 568
rect 350 526 373 560
rect 407 526 448 560
rect 350 492 448 526
rect 350 458 373 492
rect 407 458 448 492
rect 350 368 448 458
rect 478 560 548 568
rect 478 526 491 560
rect 525 526 548 560
rect 478 492 548 526
rect 478 458 491 492
rect 525 458 548 492
rect 478 424 548 458
rect 478 390 491 424
rect 525 390 548 424
rect 478 368 548 390
rect 578 560 744 568
rect 578 526 591 560
rect 625 526 687 560
rect 721 526 744 560
rect 578 492 744 526
rect 578 458 591 492
rect 625 458 687 492
rect 721 458 744 492
rect 578 368 744 458
rect 774 580 834 592
rect 774 546 787 580
rect 821 546 834 580
rect 774 497 834 546
rect 774 463 787 497
rect 821 463 834 497
rect 774 414 834 463
rect 774 380 787 414
rect 821 380 834 414
rect 774 368 834 380
rect 864 580 933 592
rect 864 546 887 580
rect 921 546 933 580
rect 864 497 933 546
rect 864 463 887 497
rect 921 463 933 497
rect 864 414 933 463
rect 864 380 887 414
rect 921 380 933 414
rect 864 368 933 380
<< ndiffc >>
rect 80 168 114 202
rect 80 86 114 120
rect 180 92 214 126
rect 294 168 328 202
rect 294 86 328 120
rect 586 176 620 210
rect 586 86 620 120
rect 712 109 746 143
rect 798 176 832 210
rect 798 86 832 120
rect 885 176 919 210
rect 885 86 919 120
<< pdiffc >>
rect 75 522 109 556
rect 75 451 109 485
rect 75 380 109 414
rect 273 522 307 556
rect 273 451 307 485
rect 273 380 307 414
rect 373 526 407 560
rect 373 458 407 492
rect 491 526 525 560
rect 491 458 525 492
rect 491 390 525 424
rect 591 526 625 560
rect 687 526 721 560
rect 591 458 625 492
rect 687 458 721 492
rect 787 546 821 580
rect 787 463 821 497
rect 787 380 821 414
rect 887 546 921 580
rect 887 463 921 497
rect 887 380 921 414
<< poly >>
rect 122 568 152 594
rect 206 568 236 594
rect 320 568 350 594
rect 448 568 478 594
rect 548 568 578 594
rect 744 592 774 618
rect 834 592 864 618
rect 122 353 152 368
rect 206 353 236 368
rect 320 353 350 368
rect 448 353 478 368
rect 548 353 578 368
rect 744 353 774 368
rect 834 353 864 368
rect 119 310 155 353
rect 21 294 155 310
rect 21 260 37 294
rect 71 260 105 294
rect 139 260 155 294
rect 21 244 155 260
rect 203 310 239 353
rect 317 310 353 353
rect 445 336 481 353
rect 545 336 581 353
rect 431 320 497 336
rect 203 294 269 310
rect 203 260 219 294
rect 253 260 269 294
rect 203 244 269 260
rect 317 294 383 310
rect 317 260 333 294
rect 367 260 383 294
rect 317 244 383 260
rect 431 286 447 320
rect 481 286 497 320
rect 431 270 497 286
rect 545 320 651 336
rect 741 326 777 353
rect 831 326 867 353
rect 545 286 601 320
rect 635 286 651 320
rect 545 270 651 286
rect 703 310 867 326
rect 703 276 719 310
rect 753 290 867 310
rect 753 276 873 290
rect 125 222 155 244
rect 239 222 269 244
rect 339 222 369 244
rect 431 222 461 270
rect 545 222 575 270
rect 703 260 873 276
rect 757 222 787 260
rect 843 222 873 260
rect 125 48 155 74
rect 239 48 269 74
rect 339 48 369 74
rect 431 48 461 74
rect 545 48 575 74
rect 757 48 787 74
rect 843 48 873 74
<< polycont >>
rect 37 260 71 294
rect 105 260 139 294
rect 219 260 253 294
rect 333 260 367 294
rect 447 286 481 320
rect 601 286 635 320
rect 719 276 753 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 59 556 125 649
rect 59 522 75 556
rect 109 522 125 556
rect 59 485 125 522
rect 59 451 75 485
rect 109 451 125 485
rect 59 414 125 451
rect 59 380 75 414
rect 109 380 125 414
rect 59 364 125 380
rect 257 556 323 572
rect 257 522 273 556
rect 307 522 323 556
rect 257 485 323 522
rect 257 451 273 485
rect 307 451 323 485
rect 357 560 423 649
rect 357 526 373 560
rect 407 526 423 560
rect 357 492 423 526
rect 357 458 373 492
rect 407 458 423 492
rect 475 560 541 576
rect 475 526 491 560
rect 525 526 541 560
rect 475 492 541 526
rect 475 458 491 492
rect 525 458 541 492
rect 575 560 737 649
rect 575 526 591 560
rect 625 526 687 560
rect 721 526 737 560
rect 575 492 737 526
rect 575 458 591 492
rect 625 458 687 492
rect 721 458 737 492
rect 771 580 837 596
rect 771 546 787 580
rect 821 546 837 580
rect 771 497 837 546
rect 771 463 787 497
rect 821 463 837 497
rect 257 424 323 451
rect 475 424 541 458
rect 257 414 491 424
rect 257 380 273 414
rect 307 390 491 414
rect 525 390 737 424
rect 307 380 323 390
rect 257 364 323 380
rect 431 320 551 356
rect 21 294 167 310
rect 21 260 37 294
rect 71 260 105 294
rect 139 260 167 294
rect 21 236 167 260
rect 203 294 269 310
rect 203 260 219 294
rect 253 260 269 294
rect 203 236 269 260
rect 313 294 383 310
rect 313 260 333 294
rect 367 260 383 294
rect 431 286 447 320
rect 481 286 551 320
rect 431 270 551 286
rect 585 320 651 356
rect 585 286 601 320
rect 635 286 651 320
rect 585 270 651 286
rect 703 326 737 390
rect 771 414 837 463
rect 771 380 787 414
rect 821 380 837 414
rect 771 364 837 380
rect 871 580 937 649
rect 871 546 887 580
rect 921 546 937 580
rect 871 497 937 546
rect 871 463 887 497
rect 921 463 937 497
rect 871 414 937 463
rect 871 380 887 414
rect 921 380 937 414
rect 871 364 937 380
rect 703 310 769 326
rect 703 276 719 310
rect 753 276 769 310
rect 313 236 383 260
rect 703 260 769 276
rect 703 236 737 260
rect 570 210 737 236
rect 803 226 837 364
rect 50 168 80 202
rect 114 168 294 202
rect 328 168 344 202
rect 50 120 116 168
rect 50 86 80 120
rect 114 86 116 120
rect 50 70 116 86
rect 150 126 244 134
rect 150 92 180 126
rect 214 92 244 126
rect 150 17 244 92
rect 278 120 344 168
rect 278 86 294 120
rect 328 86 344 120
rect 278 70 344 86
rect 570 176 586 210
rect 620 202 737 210
rect 782 210 848 226
rect 620 176 636 202
rect 570 120 636 176
rect 782 176 798 210
rect 832 176 848 210
rect 570 86 586 120
rect 620 86 636 120
rect 570 70 636 86
rect 682 143 748 165
rect 682 109 712 143
rect 746 109 748 143
rect 682 17 748 109
rect 782 120 848 176
rect 782 86 798 120
rect 832 86 848 120
rect 782 70 848 86
rect 884 210 937 226
rect 884 176 885 210
rect 919 176 937 210
rect 884 120 937 176
rect 884 86 885 120
rect 919 86 937 120
rect 884 17 937 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o2111a_2
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 127 242 161 276 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 223 242 257 276 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 319 242 353 276 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 D1
port 5 nsew
flabel corelocali s 799 94 833 128 0 FreeSans 340 0 0 0 X
port 10 nsew
flabel corelocali s 799 168 833 202 0 FreeSans 340 0 0 0 X
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 960 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1720424
string GDS_START 1712122
<< end >>
