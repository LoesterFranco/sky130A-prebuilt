magic
tech sky130A
magscale 1 2
timestamp 1604502741
<< locali >>
rect 123 424 189 547
rect 123 390 427 424
rect 25 270 217 356
rect 283 286 359 356
rect 393 330 427 390
rect 393 252 455 330
rect 601 326 743 356
rect 533 260 743 326
rect 793 270 935 356
rect 985 270 1127 356
rect 337 236 455 252
rect 123 218 455 236
rect 123 202 387 218
rect 123 80 189 202
rect 337 119 387 202
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 23 581 289 615
rect 23 390 89 581
rect 223 492 289 581
rect 323 530 427 649
rect 461 492 527 596
rect 223 458 527 492
rect 561 458 627 649
rect 461 424 527 458
rect 661 424 727 596
rect 761 458 827 649
rect 861 424 934 600
rect 968 458 1034 649
rect 1068 424 1129 600
rect 461 390 1129 424
rect 461 364 527 390
rect 23 17 89 236
rect 893 226 1129 236
rect 235 85 301 168
rect 593 184 659 216
rect 421 150 659 184
rect 705 202 1129 226
rect 705 170 927 202
rect 421 85 471 150
rect 791 116 857 136
rect 235 51 471 85
rect 507 66 857 116
rect 893 70 927 170
rect 963 17 1029 168
rect 1063 70 1129 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
rlabel locali s 283 286 359 356 6 A1
port 1 nsew signal input
rlabel locali s 601 326 743 356 6 A2
port 2 nsew signal input
rlabel locali s 533 260 743 326 6 A2
port 2 nsew signal input
rlabel locali s 793 270 935 356 6 A3
port 3 nsew signal input
rlabel locali s 985 270 1127 356 6 A4
port 4 nsew signal input
rlabel locali s 25 270 217 356 6 B1
port 5 nsew signal input
rlabel locali s 393 330 427 390 6 Y
port 6 nsew signal output
rlabel locali s 393 252 455 330 6 Y
port 6 nsew signal output
rlabel locali s 337 236 455 252 6 Y
port 6 nsew signal output
rlabel locali s 337 119 387 202 6 Y
port 6 nsew signal output
rlabel locali s 123 424 189 547 6 Y
port 6 nsew signal output
rlabel locali s 123 390 427 424 6 Y
port 6 nsew signal output
rlabel locali s 123 218 455 236 6 Y
port 6 nsew signal output
rlabel locali s 123 202 387 218 6 Y
port 6 nsew signal output
rlabel locali s 123 80 189 202 6 Y
port 6 nsew signal output
rlabel metal1 s 0 -49 1152 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 617 1152 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3088408
string GDS_START 3078574
<< end >>
