magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1380 561
rect 103 427 169 527
rect 291 439 364 527
rect 18 197 66 325
rect 103 17 169 89
rect 306 287 443 337
rect 297 17 363 181
rect 397 57 443 287
rect 680 427 740 527
rect 863 402 920 527
rect 1115 426 1185 527
rect 1042 221 1097 287
rect 1219 299 1272 491
rect 779 17 829 122
rect 1233 119 1272 299
rect 1306 297 1362 527
rect 1135 17 1169 109
rect 1212 51 1272 119
rect 1306 17 1362 177
rect 0 -17 1380 17
<< obsli1 >>
rect 35 393 69 493
rect 203 405 248 493
rect 496 451 646 485
rect 35 359 156 393
rect 122 278 156 359
rect 203 371 529 405
rect 122 212 168 278
rect 122 157 156 212
rect 35 123 156 157
rect 35 52 69 123
rect 203 52 256 371
rect 479 197 529 371
rect 612 265 646 451
rect 783 373 827 487
rect 687 368 827 373
rect 1002 379 1068 493
rect 687 307 947 368
rect 1002 345 1185 379
rect 612 231 836 265
rect 711 199 836 231
rect 870 199 947 307
rect 1151 265 1185 345
rect 479 163 645 197
rect 711 112 745 199
rect 870 123 917 199
rect 1151 187 1199 265
rect 986 153 1199 187
rect 986 124 1030 153
rect 559 78 745 112
rect 863 51 917 123
rect 967 58 1030 124
<< metal1 >>
rect 0 496 1380 592
rect 18 252 76 261
rect 1030 252 1088 261
rect 18 224 1088 252
rect 18 215 76 224
rect 1030 215 1088 224
rect 0 -48 1380 48
<< labels >>
rlabel locali s 397 57 443 287 6 GATE
port 1 nsew signal input
rlabel locali s 306 287 443 337 6 GATE
port 1 nsew signal input
rlabel locali s 1233 119 1272 299 6 GCLK
port 2 nsew signal output
rlabel locali s 1219 299 1272 491 6 GCLK
port 2 nsew signal output
rlabel locali s 1212 51 1272 119 6 GCLK
port 2 nsew signal output
rlabel locali s 18 197 66 325 6 CLK
port 3 nsew clock input
rlabel locali s 1042 221 1097 287 6 CLK
port 3 nsew clock input
rlabel metal1 s 1030 252 1088 261 6 CLK
port 3 nsew clock input
rlabel metal1 s 1030 215 1088 224 6 CLK
port 3 nsew clock input
rlabel metal1 s 18 252 76 261 6 CLK
port 3 nsew clock input
rlabel metal1 s 18 224 1088 252 6 CLK
port 3 nsew clock input
rlabel metal1 s 18 215 76 224 6 CLK
port 3 nsew clock input
rlabel locali s 1306 17 1362 177 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 1135 17 1169 109 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 779 17 829 122 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 297 17 363 181 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 103 17 169 89 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 1380 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1380 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 1306 297 1362 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 1115 426 1185 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 863 402 920 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 680 427 740 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 291 439 364 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 103 427 169 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 1380 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 1380 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1380 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2585946
string GDS_START 2575692
<< end >>
