magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 368 561
rect 31 326 75 487
rect 109 360 175 493
rect 209 326 247 487
rect 281 360 347 493
rect 31 292 351 326
rect 17 213 261 258
rect 295 179 351 292
rect 205 145 351 179
rect 112 17 171 122
rect 205 56 250 145
rect 284 17 350 111
rect 0 -17 368 17
<< metal1 >>
rect 0 496 368 592
rect 14 428 354 468
rect 108 416 166 428
rect 288 416 346 428
rect 0 -48 368 48
<< labels >>
rlabel locali s 17 213 261 258 6 A
port 1 nsew signal input
rlabel locali s 295 179 351 292 6 Y
port 2 nsew signal output
rlabel locali s 209 326 247 487 6 Y
port 2 nsew signal output
rlabel locali s 205 145 351 179 6 Y
port 2 nsew signal output
rlabel locali s 205 56 250 145 6 Y
port 2 nsew signal output
rlabel locali s 31 326 75 487 6 Y
port 2 nsew signal output
rlabel locali s 31 292 351 326 6 Y
port 2 nsew signal output
rlabel locali s 109 360 175 493 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 281 360 347 493 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 288 416 346 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 108 416 166 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 14 428 354 468 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 284 17 350 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 112 17 171 122 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 368 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 368 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 527 368 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 368 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 368 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2255326
string GDS_START 2250622
<< end >>
