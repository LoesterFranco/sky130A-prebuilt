magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 460 561
rect 32 435 86 527
rect 17 237 86 391
rect 222 367 324 527
rect 358 367 443 493
rect 188 216 254 323
rect 390 105 443 367
rect 190 17 278 105
rect 312 51 443 105
rect 0 -17 460 17
<< obsli1 >>
rect 120 427 173 493
rect 120 190 154 427
rect 37 182 154 190
rect 290 182 356 287
rect 37 139 356 182
rect 37 56 98 139
<< metal1 >>
rect 0 496 460 592
rect 0 -48 460 48
<< labels >>
rlabel locali s 17 237 86 391 6 A
port 1 nsew signal input
rlabel locali s 188 216 254 323 6 B
port 2 nsew signal input
rlabel locali s 390 105 443 367 6 X
port 3 nsew signal output
rlabel locali s 358 367 443 493 6 X
port 3 nsew signal output
rlabel locali s 312 51 443 105 6 X
port 3 nsew signal output
rlabel locali s 190 17 278 105 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 460 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 460 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 222 367 324 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 32 435 86 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 460 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 460 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 460 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3741638
string GDS_START 3737216
<< end >>
