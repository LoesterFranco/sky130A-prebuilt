magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 25 260 101 356
rect 357 405 423 471
rect 389 356 423 405
rect 389 225 461 356
rect 1561 394 1627 596
rect 1741 394 1807 596
rect 1561 360 1807 394
rect 1773 226 1807 360
rect 1564 192 1807 226
rect 1564 70 1630 192
rect 1740 70 1807 192
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 23 424 89 596
rect 129 458 163 649
rect 203 539 295 596
rect 331 573 365 649
rect 399 581 675 615
rect 743 586 809 649
rect 399 539 433 581
rect 641 552 675 581
rect 843 581 1191 615
rect 843 552 877 581
rect 203 505 433 539
rect 23 390 169 424
rect 135 310 169 390
rect 203 364 295 505
rect 261 310 295 364
rect 467 424 501 547
rect 541 497 607 547
rect 641 518 877 552
rect 563 484 607 497
rect 563 450 877 484
rect 467 390 529 424
rect 135 226 227 310
rect 23 192 227 226
rect 23 70 89 192
rect 125 17 159 158
rect 193 85 227 192
rect 261 244 353 310
rect 261 119 295 244
rect 495 248 529 390
rect 563 316 597 450
rect 631 350 775 416
rect 563 282 669 316
rect 495 214 599 248
rect 329 146 531 180
rect 329 85 363 146
rect 193 51 363 85
rect 397 17 463 112
rect 497 85 531 146
rect 565 119 599 214
rect 635 190 669 282
rect 635 124 707 190
rect 741 172 775 350
rect 811 326 877 450
rect 911 274 945 547
rect 979 308 1013 581
rect 1047 376 1081 547
rect 1125 410 1191 581
rect 1263 490 1330 649
rect 1364 378 1430 596
rect 1471 412 1521 649
rect 1667 428 1701 649
rect 1047 342 1172 376
rect 1258 362 1494 378
rect 979 274 1104 308
rect 809 240 945 274
rect 809 206 1004 240
rect 1038 230 1104 274
rect 1138 262 1172 342
rect 1226 344 1494 362
rect 1847 364 1897 649
rect 1226 296 1292 344
rect 1460 326 1494 344
rect 1360 278 1426 310
rect 1326 262 1426 278
rect 1138 244 1426 262
rect 1460 260 1733 326
rect 970 190 1004 206
rect 1138 228 1360 244
rect 1138 194 1172 228
rect 1460 210 1494 260
rect 1394 194 1494 210
rect 741 138 936 172
rect 741 85 775 138
rect 497 51 775 85
rect 818 17 868 104
rect 902 85 936 138
rect 970 119 1036 190
rect 1070 144 1172 194
rect 1133 85 1199 102
rect 902 51 1199 85
rect 1282 17 1332 194
rect 1378 176 1494 194
rect 1378 70 1428 176
rect 1464 17 1530 142
rect 1666 17 1700 158
rect 1842 17 1892 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
<< metal1 >>
rect 0 683 1920 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 0 617 1920 649
rect 0 17 1920 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
rect 0 -49 1920 -17
<< labels >>
rlabel locali s 389 356 423 405 6 D
port 1 nsew signal input
rlabel locali s 389 225 461 356 6 D
port 1 nsew signal input
rlabel locali s 357 405 423 471 6 D
port 1 nsew signal input
rlabel locali s 1773 226 1807 360 6 Q
port 2 nsew signal output
rlabel locali s 1741 394 1807 596 6 Q
port 2 nsew signal output
rlabel locali s 1740 70 1807 192 6 Q
port 2 nsew signal output
rlabel locali s 1564 192 1807 226 6 Q
port 2 nsew signal output
rlabel locali s 1564 70 1630 192 6 Q
port 2 nsew signal output
rlabel locali s 1561 394 1627 596 6 Q
port 2 nsew signal output
rlabel locali s 1561 360 1807 394 6 Q
port 2 nsew signal output
rlabel locali s 25 260 101 356 6 CLK
port 3 nsew clock input
rlabel metal1 s 0 -49 1920 49 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 617 1920 715 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1920 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3101088
string GDS_START 3086236
<< end >>
