magic
tech sky130A
magscale 1 2
timestamp 1604502705
<< nwell >>
rect -38 335 2822 704
rect -38 332 825 335
rect 1117 332 2822 335
rect 1601 311 1903 332
<< pwell >>
rect 0 0 2784 49
<< scnmos >>
rect 84 74 114 158
rect 282 81 312 165
rect 379 81 409 165
rect 515 81 545 165
rect 593 81 623 165
rect 685 81 715 165
rect 904 119 934 267
rect 1014 119 1044 267
rect 1204 119 1234 203
rect 1290 119 1320 203
rect 1367 119 1397 203
rect 1445 119 1475 203
rect 1629 74 1659 202
rect 1717 74 1747 202
rect 1936 74 1966 158
rect 2008 74 2038 158
rect 2094 74 2124 158
rect 2166 74 2196 158
rect 2378 74 2408 222
rect 2571 74 2601 184
rect 2669 74 2699 222
<< pmoshvt >>
rect 208 464 238 592
rect 308 464 338 592
rect 392 464 422 592
rect 482 464 512 592
rect 592 464 622 592
rect 706 464 736 592
rect 914 392 944 592
rect 1004 392 1034 592
rect 1212 457 1242 541
rect 1302 457 1332 541
rect 1374 457 1404 541
rect 1464 457 1494 541
rect 1694 347 1724 547
rect 1784 347 1814 547
rect 1939 489 1969 573
rect 2017 489 2047 573
rect 2144 489 2174 573
rect 2234 489 2264 573
rect 2370 368 2400 592
rect 2568 424 2598 592
rect 2672 368 2702 592
<< ndiff >>
rect 845 180 904 267
rect 27 133 84 158
rect 27 99 39 133
rect 73 99 84 133
rect 27 74 84 99
rect 114 133 171 158
rect 114 99 125 133
rect 159 99 171 133
rect 114 74 171 99
rect 225 141 282 165
rect 225 107 237 141
rect 271 107 282 141
rect 225 81 282 107
rect 312 81 379 165
rect 409 153 515 165
rect 409 119 470 153
rect 504 119 515 153
rect 409 81 515 119
rect 545 81 593 165
rect 623 130 685 165
rect 623 96 636 130
rect 670 96 685 130
rect 623 81 685 96
rect 715 130 772 165
rect 715 96 726 130
rect 760 96 772 130
rect 835 150 904 180
rect 835 116 847 150
rect 881 119 904 150
rect 934 134 1014 267
rect 934 119 957 134
rect 881 116 889 119
rect 835 98 889 116
rect 715 81 772 96
rect 949 100 957 119
rect 991 119 1014 134
rect 1044 241 1097 267
rect 1044 207 1055 241
rect 1089 207 1097 241
rect 1044 173 1097 207
rect 1044 139 1055 173
rect 1089 139 1097 173
rect 1044 119 1097 139
rect 1151 179 1204 203
rect 1151 145 1159 179
rect 1193 145 1204 179
rect 1151 119 1204 145
rect 1234 179 1290 203
rect 1234 145 1245 179
rect 1279 145 1290 179
rect 1234 119 1290 145
rect 1320 119 1367 203
rect 1397 119 1445 203
rect 1475 202 1600 203
rect 1475 119 1629 202
rect 991 100 999 119
rect 949 88 999 100
rect 1491 82 1629 119
rect 1491 48 1502 82
rect 1536 74 1629 82
rect 1659 179 1717 202
rect 1659 145 1672 179
rect 1706 145 1717 179
rect 1659 74 1717 145
rect 1747 158 1797 202
rect 1747 131 1936 158
rect 1747 97 1857 131
rect 1891 97 1936 131
rect 1747 74 1936 97
rect 1966 74 2008 158
rect 2038 133 2094 158
rect 2038 99 2049 133
rect 2083 99 2094 133
rect 2038 74 2094 99
rect 2124 74 2166 158
rect 2196 127 2253 158
rect 2196 93 2207 127
rect 2241 93 2253 127
rect 2196 74 2253 93
rect 2307 82 2378 222
rect 1536 48 1549 74
rect 2307 48 2318 82
rect 2352 74 2378 82
rect 2408 210 2464 222
rect 2408 176 2419 210
rect 2453 176 2464 210
rect 2616 210 2669 222
rect 2616 184 2624 210
rect 2408 120 2464 176
rect 2408 86 2419 120
rect 2453 86 2464 120
rect 2408 74 2464 86
rect 2518 146 2571 184
rect 2518 112 2526 146
rect 2560 112 2571 146
rect 2518 74 2571 112
rect 2601 176 2624 184
rect 2658 176 2669 210
rect 2601 120 2669 176
rect 2601 86 2624 120
rect 2658 86 2669 120
rect 2601 74 2669 86
rect 2699 210 2756 222
rect 2699 176 2710 210
rect 2744 176 2756 210
rect 2699 120 2756 176
rect 2699 86 2710 120
rect 2744 86 2756 120
rect 2699 74 2756 86
rect 2352 48 2363 74
rect 1491 36 1549 48
rect 2307 36 2363 48
<< pdiff >>
rect 27 579 208 592
rect 27 545 39 579
rect 73 545 161 579
rect 195 545 208 579
rect 27 510 208 545
rect 27 476 39 510
rect 73 476 161 510
rect 195 476 208 510
rect 27 464 208 476
rect 238 584 308 592
rect 238 550 261 584
rect 295 550 308 584
rect 238 512 308 550
rect 238 478 261 512
rect 295 478 308 512
rect 238 464 308 478
rect 338 464 392 592
rect 422 584 482 592
rect 422 550 435 584
rect 469 550 482 584
rect 422 512 482 550
rect 422 478 435 512
rect 469 478 482 512
rect 422 464 482 478
rect 512 464 592 592
rect 622 580 706 592
rect 622 546 635 580
rect 669 546 706 580
rect 622 464 706 546
rect 736 580 795 592
rect 736 546 749 580
rect 783 546 795 580
rect 736 512 795 546
rect 736 478 749 512
rect 783 478 795 512
rect 736 464 795 478
rect 855 434 914 592
rect 855 400 867 434
rect 901 400 914 434
rect 855 392 914 400
rect 944 584 1004 592
rect 944 550 957 584
rect 991 550 1004 584
rect 944 392 1004 550
rect 1034 443 1093 592
rect 1034 409 1047 443
rect 1081 409 1093 443
rect 1034 392 1093 409
rect 2065 582 2126 594
rect 2065 573 2078 582
rect 1880 547 1939 573
rect 1153 516 1212 541
rect 1153 482 1165 516
rect 1199 482 1212 516
rect 1153 457 1212 482
rect 1242 528 1302 541
rect 1242 494 1255 528
rect 1289 494 1302 528
rect 1242 457 1302 494
rect 1332 457 1374 541
rect 1404 533 1464 541
rect 1404 499 1417 533
rect 1451 499 1464 533
rect 1404 457 1464 499
rect 1494 523 1553 541
rect 1494 489 1507 523
rect 1541 489 1553 523
rect 1494 457 1553 489
rect 1637 535 1694 547
rect 1637 501 1647 535
rect 1681 501 1694 535
rect 1637 464 1694 501
rect 1637 430 1647 464
rect 1681 430 1694 464
rect 1637 393 1694 430
rect 1637 359 1647 393
rect 1681 359 1694 393
rect 1637 347 1694 359
rect 1724 535 1784 547
rect 1724 501 1737 535
rect 1771 501 1784 535
rect 1724 464 1784 501
rect 1724 430 1737 464
rect 1771 430 1784 464
rect 1724 393 1784 430
rect 1724 359 1737 393
rect 1771 359 1784 393
rect 1724 347 1784 359
rect 1814 535 1939 547
rect 1814 501 1892 535
rect 1926 501 1939 535
rect 1814 489 1939 501
rect 1969 489 2017 573
rect 2047 548 2078 573
rect 2112 573 2126 582
rect 2282 580 2370 592
rect 2282 573 2290 580
rect 2112 548 2144 573
rect 2047 489 2144 548
rect 2174 548 2234 573
rect 2174 514 2187 548
rect 2221 514 2234 548
rect 2174 489 2234 514
rect 2264 546 2290 573
rect 2324 546 2370 580
rect 2264 512 2370 546
rect 2264 489 2322 512
rect 1814 481 1869 489
rect 1814 447 1827 481
rect 1861 447 1869 481
rect 2310 478 2322 489
rect 2356 478 2370 512
rect 1814 401 1869 447
rect 1814 367 1827 401
rect 1861 367 1869 401
rect 1814 347 1869 367
rect 2310 444 2370 478
rect 2310 410 2322 444
rect 2356 410 2370 444
rect 2310 368 2370 410
rect 2400 580 2459 592
rect 2400 546 2413 580
rect 2447 546 2459 580
rect 2400 500 2459 546
rect 2400 466 2413 500
rect 2447 466 2459 500
rect 2400 428 2459 466
rect 2400 394 2413 428
rect 2447 394 2459 428
rect 2513 580 2568 592
rect 2513 546 2521 580
rect 2555 546 2568 580
rect 2513 470 2568 546
rect 2513 436 2521 470
rect 2555 436 2568 470
rect 2513 424 2568 436
rect 2598 580 2672 592
rect 2598 546 2618 580
rect 2652 546 2672 580
rect 2598 497 2672 546
rect 2598 463 2618 497
rect 2652 463 2672 497
rect 2598 424 2672 463
rect 2617 414 2672 424
rect 2400 368 2459 394
rect 2617 380 2625 414
rect 2659 380 2672 414
rect 2617 368 2672 380
rect 2702 580 2757 592
rect 2702 546 2715 580
rect 2749 546 2757 580
rect 2702 497 2757 546
rect 2702 463 2715 497
rect 2749 463 2757 497
rect 2702 414 2757 463
rect 2702 380 2715 414
rect 2749 380 2757 414
rect 2702 368 2757 380
<< ndiffc >>
rect 39 99 73 133
rect 125 99 159 133
rect 237 107 271 141
rect 470 119 504 153
rect 636 96 670 130
rect 726 96 760 130
rect 847 116 881 150
rect 957 100 991 134
rect 1055 207 1089 241
rect 1055 139 1089 173
rect 1159 145 1193 179
rect 1245 145 1279 179
rect 1502 48 1536 82
rect 1672 145 1706 179
rect 1857 97 1891 131
rect 2049 99 2083 133
rect 2207 93 2241 127
rect 2318 48 2352 82
rect 2419 176 2453 210
rect 2419 86 2453 120
rect 2526 112 2560 146
rect 2624 176 2658 210
rect 2624 86 2658 120
rect 2710 176 2744 210
rect 2710 86 2744 120
<< pdiffc >>
rect 39 545 73 579
rect 161 545 195 579
rect 39 476 73 510
rect 161 476 195 510
rect 261 550 295 584
rect 261 478 295 512
rect 435 550 469 584
rect 435 478 469 512
rect 635 546 669 580
rect 749 546 783 580
rect 749 478 783 512
rect 867 400 901 434
rect 957 550 991 584
rect 1047 409 1081 443
rect 1165 482 1199 516
rect 1255 494 1289 528
rect 1417 499 1451 533
rect 1507 489 1541 523
rect 1647 501 1681 535
rect 1647 430 1681 464
rect 1647 359 1681 393
rect 1737 501 1771 535
rect 1737 430 1771 464
rect 1737 359 1771 393
rect 1892 501 1926 535
rect 2078 548 2112 582
rect 2187 514 2221 548
rect 2290 546 2324 580
rect 1827 447 1861 481
rect 2322 478 2356 512
rect 1827 367 1861 401
rect 2322 410 2356 444
rect 2413 546 2447 580
rect 2413 466 2447 500
rect 2413 394 2447 428
rect 2521 546 2555 580
rect 2521 436 2555 470
rect 2618 546 2652 580
rect 2618 463 2652 497
rect 2625 380 2659 414
rect 2715 546 2749 580
rect 2715 463 2749 497
rect 2715 380 2749 414
<< poly >>
rect 208 592 238 618
rect 308 592 338 618
rect 392 592 422 618
rect 482 592 512 618
rect 592 592 622 618
rect 706 592 736 618
rect 914 592 944 618
rect 1004 592 1034 618
rect 1108 615 1817 645
rect 208 449 238 464
rect 308 449 338 464
rect 392 449 422 464
rect 482 449 512 464
rect 592 449 622 464
rect 706 449 736 464
rect 205 376 241 449
rect 305 376 341 449
rect 84 360 341 376
rect 84 326 137 360
rect 171 326 205 360
rect 239 326 273 360
rect 307 326 341 360
rect 84 310 341 326
rect 84 158 114 310
rect 389 262 425 449
rect 479 432 515 449
rect 467 416 533 432
rect 467 382 483 416
rect 517 382 533 416
rect 467 366 533 382
rect 577 406 643 449
rect 577 372 593 406
rect 627 372 643 406
rect 577 338 643 372
rect 213 246 279 262
rect 213 212 229 246
rect 263 226 279 246
rect 354 246 425 262
rect 469 302 535 318
rect 469 268 485 302
rect 519 268 535 302
rect 577 304 593 338
rect 627 304 643 338
rect 577 288 643 304
rect 685 432 739 449
rect 685 416 823 432
rect 685 382 773 416
rect 807 382 823 416
rect 685 370 823 382
rect 914 377 944 392
rect 685 366 819 370
rect 469 252 535 268
rect 263 212 312 226
rect 213 196 312 212
rect 354 212 370 246
rect 404 212 425 246
rect 354 196 425 212
rect 505 210 535 252
rect 282 165 312 196
rect 379 165 409 196
rect 505 180 545 210
rect 515 165 545 180
rect 593 165 623 288
rect 685 165 715 366
rect 904 324 944 377
rect 1004 375 1034 392
rect 1108 375 1138 615
rect 1212 541 1242 567
rect 1302 541 1332 615
rect 1374 541 1404 567
rect 1464 541 1494 567
rect 1694 547 1724 573
rect 1781 562 1817 615
rect 1939 573 1969 599
rect 2017 573 2047 599
rect 1784 547 1814 562
rect 1212 442 1242 457
rect 1209 375 1245 442
rect 1302 431 1332 457
rect 757 308 944 324
rect 757 274 773 308
rect 807 282 944 308
rect 990 344 1142 375
rect 990 310 1006 344
rect 1040 310 1142 344
rect 990 282 1142 310
rect 1184 359 1250 375
rect 1374 361 1404 457
rect 1464 442 1494 457
rect 1464 429 1542 442
rect 1464 409 1605 429
rect 1464 403 1555 409
rect 1504 375 1555 403
rect 1589 375 1605 409
rect 1184 325 1200 359
rect 1234 345 1250 359
rect 1367 345 1462 361
rect 1234 325 1320 345
rect 1184 309 1320 325
rect 807 274 823 282
rect 757 240 823 274
rect 904 267 934 282
rect 1014 267 1044 282
rect 1112 267 1142 282
rect 757 206 773 240
rect 807 206 823 240
rect 757 190 823 206
rect 904 93 934 119
rect 1112 223 1234 267
rect 1204 203 1234 223
rect 1290 203 1320 309
rect 1367 311 1412 345
rect 1446 311 1462 345
rect 1367 295 1462 311
rect 1504 359 1605 375
rect 1367 203 1397 295
rect 1504 253 1534 359
rect 2144 573 2174 599
rect 2234 573 2264 599
rect 2370 592 2400 618
rect 2568 592 2598 618
rect 2672 592 2702 618
rect 1939 474 1969 489
rect 2017 474 2047 489
rect 2144 474 2174 489
rect 2234 474 2264 489
rect 1936 446 1972 474
rect 1901 430 1972 446
rect 1901 396 1917 430
rect 1951 396 1972 430
rect 1901 380 1972 396
rect 2014 396 2050 474
rect 2141 444 2183 474
rect 2231 444 2285 474
rect 2153 402 2183 444
rect 2014 380 2105 396
rect 1694 332 1724 347
rect 1784 332 1814 347
rect 2014 346 2055 380
rect 2089 346 2105 380
rect 1691 319 1727 332
rect 1633 315 1727 319
rect 1445 223 1534 253
rect 1597 299 1727 315
rect 1781 302 1966 332
rect 2014 330 2105 346
rect 2147 386 2213 402
rect 2147 352 2163 386
rect 2197 352 2213 386
rect 2147 336 2213 352
rect 2255 337 2285 444
rect 2568 409 2598 424
rect 2370 353 2400 368
rect 2367 337 2403 353
rect 2565 337 2601 409
rect 2672 353 2702 368
rect 1597 265 1613 299
rect 1647 289 1727 299
rect 1647 265 1663 289
rect 1597 249 1663 265
rect 1445 203 1475 223
rect 1629 202 1659 249
rect 1717 231 1887 247
rect 1717 217 1837 231
rect 1717 202 1747 217
rect 1014 93 1044 119
rect 1204 93 1234 119
rect 1290 93 1320 119
rect 1367 93 1397 119
rect 84 48 114 74
rect 282 55 312 81
rect 379 55 409 81
rect 515 55 545 81
rect 593 55 623 81
rect 685 51 715 81
rect 1445 51 1475 119
rect 685 21 1475 51
rect 1821 197 1837 217
rect 1871 197 1887 231
rect 1821 181 1887 197
rect 1936 158 1966 302
rect 2008 300 2044 330
rect 2008 158 2038 300
rect 2147 282 2177 336
rect 2255 287 2601 337
rect 2669 326 2705 353
rect 2094 252 2177 282
rect 2219 271 2601 287
rect 2094 158 2124 252
rect 2219 237 2235 271
rect 2269 247 2408 271
rect 2269 237 2285 247
rect 2219 204 2285 237
rect 2378 222 2408 247
rect 2166 174 2285 204
rect 2166 158 2196 174
rect 1629 48 1659 74
rect 1717 48 1747 74
rect 1936 48 1966 74
rect 2008 48 2038 74
rect 2094 48 2124 74
rect 2166 48 2196 74
rect 2571 184 2601 271
rect 2643 310 2709 326
rect 2643 276 2659 310
rect 2693 276 2709 310
rect 2643 260 2709 276
rect 2669 222 2699 260
rect 2378 48 2408 74
rect 2571 48 2601 74
rect 2669 48 2699 74
<< polycont >>
rect 137 326 171 360
rect 205 326 239 360
rect 273 326 307 360
rect 483 382 517 416
rect 593 372 627 406
rect 229 212 263 246
rect 485 268 519 302
rect 593 304 627 338
rect 773 382 807 416
rect 370 212 404 246
rect 773 274 807 308
rect 1006 310 1040 344
rect 1555 375 1589 409
rect 1200 325 1234 359
rect 773 206 807 240
rect 1412 311 1446 345
rect 1917 396 1951 430
rect 2055 346 2089 380
rect 2163 352 2197 386
rect 1613 265 1647 299
rect 1837 197 1871 231
rect 2235 237 2269 271
rect 2659 276 2693 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 23 579 211 595
rect 23 545 39 579
rect 73 545 161 579
rect 195 545 211 579
rect 23 510 211 545
rect 23 476 39 510
rect 73 476 161 510
rect 195 476 211 510
rect 245 584 311 649
rect 245 550 261 584
rect 295 550 311 584
rect 245 512 311 550
rect 245 478 261 512
rect 295 478 311 512
rect 419 584 511 596
rect 419 550 435 584
rect 469 550 511 584
rect 419 520 511 550
rect 619 580 685 649
rect 619 546 635 580
rect 669 546 685 580
rect 733 580 799 596
rect 733 546 749 580
rect 783 546 799 580
rect 941 584 1007 649
rect 941 550 957 584
rect 991 550 1007 584
rect 733 524 799 546
rect 733 520 916 524
rect 419 512 589 520
rect 733 518 922 520
rect 733 517 926 518
rect 733 516 929 517
rect 1165 516 1215 545
rect 733 512 1165 516
rect 419 478 435 512
rect 469 478 749 512
rect 783 484 1165 512
rect 783 480 850 484
rect 911 483 1165 484
rect 914 482 1165 483
rect 1199 482 1215 516
rect 918 480 1215 482
rect 783 478 846 480
rect 23 444 211 476
rect 689 477 846 478
rect 923 477 1215 480
rect 1250 528 1371 545
rect 1250 494 1255 528
rect 1289 494 1371 528
rect 1250 477 1371 494
rect 689 466 757 477
rect 23 416 539 444
rect 23 410 483 416
rect 23 262 57 410
rect 473 382 483 410
rect 517 382 539 416
rect 121 360 359 376
rect 473 366 539 382
rect 587 406 653 430
rect 587 372 593 406
rect 627 372 653 406
rect 121 326 137 360
rect 171 326 205 360
rect 239 326 273 360
rect 307 332 359 360
rect 587 338 653 372
rect 307 326 545 332
rect 121 302 545 326
rect 121 298 485 302
rect 479 268 485 298
rect 519 268 545 302
rect 587 304 593 338
rect 627 304 653 338
rect 587 288 653 304
rect 23 246 279 262
rect 23 212 229 246
rect 263 212 279 246
rect 23 196 279 212
rect 313 246 420 262
rect 479 252 545 268
rect 313 212 370 246
rect 404 212 420 246
rect 689 218 723 466
rect 867 439 901 450
rect 1165 443 1215 477
rect 784 432 833 438
rect 757 424 833 432
rect 757 416 799 424
rect 757 382 773 416
rect 807 382 833 390
rect 757 366 833 382
rect 867 434 997 439
rect 901 400 997 434
rect 867 360 997 400
rect 1031 409 1047 443
rect 1081 409 1126 443
rect 1165 409 1303 443
rect 1031 391 1126 409
rect 963 355 997 360
rect 1090 375 1126 391
rect 1090 359 1235 375
rect 963 344 1056 355
rect 23 133 73 196
rect 313 162 420 212
rect 454 184 723 218
rect 757 308 929 326
rect 757 274 773 308
rect 807 274 929 308
rect 757 240 929 274
rect 757 206 773 240
rect 807 236 929 240
rect 963 310 1006 344
rect 1040 310 1056 344
rect 963 291 1056 310
rect 1090 325 1200 359
rect 1234 325 1235 359
rect 1090 309 1235 325
rect 807 206 812 236
rect 757 184 812 206
rect 963 202 1009 291
rect 1090 257 1126 309
rect 1269 274 1303 409
rect 23 99 39 133
rect 23 70 73 99
rect 109 133 175 162
rect 109 99 125 133
rect 159 99 175 133
rect 109 17 175 99
rect 221 141 271 162
rect 221 107 237 141
rect 454 153 520 184
rect 454 119 470 153
rect 504 119 520 153
rect 846 168 1009 202
rect 1043 241 1126 257
rect 1043 207 1055 241
rect 1089 214 1126 241
rect 1160 240 1303 274
rect 1337 433 1371 477
rect 1405 533 1453 649
rect 1405 499 1417 533
rect 1451 499 1453 533
rect 1405 469 1453 499
rect 1487 523 1553 549
rect 1487 489 1507 523
rect 1541 489 1553 523
rect 1487 464 1553 489
rect 1647 535 1697 649
rect 2061 582 2130 649
rect 1681 501 1697 535
rect 1647 464 1697 501
rect 1487 433 1521 464
rect 1337 397 1521 433
rect 1681 430 1697 464
rect 1089 207 1124 214
rect 1043 173 1124 207
rect 1160 199 1195 240
rect 1337 206 1371 397
rect 846 150 907 168
rect 612 130 682 150
rect 221 85 271 107
rect 612 96 636 130
rect 670 96 682 130
rect 612 85 682 96
rect 221 51 682 85
rect 718 130 776 150
rect 718 96 726 130
rect 760 96 776 130
rect 827 116 847 150
rect 881 116 907 150
rect 1043 139 1055 173
rect 1089 139 1124 173
rect 827 100 907 116
rect 941 100 957 134
rect 991 100 1007 134
rect 718 17 776 96
rect 941 17 1007 100
rect 1043 85 1124 139
rect 1159 179 1195 199
rect 1193 145 1195 179
rect 1159 119 1195 145
rect 1229 179 1371 206
rect 1405 345 1453 361
rect 1405 311 1412 345
rect 1446 311 1453 345
rect 1405 218 1453 311
rect 1487 309 1521 397
rect 1555 424 1607 430
rect 1555 409 1567 424
rect 1601 390 1607 424
rect 1589 375 1607 390
rect 1555 359 1607 375
rect 1647 393 1697 430
rect 1681 359 1697 393
rect 1647 343 1697 359
rect 1737 535 1787 551
rect 1771 501 1787 535
rect 1737 464 1787 501
rect 1771 430 1787 464
rect 1737 393 1787 430
rect 1771 359 1787 393
rect 1487 299 1663 309
rect 1487 265 1613 299
rect 1647 265 1663 299
rect 1737 283 1787 359
rect 1821 535 2019 551
rect 1821 501 1892 535
rect 1926 501 2019 535
rect 2061 548 2078 582
rect 2112 548 2130 582
rect 2274 580 2363 649
rect 2061 532 2130 548
rect 2171 548 2237 577
rect 1821 485 2019 501
rect 2171 514 2187 548
rect 2221 514 2237 548
rect 2274 546 2290 580
rect 2324 546 2363 580
rect 2274 539 2363 546
rect 2171 498 2237 514
rect 2317 512 2363 539
rect 1821 481 1865 485
rect 1821 447 1827 481
rect 1861 447 1865 481
rect 1821 401 1865 447
rect 1821 367 1827 401
rect 1861 367 1865 401
rect 1821 351 1865 367
rect 1901 430 1951 446
rect 1901 396 1917 430
rect 1901 315 1951 396
rect 1487 252 1663 265
rect 1697 249 1787 283
rect 1821 269 1951 315
rect 1985 287 2019 485
rect 2053 464 2281 498
rect 2053 380 2105 464
rect 2053 346 2055 380
rect 2089 346 2105 380
rect 2053 330 2105 346
rect 2139 424 2213 430
rect 2139 390 2143 424
rect 2177 390 2213 424
rect 2139 386 2213 390
rect 2139 352 2163 386
rect 2197 352 2213 386
rect 2139 337 2213 352
rect 2247 360 2281 464
rect 2317 478 2322 512
rect 2356 478 2363 512
rect 2317 444 2363 478
rect 2317 410 2322 444
rect 2356 410 2363 444
rect 2317 394 2363 410
rect 2403 580 2469 596
rect 2403 546 2413 580
rect 2447 546 2469 580
rect 2403 500 2469 546
rect 2403 466 2413 500
rect 2447 466 2469 500
rect 2403 428 2469 466
rect 2403 394 2413 428
rect 2447 394 2469 428
rect 2247 326 2369 360
rect 1985 271 2285 287
rect 1697 218 1731 249
rect 1405 184 1731 218
rect 1821 231 1887 269
rect 1985 237 2235 271
rect 2269 237 2285 271
rect 1985 235 2285 237
rect 1821 215 1837 231
rect 1229 145 1245 179
rect 1279 172 1371 179
rect 1654 179 1731 184
rect 1279 145 1294 172
rect 1229 119 1294 145
rect 1410 116 1620 150
rect 1654 145 1672 179
rect 1706 145 1731 179
rect 1654 119 1731 145
rect 1765 197 1837 215
rect 1871 197 1887 231
rect 1765 181 1887 197
rect 1921 201 2285 235
rect 1410 85 1444 116
rect 1043 51 1444 85
rect 1586 85 1620 116
rect 1765 85 1799 181
rect 1921 147 1955 201
rect 1486 48 1502 82
rect 1536 48 1552 82
rect 1586 51 1799 85
rect 1833 131 1955 147
rect 1833 97 1857 131
rect 1891 97 1955 131
rect 1833 81 1955 97
rect 2033 133 2099 152
rect 2335 150 2369 326
rect 2033 99 2049 133
rect 2083 99 2099 133
rect 1486 17 1552 48
rect 2033 17 2099 99
rect 2191 127 2369 150
rect 2191 93 2207 127
rect 2241 116 2369 127
rect 2403 210 2469 394
rect 2403 176 2419 210
rect 2453 176 2469 210
rect 2403 120 2469 176
rect 2241 93 2257 116
rect 2191 70 2257 93
rect 2403 86 2419 120
rect 2453 86 2469 120
rect 2514 580 2571 596
rect 2514 546 2521 580
rect 2555 546 2571 580
rect 2514 470 2571 546
rect 2514 436 2521 470
rect 2555 436 2571 470
rect 2514 326 2571 436
rect 2609 580 2665 649
rect 2609 546 2618 580
rect 2652 546 2665 580
rect 2609 497 2665 546
rect 2609 463 2618 497
rect 2652 463 2665 497
rect 2609 414 2665 463
rect 2609 380 2625 414
rect 2659 380 2665 414
rect 2609 364 2665 380
rect 2711 580 2767 596
rect 2711 546 2715 580
rect 2749 546 2767 580
rect 2711 497 2767 546
rect 2711 463 2715 497
rect 2749 463 2767 497
rect 2711 414 2767 463
rect 2711 380 2715 414
rect 2749 380 2767 414
rect 2711 364 2767 380
rect 2514 310 2697 326
rect 2514 276 2659 310
rect 2693 276 2697 310
rect 2514 260 2697 276
rect 2514 146 2571 260
rect 2733 226 2767 364
rect 2514 112 2526 146
rect 2560 112 2571 146
rect 2514 91 2571 112
rect 2624 210 2658 226
rect 2624 120 2658 176
rect 2302 48 2318 82
rect 2352 48 2368 82
rect 2403 70 2469 86
rect 2302 17 2368 48
rect 2624 17 2658 86
rect 2694 210 2767 226
rect 2694 176 2710 210
rect 2744 176 2767 210
rect 2694 120 2767 176
rect 2694 86 2710 120
rect 2744 86 2767 120
rect 2694 70 2767 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 799 416 833 424
rect 799 390 807 416
rect 807 390 833 416
rect 1567 409 1601 424
rect 1567 390 1589 409
rect 1589 390 1601 409
rect 2143 390 2177 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
<< metal1 >>
rect 0 683 2784 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 0 617 2784 649
rect 787 424 845 430
rect 787 390 799 424
rect 833 421 845 424
rect 1555 424 1613 430
rect 1555 421 1567 424
rect 833 393 1567 421
rect 833 390 845 393
rect 787 384 845 390
rect 1555 390 1567 393
rect 1601 421 1613 424
rect 2131 424 2189 430
rect 2131 421 2143 424
rect 1601 393 2143 421
rect 1601 390 1613 393
rect 1555 384 1613 390
rect 2131 390 2143 393
rect 2177 390 2189 424
rect 2131 384 2189 390
rect 0 17 2784 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
rect 0 -49 2784 -17
<< labels >>
rlabel comment s 0 0 0 0 4 sdfrbp_1
flabel comment s 1484 630 1484 630 0 FreeSans 300 0 0 0 no_jumper_check
flabel comment s 1070 36 1070 36 0 FreeSans 300 0 0 0 no_jumper_check
flabel pwell s 0 0 2784 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 0 617 2784 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 2143 390 2177 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew
flabel metal1 s 0 617 2784 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 2784 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 2431 390 2465 424 0 FreeSans 340 0 0 0 Q_N
port 11 nsew
flabel corelocali s 2431 464 2465 498 0 FreeSans 340 0 0 0 Q_N
port 11 nsew
flabel corelocali s 2431 538 2465 572 0 FreeSans 340 0 0 0 Q_N
port 11 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 799 242 833 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 SCD
port 4 nsew
flabel corelocali s 607 390 641 424 0 FreeSans 340 0 0 0 SCD
port 4 nsew
flabel corelocali s 319 168 353 202 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 2719 168 2753 202 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2719 390 2753 424 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2719 464 2753 498 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2719 538 2753 572 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2719 94 2753 128 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2431 94 2465 128 0 FreeSans 340 0 0 0 Q_N
port 11 nsew
flabel corelocali s 2431 168 2465 202 0 FreeSans 340 0 0 0 Q_N
port 11 nsew
flabel corelocali s 2431 242 2465 276 0 FreeSans 340 0 0 0 Q_N
port 11 nsew
flabel corelocali s 2431 316 2465 350 0 FreeSans 340 0 0 0 Q_N
port 11 nsew
<< properties >>
string FIXED_BBOX 0 0 2784 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 96944
string GDS_START 74194
<< end >>
