magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 25 270 110 356
rect 217 364 303 430
rect 223 226 257 364
rect 223 70 289 226
rect 409 236 505 310
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 23 498 89 540
rect 130 532 196 649
rect 327 532 452 649
rect 583 532 649 649
rect 23 464 627 498
rect 23 390 178 464
rect 144 236 178 390
rect 337 374 559 430
rect 23 202 178 236
rect 337 326 371 374
rect 593 326 627 464
rect 291 260 371 326
rect 23 70 89 202
rect 123 17 189 168
rect 337 202 371 260
rect 553 260 627 326
rect 578 202 644 226
rect 337 168 644 202
rect 323 17 480 120
rect 578 70 644 168
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel locali s 25 270 110 356 6 A_N
port 1 nsew signal input
rlabel locali s 409 236 505 310 6 B
port 2 nsew signal input
rlabel locali s 223 226 257 364 6 X
port 3 nsew signal output
rlabel locali s 223 70 289 226 6 X
port 3 nsew signal output
rlabel locali s 217 364 303 430 6 X
port 3 nsew signal output
rlabel metal1 s 0 -49 672 49 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 617 672 715 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3861426
string GDS_START 3855976
<< end >>
