magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 460 561
rect 17 299 69 527
rect 103 333 169 493
rect 203 367 237 527
rect 271 333 337 493
rect 371 367 422 527
rect 103 299 443 333
rect 17 215 169 265
rect 203 215 353 265
rect 387 181 443 299
rect 119 17 153 109
rect 271 131 443 181
rect 0 -17 460 17
<< obsli1 >>
rect 17 143 237 177
rect 17 51 85 143
rect 187 93 237 143
rect 355 93 421 97
rect 187 51 421 93
<< metal1 >>
rect 0 496 460 592
rect 0 -48 460 48
<< labels >>
rlabel locali s 203 215 353 265 6 A
port 1 nsew signal input
rlabel locali s 17 215 169 265 6 B
port 2 nsew signal input
rlabel locali s 387 181 443 299 6 Y
port 3 nsew signal output
rlabel locali s 271 333 337 493 6 Y
port 3 nsew signal output
rlabel locali s 271 131 443 181 6 Y
port 3 nsew signal output
rlabel locali s 103 333 169 493 6 Y
port 3 nsew signal output
rlabel locali s 103 299 443 333 6 Y
port 3 nsew signal output
rlabel locali s 119 17 153 109 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 460 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 460 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 371 367 422 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 203 367 237 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 17 299 69 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 460 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 460 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 460 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1604838
string GDS_START 1599858
<< end >>
