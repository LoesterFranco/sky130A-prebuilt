magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 873 323 923 425
rect 1049 323 1103 425
rect 307 289 795 323
rect 307 257 341 289
rect 20 215 341 257
rect 375 215 685 255
rect 719 215 795 289
rect 829 283 1103 323
rect 829 181 873 283
rect 1309 215 1614 255
rect 1688 215 1993 255
rect 385 145 1119 181
rect 385 129 659 145
rect 855 55 931 145
rect 1043 55 1119 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 17 325 85 493
rect 129 359 171 527
rect 215 393 263 493
rect 309 427 359 527
rect 403 393 453 493
rect 497 427 547 527
rect 591 393 641 493
rect 685 427 735 527
rect 779 459 1213 493
rect 779 393 829 459
rect 215 359 829 393
rect 215 325 263 359
rect 17 291 263 325
rect 967 359 1015 459
rect 1137 291 1213 459
rect 1251 325 1317 493
rect 1361 359 1403 527
rect 1448 325 1496 493
rect 1541 359 1591 527
rect 1635 459 2062 493
rect 1635 325 1685 459
rect 1251 291 1685 325
rect 1729 325 1779 425
rect 1823 359 1873 459
rect 1917 325 1967 425
rect 2012 359 2062 459
rect 1729 291 2092 325
rect 907 215 1265 249
rect 1231 181 1265 215
rect 2027 181 2092 291
rect 35 17 69 179
rect 103 145 351 181
rect 103 51 179 145
rect 223 17 257 111
rect 291 95 351 145
rect 1231 147 2092 181
rect 291 51 743 95
rect 787 17 821 111
rect 975 17 1009 111
rect 1335 145 1975 147
rect 1163 17 1301 111
rect 1335 51 1411 145
rect 1455 17 1489 111
rect 1523 51 1599 145
rect 1643 17 1677 111
rect 1711 51 1787 145
rect 1831 17 1865 111
rect 1899 51 1975 145
rect 2019 17 2053 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
<< metal1 >>
rect 0 561 2116 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 0 496 2116 527
rect 0 17 2116 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
rect 0 -48 2116 -17
<< labels >>
rlabel locali s 1309 215 1614 255 6 A1_N
port 1 nsew signal input
rlabel locali s 1688 215 1993 255 6 A2_N
port 2 nsew signal input
rlabel locali s 719 215 795 289 6 B1
port 3 nsew signal input
rlabel locali s 307 289 795 323 6 B1
port 3 nsew signal input
rlabel locali s 307 257 341 289 6 B1
port 3 nsew signal input
rlabel locali s 20 215 341 257 6 B1
port 3 nsew signal input
rlabel locali s 375 215 685 255 6 B2
port 4 nsew signal input
rlabel locali s 1049 323 1103 425 6 Y
port 5 nsew signal output
rlabel locali s 1043 55 1119 145 6 Y
port 5 nsew signal output
rlabel locali s 873 323 923 425 6 Y
port 5 nsew signal output
rlabel locali s 855 55 931 145 6 Y
port 5 nsew signal output
rlabel locali s 829 283 1103 323 6 Y
port 5 nsew signal output
rlabel locali s 829 181 873 283 6 Y
port 5 nsew signal output
rlabel locali s 385 145 1119 181 6 Y
port 5 nsew signal output
rlabel locali s 385 129 659 145 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -48 2116 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 2116 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2116 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1363674
string GDS_START 1348580
<< end >>
