magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 189 236 263 430
rect 365 270 455 356
rect 189 70 255 236
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 23 547 165 649
rect 23 364 84 547
rect 279 532 345 649
rect 386 498 457 576
rect 121 464 457 498
rect 121 326 155 464
rect 21 260 155 326
rect 297 236 331 464
rect 386 390 457 464
rect 103 17 153 226
rect 297 202 457 236
rect 289 17 355 168
rect 391 90 457 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< metal1 >>
rect 0 683 480 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 0 617 480 649
rect 0 17 480 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
rect 0 -49 480 -17
<< labels >>
rlabel locali s 365 270 455 356 6 A
port 1 nsew signal input
rlabel locali s 189 236 263 430 6 X
port 2 nsew signal output
rlabel locali s 189 70 255 236 6 X
port 2 nsew signal output
rlabel metal1 s 0 -49 480 49 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 617 480 715 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 480 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3225700
string GDS_START 3221008
<< end >>
