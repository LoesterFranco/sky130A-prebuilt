magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1656 561
rect 119 367 153 527
rect 831 425 865 527
rect 1193 367 1227 527
rect 1261 333 1327 493
rect 1361 367 1395 527
rect 1429 333 1495 493
rect 1529 367 1580 527
rect 1261 299 1627 333
rect 30 215 156 255
rect 214 215 340 255
rect 402 215 525 255
rect 774 215 846 255
rect 958 215 1052 255
rect 1529 181 1627 299
rect 103 17 509 93
rect 1193 17 1227 177
rect 1261 143 1627 181
rect 1261 51 1327 143
rect 1361 17 1395 109
rect 1429 51 1495 143
rect 1529 17 1580 109
rect 0 -17 1656 17
<< obsli1 >>
rect 17 333 85 493
rect 187 459 421 493
rect 187 333 253 459
rect 17 289 253 333
rect 287 338 321 409
rect 355 372 421 459
rect 459 459 693 493
rect 459 338 525 459
rect 287 289 525 338
rect 559 255 593 409
rect 627 289 693 459
rect 731 391 797 493
rect 899 457 1139 493
rect 899 391 965 457
rect 731 357 965 391
rect 731 289 797 357
rect 1005 323 1039 423
rect 880 289 1039 323
rect 1073 289 1139 457
rect 559 221 729 255
rect 17 127 593 177
rect 691 161 729 221
rect 880 161 924 289
rect 1104 249 1227 253
rect 1104 215 1495 249
rect 1104 161 1155 215
rect 691 127 1155 161
rect 17 51 69 127
rect 543 93 593 127
rect 543 51 1139 93
<< metal1 >>
rect 0 496 1656 592
rect 0 -48 1656 48
<< labels >>
rlabel locali s 30 215 156 255 6 A1
port 1 nsew signal input
rlabel locali s 214 215 340 255 6 A2
port 2 nsew signal input
rlabel locali s 402 215 525 255 6 A3
port 3 nsew signal input
rlabel locali s 774 215 846 255 6 B1
port 4 nsew signal input
rlabel locali s 958 215 1052 255 6 B2
port 5 nsew signal input
rlabel locali s 1529 181 1627 299 6 X
port 6 nsew signal output
rlabel locali s 1429 333 1495 493 6 X
port 6 nsew signal output
rlabel locali s 1429 51 1495 143 6 X
port 6 nsew signal output
rlabel locali s 1261 333 1327 493 6 X
port 6 nsew signal output
rlabel locali s 1261 299 1627 333 6 X
port 6 nsew signal output
rlabel locali s 1261 143 1627 181 6 X
port 6 nsew signal output
rlabel locali s 1261 51 1327 143 6 X
port 6 nsew signal output
rlabel locali s 1529 17 1580 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1361 17 1395 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1193 17 1227 177 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 103 17 509 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 1656 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1656 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1529 367 1580 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1361 367 1395 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1193 367 1227 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 831 425 865 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 119 367 153 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 1656 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 1656 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1656 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 924904
string GDS_START 912656
<< end >>
