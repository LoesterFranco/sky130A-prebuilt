magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 129 367 177 527
rect 18 215 94 263
rect 223 323 257 493
rect 291 367 367 527
rect 411 323 445 493
rect 223 289 445 323
rect 479 297 555 527
rect 384 181 445 289
rect 223 147 445 181
rect 105 17 163 113
rect 223 51 257 147
rect 291 17 367 113
rect 411 51 445 147
rect 479 17 555 177
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< obsli1 >>
rect 19 331 85 493
rect 19 297 172 331
rect 138 249 172 297
rect 138 215 248 249
rect 138 181 172 215
rect 35 147 172 181
rect 35 51 69 147
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 18 215 94 263 6 A
port 1 nsew signal input
rlabel locali s 411 323 445 493 6 X
port 2 nsew signal output
rlabel locali s 411 51 445 147 6 X
port 2 nsew signal output
rlabel locali s 384 181 445 289 6 X
port 2 nsew signal output
rlabel locali s 223 323 257 493 6 X
port 2 nsew signal output
rlabel locali s 223 289 445 323 6 X
port 2 nsew signal output
rlabel locali s 223 147 445 181 6 X
port 2 nsew signal output
rlabel locali s 223 51 257 147 6 X
port 2 nsew signal output
rlabel viali s 581 -17 615 17 8 VGND
port 3 nsew ground bidirectional
rlabel viali s 489 -17 523 17 8 VGND
port 3 nsew ground bidirectional
rlabel viali s 397 -17 431 17 8 VGND
port 3 nsew ground bidirectional
rlabel viali s 305 -17 339 17 8 VGND
port 3 nsew ground bidirectional
rlabel viali s 213 -17 247 17 8 VGND
port 3 nsew ground bidirectional
rlabel viali s 121 -17 155 17 8 VGND
port 3 nsew ground bidirectional
rlabel viali s 29 -17 63 17 8 VGND
port 3 nsew ground bidirectional
rlabel locali s 479 17 555 177 6 VGND
port 3 nsew ground bidirectional
rlabel locali s 291 17 367 113 6 VGND
port 3 nsew ground bidirectional
rlabel locali s 105 17 163 113 6 VGND
port 3 nsew ground bidirectional
rlabel locali s 0 -17 644 17 8 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 -48 644 48 8 VGND
port 3 nsew ground bidirectional
rlabel viali s 581 527 615 561 6 VPWR
port 4 nsew power bidirectional
rlabel viali s 489 527 523 561 6 VPWR
port 4 nsew power bidirectional
rlabel viali s 397 527 431 561 6 VPWR
port 4 nsew power bidirectional
rlabel viali s 305 527 339 561 6 VPWR
port 4 nsew power bidirectional
rlabel viali s 213 527 247 561 6 VPWR
port 4 nsew power bidirectional
rlabel viali s 121 527 155 561 6 VPWR
port 4 nsew power bidirectional
rlabel viali s 29 527 63 561 6 VPWR
port 4 nsew power bidirectional
rlabel locali s 479 297 555 527 6 VPWR
port 4 nsew power bidirectional
rlabel locali s 291 367 367 527 6 VPWR
port 4 nsew power bidirectional
rlabel locali s 129 367 177 527 6 VPWR
port 4 nsew power bidirectional
rlabel locali s 0 527 644 561 6 VPWR
port 4 nsew power bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 4 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1666920
string GDS_START 1661252
<< end >>
