magic
tech sky130A
magscale 1 2
timestamp 1599588209
<< nwell >>
rect -38 332 2726 704
rect 280 330 587 332
<< pwell >>
rect 0 0 2688 49
<< scpmos >>
rect 85 508 115 592
rect 175 508 205 592
rect 374 366 404 590
rect 464 366 494 590
rect 669 463 699 547
rect 759 463 789 547
rect 837 463 867 547
rect 959 463 989 547
rect 1230 392 1260 592
rect 1320 392 1350 592
rect 1597 493 1627 577
rect 1681 493 1711 577
rect 1789 493 1819 577
rect 1879 493 1909 577
rect 1980 409 2010 577
rect 2070 409 2100 577
rect 2171 368 2201 592
rect 2270 368 2300 592
rect 2455 368 2485 592
rect 2545 368 2575 592
<< nmoslvt >>
rect 94 78 124 162
rect 172 78 202 162
rect 370 74 400 222
rect 484 74 514 222
rect 682 138 712 222
rect 782 138 812 222
rect 860 138 890 222
rect 938 138 968 222
rect 1122 74 1152 222
rect 1407 74 1437 222
rect 1617 81 1647 165
rect 1695 81 1725 165
rect 1797 81 1827 165
rect 1875 81 1905 165
rect 2087 74 2117 222
rect 2285 74 2315 222
rect 2390 74 2420 222
rect 2490 74 2520 222
rect 2576 74 2606 222
<< ndiff >>
rect 313 210 370 222
rect 313 176 325 210
rect 359 176 370 210
rect 37 137 94 162
rect 37 103 49 137
rect 83 103 94 137
rect 37 78 94 103
rect 124 78 172 162
rect 202 137 259 162
rect 202 103 213 137
rect 247 103 259 137
rect 202 78 259 103
rect 313 120 370 176
rect 313 86 325 120
rect 359 86 370 120
rect 313 74 370 86
rect 400 132 484 222
rect 400 98 425 132
rect 459 98 484 132
rect 400 74 484 98
rect 514 132 571 222
rect 625 197 682 222
rect 625 163 637 197
rect 671 163 682 197
rect 625 138 682 163
rect 712 189 782 222
rect 712 155 737 189
rect 771 155 782 189
rect 712 138 782 155
rect 812 138 860 222
rect 890 138 938 222
rect 968 138 1122 222
rect 514 98 525 132
rect 559 98 571 132
rect 514 74 571 98
rect 983 74 1122 138
rect 1152 194 1407 222
rect 1152 160 1163 194
rect 1197 160 1255 194
rect 1289 160 1348 194
rect 1382 160 1407 194
rect 1152 74 1407 160
rect 1437 165 1487 222
rect 2016 210 2087 222
rect 2016 176 2028 210
rect 2062 176 2087 210
rect 1437 153 1617 165
rect 1437 119 1448 153
rect 1482 119 1537 153
rect 1571 119 1617 153
rect 1437 81 1617 119
rect 1647 81 1695 165
rect 1725 140 1797 165
rect 1725 106 1741 140
rect 1775 106 1797 140
rect 1725 81 1797 106
rect 1827 81 1875 165
rect 1905 140 1962 165
rect 1905 106 1916 140
rect 1950 106 1962 140
rect 1905 81 1962 106
rect 2016 120 2087 176
rect 2016 86 2028 120
rect 2062 86 2087 120
rect 1437 74 1487 81
rect 983 40 995 74
rect 1029 40 1041 74
rect 2016 74 2087 86
rect 2117 210 2174 222
rect 2117 176 2128 210
rect 2162 176 2174 210
rect 2117 120 2174 176
rect 2117 86 2128 120
rect 2162 86 2174 120
rect 2117 74 2174 86
rect 2228 210 2285 222
rect 2228 176 2240 210
rect 2274 176 2285 210
rect 2228 123 2285 176
rect 2228 89 2240 123
rect 2274 89 2285 123
rect 2228 74 2285 89
rect 2315 210 2390 222
rect 2315 176 2335 210
rect 2369 176 2390 210
rect 2315 123 2390 176
rect 2315 89 2335 123
rect 2369 89 2390 123
rect 2315 74 2390 89
rect 2420 123 2490 222
rect 2420 89 2431 123
rect 2465 89 2490 123
rect 2420 74 2490 89
rect 2520 210 2576 222
rect 2520 176 2531 210
rect 2565 176 2576 210
rect 2520 120 2576 176
rect 2520 86 2531 120
rect 2565 86 2576 120
rect 2520 74 2576 86
rect 2606 204 2661 222
rect 2606 170 2617 204
rect 2651 170 2661 204
rect 2606 120 2661 170
rect 2606 86 2617 120
rect 2651 86 2661 120
rect 2606 74 2661 86
rect 983 28 1041 40
<< pdiff >>
rect 27 567 85 592
rect 27 533 38 567
rect 72 533 85 567
rect 27 508 85 533
rect 115 567 175 592
rect 115 533 128 567
rect 162 533 175 567
rect 115 508 175 533
rect 205 580 262 592
rect 205 546 218 580
rect 252 546 262 580
rect 205 508 262 546
rect 316 412 374 590
rect 316 378 327 412
rect 361 378 374 412
rect 316 366 374 378
rect 404 574 464 590
rect 404 540 417 574
rect 451 540 464 574
rect 404 366 464 540
rect 494 415 551 590
rect 494 381 507 415
rect 541 381 551 415
rect 494 366 551 381
rect 885 582 941 594
rect 885 548 896 582
rect 930 548 941 582
rect 885 547 941 548
rect 611 522 669 547
rect 611 488 622 522
rect 656 488 669 522
rect 611 463 669 488
rect 699 532 759 547
rect 699 498 712 532
rect 746 498 759 532
rect 699 463 759 498
rect 789 463 837 547
rect 867 463 959 547
rect 989 522 1047 547
rect 989 488 1002 522
rect 1036 488 1047 522
rect 989 463 1047 488
rect 1162 583 1230 592
rect 1162 549 1182 583
rect 1216 549 1230 583
rect 1162 540 1230 549
rect 1177 392 1230 540
rect 1260 442 1320 592
rect 1260 408 1273 442
rect 1307 408 1320 442
rect 1260 392 1320 408
rect 1350 577 1403 592
rect 2118 577 2171 592
rect 1350 545 1597 577
rect 1350 511 1432 545
rect 1466 511 1550 545
rect 1584 511 1597 545
rect 1350 493 1597 511
rect 1627 493 1681 577
rect 1711 552 1789 577
rect 1711 518 1732 552
rect 1766 518 1789 552
rect 1711 493 1789 518
rect 1819 552 1879 577
rect 1819 518 1832 552
rect 1866 518 1879 552
rect 1819 493 1879 518
rect 1909 552 1980 577
rect 1909 518 1930 552
rect 1964 518 1980 552
rect 1909 493 1980 518
rect 1350 392 1403 493
rect 1927 409 1980 493
rect 2010 565 2070 577
rect 2010 531 2023 565
rect 2057 531 2070 565
rect 2010 455 2070 531
rect 2010 421 2023 455
rect 2057 421 2070 455
rect 2010 409 2070 421
rect 2100 565 2171 577
rect 2100 531 2123 565
rect 2157 531 2171 565
rect 2100 455 2171 531
rect 2100 421 2123 455
rect 2157 421 2171 455
rect 2100 409 2171 421
rect 2118 368 2171 409
rect 2201 580 2270 592
rect 2201 546 2223 580
rect 2257 546 2270 580
rect 2201 497 2270 546
rect 2201 463 2223 497
rect 2257 463 2270 497
rect 2201 414 2270 463
rect 2201 380 2223 414
rect 2257 380 2270 414
rect 2201 368 2270 380
rect 2300 580 2455 592
rect 2300 546 2314 580
rect 2348 546 2407 580
rect 2441 546 2455 580
rect 2300 478 2455 546
rect 2300 444 2314 478
rect 2348 444 2407 478
rect 2441 444 2455 478
rect 2300 368 2455 444
rect 2485 580 2545 592
rect 2485 546 2498 580
rect 2532 546 2545 580
rect 2485 497 2545 546
rect 2485 463 2498 497
rect 2532 463 2545 497
rect 2485 414 2545 463
rect 2485 380 2498 414
rect 2532 380 2545 414
rect 2485 368 2545 380
rect 2575 580 2644 592
rect 2575 546 2598 580
rect 2632 546 2644 580
rect 2575 510 2644 546
rect 2575 476 2598 510
rect 2632 476 2644 510
rect 2575 440 2644 476
rect 2575 406 2598 440
rect 2632 406 2644 440
rect 2575 368 2644 406
<< ndiffc >>
rect 325 176 359 210
rect 49 103 83 137
rect 213 103 247 137
rect 325 86 359 120
rect 425 98 459 132
rect 637 163 671 197
rect 737 155 771 189
rect 525 98 559 132
rect 1163 160 1197 194
rect 1255 160 1289 194
rect 1348 160 1382 194
rect 2028 176 2062 210
rect 1448 119 1482 153
rect 1537 119 1571 153
rect 1741 106 1775 140
rect 1916 106 1950 140
rect 2028 86 2062 120
rect 995 40 1029 74
rect 2128 176 2162 210
rect 2128 86 2162 120
rect 2240 176 2274 210
rect 2240 89 2274 123
rect 2335 176 2369 210
rect 2335 89 2369 123
rect 2431 89 2465 123
rect 2531 176 2565 210
rect 2531 86 2565 120
rect 2617 170 2651 204
rect 2617 86 2651 120
<< pdiffc >>
rect 38 533 72 567
rect 128 533 162 567
rect 218 546 252 580
rect 327 378 361 412
rect 417 540 451 574
rect 507 381 541 415
rect 896 548 930 582
rect 622 488 656 522
rect 712 498 746 532
rect 1002 488 1036 522
rect 1182 549 1216 583
rect 1273 408 1307 442
rect 1432 511 1466 545
rect 1550 511 1584 545
rect 1732 518 1766 552
rect 1832 518 1866 552
rect 1930 518 1964 552
rect 2023 531 2057 565
rect 2023 421 2057 455
rect 2123 531 2157 565
rect 2123 421 2157 455
rect 2223 546 2257 580
rect 2223 463 2257 497
rect 2223 380 2257 414
rect 2314 546 2348 580
rect 2407 546 2441 580
rect 2314 444 2348 478
rect 2407 444 2441 478
rect 2498 546 2532 580
rect 2498 463 2532 497
rect 2498 380 2532 414
rect 2598 546 2632 580
rect 2598 476 2632 510
rect 2598 406 2632 440
<< poly >>
rect 85 592 115 618
rect 175 592 205 618
rect 374 590 404 616
rect 464 590 494 616
rect 566 615 1092 645
rect 85 493 115 508
rect 175 493 205 508
rect 82 470 118 493
rect 82 402 124 470
rect 44 386 124 402
rect 44 352 60 386
rect 94 352 124 386
rect 44 318 124 352
rect 44 284 60 318
rect 94 284 124 318
rect 44 250 124 284
rect 44 216 60 250
rect 94 216 124 250
rect 44 200 124 216
rect 94 162 124 200
rect 172 428 208 493
rect 172 412 264 428
rect 172 378 214 412
rect 248 378 264 412
rect 172 344 264 378
rect 374 351 404 366
rect 464 351 494 366
rect 172 310 214 344
rect 248 310 264 344
rect 371 328 407 351
rect 461 348 497 351
rect 566 348 596 615
rect 669 547 699 573
rect 756 562 792 615
rect 759 547 789 562
rect 837 547 867 573
rect 959 547 989 573
rect 1062 508 1092 615
rect 1230 592 1260 618
rect 1320 592 1350 618
rect 1062 492 1145 508
rect 669 448 699 463
rect 666 378 702 448
rect 759 437 789 463
rect 837 448 867 463
rect 959 448 989 463
rect 1062 458 1095 492
rect 1129 458 1145 492
rect 834 421 870 448
rect 834 405 914 421
rect 172 276 264 310
rect 172 242 214 276
rect 248 242 264 276
rect 353 312 419 328
rect 353 278 369 312
rect 403 278 419 312
rect 353 262 419 278
rect 461 318 596 348
rect 638 362 704 378
rect 638 328 654 362
rect 688 348 704 362
rect 834 371 864 405
rect 898 371 914 405
rect 834 355 914 371
rect 956 400 992 448
rect 1062 442 1145 458
rect 956 384 1083 400
rect 1597 577 1627 603
rect 1681 577 1711 603
rect 1789 577 1819 603
rect 1879 577 1909 603
rect 1980 577 2010 603
rect 2070 577 2100 603
rect 2171 592 2201 618
rect 2270 592 2300 618
rect 2455 592 2485 618
rect 2545 592 2575 618
rect 1597 478 1627 493
rect 1681 478 1711 493
rect 1789 478 1819 493
rect 1879 478 1909 493
rect 1594 461 1630 478
rect 1548 445 1630 461
rect 1548 411 1564 445
rect 1598 411 1630 445
rect 1548 395 1630 411
rect 1678 425 1714 478
rect 1786 455 1822 478
rect 1762 439 1828 455
rect 1678 395 1719 425
rect 688 328 790 348
rect 638 318 790 328
rect 461 294 545 318
rect 638 312 704 318
rect 172 226 264 242
rect 172 162 202 226
rect 370 222 400 262
rect 461 260 495 294
rect 529 270 545 294
rect 760 307 790 318
rect 760 277 812 307
rect 529 260 712 270
rect 461 240 712 260
rect 484 222 514 240
rect 682 222 712 240
rect 782 222 812 277
rect 860 222 890 355
rect 956 350 1033 384
rect 1067 350 1083 384
rect 1230 377 1260 392
rect 1320 377 1350 392
rect 956 334 1083 350
rect 1227 346 1263 377
rect 1317 347 1353 377
rect 962 267 992 334
rect 1227 310 1257 346
rect 1317 318 1647 347
rect 1131 294 1257 310
rect 1131 274 1147 294
rect 938 237 992 267
rect 1122 260 1147 274
rect 1181 260 1257 294
rect 1122 244 1257 260
rect 1299 317 1647 318
rect 1299 302 1365 317
rect 1299 268 1315 302
rect 1349 268 1365 302
rect 1299 252 1365 268
rect 1407 253 1575 269
rect 938 222 968 237
rect 1122 222 1152 244
rect 1407 239 1525 253
rect 1407 222 1437 239
rect 94 52 124 78
rect 172 52 202 78
rect 682 112 712 138
rect 782 112 812 138
rect 860 112 890 138
rect 938 112 968 138
rect 1509 219 1525 239
rect 1559 219 1575 253
rect 1509 203 1575 219
rect 1617 165 1647 317
rect 1689 273 1719 395
rect 1762 405 1778 439
rect 1812 405 1828 439
rect 1762 389 1828 405
rect 1689 257 1755 273
rect 1689 223 1705 257
rect 1739 223 1755 257
rect 1689 207 1755 223
rect 1695 165 1725 207
rect 1797 165 1827 389
rect 1876 341 1912 478
rect 1980 394 2010 409
rect 2070 394 2100 409
rect 1977 341 2013 394
rect 2067 341 2103 394
rect 2171 353 2201 368
rect 2270 353 2300 368
rect 2455 353 2485 368
rect 2545 353 2575 368
rect 1869 325 2103 341
rect 1869 291 1885 325
rect 1919 311 2103 325
rect 1919 291 1935 311
rect 1869 275 1935 291
rect 1875 165 1905 275
rect 2073 267 2103 311
rect 2168 326 2204 353
rect 2267 326 2303 353
rect 2452 326 2488 353
rect 2542 326 2578 353
rect 2168 310 2606 326
rect 2168 296 2262 310
rect 2246 276 2262 296
rect 2296 276 2330 310
rect 2364 276 2398 310
rect 2432 296 2606 310
rect 2432 276 2448 296
rect 2073 237 2117 267
rect 2246 260 2448 276
rect 2087 222 2117 237
rect 2285 222 2315 260
rect 2390 222 2420 260
rect 2490 222 2520 296
rect 2576 222 2606 296
rect 370 48 400 74
rect 484 48 514 74
rect 1122 48 1152 74
rect 1407 48 1437 74
rect 1617 55 1647 81
rect 1695 55 1725 81
rect 1797 55 1827 81
rect 1875 55 1905 81
rect 2087 48 2117 74
rect 2285 48 2315 74
rect 2390 48 2420 74
rect 2490 48 2520 74
rect 2576 48 2606 74
<< polycont >>
rect 60 352 94 386
rect 60 284 94 318
rect 60 216 94 250
rect 214 378 248 412
rect 214 310 248 344
rect 1095 458 1129 492
rect 214 242 248 276
rect 369 278 403 312
rect 654 328 688 362
rect 864 371 898 405
rect 1564 411 1598 445
rect 495 260 529 294
rect 1033 350 1067 384
rect 1147 260 1181 294
rect 1315 268 1349 302
rect 1525 219 1559 253
rect 1778 405 1812 439
rect 1705 223 1739 257
rect 1885 291 1919 325
rect 2262 276 2296 310
rect 2330 276 2364 310
rect 2398 276 2432 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2688 683
rect 22 567 72 649
rect 22 533 38 567
rect 22 504 72 533
rect 112 567 178 596
rect 112 533 128 567
rect 162 533 178 567
rect 112 504 178 533
rect 218 580 268 649
rect 252 546 268 580
rect 218 530 268 546
rect 401 574 467 649
rect 401 540 417 574
rect 451 540 467 574
rect 880 582 946 649
rect 401 536 467 540
rect 137 496 178 504
rect 606 522 672 551
rect 606 502 622 522
rect 302 496 622 502
rect 137 488 622 496
rect 656 488 672 522
rect 137 468 672 488
rect 712 532 762 551
rect 880 548 896 582
rect 930 548 946 582
rect 1166 583 1233 649
rect 746 514 762 532
rect 983 522 1036 551
rect 1166 549 1182 583
rect 1216 549 1233 583
rect 983 514 1002 522
rect 746 498 1002 514
rect 712 488 1002 498
rect 1425 545 1682 561
rect 712 480 1036 488
rect 137 462 336 468
rect 25 386 103 436
rect 25 352 60 386
rect 94 352 103 386
rect 25 318 103 352
rect 25 284 60 318
rect 94 284 103 318
rect 25 250 103 284
rect 25 216 60 250
rect 94 216 103 250
rect 25 200 103 216
rect 137 166 171 462
rect 606 446 672 468
rect 205 424 257 428
rect 205 412 223 424
rect 205 378 214 412
rect 248 378 257 390
rect 205 344 257 378
rect 205 310 214 344
rect 248 310 257 344
rect 205 276 257 310
rect 205 242 214 276
rect 248 242 257 276
rect 205 226 257 242
rect 291 412 361 428
rect 291 378 327 412
rect 291 362 361 378
rect 491 415 569 434
rect 491 381 507 415
rect 541 381 569 415
rect 606 412 759 446
rect 491 378 569 381
rect 491 362 691 378
rect 291 228 325 362
rect 409 328 455 356
rect 491 344 654 362
rect 359 312 455 328
rect 359 278 369 312
rect 403 278 455 312
rect 359 262 455 278
rect 489 294 535 310
rect 489 260 495 294
rect 529 260 535 294
rect 489 228 535 260
rect 291 210 535 228
rect 291 176 325 210
rect 359 194 535 210
rect 359 176 375 194
rect 33 137 171 166
rect 33 103 49 137
rect 83 132 171 137
rect 213 137 247 166
rect 83 103 99 132
rect 33 74 99 103
rect 213 17 247 103
rect 291 120 375 176
rect 569 160 603 344
rect 638 328 654 344
rect 688 328 691 362
rect 638 312 691 328
rect 725 278 759 412
rect 291 86 325 120
rect 359 86 375 120
rect 291 70 375 86
rect 409 132 475 160
rect 409 98 425 132
rect 459 98 475 132
rect 409 17 475 98
rect 509 132 603 160
rect 637 244 759 278
rect 637 197 687 244
rect 793 210 827 480
rect 949 459 1036 480
rect 1079 492 1391 515
rect 1425 511 1432 545
rect 1466 511 1550 545
rect 1584 511 1682 545
rect 1425 495 1682 511
rect 671 163 687 197
rect 637 134 687 163
rect 721 189 827 210
rect 721 155 737 189
rect 771 176 827 189
rect 861 405 914 421
rect 861 371 864 405
rect 898 371 914 405
rect 861 210 914 371
rect 949 300 983 459
rect 1079 458 1095 492
rect 1129 481 1391 492
rect 1129 458 1145 481
rect 1231 442 1323 447
rect 1017 390 1087 424
rect 1121 390 1127 424
rect 1017 384 1127 390
rect 1017 350 1033 384
rect 1067 350 1127 384
rect 1017 334 1127 350
rect 1231 408 1273 442
rect 1307 408 1323 442
rect 1231 388 1323 408
rect 949 294 1197 300
rect 949 260 1147 294
rect 1181 260 1197 294
rect 949 244 1197 260
rect 1231 210 1265 388
rect 1357 318 1391 481
rect 1299 302 1391 318
rect 1299 268 1315 302
rect 1349 268 1391 302
rect 1299 252 1391 268
rect 861 194 1398 210
rect 861 176 1163 194
rect 771 155 787 176
rect 721 134 787 155
rect 1147 160 1163 176
rect 1197 160 1255 194
rect 1289 160 1348 194
rect 1382 160 1398 194
rect 1147 144 1398 160
rect 1432 169 1466 495
rect 1548 445 1614 461
rect 1548 411 1564 445
rect 1598 411 1614 445
rect 1548 269 1614 411
rect 1648 341 1682 495
rect 1716 552 1782 649
rect 1716 518 1732 552
rect 1766 518 1782 552
rect 1716 489 1782 518
rect 1816 552 1896 581
rect 1816 518 1832 552
rect 1866 518 1896 552
rect 1816 489 1896 518
rect 1930 552 1980 649
rect 1964 518 1980 552
rect 1930 489 1980 518
rect 2023 565 2073 581
rect 2057 531 2073 565
rect 1753 439 1828 455
rect 1753 424 1778 439
rect 1753 390 1759 424
rect 1812 405 1828 439
rect 1793 390 1828 405
rect 1753 384 1828 390
rect 1862 409 1896 489
rect 2023 455 2073 531
rect 2057 421 2073 455
rect 1862 375 1989 409
rect 1648 325 1921 341
rect 1648 307 1885 325
rect 1869 291 1885 307
rect 1919 291 1921 325
rect 1869 275 1921 291
rect 1509 253 1655 269
rect 1509 219 1525 253
rect 1559 219 1655 253
rect 1509 203 1655 219
rect 1689 257 1755 273
rect 1689 223 1705 257
rect 1739 241 1755 257
rect 1955 241 1989 375
rect 2023 326 2073 421
rect 2107 565 2173 649
rect 2107 531 2123 565
rect 2157 531 2173 565
rect 2107 455 2173 531
rect 2107 421 2123 455
rect 2157 421 2173 455
rect 2107 405 2173 421
rect 2207 580 2273 596
rect 2207 546 2223 580
rect 2257 546 2273 580
rect 2207 497 2273 546
rect 2207 463 2223 497
rect 2257 463 2273 497
rect 2207 414 2273 463
rect 2307 580 2448 649
rect 2307 546 2314 580
rect 2348 546 2407 580
rect 2441 546 2448 580
rect 2307 478 2448 546
rect 2307 444 2314 478
rect 2348 444 2407 478
rect 2441 444 2448 478
rect 2307 428 2448 444
rect 2482 580 2548 596
rect 2482 546 2498 580
rect 2532 546 2548 580
rect 2482 497 2548 546
rect 2482 463 2498 497
rect 2532 463 2548 497
rect 2207 380 2223 414
rect 2257 394 2273 414
rect 2482 414 2548 463
rect 2482 394 2498 414
rect 2257 380 2498 394
rect 2532 380 2548 414
rect 2582 580 2648 649
rect 2582 546 2598 580
rect 2632 546 2648 580
rect 2582 510 2648 546
rect 2582 476 2598 510
rect 2632 476 2648 510
rect 2582 440 2648 476
rect 2582 406 2598 440
rect 2632 406 2648 440
rect 2582 390 2648 406
rect 2207 360 2548 380
rect 2482 356 2548 360
rect 2023 310 2448 326
rect 2482 322 2663 356
rect 2023 292 2262 310
rect 1739 223 1989 241
rect 2112 276 2262 292
rect 2296 276 2330 310
rect 2364 276 2398 310
rect 2432 276 2448 310
rect 2112 260 2448 276
rect 1689 207 1989 223
rect 2023 210 2078 226
rect 1432 153 1587 169
rect 509 98 525 132
rect 559 100 603 132
rect 861 108 1113 142
rect 1432 119 1448 153
rect 1482 119 1537 153
rect 1571 119 1587 153
rect 861 100 895 108
rect 559 98 895 100
rect 509 66 895 98
rect 1079 85 1113 108
rect 1621 85 1655 203
rect 979 40 995 74
rect 1029 40 1045 74
rect 1079 51 1655 85
rect 1725 140 1791 169
rect 1725 106 1741 140
rect 1775 106 1791 140
rect 979 17 1045 40
rect 1725 17 1791 106
rect 1900 140 1966 207
rect 1900 106 1916 140
rect 1950 106 1966 140
rect 1900 77 1966 106
rect 2023 176 2028 210
rect 2062 176 2078 210
rect 2023 120 2078 176
rect 2023 86 2028 120
rect 2062 86 2078 120
rect 2023 17 2078 86
rect 2112 210 2178 260
rect 2515 254 2663 322
rect 2515 226 2565 254
rect 2112 176 2128 210
rect 2162 176 2178 210
rect 2112 120 2178 176
rect 2112 86 2128 120
rect 2162 86 2178 120
rect 2112 70 2178 86
rect 2224 210 2282 226
rect 2224 176 2240 210
rect 2274 176 2282 210
rect 2224 123 2282 176
rect 2224 89 2240 123
rect 2274 89 2282 123
rect 2224 17 2282 89
rect 2319 210 2565 226
rect 2319 176 2335 210
rect 2369 176 2531 210
rect 2319 123 2382 176
rect 2319 89 2335 123
rect 2369 89 2382 123
rect 2319 73 2382 89
rect 2416 123 2481 142
rect 2416 89 2431 123
rect 2465 89 2481 123
rect 2416 17 2481 89
rect 2515 120 2565 176
rect 2515 86 2531 120
rect 2515 70 2565 86
rect 2601 204 2667 220
rect 2601 170 2617 204
rect 2651 170 2667 204
rect 2601 120 2667 170
rect 2601 86 2617 120
rect 2651 86 2667 120
rect 2601 17 2667 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2688 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 223 412 257 424
rect 223 390 248 412
rect 248 390 257 412
rect 1087 390 1121 424
rect 1759 405 1778 424
rect 1778 405 1793 424
rect 1759 390 1793 405
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
<< metal1 >>
rect 0 683 2688 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2688 683
rect 0 617 2688 649
rect 211 424 269 430
rect 211 390 223 424
rect 257 421 269 424
rect 1075 424 1133 430
rect 1075 421 1087 424
rect 257 393 1087 421
rect 257 390 269 393
rect 211 384 269 390
rect 1075 390 1087 393
rect 1121 421 1133 424
rect 1747 424 1805 430
rect 1747 421 1759 424
rect 1121 393 1759 421
rect 1121 390 1133 393
rect 1075 384 1133 390
rect 1747 390 1759 393
rect 1793 390 1805 424
rect 1747 384 1805 390
rect 0 17 2688 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2688 17
rect 0 -49 2688 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dfrtp_4
flabel comment s 731 633 731 633 0 FreeSans 200 0 0 0 no_jumper_check
flabel pwell s 0 0 2688 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 0 617 2688 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 223 390 257 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew
flabel metal1 s 0 617 2688 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 2688 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 31 390 65 424 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 2623 316 2657 350 0 FreeSans 340 0 0 0 Q
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 2688 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 2926364
string GDS_START 2907590
<< end >>
