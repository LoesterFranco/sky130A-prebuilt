magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 710 704
<< pwell >>
rect 0 0 672 49
<< scnmos >>
rect 98 74 128 222
rect 184 74 214 222
rect 298 74 328 222
rect 384 74 414 222
rect 558 74 588 222
<< pmoshvt >>
rect 89 368 119 592
rect 179 368 209 592
rect 269 368 299 592
rect 359 368 389 592
rect 466 368 496 536
rect 556 368 586 536
<< ndiff >>
rect 27 153 98 222
rect 27 119 39 153
rect 73 119 98 153
rect 27 74 98 119
rect 128 210 184 222
rect 128 176 139 210
rect 173 176 184 210
rect 128 120 184 176
rect 128 86 139 120
rect 173 86 184 120
rect 128 74 184 86
rect 214 131 298 222
rect 214 97 239 131
rect 273 97 298 131
rect 214 74 298 97
rect 328 210 384 222
rect 328 176 339 210
rect 373 176 384 210
rect 328 120 384 176
rect 328 86 339 120
rect 373 86 384 120
rect 328 74 384 86
rect 414 120 558 222
rect 414 86 469 120
rect 503 86 558 120
rect 414 74 558 86
rect 588 210 645 222
rect 588 176 599 210
rect 633 176 645 210
rect 588 120 645 176
rect 588 86 599 120
rect 633 86 645 120
rect 588 74 645 86
<< pdiff >>
rect 30 580 89 592
rect 30 546 42 580
rect 76 546 89 580
rect 30 497 89 546
rect 30 463 42 497
rect 76 463 89 497
rect 30 414 89 463
rect 30 380 42 414
rect 76 380 89 414
rect 30 368 89 380
rect 119 580 179 592
rect 119 546 132 580
rect 166 546 179 580
rect 119 497 179 546
rect 119 463 132 497
rect 166 463 179 497
rect 119 414 179 463
rect 119 380 132 414
rect 166 380 179 414
rect 119 368 179 380
rect 209 580 269 592
rect 209 546 222 580
rect 256 546 269 580
rect 209 462 269 546
rect 209 428 222 462
rect 256 428 269 462
rect 209 368 269 428
rect 299 580 359 592
rect 299 546 312 580
rect 346 546 359 580
rect 299 497 359 546
rect 299 463 312 497
rect 346 463 359 497
rect 299 414 359 463
rect 299 380 312 414
rect 346 380 359 414
rect 299 368 359 380
rect 389 580 448 592
rect 389 546 402 580
rect 436 546 448 580
rect 389 536 448 546
rect 389 497 466 536
rect 389 463 402 497
rect 436 463 466 497
rect 389 414 466 463
rect 389 380 402 414
rect 436 380 466 414
rect 389 368 466 380
rect 496 440 556 536
rect 496 406 509 440
rect 543 406 556 440
rect 496 368 556 406
rect 586 524 645 536
rect 586 490 599 524
rect 633 490 645 524
rect 586 368 645 490
<< ndiffc >>
rect 39 119 73 153
rect 139 176 173 210
rect 139 86 173 120
rect 239 97 273 131
rect 339 176 373 210
rect 339 86 373 120
rect 469 86 503 120
rect 599 176 633 210
rect 599 86 633 120
<< pdiffc >>
rect 42 546 76 580
rect 42 463 76 497
rect 42 380 76 414
rect 132 546 166 580
rect 132 463 166 497
rect 132 380 166 414
rect 222 546 256 580
rect 222 428 256 462
rect 312 546 346 580
rect 312 463 346 497
rect 312 380 346 414
rect 402 546 436 580
rect 402 463 436 497
rect 402 380 436 414
rect 509 406 543 440
rect 599 490 633 524
<< poly >>
rect 89 592 119 618
rect 179 592 209 618
rect 269 592 299 618
rect 359 592 389 618
rect 466 536 496 562
rect 556 536 586 562
rect 89 353 119 368
rect 179 353 209 368
rect 269 353 299 368
rect 359 353 389 368
rect 466 353 496 368
rect 556 353 586 368
rect 86 290 122 353
rect 176 326 212 353
rect 266 326 302 353
rect 356 326 392 353
rect 463 336 499 353
rect 553 336 589 353
rect 176 310 414 326
rect 176 290 228 310
rect 86 276 228 290
rect 262 276 296 310
rect 330 276 364 310
rect 398 276 414 310
rect 463 320 589 336
rect 463 306 531 320
rect 86 260 414 276
rect 515 286 531 306
rect 565 286 589 320
rect 515 270 589 286
rect 98 222 128 260
rect 184 222 214 260
rect 298 222 328 260
rect 384 222 414 260
rect 558 222 588 270
rect 98 48 128 74
rect 184 48 214 74
rect 298 48 328 74
rect 384 48 414 74
rect 558 48 588 74
<< polycont >>
rect 228 276 262 310
rect 296 276 330 310
rect 364 276 398 310
rect 531 286 565 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 26 580 92 649
rect 26 546 42 580
rect 76 546 92 580
rect 26 497 92 546
rect 26 463 42 497
rect 76 463 92 497
rect 26 414 92 463
rect 26 380 42 414
rect 76 380 92 414
rect 26 364 92 380
rect 132 580 167 596
rect 166 546 167 580
rect 132 497 167 546
rect 166 463 167 497
rect 132 414 167 463
rect 206 580 272 649
rect 206 546 222 580
rect 256 546 272 580
rect 206 462 272 546
rect 206 428 222 462
rect 256 428 272 462
rect 312 580 346 596
rect 312 497 346 546
rect 166 394 167 414
rect 312 414 346 463
rect 166 380 312 394
rect 132 360 346 380
rect 386 580 452 649
rect 386 546 402 580
rect 436 546 452 580
rect 386 497 452 546
rect 386 463 402 497
rect 436 463 452 497
rect 583 524 649 649
rect 583 490 599 524
rect 633 490 649 524
rect 583 474 649 490
rect 386 414 452 463
rect 386 380 402 414
rect 436 380 452 414
rect 493 406 509 440
rect 543 406 649 440
rect 493 390 649 406
rect 386 364 452 380
rect 132 282 167 360
rect 121 236 167 282
rect 212 310 457 326
rect 212 276 228 310
rect 262 276 296 310
rect 330 276 364 310
rect 398 276 457 310
rect 212 260 457 276
rect 505 320 581 356
rect 505 286 531 320
rect 565 286 581 320
rect 505 270 581 286
rect 123 226 167 236
rect 423 226 457 260
rect 615 226 649 390
rect 123 210 389 226
rect 23 153 89 202
rect 23 119 39 153
rect 73 119 89 153
rect 23 17 89 119
rect 123 176 139 210
rect 173 192 339 210
rect 173 176 189 192
rect 123 120 189 176
rect 323 176 339 192
rect 373 176 389 210
rect 423 210 649 226
rect 423 192 599 210
rect 123 86 139 120
rect 173 86 189 120
rect 123 70 189 86
rect 223 131 289 158
rect 223 97 239 131
rect 273 97 289 131
rect 223 17 289 97
rect 323 120 389 176
rect 583 176 599 192
rect 633 176 649 210
rect 323 86 339 120
rect 373 86 389 120
rect 323 70 389 86
rect 423 120 549 136
rect 423 86 469 120
rect 503 86 549 120
rect 423 17 549 86
rect 583 120 649 176
rect 583 86 599 120
rect 633 86 649 120
rect 583 70 649 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel comment s 0 0 0 0 4 buf_4
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew
flabel nbase s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 127 242 161 276 0 FreeSans 340 0 0 0 X
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 672 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3231474
string GDS_START 3225754
<< end >>
