magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 460 561
rect 229 367 295 527
rect 329 369 436 493
rect 29 153 100 265
rect 202 153 255 265
rect 373 165 436 369
rect 50 17 98 119
rect 236 17 279 119
rect 313 51 436 165
rect 0 -17 460 17
<< obsli1 >>
rect 54 333 132 368
rect 54 299 339 333
rect 134 119 168 299
rect 305 199 339 299
rect 134 53 190 119
<< metal1 >>
rect 0 496 460 592
rect 0 -48 460 48
<< labels >>
rlabel locali s 202 153 255 265 6 A
port 1 nsew signal input
rlabel locali s 29 153 100 265 6 B
port 2 nsew signal input
rlabel locali s 373 165 436 369 6 X
port 3 nsew signal output
rlabel locali s 329 369 436 493 6 X
port 3 nsew signal output
rlabel locali s 313 51 436 165 6 X
port 3 nsew signal output
rlabel locali s 236 17 279 119 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 50 17 98 119 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 460 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 460 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 229 367 295 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 460 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 460 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 460 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 999018
string GDS_START 994852
<< end >>
