magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 552 561
rect 113 367 175 527
rect 209 401 261 493
rect 295 435 346 527
rect 381 401 433 493
rect 209 367 433 401
rect 85 151 155 265
rect 381 317 433 367
rect 467 353 524 527
rect 381 283 532 317
rect 451 181 532 283
rect 202 147 532 181
rect 111 17 166 113
rect 202 69 261 147
rect 295 17 346 113
rect 381 69 433 147
rect 467 17 523 113
rect 0 -17 552 17
<< obsli1 >>
rect 17 333 79 493
rect 17 299 223 333
rect 17 117 51 299
rect 189 249 223 299
rect 189 215 417 249
rect 17 51 77 117
<< metal1 >>
rect 0 496 552 592
rect 0 -48 552 48
<< labels >>
rlabel locali s 85 151 155 265 6 A
port 1 nsew signal input
rlabel locali s 451 181 532 283 6 X
port 2 nsew signal output
rlabel locali s 381 401 433 493 6 X
port 2 nsew signal output
rlabel locali s 381 317 433 367 6 X
port 2 nsew signal output
rlabel locali s 381 283 532 317 6 X
port 2 nsew signal output
rlabel locali s 381 69 433 147 6 X
port 2 nsew signal output
rlabel locali s 209 401 261 493 6 X
port 2 nsew signal output
rlabel locali s 209 367 433 401 6 X
port 2 nsew signal output
rlabel locali s 202 147 532 181 6 X
port 2 nsew signal output
rlabel locali s 202 69 261 147 6 X
port 2 nsew signal output
rlabel locali s 467 17 523 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 295 17 346 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 111 17 166 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 0 -17 552 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 552 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 467 353 524 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 295 435 346 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 113 367 175 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 0 527 552 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 496 552 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 552 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3168094
string GDS_START 3162938
<< end >>
