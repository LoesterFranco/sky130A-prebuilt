magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< obsli1 >>
rect 0 1071 46920 1105
rect 388424 1071 412804 1105
rect 41 911 107 1071
rect 207 953 273 1033
rect 389 987 455 1071
rect 489 953 549 1037
rect 583 987 747 1071
rect 207 911 747 953
rect 781 949 847 1037
rect 881 983 935 1071
rect 969 949 1035 1037
rect 1069 983 1123 1071
rect 1157 949 1223 1037
rect 781 915 1223 949
rect 19 830 139 877
rect 173 830 307 877
rect 341 830 409 877
rect 105 796 139 830
rect 341 796 375 830
rect 19 728 71 796
rect 105 762 375 796
rect 409 728 455 796
rect 19 694 455 728
rect 19 595 85 694
rect 119 561 173 660
rect 207 595 273 694
rect 307 561 361 660
rect 395 629 455 694
rect 489 730 539 911
rect 713 881 747 911
rect 573 765 639 877
rect 713 833 1091 881
rect 1125 799 1175 915
rect 1257 907 1307 1071
rect 1397 926 1455 1071
rect 1513 911 1579 1071
rect 1679 953 1745 1033
rect 1861 987 1927 1071
rect 1961 953 2021 1037
rect 2055 987 2219 1071
rect 1679 911 2219 953
rect 2253 949 2319 1037
rect 2353 983 2407 1071
rect 2441 949 2507 1037
rect 2541 983 2595 1071
rect 2629 949 2695 1037
rect 2729 983 2783 1071
rect 2817 949 2883 1037
rect 2253 915 2883 949
rect 1491 830 1611 877
rect 1645 830 1779 877
rect 1813 830 1881 877
rect 489 663 549 730
rect 583 629 649 731
rect 395 595 649 629
rect 697 561 747 789
rect 787 765 1217 799
rect 787 595 841 765
rect 875 561 941 731
rect 975 595 1029 765
rect 1063 561 1129 731
rect 1163 595 1217 765
rect 1253 561 1319 799
rect 1577 796 1611 830
rect 1813 796 1847 830
rect 1397 561 1455 794
rect 1491 728 1543 796
rect 1577 762 1847 796
rect 1881 728 1927 796
rect 1491 694 1927 728
rect 1491 595 1557 694
rect 1591 561 1645 660
rect 1679 595 1745 694
rect 1779 561 1833 660
rect 1867 629 1927 694
rect 1961 730 2011 911
rect 2185 881 2219 911
rect 2045 765 2111 877
rect 2185 833 2699 881
rect 2781 799 2831 915
rect 2917 907 2967 1071
rect 3053 926 3111 1071
rect 3147 923 3213 1071
rect 3331 957 3397 1037
rect 3516 991 3582 1071
rect 3331 923 3589 957
rect 3145 823 3251 889
rect 3301 829 3435 889
rect 1961 663 2021 730
rect 2055 629 2121 731
rect 1867 595 2121 629
rect 2169 561 2219 789
rect 2259 765 2877 799
rect 2259 595 2313 765
rect 2347 561 2413 731
rect 2447 595 2501 765
rect 2535 561 2601 731
rect 2635 595 2689 765
rect 2723 561 2789 731
rect 2823 595 2877 765
rect 2915 561 2977 799
rect 3215 795 3251 823
rect 3469 823 3521 889
rect 3555 877 3589 923
rect 3623 945 3677 1037
rect 3711 979 3777 1071
rect 3811 945 3865 1037
rect 3899 979 3965 1071
rect 3999 945 4053 1037
rect 4087 979 4153 1071
rect 3623 911 4123 945
rect 4249 926 4307 1071
rect 4343 923 4409 1071
rect 4527 957 4593 1037
rect 4712 991 4778 1071
rect 4527 923 4785 957
rect 3555 835 3989 877
rect 3469 795 3505 823
rect 3053 561 3111 794
rect 3215 761 3505 795
rect 3555 727 3589 835
rect 4023 799 4123 911
rect 4341 823 4447 889
rect 4497 829 4631 889
rect 3147 561 3207 727
rect 3241 693 3589 727
rect 3623 765 4123 799
rect 4411 795 4447 823
rect 4665 823 4717 889
rect 4751 877 4785 923
rect 4819 945 4873 1037
rect 4907 979 4973 1071
rect 5007 945 5061 1037
rect 5095 979 5161 1071
rect 5195 945 5249 1037
rect 5283 979 5349 1071
rect 5383 945 5437 1037
rect 5471 979 5537 1071
rect 4819 911 5507 945
rect 5629 926 5687 1071
rect 5733 979 5783 1071
rect 4751 835 5389 877
rect 4665 795 4701 823
rect 3241 595 3301 693
rect 3335 561 3401 659
rect 3435 595 3489 693
rect 3523 561 3589 656
rect 3623 595 3677 765
rect 3711 561 3777 731
rect 3811 595 3865 765
rect 3899 561 3965 731
rect 3999 595 4053 765
rect 4087 561 4153 731
rect 4249 561 4307 794
rect 4411 761 4701 795
rect 4751 727 4785 835
rect 5423 799 5507 911
rect 5721 823 5783 945
rect 5817 873 5883 1035
rect 5917 966 5971 1071
rect 6005 941 6071 1037
rect 6105 975 6159 1071
rect 6193 941 6259 1037
rect 6293 975 6347 1071
rect 6381 941 6447 1037
rect 6481 975 6535 1071
rect 6005 907 6519 941
rect 6641 926 6699 1071
rect 6735 966 6801 1071
rect 6835 945 6889 1032
rect 6923 979 6989 1071
rect 7023 945 7077 1032
rect 7111 979 7177 1071
rect 6835 907 7077 945
rect 7211 945 7265 1032
rect 7299 979 7365 1071
rect 7399 945 7453 1032
rect 7487 979 7553 1071
rect 7587 945 7641 1032
rect 7675 979 7741 1071
rect 7775 945 7829 1032
rect 7863 979 7929 1071
rect 7963 945 8017 1032
rect 8051 979 8117 1071
rect 8151 945 8205 1032
rect 8239 966 8305 1071
rect 7211 907 8205 945
rect 8389 926 8447 1071
rect 8697 983 8831 1071
rect 8865 949 8919 1037
rect 8953 983 9019 1071
rect 9053 949 9107 1037
rect 9141 983 9207 1071
rect 9241 949 9295 1037
rect 9329 983 9395 1071
rect 9429 949 9483 1037
rect 9517 983 9583 1071
rect 9617 949 9671 1037
rect 9705 983 9771 1071
rect 9805 949 9859 1037
rect 9893 983 10027 1071
rect 5817 823 6382 873
rect 4343 561 4403 727
rect 4437 693 4785 727
rect 4819 765 5507 799
rect 4437 595 4497 693
rect 4531 561 4597 659
rect 4631 595 4685 693
rect 4719 561 4785 656
rect 4819 595 4873 765
rect 4907 561 4973 731
rect 5007 595 5061 765
rect 5095 561 5161 731
rect 5195 595 5249 765
rect 5283 561 5349 731
rect 5383 595 5437 765
rect 5471 561 5537 731
rect 5629 561 5687 794
rect 5723 561 5783 789
rect 5817 595 5883 823
rect 6453 789 6519 907
rect 7023 873 7077 907
rect 6821 827 6980 873
rect 7023 827 8053 873
rect 5917 561 5971 789
rect 6005 755 6519 789
rect 6005 596 6071 755
rect 6105 561 6159 721
rect 6193 596 6259 755
rect 6293 561 6347 721
rect 6381 596 6447 755
rect 6481 561 6535 721
rect 6641 561 6699 794
rect 7023 793 7077 827
rect 8108 793 8205 907
rect 8487 915 10195 949
rect 10321 926 10379 1071
rect 10415 1003 10857 1037
rect 8487 796 8521 915
rect 8555 830 10049 881
rect 10084 796 10195 915
rect 6830 789 7077 793
rect 6735 561 6795 789
rect 6829 755 7077 789
rect 6829 595 6895 755
rect 6929 561 6983 721
rect 7023 595 7077 755
rect 7111 561 7171 793
rect 7205 755 8205 793
rect 7205 595 7265 755
rect 7299 561 7365 721
rect 7399 595 7453 755
rect 7487 561 7553 721
rect 7587 595 7641 755
rect 7675 561 7741 721
rect 7775 595 7829 755
rect 7863 561 7929 721
rect 7963 595 8017 755
rect 8051 561 8117 721
rect 8151 595 8205 755
rect 8239 561 8305 795
rect 8389 561 8447 794
rect 8487 762 10195 796
rect 8483 561 8549 728
rect 8583 595 8637 762
rect 8671 561 8737 728
rect 8771 595 8825 762
rect 8859 561 8925 728
rect 8959 595 9013 762
rect 9047 561 9113 728
rect 9147 595 9201 762
rect 9235 561 9301 728
rect 9335 595 9389 762
rect 9423 561 9489 728
rect 9523 595 9577 762
rect 9611 561 9677 728
rect 9711 595 9765 762
rect 9799 561 9865 728
rect 9899 595 9953 762
rect 9987 561 10053 728
rect 10087 595 10141 762
rect 10175 561 10241 728
rect 10321 561 10379 794
rect 10415 629 10475 1003
rect 10609 979 10663 1003
rect 10797 978 10857 1003
rect 10901 978 10955 1071
rect 10509 943 10575 969
rect 10697 943 10763 969
rect 10989 943 11055 1037
rect 11089 979 11143 1071
rect 11177 943 11243 1037
rect 10509 907 11243 943
rect 11277 907 11331 1071
rect 11365 873 11431 1037
rect 11465 907 11519 1071
rect 11553 943 11619 1037
rect 11653 979 11707 1071
rect 11741 943 11807 1037
rect 11841 978 11895 1071
rect 11939 1003 12381 1037
rect 11939 978 11999 1003
rect 12133 979 12187 1003
rect 12033 943 12099 969
rect 12221 943 12287 969
rect 11553 907 12287 943
rect 12321 873 12381 1003
rect 12425 907 12479 1071
rect 12513 943 12579 1037
rect 12613 979 12667 1071
rect 12701 943 12767 1037
rect 12801 979 12855 1071
rect 12889 943 12955 1037
rect 12989 979 13043 1071
rect 13077 943 13143 1037
rect 13177 978 13231 1071
rect 13265 943 13331 1037
rect 13365 979 13419 1071
rect 13453 943 13519 1037
rect 12513 907 13519 943
rect 13553 907 13607 1071
rect 13725 926 13783 1071
rect 13819 1003 14261 1037
rect 10509 823 10779 873
rect 10981 823 11251 873
rect 11365 823 11815 873
rect 12017 823 12287 873
rect 12321 823 13361 873
rect 10509 755 10763 789
rect 10509 663 10575 755
rect 10609 629 10663 721
rect 10697 663 10763 755
rect 10797 629 10857 789
rect 10415 595 10857 629
rect 10901 561 10955 789
rect 10989 755 11243 789
rect 10989 595 11055 755
rect 11089 561 11143 721
rect 11177 595 11243 755
rect 11277 561 11331 789
rect 11365 595 11431 823
rect 11465 561 11519 789
rect 11553 755 11807 789
rect 11553 595 11619 755
rect 11653 561 11707 721
rect 11741 595 11807 755
rect 11841 561 11895 789
rect 11939 629 11999 789
rect 12033 755 12287 789
rect 12033 663 12099 755
rect 12133 629 12187 721
rect 12221 663 12287 755
rect 12321 629 12381 823
rect 13453 789 13519 907
rect 11939 595 12381 629
rect 12425 561 12479 789
rect 12513 755 13519 789
rect 12513 595 12579 755
rect 12613 561 12667 721
rect 12701 595 12767 755
rect 12801 561 12855 721
rect 12889 595 12955 755
rect 12989 561 13043 721
rect 13077 595 13143 755
rect 13177 561 13231 721
rect 13265 595 13331 755
rect 13365 561 13419 721
rect 13453 595 13519 755
rect 13553 561 13607 789
rect 13725 561 13783 794
rect 13819 629 13879 1003
rect 14013 979 14067 1003
rect 14201 978 14261 1003
rect 14305 978 14359 1071
rect 13913 943 13979 969
rect 14101 943 14167 969
rect 14393 943 14459 1037
rect 14493 979 14547 1071
rect 14581 943 14647 1037
rect 13913 907 14647 943
rect 14681 907 14735 1071
rect 14769 873 14835 1037
rect 14869 907 14923 1071
rect 14957 943 15023 1037
rect 15057 979 15111 1071
rect 15145 943 15211 1037
rect 15245 978 15299 1071
rect 15343 1003 15785 1037
rect 15343 978 15403 1003
rect 15537 979 15591 1003
rect 15437 943 15503 969
rect 15625 943 15691 969
rect 14957 907 15691 943
rect 15725 873 15785 1003
rect 15829 907 15883 1071
rect 15917 943 15983 1037
rect 16017 979 16071 1071
rect 16105 943 16171 1037
rect 16205 979 16259 1071
rect 16293 943 16359 1037
rect 16393 979 16447 1071
rect 16481 943 16547 1037
rect 16581 978 16635 1071
rect 16669 943 16735 1037
rect 16769 979 16823 1071
rect 16857 943 16923 1037
rect 16957 979 17011 1071
rect 17045 943 17111 1037
rect 17145 979 17199 1071
rect 17233 943 17299 1037
rect 15917 907 17299 943
rect 17333 907 17387 1071
rect 17497 926 17555 1071
rect 17590 945 17657 1037
rect 17691 979 17745 1071
rect 17779 945 17845 1037
rect 17879 979 17933 1071
rect 17967 945 18033 1037
rect 18067 979 18121 1071
rect 18155 995 18785 1037
rect 18155 945 18205 995
rect 17590 911 18205 945
rect 18239 911 18691 961
rect 18725 911 18785 995
rect 18877 926 18935 1071
rect 18970 945 19037 1037
rect 19071 979 19125 1071
rect 19159 945 19225 1037
rect 19259 979 19313 1071
rect 19347 945 19413 1037
rect 19447 979 19501 1071
rect 19535 945 19601 1037
rect 19635 979 19689 1071
rect 19723 945 19789 1037
rect 19823 979 19877 1071
rect 19911 945 19977 1037
rect 20011 979 20065 1071
rect 20099 995 21293 1037
rect 20099 945 20149 995
rect 18970 911 20149 945
rect 20183 911 21199 961
rect 21243 911 21293 995
rect 21361 926 21419 1071
rect 21455 945 21521 1037
rect 21555 979 21609 1071
rect 21643 945 21709 1037
rect 21743 979 21797 1071
rect 21831 945 21897 1037
rect 21931 979 21985 1071
rect 22019 945 22085 1037
rect 22119 979 22173 1071
rect 22207 945 22273 1037
rect 22307 979 22361 1071
rect 22395 945 22461 1037
rect 22495 979 22549 1071
rect 22583 945 22649 1037
rect 22683 979 22737 1071
rect 22771 945 22837 1037
rect 22871 979 22925 1071
rect 22959 995 24529 1037
rect 22959 945 23009 995
rect 21455 911 23009 945
rect 23043 911 24435 961
rect 24479 911 24529 995
rect 24581 926 24639 1071
rect 13913 823 14183 873
rect 14385 823 14655 873
rect 14769 823 15219 873
rect 15421 823 15691 873
rect 15725 823 17173 873
rect 13913 755 14167 789
rect 13913 663 13979 755
rect 14013 629 14067 721
rect 14101 663 14167 755
rect 14201 629 14261 789
rect 13819 595 14261 629
rect 14305 561 14359 789
rect 14393 755 14647 789
rect 14393 595 14459 755
rect 14493 561 14547 721
rect 14581 595 14647 755
rect 14681 561 14735 789
rect 14769 595 14835 823
rect 14869 561 14923 789
rect 14957 755 15211 789
rect 14957 595 15023 755
rect 15057 561 15111 721
rect 15145 595 15211 755
rect 15245 561 15299 789
rect 15343 629 15403 789
rect 15437 755 15691 789
rect 15437 663 15503 755
rect 15537 629 15591 721
rect 15625 663 15691 755
rect 15725 629 15785 823
rect 17217 789 17299 907
rect 17651 823 18125 877
rect 15343 595 15785 629
rect 15829 561 15883 789
rect 15917 755 17299 789
rect 15917 595 15983 755
rect 16017 561 16071 721
rect 16105 595 16171 755
rect 16205 561 16259 721
rect 16293 595 16359 755
rect 16393 561 16447 721
rect 16481 595 16547 755
rect 16581 561 16635 721
rect 16669 595 16735 755
rect 16769 561 16823 721
rect 16857 595 16923 755
rect 16957 561 17011 721
rect 17045 595 17111 755
rect 17145 561 17199 721
rect 17233 595 17299 755
rect 17333 561 17387 789
rect 17497 561 17555 794
rect 18239 789 18299 911
rect 18637 877 18691 911
rect 20183 877 20243 911
rect 21145 877 21199 911
rect 23043 877 23103 911
rect 24381 877 24435 911
rect 24679 907 24739 1071
rect 24773 943 24839 1037
rect 24873 977 24927 1071
rect 24961 943 25027 1037
rect 25061 977 25115 1071
rect 25149 943 25215 1037
rect 25249 977 25303 1071
rect 25337 943 25403 1037
rect 25437 977 25491 1071
rect 25525 943 25591 1037
rect 25625 977 25679 1071
rect 25713 943 25779 1037
rect 25813 977 25971 1071
rect 26005 943 26071 1037
rect 26105 977 26159 1071
rect 26193 943 26259 1037
rect 26293 977 26347 1071
rect 26381 943 26447 1037
rect 26481 977 26535 1071
rect 26569 943 26635 1037
rect 26669 977 26723 1071
rect 26757 943 26823 1037
rect 26857 977 26911 1071
rect 26945 943 27023 1037
rect 24773 907 27023 943
rect 27057 907 27107 1071
rect 27157 926 27215 1071
rect 27259 907 27311 1071
rect 27345 943 27411 1037
rect 27445 977 27499 1071
rect 27533 943 27599 1037
rect 27633 977 27687 1071
rect 27721 943 27787 1037
rect 27821 977 27875 1071
rect 27909 943 27975 1037
rect 28009 977 28063 1071
rect 28097 943 28163 1037
rect 28197 977 28251 1071
rect 28285 943 28351 1037
rect 28385 977 28439 1071
rect 28473 943 28539 1037
rect 28573 977 28627 1071
rect 28661 943 28727 1037
rect 28761 977 28919 1071
rect 28953 943 29019 1037
rect 29053 977 29107 1071
rect 29141 943 29207 1037
rect 29241 977 29295 1071
rect 29329 943 29395 1037
rect 29429 977 29483 1071
rect 29517 943 29583 1037
rect 29617 977 29671 1071
rect 29705 943 29771 1037
rect 29805 977 29859 1071
rect 29893 943 29959 1037
rect 29993 977 30047 1071
rect 30081 943 30147 1037
rect 30181 977 30235 1071
rect 30269 943 30335 1037
rect 27345 907 30335 943
rect 30369 907 30425 1071
rect 30469 926 30527 1071
rect 30573 941 30633 1037
rect 30667 975 30723 1071
rect 30757 941 30811 1037
rect 30845 975 30905 1071
rect 30939 941 31005 1037
rect 31039 975 31093 1071
rect 31127 941 31193 1037
rect 31227 975 31281 1071
rect 31315 941 31381 1037
rect 31415 975 31469 1071
rect 31503 941 31569 1037
rect 30573 907 30863 941
rect 30939 907 31569 941
rect 31603 911 31653 1071
rect 31757 926 31815 1071
rect 31861 907 31915 1071
rect 31949 943 32015 1037
rect 32049 977 32103 1071
rect 32137 943 32203 1037
rect 32237 977 32395 1071
rect 31949 941 32203 943
rect 31949 907 32307 941
rect 32341 907 32395 977
rect 32429 943 32489 1037
rect 32523 977 32589 1071
rect 32623 943 32677 1037
rect 32711 977 32777 1071
rect 32811 943 32865 1037
rect 32899 977 32965 1071
rect 32999 943 33053 1037
rect 33087 977 33153 1071
rect 32429 907 33099 943
rect 33229 926 33287 1071
rect 33321 926 33379 1071
rect 33425 907 33479 1071
rect 33513 943 33579 1037
rect 33613 977 33667 1071
rect 33701 943 33767 1037
rect 33801 977 33959 1071
rect 33513 941 33767 943
rect 33513 907 33871 941
rect 33905 907 33959 977
rect 33993 943 34053 1037
rect 34087 977 34153 1071
rect 34187 943 34241 1037
rect 34275 977 34341 1071
rect 34375 943 34429 1037
rect 34463 977 34529 1071
rect 33993 907 34479 943
rect 34609 926 34667 1071
rect 34713 941 34773 1037
rect 34807 975 34863 1071
rect 34897 941 34951 1037
rect 34985 975 35045 1071
rect 35079 941 35145 1037
rect 35179 975 35233 1071
rect 35267 941 35333 1037
rect 35367 975 35421 1071
rect 35455 941 35521 1037
rect 35555 975 35609 1071
rect 35643 941 35709 1037
rect 34713 907 35003 941
rect 35079 907 35709 941
rect 35743 911 35793 1071
rect 35897 926 35955 1071
rect 36017 961 36051 1032
rect 36085 995 36151 1071
rect 36017 927 36127 961
rect 18333 823 18603 877
rect 18637 823 18755 877
rect 19019 823 20105 877
rect 18637 789 18691 823
rect 17597 561 17651 789
rect 17685 755 18691 789
rect 17685 595 17751 755
rect 17785 561 17839 721
rect 17873 595 17939 755
rect 17973 561 18027 721
rect 18061 595 18127 755
rect 18161 561 18215 721
rect 18249 595 18315 755
rect 18349 561 18403 721
rect 18437 595 18503 755
rect 18537 561 18591 721
rect 18625 595 18691 755
rect 18725 561 18779 789
rect 18877 561 18935 794
rect 20161 789 20243 877
rect 20277 823 21091 877
rect 21145 823 21239 877
rect 21515 823 22941 877
rect 21145 789 21199 823
rect 18977 561 19031 789
rect 19065 755 21199 789
rect 19065 595 19131 755
rect 19165 561 19219 721
rect 19253 595 19319 755
rect 19353 561 19407 721
rect 19441 595 19507 755
rect 19541 561 19595 721
rect 19629 595 19695 755
rect 19729 561 19783 721
rect 19817 595 19883 755
rect 19917 561 19971 721
rect 20005 595 20071 755
rect 20105 561 20159 721
rect 20193 595 20259 755
rect 20293 561 20347 721
rect 20381 595 20447 755
rect 20481 561 20535 721
rect 20569 595 20635 755
rect 20669 561 20723 721
rect 20757 595 20823 755
rect 20857 561 20911 721
rect 20945 595 21011 755
rect 21045 561 21099 721
rect 21133 595 21199 755
rect 21233 561 21287 789
rect 21361 561 21419 794
rect 23021 789 23103 877
rect 23137 823 24291 877
rect 24381 823 24459 877
rect 24757 831 25231 873
rect 25321 831 25795 873
rect 25989 831 26463 873
rect 26535 831 26873 873
rect 24381 789 24435 823
rect 26945 797 27023 907
rect 27313 831 27991 873
rect 28081 831 28759 873
rect 28921 831 29599 873
rect 29713 797 29795 907
rect 30828 873 30863 907
rect 29829 831 30303 873
rect 30572 833 30792 873
rect 30828 839 31353 873
rect 30828 799 30863 839
rect 31402 799 31569 907
rect 32271 873 32307 907
rect 31915 833 32049 873
rect 32103 833 32237 873
rect 32271 833 32937 873
rect 32271 799 32307 833
rect 21461 561 21515 789
rect 21549 755 24435 789
rect 21549 595 21615 755
rect 21649 561 21703 721
rect 21737 595 21803 755
rect 21837 561 21891 721
rect 21925 595 21991 755
rect 22025 561 22079 721
rect 22113 595 22179 755
rect 22213 561 22267 721
rect 22301 595 22367 755
rect 22401 561 22455 721
rect 22489 595 22555 755
rect 22589 561 22643 721
rect 22677 595 22743 755
rect 22777 561 22831 721
rect 22865 595 22931 755
rect 22965 561 23019 721
rect 23053 595 23119 755
rect 23153 561 23207 721
rect 23241 595 23307 755
rect 23341 561 23395 721
rect 23429 595 23495 755
rect 23529 561 23583 721
rect 23617 595 23683 755
rect 23717 561 23771 721
rect 23805 595 23871 755
rect 23905 561 23959 721
rect 23993 595 24059 755
rect 24093 561 24147 721
rect 24181 595 24247 755
rect 24281 561 24335 721
rect 24369 595 24435 755
rect 24469 561 24523 789
rect 24581 561 24639 794
rect 24679 763 25301 797
rect 24679 595 24737 763
rect 24781 561 24831 729
rect 24875 595 24925 763
rect 24969 561 25019 729
rect 25063 595 25113 763
rect 25157 561 25207 729
rect 25251 629 25301 763
rect 25345 763 26439 797
rect 25345 663 25395 763
rect 25439 629 25489 729
rect 25533 663 25583 763
rect 25627 629 25677 729
rect 25721 663 25771 763
rect 25815 629 25873 729
rect 25251 595 25873 629
rect 25911 629 25969 729
rect 26013 663 26063 763
rect 26107 629 26157 729
rect 26201 663 26251 763
rect 26295 629 26345 729
rect 26389 663 26439 763
rect 26483 629 26533 797
rect 26577 763 27023 797
rect 26577 663 26627 763
rect 26671 629 26721 729
rect 26765 663 26815 763
rect 26859 629 26909 729
rect 26945 663 27023 763
rect 27057 629 27107 797
rect 25911 595 27107 629
rect 27157 561 27215 794
rect 27251 763 28061 797
rect 27251 595 27317 763
rect 27353 561 27403 729
rect 27447 595 27497 763
rect 27541 561 27591 729
rect 27635 595 27685 763
rect 27729 561 27779 729
rect 27823 595 27873 763
rect 27917 561 27967 729
rect 28011 629 28061 763
rect 28105 763 29575 797
rect 28105 663 28155 763
rect 28199 629 28249 729
rect 28293 663 28343 763
rect 28387 629 28437 729
rect 28481 663 28531 763
rect 28575 629 28625 729
rect 28669 663 28719 763
rect 28763 629 28821 729
rect 28011 595 28821 629
rect 28859 629 28917 729
rect 28961 663 29011 763
rect 29047 629 29105 729
rect 29149 663 29199 763
rect 29243 629 29293 729
rect 29337 663 29387 763
rect 29431 629 29481 729
rect 29525 663 29575 763
rect 29619 629 29669 797
rect 29713 763 30327 797
rect 29713 663 29763 763
rect 29807 629 29857 729
rect 29901 663 29951 763
rect 29995 629 30045 729
rect 30089 663 30139 763
rect 30183 629 30233 729
rect 30277 663 30327 763
rect 30371 629 30431 795
rect 28859 595 30431 629
rect 30469 561 30527 794
rect 30563 765 30863 799
rect 30939 765 31569 799
rect 30563 595 30629 765
rect 30663 561 30717 721
rect 30751 595 30817 765
rect 30851 561 30905 721
rect 30939 595 31005 765
rect 31039 561 31093 721
rect 31127 595 31193 765
rect 31227 561 31281 721
rect 31315 595 31381 765
rect 31415 561 31469 721
rect 31503 595 31569 765
rect 31603 561 31663 791
rect 31757 561 31815 794
rect 31850 755 32103 797
rect 31850 595 31915 755
rect 31949 561 32015 721
rect 32049 629 32103 755
rect 32137 755 32307 799
rect 33019 789 33099 907
rect 33835 873 33871 907
rect 33479 833 33613 873
rect 33667 833 33801 873
rect 33835 833 34365 873
rect 33835 799 33871 833
rect 32137 663 32203 755
rect 32237 629 32297 721
rect 32049 595 32297 629
rect 32341 561 32395 789
rect 32429 755 33099 789
rect 32429 595 32495 755
rect 32529 561 32583 721
rect 32617 595 32683 755
rect 32717 561 32771 721
rect 32805 595 32871 755
rect 32905 561 32959 721
rect 32993 595 33059 755
rect 33093 561 33147 721
rect 33229 597 33287 794
rect 33321 597 33379 794
rect 33414 755 33667 797
rect 33414 595 33479 755
rect 33513 561 33579 721
rect 33613 629 33667 755
rect 33701 755 33871 799
rect 34399 789 34479 907
rect 34968 873 35003 907
rect 34712 833 34932 873
rect 34968 839 35493 873
rect 34968 799 35003 839
rect 35542 799 35709 907
rect 33701 663 33767 755
rect 33801 629 33861 721
rect 33613 595 33861 629
rect 33905 561 33959 789
rect 33993 755 34479 789
rect 33993 595 34059 755
rect 34093 561 34147 721
rect 34181 595 34247 755
rect 34281 561 34335 721
rect 34369 595 34435 755
rect 34469 561 34523 721
rect 34609 561 34667 794
rect 34703 765 35003 799
rect 35079 765 35709 799
rect 34703 595 34769 765
rect 34803 561 34857 721
rect 34891 595 34957 765
rect 34991 561 35045 721
rect 35079 595 35145 765
rect 35179 561 35233 721
rect 35267 595 35333 765
rect 35367 561 35421 721
rect 35455 595 35521 765
rect 35555 561 35609 721
rect 35643 595 35709 765
rect 35743 561 35803 791
rect 35897 561 35955 794
rect 35989 763 36059 891
rect 36093 874 36127 927
rect 36093 729 36151 874
rect 35989 695 36151 729
rect 36185 799 36219 1032
rect 36304 965 36343 1019
rect 36377 999 36443 1071
rect 36580 975 36704 1032
rect 36304 935 36395 965
rect 36304 931 36479 935
rect 36259 828 36325 897
rect 36361 869 36479 931
rect 36528 869 36631 941
rect 35989 595 36051 695
rect 36085 561 36151 661
rect 36185 595 36239 799
rect 36361 789 36395 869
rect 36283 755 36395 789
rect 36283 595 36349 755
rect 36461 751 36563 835
rect 36597 773 36631 869
rect 36670 889 36704 975
rect 36746 966 36812 1071
rect 36863 923 36929 1037
rect 37036 963 37091 1071
rect 37125 989 37231 1037
rect 37036 923 37102 963
rect 36670 855 36848 889
rect 36708 823 36848 855
rect 36383 561 36437 721
rect 36597 689 36674 773
rect 36708 655 36742 823
rect 36882 781 36916 923
rect 37136 911 37231 989
rect 37277 926 37335 1071
rect 37397 961 37431 1032
rect 37465 995 37531 1071
rect 37397 927 37507 961
rect 36950 823 37049 889
rect 37083 823 37151 877
rect 37083 781 37117 823
rect 37185 789 37231 911
rect 36776 747 37117 781
rect 36776 715 37006 747
rect 36576 611 36742 655
rect 36782 561 36899 661
rect 36949 595 37006 715
rect 37041 658 37107 711
rect 37041 561 37101 658
rect 37151 637 37231 789
rect 37135 595 37231 637
rect 37277 561 37335 794
rect 37369 763 37439 891
rect 37473 874 37507 927
rect 37473 808 37531 874
rect 37473 729 37507 808
rect 37369 695 37507 729
rect 37565 751 37599 1032
rect 37684 965 37723 1019
rect 37757 999 37823 1071
rect 37960 975 38084 1032
rect 37684 935 37775 965
rect 37684 931 37859 935
rect 37639 823 37705 897
rect 37741 869 37859 931
rect 37908 869 38011 941
rect 37741 789 37775 869
rect 37663 755 37775 789
rect 37369 595 37431 695
rect 37465 561 37531 661
rect 37565 595 37619 751
rect 37663 595 37729 755
rect 37841 751 37943 835
rect 37977 773 38011 869
rect 38050 889 38084 975
rect 38126 966 38192 1071
rect 38243 923 38309 1037
rect 38416 963 38471 1071
rect 38505 989 38611 1037
rect 38416 923 38482 963
rect 38050 855 38228 889
rect 38088 823 38228 855
rect 37763 561 37817 721
rect 37977 689 38054 773
rect 38088 655 38122 823
rect 38262 781 38296 923
rect 38516 911 38611 989
rect 38657 926 38715 1071
rect 38777 961 38811 1032
rect 38845 995 38911 1071
rect 38777 927 38887 961
rect 38330 823 38429 889
rect 38463 823 38531 877
rect 38463 781 38497 823
rect 38565 789 38611 911
rect 38156 747 38497 781
rect 38156 715 38386 747
rect 37956 611 38122 655
rect 38162 561 38279 661
rect 38329 595 38386 715
rect 38421 658 38487 711
rect 38421 561 38481 658
rect 38531 637 38611 789
rect 38515 595 38611 637
rect 38657 561 38715 794
rect 38749 763 38819 891
rect 38853 874 38887 927
rect 38853 729 38911 874
rect 38749 695 38911 729
rect 38945 799 38979 1032
rect 39064 965 39103 1019
rect 39137 999 39203 1071
rect 39340 975 39464 1032
rect 39064 935 39155 965
rect 39064 931 39239 935
rect 39019 828 39085 897
rect 39121 869 39239 931
rect 39288 869 39391 941
rect 38749 595 38811 695
rect 38845 561 38911 661
rect 38945 595 38999 799
rect 39121 789 39155 869
rect 39043 755 39155 789
rect 39043 595 39109 755
rect 39221 751 39323 835
rect 39357 773 39391 869
rect 39430 889 39464 975
rect 39506 966 39572 1071
rect 39623 923 39689 1037
rect 39795 923 39861 1071
rect 39895 923 39973 1037
rect 39430 855 39608 889
rect 39468 823 39608 855
rect 39143 561 39197 721
rect 39357 689 39434 773
rect 39468 655 39502 823
rect 39642 781 39676 923
rect 39710 823 39809 889
rect 39843 823 39905 889
rect 39939 877 39973 923
rect 40007 911 40049 1071
rect 40129 926 40187 1071
rect 40249 961 40283 1032
rect 40317 995 40383 1071
rect 40249 927 40359 961
rect 39939 823 40019 877
rect 39843 781 39877 823
rect 39939 789 39973 823
rect 39536 747 39877 781
rect 39536 715 39766 747
rect 39336 611 39502 655
rect 39542 561 39659 661
rect 39709 595 39766 715
rect 39801 658 39867 711
rect 39801 561 39861 658
rect 39911 637 39973 789
rect 39895 597 39973 637
rect 40007 561 40048 789
rect 40129 561 40187 794
rect 40221 763 40291 891
rect 40325 874 40359 927
rect 40325 808 40383 874
rect 40325 729 40359 808
rect 40221 695 40359 729
rect 40417 751 40451 1032
rect 40536 965 40575 1019
rect 40609 999 40675 1071
rect 40812 975 40936 1032
rect 40536 935 40627 965
rect 40536 931 40711 935
rect 40491 823 40557 897
rect 40593 869 40711 931
rect 40760 869 40863 941
rect 40593 789 40627 869
rect 40515 755 40627 789
rect 40221 595 40283 695
rect 40317 561 40383 661
rect 40417 595 40471 751
rect 40515 595 40581 755
rect 40693 751 40795 835
rect 40829 773 40863 869
rect 40902 889 40936 975
rect 40978 966 41044 1071
rect 41095 923 41161 1037
rect 41267 923 41333 1071
rect 41367 923 41445 1037
rect 40902 855 41080 889
rect 40940 823 41080 855
rect 40615 561 40669 721
rect 40829 689 40906 773
rect 40940 655 40974 823
rect 41114 781 41148 923
rect 41182 823 41281 889
rect 41315 823 41377 889
rect 41411 877 41445 923
rect 41479 911 41521 1071
rect 41601 926 41659 1071
rect 41721 961 41755 1032
rect 41789 995 41855 1071
rect 41721 927 41831 961
rect 41411 823 41491 877
rect 41315 781 41349 823
rect 41411 789 41445 823
rect 41008 747 41349 781
rect 41008 715 41238 747
rect 40808 611 40974 655
rect 41014 561 41131 661
rect 41181 595 41238 715
rect 41273 658 41339 711
rect 41273 561 41333 658
rect 41383 637 41445 789
rect 41367 597 41445 637
rect 41479 561 41520 789
rect 41601 561 41659 794
rect 41693 763 41763 891
rect 41797 874 41831 927
rect 41797 729 41855 874
rect 41693 695 41855 729
rect 41889 799 41923 1032
rect 42008 965 42047 1019
rect 42081 999 42147 1071
rect 42284 975 42408 1032
rect 42008 935 42099 965
rect 42008 931 42183 935
rect 41963 828 42029 897
rect 42065 869 42183 931
rect 42232 869 42335 941
rect 41693 595 41755 695
rect 41789 561 41855 661
rect 41889 595 41943 799
rect 42065 789 42099 869
rect 41987 755 42099 789
rect 41987 595 42053 755
rect 42165 751 42267 835
rect 42301 773 42335 869
rect 42374 889 42408 975
rect 42450 966 42516 1071
rect 42567 923 42633 1037
rect 42739 923 42805 1071
rect 42839 941 42915 1037
rect 42951 975 42993 1071
rect 43027 941 43093 1037
rect 42374 855 42552 889
rect 42412 823 42552 855
rect 42087 561 42141 721
rect 42301 689 42378 773
rect 42412 655 42446 823
rect 42586 781 42620 923
rect 42839 907 43093 941
rect 43127 911 43169 1071
rect 43257 926 43315 1071
rect 43377 961 43411 1032
rect 43445 995 43511 1071
rect 43377 927 43487 961
rect 42654 823 42753 889
rect 42957 877 43093 907
rect 42787 823 42923 873
rect 42957 823 43129 877
rect 42787 781 42821 823
rect 42957 789 43093 823
rect 42480 747 42821 781
rect 42855 755 43093 789
rect 42480 715 42711 747
rect 42280 611 42446 655
rect 42480 561 42617 661
rect 42651 601 42711 715
rect 42855 713 42905 755
rect 42745 658 42811 713
rect 42745 561 42805 658
rect 42845 637 42905 713
rect 42839 595 42905 637
rect 42939 561 42993 721
rect 43027 595 43093 755
rect 43127 561 43178 789
rect 43257 561 43315 794
rect 43349 763 43419 891
rect 43453 874 43487 927
rect 43453 808 43511 874
rect 43453 729 43487 808
rect 43349 695 43487 729
rect 43545 751 43579 1032
rect 43664 965 43703 1019
rect 43737 999 43803 1071
rect 43940 975 44064 1032
rect 43664 935 43755 965
rect 43664 931 43839 935
rect 43619 823 43685 897
rect 43721 869 43839 931
rect 43888 869 43991 941
rect 43721 789 43755 869
rect 43643 755 43755 789
rect 43349 595 43411 695
rect 43445 561 43511 661
rect 43545 595 43599 751
rect 43643 595 43709 755
rect 43821 751 43923 835
rect 43957 773 43991 869
rect 44030 889 44064 975
rect 44106 966 44172 1071
rect 44223 923 44289 1037
rect 44395 923 44461 1071
rect 44495 941 44571 1037
rect 44607 975 44649 1071
rect 44683 941 44749 1037
rect 44030 855 44208 889
rect 44068 823 44208 855
rect 43743 561 43797 721
rect 43957 689 44034 773
rect 44068 655 44102 823
rect 44242 781 44276 923
rect 44495 907 44749 941
rect 44783 911 44825 1071
rect 44913 926 44971 1071
rect 44310 823 44409 889
rect 44613 877 44749 907
rect 44443 823 44579 873
rect 44613 823 44785 877
rect 44443 781 44477 823
rect 44613 789 44749 823
rect 44136 747 44477 781
rect 44511 755 44749 789
rect 44136 715 44367 747
rect 43936 611 44102 655
rect 44136 561 44273 661
rect 44307 601 44367 715
rect 44511 713 44561 755
rect 44401 658 44467 713
rect 44401 561 44461 658
rect 44501 637 44561 713
rect 44495 595 44561 637
rect 44595 561 44649 721
rect 44683 595 44749 755
rect 44783 561 44834 789
rect 44913 561 44971 794
rect 45005 595 45155 1037
rect 45189 595 45523 1037
rect 45557 595 46075 1037
rect 46109 595 46811 1037
rect 46845 926 46903 1071
rect 388441 926 388499 1071
rect 388570 966 388628 1071
rect 388670 923 388720 1032
rect 388754 966 388812 1071
rect 388913 1003 389319 1037
rect 388913 934 388963 1003
rect 388533 823 388652 889
rect 388686 875 388720 923
rect 388997 875 389063 969
rect 389097 934 389131 1003
rect 389165 911 389231 969
rect 389265 945 389319 1003
rect 389353 979 389403 1071
rect 389437 945 389503 1037
rect 389537 979 389591 1071
rect 389625 945 389691 1037
rect 389265 911 389691 945
rect 389725 911 389791 1071
rect 389825 945 389891 1037
rect 389925 979 389979 1071
rect 390013 945 390079 1037
rect 390113 979 390163 1071
rect 390197 1003 390603 1037
rect 390197 945 390251 1003
rect 389825 911 390251 945
rect 390285 911 390351 969
rect 390385 934 390419 1003
rect 389165 875 389211 911
rect 388686 809 388923 875
rect 388957 815 389211 875
rect 389447 823 389725 877
rect 389791 823 390069 877
rect 390305 875 390351 911
rect 390453 875 390519 969
rect 390553 934 390603 1003
rect 390704 966 390762 1071
rect 390796 923 390846 1032
rect 390888 966 390946 1071
rect 391054 966 391112 1071
rect 391154 923 391204 1032
rect 391238 966 391296 1071
rect 391397 1003 391803 1037
rect 391397 934 391447 1003
rect 390796 875 390830 923
rect 46845 561 46903 794
rect 388441 561 388499 794
rect 388686 767 388720 809
rect 388560 561 388620 767
rect 388654 595 388720 767
rect 388759 561 388814 767
rect 388863 595 388923 775
rect 0 527 388923 561
rect 18 337 71 491
rect 105 383 181 527
rect 219 419 271 491
rect 305 453 417 527
rect 461 419 513 491
rect 219 373 513 419
rect 641 337 709 491
rect 18 53 85 337
rect 121 301 709 337
rect 121 163 169 301
rect 753 294 811 527
rect 846 298 905 527
rect 203 199 339 265
rect 373 199 478 265
rect 518 199 615 265
rect 661 199 717 265
rect 121 125 707 163
rect 131 17 280 91
rect 439 53 504 125
rect 540 17 616 91
rect 662 53 707 125
rect 753 17 811 162
rect 846 17 905 181
rect 949 51 995 467
rect 1048 366 1099 527
rect 1139 404 1215 493
rect 1259 438 1314 527
rect 1371 404 1437 493
rect 1139 368 1437 404
rect 1539 332 1615 465
rect 1048 298 1615 332
rect 1048 175 1099 298
rect 1673 294 1731 527
rect 1766 375 1833 527
rect 1877 341 1914 493
rect 1958 375 2024 527
rect 2068 341 2106 493
rect 2150 367 2200 527
rect 2262 442 2728 493
rect 2762 455 2838 527
rect 2662 421 2728 442
rect 2880 421 2942 493
rect 2976 455 3052 527
rect 3096 421 3147 493
rect 2254 374 2520 408
rect 2662 376 3147 421
rect 1765 299 2106 341
rect 2254 335 2289 374
rect 2225 301 2289 335
rect 1133 209 1220 255
rect 1286 209 1367 255
rect 1401 209 1467 255
rect 1501 209 1575 255
rect 1765 175 1816 299
rect 2225 265 2272 301
rect 2323 289 2673 340
rect 2323 265 2369 289
rect 1853 209 2272 265
rect 1048 139 1615 175
rect 1029 17 1182 89
rect 1323 55 1399 139
rect 1450 17 1505 105
rect 1539 55 1615 139
rect 1673 17 1731 162
rect 1765 127 2193 175
rect 1965 123 2193 127
rect 2227 161 2272 209
rect 2306 197 2369 265
rect 2403 197 2557 255
rect 2597 197 2673 289
rect 2737 302 3037 340
rect 3071 307 3147 376
rect 2737 204 2813 302
rect 2855 204 2934 266
rect 2973 264 3037 302
rect 3237 294 3295 527
rect 3337 345 3387 491
rect 3421 381 3497 527
rect 3541 345 3578 491
rect 3337 305 3578 345
rect 2973 204 3123 264
rect 2227 123 2956 161
rect 1845 17 1921 93
rect 1965 51 2003 123
rect 2037 17 2113 89
rect 2157 51 2193 123
rect 2232 17 2309 89
rect 2353 51 2402 123
rect 2436 17 2512 89
rect 2556 51 2632 123
rect 2676 17 2750 89
rect 2880 55 2956 123
rect 3071 17 3147 161
rect 3237 17 3295 162
rect 3331 153 3399 265
rect 3433 199 3568 265
rect 3612 199 3671 491
rect 3705 357 3842 491
rect 3708 199 3765 323
rect 3329 17 3397 119
rect 3433 53 3493 199
rect 3799 163 3842 357
rect 3881 294 3939 527
rect 3985 457 4439 491
rect 3985 357 4037 457
rect 4191 451 4439 457
rect 3976 199 4037 323
rect 4071 171 4135 423
rect 4191 357 4229 451
rect 4263 331 4339 415
rect 4383 367 4439 451
rect 4483 367 4529 527
rect 4575 331 4629 493
rect 4675 367 4721 527
rect 4767 331 4821 493
rect 4867 367 4913 527
rect 4169 257 4213 323
rect 4263 291 4821 331
rect 4893 257 4939 331
rect 4985 294 5043 527
rect 5079 417 5129 493
rect 5163 451 5239 527
rect 5283 421 5317 493
rect 5351 455 5427 527
rect 5471 421 5505 493
rect 5539 455 5615 527
rect 5659 421 5693 493
rect 5727 455 5803 527
rect 5847 451 6674 493
rect 5847 421 5881 451
rect 5283 417 5881 421
rect 5079 359 5881 417
rect 5915 357 6152 417
rect 6204 373 6692 417
rect 6086 339 6152 357
rect 4169 207 4343 257
rect 4518 207 4670 257
rect 4734 207 4939 257
rect 5080 289 5855 325
rect 5080 207 5367 289
rect 5421 207 5721 255
rect 5779 207 5855 289
rect 5889 255 6052 323
rect 6086 289 6382 339
rect 6426 255 6470 339
rect 5889 207 6121 255
rect 6170 207 6470 255
rect 6520 265 6562 331
rect 6596 299 6692 373
rect 6520 199 6607 265
rect 3543 125 3842 163
rect 3543 53 3580 125
rect 3622 17 3698 91
rect 3763 53 3808 125
rect 3881 17 3939 162
rect 3985 17 4035 163
rect 4071 131 4635 171
rect 4071 51 4133 131
rect 4681 127 4923 171
rect 4681 95 4715 127
rect 4167 17 4243 95
rect 4359 17 4435 95
rect 4473 53 4715 95
rect 4751 17 4827 91
rect 4873 53 4923 127
rect 4985 17 5043 162
rect 5183 139 5411 173
rect 5079 17 5139 117
rect 5183 106 5225 139
rect 5260 17 5317 105
rect 5351 101 5411 139
rect 5445 165 6471 173
rect 6641 165 6692 299
rect 6733 294 6791 527
rect 6829 409 6877 487
rect 6911 445 6991 527
rect 6829 369 7001 409
rect 5445 139 6692 165
rect 5445 135 5796 139
rect 5915 125 6692 139
rect 5915 123 6179 125
rect 5351 51 5803 101
rect 5847 17 5881 105
rect 5915 51 5989 123
rect 6033 17 6099 89
rect 6145 51 6179 123
rect 6333 123 6692 125
rect 6223 17 6289 89
rect 6333 51 6367 123
rect 6411 17 6477 89
rect 6593 17 6674 89
rect 6733 17 6791 162
rect 6829 65 6875 333
rect 6911 233 7001 369
rect 7035 269 7101 491
rect 7145 397 7181 491
rect 7215 431 7291 527
rect 7336 397 7370 491
rect 7145 357 7370 397
rect 6911 53 6967 233
rect 7035 209 7154 269
rect 7017 17 7066 173
rect 7100 163 7154 209
rect 7188 199 7263 323
rect 7297 199 7349 323
rect 7423 299 7480 527
rect 7465 163 7517 265
rect 7100 125 7517 163
rect 7100 53 7196 125
rect 7332 17 7478 91
rect 7551 53 7607 491
rect 7653 294 7711 527
rect 7746 451 7813 527
rect 7857 401 7908 485
rect 7956 455 8022 527
rect 8153 421 8203 493
rect 7750 367 7908 401
rect 7971 379 8203 421
rect 7750 177 7804 367
rect 7971 333 8005 379
rect 7852 299 8005 333
rect 8039 311 8135 345
rect 7852 215 7918 299
rect 8101 265 8135 311
rect 8169 335 8203 379
rect 8237 403 8313 493
rect 8359 437 8393 527
rect 8427 403 8503 493
rect 8237 369 8503 403
rect 8169 301 8271 335
rect 7973 199 8067 265
rect 8101 199 8193 265
rect 7653 17 7711 162
rect 7750 143 7908 177
rect 8101 165 8135 199
rect 7746 17 7797 109
rect 7832 63 7908 143
rect 7942 17 8008 157
rect 8049 131 8135 165
rect 8227 165 8271 301
rect 8305 199 8345 323
rect 8403 199 8461 323
rect 8573 294 8631 527
rect 8669 421 8752 493
rect 8786 455 8862 527
rect 8978 455 9054 527
rect 9169 455 9246 527
rect 9303 442 9525 476
rect 9559 455 9635 527
rect 9747 455 9823 527
rect 8669 387 9266 421
rect 8669 359 8755 387
rect 8669 168 8708 359
rect 8742 202 8818 325
rect 8858 319 9164 353
rect 8227 127 8316 165
rect 8153 17 8219 93
rect 8427 17 8503 165
rect 8573 17 8631 162
rect 8669 51 8750 168
rect 8858 157 8956 319
rect 9232 305 9266 387
rect 9303 339 9337 442
rect 9489 421 9525 442
rect 9489 387 9917 421
rect 9232 271 9353 305
rect 8990 237 9198 265
rect 8990 199 9254 237
rect 9291 199 9353 271
rect 9220 157 9254 199
rect 9397 168 9431 361
rect 9489 289 9525 387
rect 9561 319 9820 353
rect 9561 255 9606 319
rect 9517 202 9606 255
rect 9640 202 9723 272
rect 9774 258 9820 319
rect 9866 292 9917 387
rect 9953 294 10011 527
rect 10047 401 10099 487
rect 10133 435 10207 527
rect 10047 367 10199 401
rect 9774 211 9892 258
rect 10049 195 10095 333
rect 9397 157 9725 168
rect 8858 123 9150 157
rect 9220 134 9725 157
rect 9220 123 9431 134
rect 8784 17 8862 89
rect 8978 17 9054 89
rect 9195 17 9349 89
rect 9397 51 9431 123
rect 9483 17 9549 89
rect 9669 81 9725 134
rect 9861 17 9917 177
rect 9953 17 10011 162
rect 10131 143 10199 367
rect 10241 269 10333 491
rect 10377 345 10415 491
rect 10449 381 10525 527
rect 10595 345 10629 491
rect 10377 305 10629 345
rect 10689 294 10747 527
rect 10783 416 10849 527
rect 10984 457 11247 493
rect 10241 209 10384 269
rect 10101 53 10199 143
rect 10233 17 10279 173
rect 10316 53 10384 209
rect 10425 75 10476 269
rect 10558 199 10653 269
rect 10571 17 10643 163
rect 10689 17 10747 162
rect 10788 153 10849 361
rect 10893 257 10929 453
rect 10984 359 11034 457
rect 10893 214 11035 257
rect 10893 106 10929 214
rect 10817 72 10929 106
rect 10981 17 11029 177
rect 11069 157 11137 423
rect 11171 405 11247 457
rect 11291 439 11325 527
rect 11386 421 11420 493
rect 11456 455 11532 527
rect 11576 421 11628 493
rect 11386 405 11628 421
rect 11171 371 11628 405
rect 11224 299 11581 335
rect 11224 249 11299 299
rect 11223 215 11299 249
rect 11335 199 11477 265
rect 11511 199 11581 299
rect 11701 294 11759 527
rect 11795 401 11861 493
rect 11905 435 11957 527
rect 12012 443 12449 493
rect 12483 455 12559 527
rect 12675 455 12751 527
rect 11795 357 11978 401
rect 12012 359 12061 443
rect 12187 441 12449 443
rect 12409 421 12449 441
rect 12795 421 12833 493
rect 12867 455 12943 527
rect 12986 421 13023 493
rect 13059 455 13135 527
rect 13174 421 13224 493
rect 11799 215 11910 323
rect 11866 199 11910 215
rect 11944 269 11978 357
rect 12112 341 12365 407
rect 12409 375 13224 421
rect 12112 317 12402 341
rect 11944 207 12300 269
rect 11069 123 11436 157
rect 11069 51 11138 123
rect 11192 17 11258 89
rect 11360 51 11436 123
rect 11562 17 11630 157
rect 11701 17 11759 162
rect 11944 159 12007 207
rect 12340 179 12402 317
rect 12436 296 13200 341
rect 12436 213 12515 296
rect 12549 213 12864 262
rect 12921 215 13200 296
rect 13265 294 13323 527
rect 12340 173 12853 179
rect 11794 123 12007 159
rect 12051 139 12853 173
rect 12051 123 12281 139
rect 12487 135 12853 139
rect 12897 147 13141 181
rect 11794 51 11865 123
rect 11930 17 12007 89
rect 12051 74 12089 123
rect 12133 17 12209 89
rect 12243 51 12281 123
rect 12325 17 12453 105
rect 12897 101 12949 147
rect 12489 51 12949 101
rect 12993 17 13031 113
rect 13065 51 13141 147
rect 13176 17 13224 177
rect 13265 17 13323 162
rect 13359 53 13411 491
rect 13445 381 13523 527
rect 13559 345 13613 491
rect 13449 301 13613 345
rect 13659 349 13705 491
rect 13741 385 13817 527
rect 13861 349 13913 491
rect 13659 301 13913 349
rect 13449 167 13517 301
rect 14001 294 14059 527
rect 14095 333 14151 527
rect 13553 203 13662 265
rect 13696 203 13783 265
rect 13449 127 13703 167
rect 13473 17 13607 91
rect 13643 53 13703 127
rect 13737 75 13783 203
rect 13822 199 13872 265
rect 13855 17 13913 163
rect 14001 17 14059 162
rect 14111 17 14145 111
rect 14185 51 14241 493
rect 14287 444 14373 527
rect 14411 384 14484 493
rect 14275 338 14484 384
rect 14528 387 14573 493
rect 14617 425 14683 527
rect 14727 387 14771 493
rect 14275 165 14362 338
rect 14528 334 14771 387
rect 14829 294 14887 527
rect 14927 387 14993 527
rect 15039 351 15073 437
rect 15109 387 15185 527
rect 15231 351 15281 437
rect 14933 317 15281 351
rect 14449 199 14524 282
rect 14275 131 14524 165
rect 14331 17 14407 89
rect 14486 51 14524 131
rect 14558 73 14622 265
rect 14708 150 14783 265
rect 14707 17 14783 113
rect 14829 17 14887 162
rect 14933 157 15040 317
rect 15317 303 15367 527
rect 15435 459 15657 493
rect 15435 339 15469 459
rect 15074 199 15364 265
rect 15404 199 15485 305
rect 15330 157 15364 199
rect 15529 168 15563 425
rect 15621 404 15657 459
rect 15691 455 15767 527
rect 15811 404 15845 493
rect 15879 455 15955 527
rect 16010 404 16076 479
rect 15621 370 16076 404
rect 15621 289 15657 370
rect 15693 302 15991 336
rect 15693 255 15738 302
rect 15931 258 15991 302
rect 16025 292 16076 370
rect 16117 294 16175 527
rect 16211 337 16266 491
rect 16300 405 16376 491
rect 16420 439 16459 527
rect 16495 405 16571 491
rect 16300 371 16571 405
rect 16211 299 16338 337
rect 16372 305 16571 371
rect 15649 202 15738 255
rect 15772 202 15897 255
rect 15931 211 16024 258
rect 15529 157 15857 168
rect 14933 123 15281 157
rect 15330 134 15857 157
rect 15330 123 15563 134
rect 14925 17 14993 89
rect 15109 17 15185 89
rect 15326 17 15481 89
rect 15529 51 15563 123
rect 15615 17 15681 89
rect 15801 81 15857 134
rect 15993 17 16049 177
rect 16117 17 16175 162
rect 16211 135 16259 265
rect 16293 165 16338 299
rect 16669 294 16727 527
rect 16766 421 16818 493
rect 16852 455 16928 527
rect 16974 421 17008 493
rect 17069 439 17103 527
rect 17147 457 17422 493
rect 16766 405 17008 421
rect 17147 405 17213 457
rect 16766 371 17213 405
rect 16773 299 17170 335
rect 16372 199 16451 265
rect 16497 199 16556 265
rect 16773 207 16883 299
rect 16923 199 17059 265
rect 17095 215 17170 299
rect 17247 266 17317 423
rect 17361 359 17422 457
rect 16293 129 16369 165
rect 16214 17 16280 95
rect 16324 53 16369 129
rect 16405 75 16451 199
rect 16511 17 16571 163
rect 16669 17 16727 162
rect 16764 17 16823 173
rect 17226 157 17317 266
rect 17351 199 17451 325
rect 17497 294 17555 527
rect 17608 443 18035 493
rect 18069 455 18145 527
rect 17608 359 17647 443
rect 17773 441 18035 443
rect 17995 421 18035 441
rect 18189 421 18227 493
rect 18261 455 18337 527
rect 18381 421 18419 493
rect 18453 455 18529 527
rect 18573 421 18609 493
rect 18645 455 18721 527
rect 18765 421 18817 493
rect 17698 341 17951 407
rect 17995 375 18817 421
rect 17698 317 17988 341
rect 17590 207 17888 283
rect 17590 199 17652 207
rect 17922 179 17988 317
rect 18022 296 18786 341
rect 18022 213 18101 296
rect 18135 213 18452 262
rect 18507 215 18786 296
rect 18877 294 18935 527
rect 18987 325 19021 493
rect 19055 459 19319 493
rect 19055 359 19115 459
rect 19243 451 19319 459
rect 19357 443 19423 527
rect 19175 409 19220 425
rect 19467 409 19517 493
rect 19175 367 19517 409
rect 19561 375 19627 527
rect 19175 359 19387 367
rect 19412 325 19659 333
rect 18987 299 19659 325
rect 18987 291 19442 299
rect 18969 215 19039 257
rect 19073 215 19183 257
rect 19217 215 19315 257
rect 17922 173 18433 179
rect 16945 123 17317 157
rect 16945 51 17024 123
rect 17126 17 17202 89
rect 17253 51 17317 123
rect 17363 17 17429 165
rect 17497 17 17555 162
rect 17590 17 17657 161
rect 17701 139 18433 173
rect 17701 123 17931 139
rect 18067 135 18433 139
rect 18477 147 18721 181
rect 17701 74 17739 123
rect 17773 17 17849 89
rect 17893 51 17931 123
rect 17969 17 18035 105
rect 18477 101 18529 147
rect 18069 51 18529 101
rect 18573 17 18611 113
rect 18645 51 18721 147
rect 18765 17 18817 177
rect 18877 17 18935 162
rect 18986 147 19219 181
rect 18986 51 19021 147
rect 19055 17 19131 113
rect 19185 101 19219 147
rect 19257 135 19315 215
rect 19349 215 19437 257
rect 19349 135 19422 215
rect 19486 199 19567 265
rect 19603 165 19659 299
rect 19705 294 19763 527
rect 19798 459 20055 493
rect 19798 359 19867 459
rect 19798 215 19864 323
rect 19901 181 19961 425
rect 20005 391 20055 459
rect 20101 459 20535 493
rect 20101 425 20151 459
rect 20289 425 20339 459
rect 20195 391 20245 425
rect 20383 391 20433 425
rect 20005 357 20433 391
rect 20485 391 20535 459
rect 20587 425 20637 527
rect 20681 391 20731 493
rect 20775 425 20825 527
rect 20878 391 20919 493
rect 20485 357 20919 391
rect 20005 299 20055 357
rect 20126 289 20493 323
rect 20126 215 20218 289
rect 20252 215 20383 255
rect 20417 215 20493 289
rect 20527 289 20834 323
rect 20878 291 20919 357
rect 20993 294 21051 527
rect 21086 459 21533 493
rect 21086 289 21149 459
rect 21193 323 21243 425
rect 21287 357 21337 459
rect 21381 323 21431 425
rect 21483 323 21533 459
rect 21581 443 22399 493
rect 22433 443 22885 527
rect 21581 359 21631 443
rect 22349 409 22399 443
rect 22923 409 22957 493
rect 21675 367 22305 409
rect 21675 323 21734 367
rect 22349 357 22973 409
rect 23017 359 23051 527
rect 22939 323 22973 357
rect 23103 323 23153 493
rect 21193 289 21439 323
rect 21483 289 21734 323
rect 21857 289 22350 323
rect 20527 215 20593 289
rect 20800 255 20834 289
rect 21399 255 21439 289
rect 21857 265 21901 289
rect 20627 215 20763 255
rect 20800 215 20957 255
rect 21086 215 21355 255
rect 21399 219 21787 255
rect 21399 181 21439 219
rect 19468 131 19659 165
rect 19468 101 19508 131
rect 19185 51 19508 101
rect 19558 17 19624 97
rect 19705 17 19763 162
rect 19801 17 19851 179
rect 19901 173 20739 181
rect 19885 145 20739 173
rect 19885 61 19961 145
rect 20267 129 20347 145
rect 20663 129 20739 145
rect 20005 17 20143 111
rect 20177 51 20441 95
rect 20494 17 20528 111
rect 20783 95 20833 181
rect 20569 51 20833 95
rect 20877 17 20911 181
rect 20993 17 21051 162
rect 21091 17 21141 179
rect 21175 145 21439 181
rect 21175 51 21251 145
rect 21295 17 21329 111
rect 21363 51 21439 145
rect 21483 129 21709 185
rect 21743 164 21787 219
rect 21821 199 21901 265
rect 21935 199 22245 255
rect 22281 215 22350 289
rect 22385 289 22895 323
rect 22939 289 23153 323
rect 23201 294 23259 527
rect 23389 459 23769 493
rect 23295 359 23345 459
rect 23389 411 23455 459
rect 23710 427 23769 459
rect 23813 366 23863 450
rect 23907 381 23973 527
rect 23295 297 23607 359
rect 23641 347 23863 366
rect 24029 347 24081 450
rect 23641 300 24081 347
rect 22385 215 22461 289
rect 22861 255 22895 289
rect 22497 215 22819 255
rect 22861 215 23148 255
rect 23293 200 23395 263
rect 23429 200 23523 263
rect 22290 164 22494 181
rect 21743 147 22785 164
rect 21743 129 22324 147
rect 22460 129 22785 147
rect 22829 145 23067 181
rect 21483 17 21517 129
rect 21675 119 21709 129
rect 21555 85 21640 95
rect 21735 85 22305 95
rect 21555 51 22305 85
rect 22359 17 22393 111
rect 22829 95 22879 145
rect 22427 51 22879 95
rect 22923 17 22957 111
rect 22991 51 23067 145
rect 23101 17 23135 181
rect 23557 163 23607 297
rect 24121 294 24179 527
rect 24214 449 24281 493
rect 24504 451 24575 527
rect 24214 343 24265 449
rect 24609 417 24675 493
rect 24309 377 24675 417
rect 24713 387 24779 527
rect 24851 357 24903 493
rect 24214 299 24803 343
rect 23653 200 23725 266
rect 23759 200 23823 266
rect 23857 200 23937 266
rect 23971 200 24075 266
rect 24213 215 24321 255
rect 24359 215 24453 257
rect 23201 17 23259 162
rect 23295 129 23871 163
rect 23295 51 23361 129
rect 23461 17 23617 93
rect 23758 59 23871 129
rect 23987 17 24069 163
rect 24121 17 24179 162
rect 24214 17 24315 170
rect 24409 135 24453 215
rect 24501 213 24613 257
rect 24501 135 24545 213
rect 24651 196 24721 257
rect 24769 157 24803 299
rect 24618 123 24803 157
rect 24618 93 24652 123
rect 24869 117 24903 357
rect 24949 294 25007 527
rect 25043 459 25297 493
rect 25043 325 25109 459
rect 25231 451 25297 459
rect 25335 443 25406 527
rect 25153 407 25199 425
rect 25450 407 25500 493
rect 25153 359 25500 407
rect 25544 375 25610 527
rect 25654 357 25736 493
rect 25043 291 25627 325
rect 25042 215 25149 255
rect 25187 215 25292 257
rect 24370 51 24652 93
rect 24713 17 24779 89
rect 24851 51 24903 117
rect 24949 17 25007 162
rect 25043 17 25143 170
rect 25237 135 25292 215
rect 25329 215 25412 257
rect 25456 215 25547 255
rect 25329 135 25388 215
rect 25593 181 25627 291
rect 25449 147 25627 181
rect 25449 101 25483 147
rect 25672 117 25736 357
rect 25775 289 25809 527
rect 25869 294 25927 527
rect 25988 365 26038 527
rect 26082 323 26132 493
rect 26176 359 26226 527
rect 26270 323 26320 493
rect 26364 425 26414 527
rect 26468 459 26910 493
rect 26468 425 26518 459
rect 26656 425 26706 459
rect 26562 391 26612 425
rect 26750 391 26800 425
rect 25961 289 26320 323
rect 26364 357 26800 391
rect 26844 391 26910 459
rect 26954 425 27004 527
rect 27048 391 27098 493
rect 27142 425 27192 527
rect 27245 391 27286 493
rect 26844 357 27286 391
rect 25198 51 25483 101
rect 25525 17 25601 113
rect 25654 51 25736 117
rect 25775 17 25809 197
rect 25961 181 26018 289
rect 26364 255 26430 357
rect 26052 215 26430 255
rect 26468 289 26860 323
rect 26468 215 26585 289
rect 26619 215 26750 255
rect 26784 215 26860 289
rect 26894 289 27201 323
rect 27245 291 27286 357
rect 27341 294 27399 527
rect 27435 459 27691 493
rect 27435 323 27501 459
rect 27623 439 27691 459
rect 27727 451 27798 527
rect 27545 396 27579 423
rect 27837 396 27871 433
rect 27545 357 27871 396
rect 27928 371 27981 527
rect 27435 289 28043 323
rect 28077 294 28135 527
rect 28171 331 28221 493
rect 28255 459 28717 493
rect 28255 365 28315 459
rect 28349 331 28425 425
rect 28469 365 28503 459
rect 28537 331 28624 425
rect 28171 297 28624 331
rect 28667 331 28717 459
rect 28761 365 28795 527
rect 28829 331 28925 493
rect 28969 365 29003 527
rect 29037 331 29113 493
rect 28667 297 29113 331
rect 26894 215 26970 289
rect 27167 255 27201 289
rect 27014 215 27123 255
rect 27167 215 27307 255
rect 26372 181 26430 215
rect 25869 17 25927 162
rect 25961 145 26328 181
rect 26372 147 27106 181
rect 25996 17 26030 111
rect 26064 53 26140 145
rect 26184 17 26218 111
rect 26252 51 26328 145
rect 26628 129 26725 147
rect 27021 129 27106 147
rect 26372 17 26510 111
rect 26544 51 26808 95
rect 26861 17 26895 111
rect 27150 95 27200 179
rect 26936 51 27200 95
rect 27244 17 27278 179
rect 27341 17 27399 162
rect 27441 153 27541 255
rect 27579 215 27679 255
rect 27629 135 27679 215
rect 27721 211 27833 255
rect 27721 135 27763 211
rect 27869 199 27941 255
rect 27975 165 28043 289
rect 28182 215 28318 255
rect 28358 215 28501 255
rect 27835 131 28043 165
rect 27435 17 27535 119
rect 27835 101 27871 131
rect 27590 51 27871 101
rect 27917 17 27983 97
rect 28077 17 28135 162
rect 28171 136 28409 170
rect 28538 169 28624 297
rect 29181 294 29239 527
rect 29274 459 30189 493
rect 29274 291 29341 459
rect 29385 325 29427 425
rect 29471 359 29521 459
rect 29565 325 29615 425
rect 29659 359 29709 459
rect 29753 325 29803 425
rect 29847 359 29897 459
rect 29941 325 29991 425
rect 29385 289 29991 325
rect 30035 325 30189 459
rect 30233 359 30283 527
rect 30327 325 30377 493
rect 30421 359 30471 527
rect 30515 325 30565 493
rect 30609 359 30659 527
rect 30703 325 30753 493
rect 30797 359 30847 527
rect 30891 325 30941 493
rect 30035 291 30941 325
rect 31021 294 31079 527
rect 28681 215 28859 255
rect 28906 215 29076 255
rect 29274 215 29675 255
rect 28171 51 28221 136
rect 28255 17 28331 102
rect 28375 101 28409 136
rect 28443 135 28811 169
rect 28875 136 29127 170
rect 28875 101 28909 136
rect 28375 51 28613 101
rect 28651 51 28909 101
rect 28948 17 29024 102
rect 29063 51 29127 136
rect 29181 17 29239 162
rect 29275 145 29701 181
rect 29275 51 29341 145
rect 29385 17 29419 111
rect 29453 51 29529 145
rect 29573 17 29607 111
rect 29641 95 29701 145
rect 29735 177 29795 289
rect 29829 215 30144 255
rect 30191 215 30513 257
rect 30558 215 30963 257
rect 29735 129 30479 177
rect 30523 145 30949 181
rect 30523 95 30573 145
rect 29641 51 30093 95
rect 30131 51 30573 95
rect 30617 17 30651 111
rect 30685 51 30761 145
rect 30805 17 30839 111
rect 30873 51 30949 145
rect 31021 17 31079 162
rect 31113 51 31165 493
rect 31199 447 31275 527
rect 31522 474 31573 493
rect 31327 440 31573 474
rect 31617 451 31685 485
rect 31327 395 31371 440
rect 31199 361 31371 395
rect 31522 413 31573 440
rect 31199 199 31233 361
rect 31434 343 31468 381
rect 31522 379 31616 413
rect 31285 199 31361 323
rect 31434 309 31538 343
rect 31395 199 31442 275
rect 31504 165 31538 309
rect 31349 131 31538 165
rect 31572 174 31616 379
rect 31651 401 31685 451
rect 31727 435 31779 527
rect 31823 401 31859 493
rect 31651 367 31859 401
rect 31675 208 31727 331
rect 31572 140 31667 174
rect 31769 153 31821 331
rect 31941 294 31999 527
rect 32053 289 32087 527
rect 32121 305 32182 493
rect 32216 447 32292 527
rect 32556 474 32590 493
rect 32344 440 32590 474
rect 32641 451 32707 485
rect 32344 395 32388 440
rect 32216 361 32388 395
rect 32544 413 32590 440
rect 31199 17 31295 106
rect 31349 51 31383 131
rect 31430 17 31574 97
rect 31633 51 31667 140
rect 31794 17 31884 119
rect 31941 17 31999 162
rect 32053 17 32087 186
rect 32121 162 32165 305
rect 32216 265 32260 361
rect 32451 343 32485 381
rect 32544 379 32636 413
rect 32199 199 32260 265
rect 32305 199 32379 323
rect 32451 309 32558 343
rect 32413 199 32483 275
rect 32524 165 32558 309
rect 32121 51 32182 162
rect 32369 131 32558 165
rect 32592 174 32636 379
rect 32673 401 32707 451
rect 32751 435 32801 527
rect 32845 401 32879 493
rect 32673 367 32879 401
rect 32676 210 32768 331
rect 32592 140 32672 174
rect 32832 153 32907 331
rect 32953 294 33011 527
rect 33055 391 33105 493
rect 33149 425 33199 527
rect 33243 391 33293 493
rect 33337 425 33387 527
rect 33431 459 33669 493
rect 33431 391 33481 459
rect 33619 427 33669 459
rect 33723 427 33773 527
rect 33817 459 34055 493
rect 33817 427 33867 459
rect 33055 357 33481 391
rect 33045 289 33395 323
rect 33439 291 33481 357
rect 33525 393 33575 425
rect 33911 393 33961 425
rect 33045 215 33153 289
rect 33199 215 33317 255
rect 33361 249 33395 289
rect 33525 283 33602 393
rect 33715 357 33961 393
rect 34005 357 34055 459
rect 34099 359 34149 527
rect 34193 391 34243 493
rect 34287 433 34337 527
rect 34381 391 34431 493
rect 34193 357 34431 391
rect 34475 365 34525 527
rect 33715 333 33749 357
rect 33679 299 33749 333
rect 34381 331 34431 357
rect 33361 215 33447 249
rect 33525 181 33567 283
rect 33679 249 33717 299
rect 33783 289 34121 323
rect 33783 265 33829 289
rect 33601 215 33717 249
rect 33751 215 33829 265
rect 33869 215 34011 255
rect 34045 215 34121 289
rect 34155 249 34230 323
rect 34381 283 34563 331
rect 34609 294 34667 527
rect 34703 361 34769 527
rect 34869 323 34945 493
rect 34988 391 35061 493
rect 35095 447 35183 493
rect 35149 391 35183 447
rect 35217 427 35267 527
rect 35311 391 35362 493
rect 34988 357 35115 391
rect 35149 357 35362 391
rect 34155 215 34446 249
rect 33679 181 33717 215
rect 34490 181 34563 283
rect 34714 199 34788 323
rect 34869 289 35047 323
rect 34839 202 34952 255
rect 32216 17 32312 106
rect 32369 51 32403 131
rect 32447 17 32594 97
rect 32638 51 32672 140
rect 32797 17 32887 119
rect 32953 17 33011 162
rect 33063 17 33097 179
rect 33131 95 33191 181
rect 33225 147 33583 181
rect 33225 129 33302 147
rect 33131 51 33395 95
rect 33439 17 33473 111
rect 33507 51 33583 147
rect 33679 145 34063 181
rect 33627 17 33765 111
rect 33799 51 33875 145
rect 33919 17 33953 111
rect 33987 51 34063 145
rect 34107 17 34141 179
rect 34175 145 34563 181
rect 35013 166 35047 289
rect 34175 55 34251 145
rect 34295 17 34329 111
rect 34363 55 34439 145
rect 34483 17 34517 111
rect 34609 17 34667 162
rect 34703 17 34769 165
rect 34813 132 35047 166
rect 35081 165 35115 357
rect 35161 199 35207 323
rect 35261 199 35329 323
rect 35437 294 35495 527
rect 35539 391 35589 493
rect 35633 427 35683 527
rect 35727 391 35777 493
rect 35821 427 35871 527
rect 35915 459 36153 493
rect 35915 391 35965 459
rect 35539 357 35965 391
rect 35534 289 35931 323
rect 35534 215 35640 289
rect 35683 215 35801 255
rect 35855 215 35931 289
rect 34813 51 34847 132
rect 34893 17 35027 98
rect 35081 51 35139 165
rect 35173 85 35207 199
rect 36001 181 36067 425
rect 36103 359 36153 459
rect 36207 393 36257 493
rect 36301 427 36351 527
rect 36395 459 36633 493
rect 36395 393 36445 459
rect 36207 357 36445 393
rect 36489 323 36539 425
rect 36135 289 36539 323
rect 36583 291 36633 459
rect 36725 294 36783 527
rect 36817 325 36885 493
rect 36929 359 36971 527
rect 37015 393 37063 493
rect 37109 427 37159 527
rect 37203 393 37253 493
rect 37297 427 37347 527
rect 37391 393 37441 493
rect 37485 427 37535 527
rect 37579 459 38013 493
rect 37579 393 37629 459
rect 37015 359 37629 393
rect 37015 325 37063 359
rect 36817 291 37063 325
rect 37673 323 37723 425
rect 37767 359 37815 459
rect 37849 323 37903 425
rect 37107 289 37595 323
rect 36135 265 36169 289
rect 36111 199 36169 265
rect 37107 257 37141 289
rect 36207 215 36406 255
rect 36456 215 36599 255
rect 36820 215 37141 257
rect 37175 215 37485 255
rect 37519 215 37595 289
rect 37629 283 37903 323
rect 37937 291 38013 459
rect 38051 325 38117 493
rect 38161 359 38203 527
rect 38248 325 38296 493
rect 38341 359 38391 527
rect 38435 459 38862 493
rect 38435 325 38485 459
rect 38051 291 38485 325
rect 38529 325 38579 425
rect 38623 359 38673 459
rect 38717 325 38767 425
rect 38812 359 38862 459
rect 38529 291 38892 325
rect 38933 294 38991 527
rect 39027 315 39093 485
rect 35285 17 35361 165
rect 35437 17 35495 162
rect 35547 17 35581 179
rect 35615 95 35675 179
rect 35709 145 36067 181
rect 36135 181 36169 199
rect 37629 181 37673 283
rect 37707 215 38065 249
rect 38109 215 38414 255
rect 38488 215 38793 255
rect 38031 181 38065 215
rect 38827 181 38892 291
rect 36135 145 36547 181
rect 35709 129 35785 145
rect 35615 51 35879 95
rect 35923 17 35957 111
rect 35991 51 36067 145
rect 36111 17 36249 111
rect 36283 51 36359 145
rect 36403 17 36437 111
rect 36471 51 36547 145
rect 36591 17 36625 181
rect 36725 17 36783 162
rect 36835 17 36869 179
rect 36903 145 37151 181
rect 36903 51 36979 145
rect 37023 17 37057 111
rect 37091 95 37151 145
rect 37185 145 37919 181
rect 38031 147 38892 181
rect 39027 162 39065 315
rect 39137 299 39187 527
rect 39225 399 39285 483
rect 39341 433 39407 527
rect 39463 399 39513 483
rect 39225 365 39513 399
rect 39559 365 39625 485
rect 39223 265 39276 331
rect 39099 199 39171 265
rect 39205 199 39276 265
rect 39311 199 39371 331
rect 39405 199 39463 331
rect 39497 199 39557 331
rect 39137 165 39171 199
rect 39591 165 39625 365
rect 39669 294 39727 527
rect 39771 435 39821 527
rect 39873 401 39907 493
rect 39762 367 39907 401
rect 39941 367 40001 527
rect 40035 401 40095 485
rect 40147 435 40213 527
rect 40261 401 40323 485
rect 40035 367 40323 401
rect 37185 129 37459 145
rect 37091 51 37543 95
rect 37587 17 37621 111
rect 37655 55 37731 145
rect 37775 17 37809 111
rect 37843 55 37919 145
rect 38135 145 38775 147
rect 37963 17 38101 111
rect 38135 51 38211 145
rect 38255 17 38289 111
rect 38323 51 38399 145
rect 38443 17 38477 111
rect 38511 51 38587 145
rect 38631 17 38665 111
rect 38699 51 38775 145
rect 38819 17 38853 111
rect 38933 17 38991 162
rect 39027 60 39093 162
rect 39137 131 39625 165
rect 39762 177 39813 367
rect 40379 333 40413 493
rect 39847 299 40413 333
rect 39847 249 39881 299
rect 39847 215 39913 249
rect 39950 199 40053 265
rect 39129 17 39195 97
rect 39433 63 39509 131
rect 39553 17 39619 97
rect 39669 17 39727 162
rect 39762 143 39907 177
rect 39950 152 40018 199
rect 39762 17 39829 93
rect 39873 51 39907 143
rect 39945 17 40021 93
rect 40125 80 40175 265
rect 40221 83 40267 265
rect 40301 51 40335 299
rect 40497 294 40555 527
rect 40607 391 40641 493
rect 40675 425 40751 527
rect 40795 391 40829 493
rect 40863 425 40939 527
rect 40983 391 41017 493
rect 41051 425 41127 527
rect 41195 459 41417 493
rect 41195 391 41229 459
rect 40607 357 41229 391
rect 41263 325 41339 423
rect 41383 359 41417 459
rect 41471 425 41537 527
rect 41581 391 41615 493
rect 41649 425 41725 527
rect 41769 391 41803 493
rect 41837 425 41913 527
rect 41559 357 41928 391
rect 40601 289 41203 323
rect 40383 151 40451 265
rect 40601 215 40677 289
rect 40727 181 40823 255
rect 40863 215 40943 255
rect 41009 215 41085 255
rect 41127 215 41203 289
rect 41263 291 41536 325
rect 41009 181 41046 215
rect 40379 17 40437 113
rect 40497 17 40555 162
rect 40607 17 40641 181
rect 40727 147 41046 181
rect 41263 174 41311 291
rect 41502 265 41536 291
rect 41357 215 41463 257
rect 41092 161 41311 174
rect 41092 140 41339 161
rect 41415 149 41463 215
rect 41502 199 41843 265
rect 41889 165 41928 357
rect 41969 294 42027 527
rect 42062 299 42128 527
rect 42172 401 42207 483
rect 42251 435 42317 527
rect 42368 401 42407 483
rect 42172 367 42407 401
rect 42257 289 42383 333
rect 42061 199 42131 265
rect 41092 113 41126 140
rect 40863 79 41126 113
rect 41162 17 41229 106
rect 41263 59 41339 140
rect 41553 131 41928 165
rect 41399 17 41505 113
rect 41649 17 41725 97
rect 41837 17 41913 97
rect 41969 17 42027 162
rect 42062 17 42130 163
rect 42165 67 42277 255
rect 42318 199 42383 289
rect 42441 299 42526 489
rect 42441 165 42475 299
rect 42613 294 42671 527
rect 42723 391 42757 493
rect 42791 425 42867 527
rect 42911 391 42945 493
rect 42979 425 43055 527
rect 43099 391 43133 493
rect 43200 425 43344 527
rect 43425 459 43663 493
rect 43425 391 43459 459
rect 42723 357 43459 391
rect 43519 323 43585 423
rect 43629 359 43663 459
rect 42509 199 42574 265
rect 42717 199 42862 323
rect 42918 199 43069 323
rect 43154 199 43306 323
rect 43354 289 43585 323
rect 43354 169 43417 289
rect 43631 255 43676 325
rect 43717 294 43775 527
rect 43827 333 43861 493
rect 43895 383 43971 527
rect 44015 333 44049 493
rect 44083 383 44159 527
rect 44203 333 44237 493
rect 44271 383 44347 527
rect 44391 333 44425 493
rect 44459 383 44535 527
rect 44579 333 44613 493
rect 44651 383 44727 527
rect 44771 333 44805 493
rect 44839 451 44915 527
rect 44959 485 44993 493
rect 44959 451 45495 485
rect 44959 333 44993 451
rect 45137 383 45409 417
rect 43827 299 44993 333
rect 43532 215 43676 255
rect 43816 199 44169 265
rect 44219 199 44582 265
rect 44637 199 44996 265
rect 45046 199 45313 326
rect 43354 165 43679 169
rect 42340 59 42475 165
rect 42509 17 42561 113
rect 42613 17 42671 162
rect 42707 131 43149 165
rect 43197 131 43679 165
rect 42791 17 42867 93
rect 42979 59 43363 93
rect 43409 51 43443 131
rect 43493 17 43569 93
rect 43603 59 43679 131
rect 43717 17 43775 162
rect 45361 161 45409 383
rect 45445 299 45495 451
rect 45557 294 45615 527
rect 45650 383 45717 485
rect 43827 127 44629 161
rect 44677 127 45479 161
rect 43827 51 43861 127
rect 43895 17 43971 93
rect 44015 51 44049 127
rect 44083 17 44159 93
rect 44203 51 44237 127
rect 44271 59 45025 93
rect 45137 17 45213 93
rect 45257 51 45291 127
rect 45325 17 45401 93
rect 45445 51 45479 127
rect 45557 17 45615 162
rect 45650 112 45701 383
rect 45777 367 45843 527
rect 45902 409 45959 493
rect 46020 443 46086 527
rect 46141 459 46411 493
rect 46141 409 46207 459
rect 45902 375 46207 409
rect 46263 333 46297 425
rect 46359 359 46411 459
rect 45767 299 46297 333
rect 45767 265 45801 299
rect 46390 265 46438 323
rect 46477 294 46535 527
rect 46579 391 46621 493
rect 46655 425 46731 527
rect 46775 391 46809 493
rect 46579 357 46809 391
rect 46879 459 47101 493
rect 46879 357 46913 459
rect 46957 389 47023 423
rect 47067 393 47101 459
rect 47135 428 47211 527
rect 47287 393 47321 493
rect 45746 199 45801 265
rect 45835 199 45903 265
rect 45767 165 45801 199
rect 45767 131 45895 165
rect 45937 133 46022 265
rect 46084 191 46165 265
rect 46108 133 46165 191
rect 46199 132 46259 265
rect 46318 199 46438 265
rect 46579 165 46621 357
rect 46957 323 47007 389
rect 47067 359 47321 393
rect 47355 383 47432 527
rect 46659 289 47007 323
rect 46659 199 46703 289
rect 45650 60 45717 112
rect 45861 97 45895 131
rect 45751 17 45827 97
rect 45861 63 46214 97
rect 46333 17 46409 161
rect 46477 17 46535 162
rect 46579 131 46731 165
rect 46765 149 46878 255
rect 46912 169 46960 289
rect 47041 249 47086 323
rect 46999 215 47086 249
rect 46912 135 47093 169
rect 46570 17 46637 93
rect 46749 17 46900 89
rect 47033 59 47093 135
rect 47127 83 47181 265
rect 47215 85 47282 325
rect 47385 199 47453 326
rect 47489 294 47547 527
rect 47583 383 47649 527
rect 47693 333 47727 493
rect 47761 383 47837 527
rect 47881 333 47915 493
rect 47949 383 48025 527
rect 48069 417 48103 493
rect 48137 451 48213 527
rect 48267 417 48301 493
rect 48335 451 48411 527
rect 48455 417 48489 493
rect 48523 451 48599 527
rect 48643 451 49201 485
rect 48643 417 48677 451
rect 48069 383 48677 417
rect 48853 415 49107 417
rect 48720 383 49107 415
rect 48720 381 48866 383
rect 48720 333 48754 381
rect 49151 351 49201 451
rect 47588 299 47915 333
rect 47954 299 48754 333
rect 47355 17 47432 161
rect 47489 17 47547 162
rect 47588 161 47632 299
rect 47954 265 47998 299
rect 47688 199 47998 265
rect 48046 215 48245 259
rect 48291 215 48450 265
rect 48500 215 48679 265
rect 47588 127 47915 161
rect 47583 17 47649 93
rect 47693 51 47727 127
rect 47761 17 47837 93
rect 47881 51 47915 127
rect 48069 131 48411 165
rect 48720 161 48754 299
rect 48788 215 48992 325
rect 49052 259 49091 327
rect 49237 294 49295 527
rect 49329 451 49601 493
rect 49329 367 49381 451
rect 49415 357 49495 417
rect 49551 391 49601 451
rect 49653 427 49703 527
rect 49755 391 49789 493
rect 49551 357 49789 391
rect 49052 215 49198 259
rect 49329 199 49381 265
rect 47949 17 48025 93
rect 48069 51 48103 131
rect 48523 127 48911 161
rect 48963 129 49185 163
rect 48963 93 48997 129
rect 48137 17 48213 93
rect 48251 59 48693 93
rect 48750 59 48997 93
rect 48963 51 48997 59
rect 49031 17 49107 93
rect 49151 51 49185 129
rect 49237 17 49295 162
rect 49415 161 49467 357
rect 49755 349 49789 357
rect 49501 199 49559 323
rect 49823 299 49901 527
rect 49973 294 50031 527
rect 50083 459 50493 493
rect 50083 359 50117 459
rect 50161 325 50227 425
rect 50271 359 50305 459
rect 50365 325 50399 425
rect 50459 393 50493 459
rect 50537 451 50681 527
rect 50731 393 50765 493
rect 50802 451 50953 527
rect 50987 393 51021 493
rect 51073 451 51217 527
rect 51267 393 51301 493
rect 50459 359 51301 393
rect 49415 127 49565 161
rect 49334 17 49400 93
rect 49505 59 49565 127
rect 49607 69 49651 265
rect 49709 83 49749 265
rect 49790 203 49883 265
rect 50077 257 50113 325
rect 50161 291 50487 325
rect 50077 215 50223 257
rect 50261 215 50407 257
rect 49826 17 49904 161
rect 49973 17 50031 162
rect 50067 143 50305 177
rect 50441 165 50487 291
rect 50523 215 50699 325
rect 50792 215 50963 325
rect 51053 215 51312 325
rect 51353 294 51411 527
rect 51447 451 52249 485
rect 51450 261 51494 393
rect 51531 349 51607 417
rect 51719 349 51795 417
rect 51863 349 51983 417
rect 52095 349 52171 417
rect 51531 315 52171 349
rect 52215 349 52249 451
rect 52287 383 52363 527
rect 52407 349 52441 493
rect 52492 383 52636 527
rect 52686 349 52720 493
rect 52801 383 52877 527
rect 52921 349 52955 493
rect 52989 383 53065 527
rect 53109 349 53143 493
rect 53281 383 53357 527
rect 53401 349 53435 493
rect 53469 383 53545 527
rect 53589 349 53623 493
rect 52215 315 53623 349
rect 51450 215 51808 261
rect 51863 198 51951 315
rect 53745 294 53803 527
rect 53845 393 53901 527
rect 53945 349 54005 459
rect 54039 383 54105 527
rect 54166 383 54251 493
rect 53840 265 53911 337
rect 53945 315 54135 349
rect 54101 265 54135 315
rect 51995 199 52219 265
rect 52263 215 52641 257
rect 52777 215 53137 260
rect 53257 215 53635 256
rect 53840 215 53953 265
rect 53997 215 54067 265
rect 50067 59 50133 143
rect 50177 17 50211 109
rect 50255 93 50305 143
rect 50339 131 50697 165
rect 50799 127 51208 161
rect 50255 59 50509 93
rect 50547 59 50969 93
rect 51021 17 51098 93
rect 51132 55 51208 127
rect 51267 17 51301 177
rect 51353 17 51411 162
rect 51907 161 51951 198
rect 51463 127 51873 161
rect 51907 127 52661 161
rect 52801 127 53529 161
rect 53579 151 53635 215
rect 54101 199 54152 265
rect 54101 181 54135 199
rect 51463 51 51497 127
rect 51531 17 51607 93
rect 51651 51 51685 127
rect 51839 93 51873 127
rect 51719 17 51795 93
rect 51839 59 52265 93
rect 52313 59 53159 93
rect 53197 17 53263 93
rect 53307 51 53341 127
rect 53375 17 53451 93
rect 53495 51 53529 127
rect 53565 17 53643 93
rect 53745 17 53803 162
rect 53845 143 54135 181
rect 53845 71 53911 143
rect 54192 109 54251 383
rect 54297 294 54355 527
rect 54395 393 54451 527
rect 54391 265 54442 353
rect 54495 349 54555 459
rect 54605 383 54673 527
rect 54721 383 54813 493
rect 54495 315 54693 349
rect 54659 265 54693 315
rect 54391 215 54515 265
rect 54549 215 54625 265
rect 54659 199 54725 265
rect 54659 181 54693 199
rect 54041 17 54091 109
rect 54125 51 54251 109
rect 54297 17 54355 162
rect 54395 143 54693 181
rect 54395 71 54461 143
rect 54759 109 54813 383
rect 54847 299 54905 527
rect 54941 294 54999 527
rect 55035 376 55101 527
rect 55147 350 55183 493
rect 55234 387 55300 527
rect 55352 352 55390 493
rect 55424 387 55500 527
rect 55544 353 55582 493
rect 55616 387 55692 527
rect 55544 352 55730 353
rect 55041 199 55103 323
rect 55147 316 55308 350
rect 55266 271 55308 316
rect 55352 307 55730 352
rect 55137 199 55232 265
rect 55266 204 55603 271
rect 54607 17 54657 109
rect 54691 51 54813 109
rect 54847 17 54905 177
rect 54941 17 54999 162
rect 55266 161 55308 204
rect 55674 169 55730 307
rect 55769 294 55827 527
rect 55879 403 55913 489
rect 55947 437 56023 527
rect 55879 357 56024 403
rect 55035 123 55308 161
rect 55352 123 55730 169
rect 55035 51 55101 123
rect 55352 103 55390 123
rect 55227 17 55293 89
rect 55424 17 55500 89
rect 55544 51 55582 123
rect 55616 17 55692 89
rect 55769 17 55827 162
rect 55873 153 55933 323
rect 55977 227 56024 357
rect 56058 295 56125 484
rect 56171 433 56299 527
rect 56170 329 56299 391
rect 56333 316 56460 473
rect 56058 265 56260 295
rect 56058 261 56345 265
rect 55977 161 56094 227
rect 56128 189 56345 261
rect 55977 131 56021 161
rect 55862 17 55929 118
rect 55973 56 56021 131
rect 56128 122 56172 189
rect 56398 155 56460 316
rect 56505 294 56563 527
rect 56615 403 56649 489
rect 56683 437 56759 527
rect 56615 357 56761 403
rect 56087 83 56172 122
rect 56087 54 56121 83
rect 56244 17 56333 116
rect 56385 51 56460 155
rect 56505 17 56563 162
rect 56609 153 56670 323
rect 56714 227 56761 357
rect 56799 295 56866 484
rect 56912 433 57059 527
rect 56911 329 57060 391
rect 57095 316 57198 473
rect 57245 336 57299 527
rect 56799 265 57001 295
rect 56799 261 57087 265
rect 56714 161 56835 227
rect 56869 189 57087 261
rect 56714 131 56757 161
rect 56599 17 56665 118
rect 56709 56 56757 131
rect 56869 122 56913 189
rect 57131 155 57198 316
rect 57333 294 57391 527
rect 57426 451 57493 527
rect 57626 455 57692 527
rect 57819 455 57895 527
rect 58007 455 58083 527
rect 57441 383 58196 417
rect 57441 265 57475 383
rect 57511 300 57691 349
rect 57735 307 58004 349
rect 57657 297 57691 300
rect 57657 271 57692 297
rect 57441 199 57493 265
rect 57529 199 57623 265
rect 57657 199 57843 271
rect 56823 83 56913 122
rect 56823 54 56857 83
rect 57001 17 57075 116
rect 57119 51 57198 155
rect 57245 17 57299 144
rect 57333 17 57391 162
rect 57657 161 57699 199
rect 57897 165 58004 307
rect 57426 123 57699 161
rect 57743 123 58004 165
rect 58048 125 58117 349
rect 57426 51 57493 123
rect 57743 99 57781 123
rect 58153 99 58196 383
rect 58253 294 58311 527
rect 58345 416 58476 527
rect 58511 425 58627 493
rect 58710 418 58761 527
rect 58345 396 58478 416
rect 58431 391 58478 396
rect 58345 272 58397 362
rect 58431 342 58507 391
rect 58560 318 58761 377
rect 58805 353 58860 493
rect 58560 308 58782 318
rect 58507 274 58782 308
rect 58507 272 58543 274
rect 58345 238 58543 272
rect 57619 17 57685 89
rect 57815 17 57891 89
rect 58007 17 58083 89
rect 58253 17 58311 162
rect 58345 127 58465 204
rect 58499 93 58543 238
rect 58345 59 58543 93
rect 58606 61 58680 240
rect 58736 198 58782 274
rect 58826 147 58860 353
rect 58897 294 58955 527
rect 58989 426 59125 527
rect 58992 319 59043 392
rect 59077 391 59125 426
rect 59161 425 59276 493
rect 59077 353 59153 391
rect 59208 319 59268 378
rect 59313 358 59356 527
rect 59406 359 59496 493
rect 58992 285 59380 319
rect 58714 17 58748 125
rect 58808 51 58860 147
rect 58897 17 58955 162
rect 58989 153 59066 249
rect 59110 114 59151 285
rect 58993 61 59151 114
rect 59185 150 59297 249
rect 59334 199 59380 285
rect 59424 289 59496 359
rect 59530 325 59582 527
rect 59633 294 59691 527
rect 59424 185 59557 289
rect 59731 268 59774 467
rect 59808 350 59844 493
rect 59887 387 59987 527
rect 60032 350 60068 493
rect 60120 387 60186 527
rect 60238 352 60276 493
rect 60310 387 60386 527
rect 60430 353 60468 493
rect 60502 387 60578 527
rect 60430 352 60606 353
rect 59808 316 60194 350
rect 60152 271 60194 316
rect 60238 307 60606 352
rect 59731 199 59883 268
rect 59185 61 59235 150
rect 59424 143 59458 185
rect 59269 17 59335 116
rect 59369 51 59458 143
rect 59511 17 59566 149
rect 59633 17 59691 162
rect 59801 89 59868 161
rect 59917 149 59979 268
rect 60013 199 60118 265
rect 60152 204 60489 271
rect 60152 161 60194 204
rect 60550 169 60606 307
rect 60645 294 60703 527
rect 60737 425 60789 527
rect 60737 215 60805 391
rect 60849 249 60883 493
rect 60937 426 61070 527
rect 61021 391 61070 426
rect 61104 425 61219 493
rect 61279 418 61322 527
rect 60937 319 60987 388
rect 61021 353 61097 391
rect 61151 319 61330 378
rect 61374 353 61427 493
rect 60937 315 61330 319
rect 60937 285 61357 315
rect 60849 199 61024 249
rect 60849 181 60899 199
rect 60035 123 60194 161
rect 60238 123 60606 169
rect 60035 89 60073 123
rect 60238 103 60276 123
rect 59801 51 60073 89
rect 60119 17 60185 89
rect 60310 17 60386 89
rect 60430 51 60468 123
rect 60502 17 60578 89
rect 60645 17 60703 162
rect 60737 17 60789 181
rect 60823 97 60899 181
rect 61058 110 61109 285
rect 60941 57 61109 110
rect 61176 61 61249 251
rect 61313 195 61357 285
rect 61393 147 61427 353
rect 61473 294 61531 527
rect 61565 315 61628 527
rect 61764 426 61897 527
rect 61283 17 61341 125
rect 61375 51 61427 147
rect 61473 17 61531 162
rect 61577 149 61630 265
rect 61674 249 61729 381
rect 61768 319 61815 392
rect 61849 391 61897 426
rect 61931 425 62046 493
rect 61849 353 61925 391
rect 61980 319 62018 378
rect 62080 358 62123 527
rect 62173 359 62266 493
rect 61768 285 62152 319
rect 61674 203 61841 249
rect 61565 17 61619 115
rect 61674 61 61729 203
rect 61877 114 61911 285
rect 61769 61 61911 114
rect 61945 153 62072 249
rect 62106 199 62152 285
rect 62196 289 62266 359
rect 62300 325 62353 527
rect 62393 294 62451 527
rect 62614 455 62714 527
rect 62847 455 62913 527
rect 63037 455 63114 527
rect 63229 455 63305 527
rect 62498 299 62570 433
rect 62604 375 63449 421
rect 62196 185 62356 289
rect 61945 61 62022 153
rect 62196 143 62262 185
rect 62070 17 62136 116
rect 62181 51 62262 143
rect 62300 17 62353 149
rect 62393 17 62451 162
rect 62498 161 62542 299
rect 62604 265 62641 375
rect 62734 305 62909 339
rect 62943 307 63267 341
rect 62875 271 62909 305
rect 62576 199 62641 265
rect 62498 109 62595 161
rect 62675 145 62725 268
rect 62766 199 62841 268
rect 62875 204 63148 271
rect 62875 161 62921 204
rect 63182 169 63267 307
rect 62772 123 62921 161
rect 62965 123 63267 169
rect 63301 123 63359 341
rect 62772 109 62808 123
rect 62498 71 62808 109
rect 62965 103 63003 123
rect 62498 51 62595 71
rect 62854 17 62920 89
rect 63037 17 63107 89
rect 63141 51 63195 123
rect 63229 17 63305 89
rect 63393 85 63449 375
rect 63497 294 63555 527
rect 63590 451 63657 527
rect 63497 17 63555 162
rect 63589 153 63637 415
rect 63693 333 63743 493
rect 63779 383 63845 527
rect 63884 333 63934 493
rect 63973 367 64047 527
rect 64111 441 64189 493
rect 63671 299 64079 333
rect 63671 117 63709 299
rect 63606 51 63709 117
rect 63743 72 63819 265
rect 63853 71 63911 265
rect 63949 143 64005 265
rect 64039 199 64079 299
rect 64137 161 64189 441
rect 64233 294 64291 527
rect 64327 451 64393 527
rect 63985 17 64039 109
rect 64111 59 64189 161
rect 64233 17 64291 162
rect 64333 151 64374 415
rect 64437 333 64471 493
rect 64515 383 64581 527
rect 64622 333 64672 493
rect 64741 367 64791 527
rect 64833 367 64923 493
rect 64957 367 65021 527
rect 64408 299 64841 333
rect 64408 117 64442 299
rect 64343 51 64442 117
rect 64479 84 64555 265
rect 64589 83 64649 265
rect 64685 148 64739 265
rect 64807 199 64841 299
rect 64875 161 64923 367
rect 65061 294 65119 527
rect 65157 367 65213 527
rect 65257 333 65299 493
rect 65347 387 65413 527
rect 65457 333 65495 493
rect 65581 371 65647 527
rect 64765 17 64799 110
rect 64833 59 64923 161
rect 64957 17 65023 162
rect 65061 17 65119 162
rect 65161 153 65202 331
rect 65236 299 65659 333
rect 65236 117 65280 299
rect 65171 51 65280 117
rect 65314 84 65405 265
rect 65439 85 65492 265
rect 65533 146 65591 265
rect 65625 261 65659 299
rect 65693 331 65743 493
rect 65787 367 65837 527
rect 65881 349 65915 493
rect 65949 383 66025 527
rect 65881 331 66027 349
rect 65693 297 66027 331
rect 65625 215 65923 261
rect 65976 162 66027 297
rect 66073 294 66131 527
rect 66182 403 66217 493
rect 66251 439 66327 527
rect 66388 409 66422 493
rect 66479 445 66623 527
rect 66674 409 66708 493
rect 66760 445 66826 527
rect 66182 369 66318 403
rect 66165 199 66238 335
rect 66284 265 66318 369
rect 66388 375 66831 409
rect 66284 199 66353 265
rect 66284 165 66318 199
rect 65693 128 66027 162
rect 65581 17 65643 110
rect 65693 51 65727 128
rect 65761 17 65837 94
rect 65881 51 65915 128
rect 65949 17 66025 94
rect 66073 17 66131 162
rect 66182 131 66318 165
rect 66182 51 66217 131
rect 66388 117 66422 375
rect 66251 17 66327 93
rect 66376 51 66422 117
rect 66483 84 66579 339
rect 66613 84 66671 339
rect 66705 133 66763 339
rect 66797 265 66831 375
rect 66875 299 66947 493
rect 66797 199 66855 265
rect 66893 161 66947 299
rect 66993 294 67051 527
rect 67103 400 67137 493
rect 67171 439 67247 527
rect 67291 417 67325 493
rect 67409 451 67553 527
rect 67602 417 67640 493
rect 67696 439 67762 527
rect 67103 366 67239 400
rect 66739 17 66818 93
rect 66852 59 66947 161
rect 66993 17 67051 162
rect 67095 148 67135 326
rect 67205 265 67239 366
rect 67291 393 67640 417
rect 67291 383 67761 393
rect 67291 332 67351 383
rect 67606 359 67761 383
rect 67205 199 67283 265
rect 67205 117 67239 199
rect 67317 117 67351 332
rect 67087 17 67153 93
rect 67197 51 67239 117
rect 67307 51 67351 117
rect 67447 84 67499 349
rect 67543 84 67591 323
rect 67625 129 67691 323
rect 67727 265 67761 359
rect 67806 333 67867 493
rect 67907 367 67958 527
rect 67806 307 67959 333
rect 67727 199 67779 265
rect 67823 165 67959 307
rect 68005 294 68063 527
rect 68097 417 68149 493
rect 68183 451 68259 527
rect 68382 451 68458 527
rect 68570 451 68646 527
rect 68782 451 68858 527
rect 68994 451 69070 527
rect 68097 383 69057 417
rect 67780 128 67959 165
rect 67670 17 67746 93
rect 67780 51 67847 128
rect 67881 17 67958 93
rect 68005 17 68063 162
rect 68097 117 68132 383
rect 68168 153 68248 327
rect 68286 309 68552 343
rect 68586 309 68986 343
rect 68286 164 68352 309
rect 68586 265 68620 309
rect 68386 199 68620 265
rect 68654 199 68704 265
rect 68286 130 68536 164
rect 68746 151 68808 265
rect 68842 147 68918 265
rect 68952 162 68986 309
rect 69023 199 69057 383
rect 69109 294 69167 527
rect 69201 427 69253 493
rect 69299 451 69375 527
rect 69201 291 69235 427
rect 69417 417 69459 493
rect 69509 451 69575 527
rect 69621 417 69655 493
rect 69694 451 69770 527
rect 69826 417 69860 493
rect 69924 451 69990 527
rect 69269 325 69347 391
rect 69417 383 69581 417
rect 69387 315 69513 349
rect 69387 291 69431 315
rect 69201 257 69431 291
rect 69547 281 69581 383
rect 68097 51 68149 117
rect 68193 17 68243 109
rect 68286 51 68348 130
rect 68382 17 68458 94
rect 68502 51 68536 130
rect 68952 128 69060 162
rect 68587 17 68653 89
rect 69109 17 69167 162
rect 69201 117 69235 257
rect 69467 247 69581 281
rect 69615 383 69980 417
rect 69289 189 69417 223
rect 69289 153 69341 189
rect 69467 151 69501 247
rect 69615 185 69649 383
rect 69201 51 69253 117
rect 69299 17 69375 93
rect 69421 85 69501 151
rect 69535 119 69649 185
rect 69683 85 69717 265
rect 69421 51 69717 85
rect 69759 83 69819 327
rect 69853 84 69912 327
rect 69946 265 69980 383
rect 70034 289 70086 493
rect 70121 294 70179 527
rect 70231 411 70265 493
rect 70299 451 70375 527
rect 70524 451 70658 527
rect 70715 417 70749 493
rect 70783 451 70861 527
rect 70905 417 70939 493
rect 71017 451 71083 527
rect 71127 417 71179 493
rect 70231 377 70611 411
rect 69946 199 70007 265
rect 70041 165 70086 289
rect 70226 199 70262 327
rect 69946 17 69980 109
rect 70034 51 70086 165
rect 70121 17 70179 162
rect 70296 161 70340 377
rect 70231 127 70340 161
rect 70409 309 70480 343
rect 70231 51 70265 127
rect 70299 17 70375 93
rect 70409 51 70464 309
rect 70577 265 70611 377
rect 70673 383 70939 417
rect 70973 383 71179 417
rect 70499 161 70543 265
rect 70577 199 70639 265
rect 70673 161 70717 383
rect 70973 349 71017 383
rect 70755 315 71017 349
rect 70755 280 70799 315
rect 70499 127 70717 161
rect 70498 17 70574 93
rect 70625 51 70659 127
rect 70850 84 70903 255
rect 70937 85 70997 281
rect 71031 153 71101 261
rect 71145 117 71179 383
rect 71225 294 71283 527
rect 71317 417 71369 493
rect 71403 451 71479 527
rect 71602 451 71678 527
rect 71790 451 71866 527
rect 72036 451 72102 527
rect 72262 451 72464 527
rect 72519 417 72553 493
rect 71317 383 72288 417
rect 71033 17 71083 117
rect 71127 51 71179 117
rect 71225 17 71283 162
rect 71317 117 71352 383
rect 71386 153 71466 327
rect 71502 309 71772 343
rect 71806 309 72210 343
rect 71502 164 71568 309
rect 71806 249 71840 309
rect 72254 275 72288 383
rect 71602 215 71840 249
rect 71502 130 71756 164
rect 71317 51 71369 117
rect 71424 17 71490 94
rect 71534 51 71568 130
rect 71602 17 71678 94
rect 71722 51 71756 130
rect 71806 157 71840 215
rect 71881 199 71939 265
rect 71806 123 71939 157
rect 71973 128 72068 265
rect 72116 241 72288 275
rect 72372 383 72553 417
rect 72116 199 72160 241
rect 72372 165 72406 383
rect 72487 199 72569 324
rect 72605 294 72663 527
rect 72713 341 72749 493
rect 72785 375 72859 527
rect 72713 307 72858 341
rect 72893 312 72959 493
rect 72824 278 72858 307
rect 72701 197 72789 271
rect 72824 212 72887 278
rect 71895 94 71939 123
rect 72242 94 72312 162
rect 72372 131 72553 165
rect 71794 17 71860 89
rect 71895 60 72312 94
rect 72377 17 72443 93
rect 72519 51 72553 131
rect 72605 17 72663 162
rect 72824 161 72858 212
rect 72715 127 72858 161
rect 72923 152 72959 312
rect 73065 294 73123 527
rect 73175 367 73209 527
rect 73243 323 73319 493
rect 73363 367 73397 527
rect 73431 323 73507 493
rect 73551 367 73585 527
rect 73645 323 73679 493
rect 73713 367 73789 527
rect 73833 323 73867 493
rect 73901 367 73977 527
rect 74021 323 74055 493
rect 74089 367 74165 527
rect 74209 323 74243 493
rect 74277 367 74353 527
rect 74397 323 74431 493
rect 74465 367 74541 527
rect 74585 323 74619 493
rect 73243 289 73583 323
rect 73645 289 74619 323
rect 74653 297 74729 527
rect 74813 294 74871 527
rect 74923 289 74957 527
rect 74991 323 75067 493
rect 75111 367 75145 527
rect 75179 323 75255 493
rect 75299 367 75333 527
rect 75367 323 75443 493
rect 75487 367 75521 527
rect 75555 323 75631 493
rect 75675 367 75709 527
rect 75743 323 75819 493
rect 75863 367 75897 527
rect 75931 323 76007 493
rect 76051 367 76085 527
rect 76119 323 76195 493
rect 76239 367 76273 527
rect 76307 323 76383 493
rect 76427 367 76461 527
rect 76495 323 76571 493
rect 76615 367 76649 527
rect 76683 323 76759 493
rect 76803 367 76837 527
rect 76871 323 76947 493
rect 76991 367 77025 527
rect 77060 323 77115 472
rect 74991 289 75521 323
rect 75555 289 77115 323
rect 77205 294 77263 527
rect 77315 341 77349 493
rect 77400 375 77466 527
rect 77315 307 77459 341
rect 73167 215 73502 255
rect 73548 249 73583 289
rect 73548 215 74133 249
rect 73548 181 73583 215
rect 74182 181 74619 289
rect 75486 255 75521 289
rect 74905 215 75435 255
rect 75486 215 76923 255
rect 75486 181 75521 215
rect 77015 181 77115 289
rect 77297 197 77368 271
rect 77425 265 77459 307
rect 77425 199 77485 265
rect 72715 51 72749 127
rect 72785 17 72859 93
rect 72893 51 72959 152
rect 73065 17 73123 162
rect 73269 147 73583 181
rect 73645 147 74619 181
rect 73159 17 73225 113
rect 73269 51 73303 147
rect 73337 17 73413 113
rect 73457 52 73491 147
rect 73525 17 73601 113
rect 73645 51 73679 147
rect 73713 17 73789 113
rect 73833 51 73867 147
rect 73901 17 73977 113
rect 74021 51 74055 147
rect 74089 17 74165 113
rect 74209 51 74243 147
rect 74277 17 74353 113
rect 74397 51 74431 147
rect 74465 17 74541 113
rect 74585 51 74619 147
rect 74653 17 74729 177
rect 74813 17 74871 162
rect 74923 17 74957 181
rect 74991 147 75521 181
rect 75555 147 77115 181
rect 74991 52 75067 147
rect 75111 17 75145 113
rect 75179 52 75255 147
rect 75299 17 75333 113
rect 75367 52 75443 147
rect 75487 17 75521 113
rect 75555 52 75631 147
rect 75555 51 75615 52
rect 75675 17 75709 113
rect 75743 52 75819 147
rect 75769 51 75803 52
rect 75863 17 75897 113
rect 75931 52 76007 147
rect 75957 51 75991 52
rect 76051 17 76085 113
rect 76119 52 76195 147
rect 76239 17 76273 113
rect 76307 52 76383 147
rect 76427 17 76461 113
rect 76495 52 76571 147
rect 76615 17 76649 113
rect 76683 52 76759 147
rect 76803 17 76837 113
rect 76871 52 76947 147
rect 76991 17 77025 113
rect 77060 73 77115 147
rect 77205 17 77263 162
rect 77425 161 77468 199
rect 77315 127 77468 161
rect 77315 51 77349 127
rect 77402 17 77468 93
rect 77534 51 77619 493
rect 77653 297 77705 527
rect 77757 294 77815 527
rect 77851 331 77917 493
rect 77961 367 78009 527
rect 77851 297 78004 331
rect 77850 215 77926 263
rect 77970 249 78004 297
rect 78055 323 78089 493
rect 78123 367 78199 527
rect 78243 323 78277 493
rect 78055 289 78277 323
rect 78311 297 78387 527
rect 78493 294 78551 527
rect 78655 297 78689 527
rect 78723 331 78799 493
rect 78843 367 78891 527
rect 78723 297 78893 331
rect 77970 215 78080 249
rect 77653 17 77705 185
rect 77970 181 78004 215
rect 78216 181 78277 289
rect 78624 215 78821 263
rect 78859 249 78893 297
rect 78937 323 78971 493
rect 79005 367 79081 527
rect 79125 323 79159 493
rect 79193 367 79269 527
rect 79313 323 79347 493
rect 78937 289 79347 323
rect 79381 297 79457 527
rect 79505 294 79563 527
rect 79599 323 79665 493
rect 79709 367 79743 527
rect 79777 323 79853 493
rect 79897 367 79931 527
rect 79991 323 80025 493
rect 80059 367 80135 527
rect 80179 323 80213 493
rect 80247 367 80323 527
rect 80367 323 80401 493
rect 80435 367 80511 527
rect 80555 323 80589 493
rect 79599 289 79929 323
rect 79991 289 80589 323
rect 80623 297 80699 527
rect 80793 294 80851 527
rect 80903 289 80937 527
rect 80971 289 81047 493
rect 81085 323 81151 493
rect 81195 357 81229 527
rect 81263 323 81339 493
rect 81383 357 81417 527
rect 81451 323 81527 493
rect 81571 367 81605 527
rect 81639 323 81715 493
rect 81759 367 81793 527
rect 81827 323 81903 493
rect 81947 367 81981 527
rect 82015 323 82091 493
rect 82135 367 82169 527
rect 82203 323 82279 493
rect 82323 367 82357 527
rect 82391 323 82467 493
rect 82511 367 82545 527
rect 82579 323 82655 493
rect 82699 367 82733 527
rect 82767 323 82843 493
rect 82887 367 82921 527
rect 82955 323 83031 493
rect 83075 367 83109 527
rect 83143 323 83219 493
rect 83263 367 83297 527
rect 83331 323 83407 493
rect 83451 367 83485 527
rect 81085 289 81417 323
rect 81451 289 81981 323
rect 82015 289 83512 323
rect 83553 294 83611 527
rect 83647 323 83713 432
rect 83757 357 83791 527
rect 83647 289 83794 323
rect 83838 309 83924 493
rect 78859 215 78963 249
rect 78859 181 78893 215
rect 79050 181 79347 289
rect 79608 215 79848 255
rect 79894 249 79929 289
rect 79894 215 80479 249
rect 79894 181 79929 215
rect 80518 181 80589 289
rect 81000 255 81047 289
rect 81383 255 81417 289
rect 81946 255 81981 289
rect 80890 215 80956 255
rect 81000 215 81339 255
rect 81383 215 81895 255
rect 81946 215 83408 255
rect 81000 181 81047 215
rect 81383 181 81417 215
rect 81946 181 81981 215
rect 83452 181 83512 289
rect 83760 265 83794 289
rect 83650 215 83716 255
rect 83760 199 83856 265
rect 83890 255 83924 309
rect 83958 323 84024 493
rect 84068 357 84102 527
rect 84136 323 84212 493
rect 84256 357 84290 527
rect 84324 323 84400 493
rect 84444 367 84478 527
rect 84512 323 84588 493
rect 84632 367 84666 527
rect 84700 323 84776 493
rect 84820 367 84854 527
rect 84888 323 84964 493
rect 85008 367 85042 527
rect 83958 289 84290 323
rect 84324 289 85076 323
rect 85117 294 85175 527
rect 85211 323 85277 493
rect 85321 357 85355 527
rect 85389 323 85465 493
rect 85509 357 85543 527
rect 85577 323 85653 493
rect 85697 367 85731 527
rect 85765 323 85841 493
rect 85885 367 85919 527
rect 85953 323 86029 493
rect 86073 367 86107 527
rect 86141 323 86217 493
rect 86261 367 86295 527
rect 86329 323 86405 493
rect 86449 367 86483 527
rect 86517 323 86593 493
rect 86637 367 86671 527
rect 86705 323 86781 493
rect 86825 367 86859 527
rect 86893 323 86969 493
rect 87013 367 87047 527
rect 87081 323 87157 493
rect 87201 367 87235 527
rect 87269 323 87345 493
rect 87389 367 87423 527
rect 87457 323 87533 493
rect 87577 367 87611 527
rect 85211 289 85543 323
rect 85577 289 86107 323
rect 86141 289 87633 323
rect 87693 294 87751 527
rect 87803 289 87837 527
rect 87871 309 87947 493
rect 84256 255 84290 289
rect 83890 215 84212 255
rect 84256 215 84810 255
rect 83760 181 83794 199
rect 77757 17 77815 162
rect 77867 147 78004 181
rect 78055 147 78277 181
rect 77867 51 77901 147
rect 77937 17 77995 113
rect 78055 51 78089 147
rect 78123 17 78199 113
rect 78243 51 78277 147
rect 78311 17 78387 177
rect 78493 17 78551 162
rect 78723 147 78893 181
rect 78937 147 79347 181
rect 78655 17 78689 113
rect 78723 51 78799 147
rect 78843 17 78877 113
rect 78937 51 78971 147
rect 79005 17 79081 113
rect 79125 51 79159 147
rect 79193 17 79269 113
rect 79313 51 79347 147
rect 79381 17 79457 177
rect 79505 17 79563 162
rect 79615 147 79929 181
rect 79991 147 80589 181
rect 79615 51 79649 147
rect 79683 17 79759 113
rect 79803 52 79837 147
rect 79871 17 79947 113
rect 79991 51 80025 147
rect 80059 17 80135 113
rect 80179 51 80213 147
rect 80247 17 80323 113
rect 80367 51 80401 147
rect 80435 17 80511 113
rect 80555 51 80589 147
rect 80623 17 80699 177
rect 80793 17 80851 162
rect 80903 17 80937 181
rect 80971 52 81047 181
rect 81085 147 81417 181
rect 81451 147 81981 181
rect 82015 147 83512 181
rect 81085 52 81151 147
rect 81195 17 81229 113
rect 81263 52 81339 147
rect 81383 17 81417 113
rect 81451 52 81527 147
rect 81571 17 81605 113
rect 81639 52 81715 147
rect 81759 17 81793 113
rect 81827 52 81903 147
rect 81947 17 81981 113
rect 82015 52 82091 147
rect 82015 51 82075 52
rect 82135 17 82169 113
rect 82203 52 82279 147
rect 82229 51 82263 52
rect 82323 17 82357 113
rect 82391 52 82467 147
rect 82417 51 82451 52
rect 82511 17 82545 113
rect 82579 52 82655 147
rect 82699 17 82733 113
rect 82767 52 82843 147
rect 82887 17 82921 113
rect 82955 52 83031 147
rect 83075 17 83109 113
rect 83143 52 83219 147
rect 83263 17 83297 113
rect 83331 52 83407 147
rect 83451 17 83485 113
rect 83553 17 83611 162
rect 83647 147 83794 181
rect 83890 165 83924 215
rect 84256 181 84290 215
rect 85000 181 85076 289
rect 85509 255 85543 289
rect 86072 255 86107 289
rect 85210 215 85465 255
rect 85509 215 86021 255
rect 86072 215 87534 255
rect 85509 181 85543 215
rect 86072 181 86107 215
rect 87578 181 87633 289
rect 87913 255 87947 309
rect 87985 323 88051 493
rect 88095 357 88129 527
rect 88163 323 88239 493
rect 88283 357 88317 527
rect 88351 323 88427 493
rect 88471 367 88505 527
rect 88539 323 88615 493
rect 88659 367 88693 527
rect 88727 323 88803 493
rect 88847 367 88881 527
rect 88915 323 88991 493
rect 89035 367 89069 527
rect 87985 289 88317 323
rect 88351 289 89129 323
rect 89165 294 89223 527
rect 89257 312 89311 493
rect 89345 375 89495 527
rect 89539 341 89573 493
rect 88283 255 88317 289
rect 87785 215 87869 255
rect 87913 215 88239 255
rect 88283 215 89017 255
rect 87913 181 87947 215
rect 88283 181 88317 215
rect 89051 181 89129 289
rect 83647 52 83713 147
rect 83757 17 83791 113
rect 83838 52 83924 165
rect 83958 147 84290 181
rect 84324 147 85076 181
rect 83958 52 84024 147
rect 84068 17 84102 113
rect 84136 52 84212 147
rect 84256 17 84290 113
rect 84324 52 84400 147
rect 84444 17 84478 113
rect 84512 52 84588 147
rect 84632 17 84666 113
rect 84700 52 84776 147
rect 84820 17 84854 113
rect 84888 52 84964 147
rect 85008 17 85042 113
rect 85117 17 85175 162
rect 85211 147 85543 181
rect 85577 147 86107 181
rect 86141 147 87633 181
rect 85211 52 85277 147
rect 85321 17 85355 113
rect 85389 52 85465 147
rect 85509 17 85543 113
rect 85577 52 85653 147
rect 85697 17 85731 113
rect 85765 52 85841 147
rect 85885 17 85919 113
rect 85953 52 86029 147
rect 86073 17 86107 113
rect 86141 52 86217 147
rect 86141 51 86201 52
rect 86261 17 86295 113
rect 86329 52 86405 147
rect 86355 51 86389 52
rect 86449 17 86483 113
rect 86517 52 86593 147
rect 86543 51 86577 52
rect 86637 17 86671 113
rect 86705 52 86781 147
rect 86825 17 86859 113
rect 86893 52 86969 147
rect 87013 17 87047 113
rect 87081 52 87157 147
rect 87201 17 87235 113
rect 87269 52 87345 147
rect 87389 17 87423 113
rect 87457 52 87533 147
rect 87577 17 87611 113
rect 87693 17 87751 162
rect 87803 17 87837 181
rect 87871 52 87947 181
rect 87985 147 88317 181
rect 88351 147 89129 181
rect 87985 52 88051 147
rect 88095 17 88129 113
rect 88163 52 88239 147
rect 88283 17 88317 113
rect 88351 52 88427 147
rect 88471 17 88505 113
rect 88539 52 88615 147
rect 88659 17 88693 113
rect 88727 52 88803 147
rect 88847 17 88881 113
rect 88915 52 88991 147
rect 89035 17 89069 113
rect 89165 17 89223 162
rect 89257 152 89291 312
rect 89348 307 89573 341
rect 89348 278 89392 307
rect 89625 294 89683 527
rect 89719 365 89778 527
rect 89325 212 89392 278
rect 89348 161 89392 212
rect 89513 197 89589 271
rect 89824 265 89873 493
rect 89918 365 89970 527
rect 90110 526 91505 527
rect 90016 265 90066 492
rect 90110 367 90162 526
rect 90206 347 90258 492
rect 90302 381 90354 526
rect 90398 347 90450 492
rect 90494 381 90546 526
rect 90590 347 90642 492
rect 90686 381 90738 526
rect 90782 347 90834 492
rect 90878 381 90927 526
rect 90971 347 91023 492
rect 91070 381 91119 526
rect 91163 347 91215 492
rect 91262 381 91311 526
rect 91355 347 91407 492
rect 91454 381 91505 526
rect 90206 344 91407 347
rect 91549 344 91607 492
rect 91651 378 91705 527
rect 90206 299 91705 344
rect 89257 51 89309 152
rect 89348 127 89565 161
rect 89345 17 89495 93
rect 89531 51 89565 127
rect 89625 17 89683 162
rect 89717 153 89780 265
rect 89824 215 91408 265
rect 89717 17 89778 119
rect 89824 53 89874 215
rect 89918 17 89970 122
rect 90016 53 90066 215
rect 91452 181 91705 299
rect 91741 294 91799 527
rect 91833 333 91887 487
rect 91921 371 91997 527
rect 92048 406 92085 487
rect 92119 442 92196 527
rect 92048 371 92191 406
rect 91833 299 92079 333
rect 90206 147 91705 181
rect 90110 17 90162 129
rect 90206 56 90258 147
rect 90302 17 90354 113
rect 90398 56 90450 147
rect 90494 17 90546 113
rect 90590 56 90642 147
rect 90686 17 90735 113
rect 90769 56 90834 147
rect 90878 17 90927 113
rect 90971 56 91023 147
rect 91069 17 91119 113
rect 91163 56 91215 147
rect 91261 17 91311 113
rect 91355 56 91407 147
rect 91453 17 91505 113
rect 91549 56 91601 147
rect 91645 17 91705 113
rect 91741 17 91799 162
rect 91833 117 91867 299
rect 91901 149 91983 265
rect 92019 199 92079 299
rect 92113 165 92191 371
rect 92293 294 92351 527
rect 92385 333 92447 493
rect 92491 367 92553 527
rect 92597 401 92649 493
rect 92693 435 92744 527
rect 92789 401 92841 493
rect 92597 367 92841 401
rect 92877 369 92943 527
rect 92385 299 92611 333
rect 92044 131 92191 165
rect 91833 51 91885 117
rect 91937 17 91992 113
rect 92044 51 92085 131
rect 92119 17 92196 97
rect 92293 17 92351 162
rect 92385 117 92419 299
rect 92453 151 92533 265
rect 92567 249 92611 299
rect 92789 330 92841 367
rect 92789 283 92950 330
rect 93029 294 93087 527
rect 93123 305 93182 527
rect 92567 215 92816 249
rect 92850 181 92950 283
rect 93228 265 93278 492
rect 93322 305 93374 527
rect 93418 347 93470 492
rect 93514 381 93566 527
rect 93610 347 93662 492
rect 93706 381 93758 527
rect 93802 347 93854 492
rect 93898 381 93950 527
rect 93994 347 94046 492
rect 94090 381 94149 527
rect 93418 299 94150 347
rect 92578 147 92950 181
rect 92385 51 92445 117
rect 92489 17 92544 113
rect 92578 69 92649 147
rect 92693 17 92744 113
rect 92789 69 92841 147
rect 92885 17 92941 113
rect 93029 17 93087 162
rect 93121 143 93184 265
rect 93228 215 93902 265
rect 93133 17 93182 109
rect 93228 53 93278 215
rect 93936 181 94150 299
rect 94225 294 94283 527
rect 94317 333 94369 527
rect 93418 147 94150 181
rect 93322 17 93374 122
rect 93418 56 93470 147
rect 93514 17 93566 113
rect 93610 56 93662 147
rect 93706 17 93758 113
rect 93802 56 93854 147
rect 93898 17 93950 113
rect 93994 56 94046 147
rect 94090 17 94150 113
rect 94225 17 94283 162
rect 94317 75 94365 265
rect 94403 258 94479 493
rect 94523 333 94579 527
rect 94685 294 94743 527
rect 94788 299 94841 527
rect 94885 333 94936 493
rect 94980 367 95032 527
rect 95077 333 95128 490
rect 95173 367 95224 527
rect 95275 333 95320 493
rect 95364 367 95416 527
rect 95461 333 95512 490
rect 95557 367 95608 527
rect 95653 333 95701 490
rect 95753 367 95804 527
rect 95851 333 95926 490
rect 95978 424 96030 527
rect 95978 367 96029 424
rect 96075 333 96125 490
rect 96171 367 96222 527
rect 96267 333 96317 490
rect 96363 367 96414 527
rect 96459 333 96509 490
rect 96555 367 96606 527
rect 96651 333 96701 490
rect 96747 367 96798 527
rect 96843 333 96891 490
rect 96939 367 96990 527
rect 97035 333 97086 490
rect 97130 367 97182 527
rect 94885 291 97086 333
rect 97261 294 97319 527
rect 97367 326 97418 487
rect 97462 360 97514 527
rect 97558 326 97610 487
rect 97657 360 97708 527
rect 97367 292 97767 326
rect 97813 294 97871 527
rect 97905 360 97974 527
rect 98019 326 98070 487
rect 98114 360 98166 527
rect 98211 326 98262 487
rect 98306 360 98358 527
rect 98402 326 98454 487
rect 98498 360 98575 527
rect 95275 283 96701 291
rect 94403 152 94579 258
rect 94829 179 95231 255
rect 94403 51 94478 152
rect 94523 17 94579 118
rect 94685 17 94743 162
rect 95171 17 95225 122
rect 95275 56 95320 283
rect 95364 17 95417 122
rect 95461 56 95512 283
rect 95556 17 95609 122
rect 95653 56 95701 283
rect 95753 17 95806 122
rect 95851 56 95921 283
rect 95978 17 96031 122
rect 96075 56 96125 283
rect 96170 17 96215 122
rect 96267 56 96317 283
rect 96362 17 96415 122
rect 96459 56 96509 283
rect 96554 17 96607 122
rect 96651 56 96701 283
rect 96746 179 97142 255
rect 97353 213 97603 258
rect 97640 179 97767 292
rect 96746 17 96799 122
rect 97261 17 97319 162
rect 97561 145 97767 179
rect 97909 292 98602 326
rect 98641 294 98699 527
rect 98743 360 98795 527
rect 98839 326 98887 487
rect 98931 360 98983 527
rect 99027 326 99075 487
rect 99119 360 99171 527
rect 99215 326 99265 487
rect 99309 360 99358 527
rect 99402 326 99451 487
rect 99495 360 99556 527
rect 99600 326 99661 487
rect 99705 360 99765 527
rect 99809 326 99857 487
rect 99901 360 99952 527
rect 97909 179 97943 292
rect 97977 213 98470 258
rect 98542 179 98602 292
rect 97448 17 97517 122
rect 97561 56 97606 145
rect 97640 17 97716 111
rect 97813 17 97871 162
rect 97909 145 98602 179
rect 98739 292 99982 326
rect 100021 294 100079 527
rect 100141 525 100429 527
rect 100141 367 100207 525
rect 98739 173 98773 292
rect 98807 207 99829 258
rect 99928 173 99982 292
rect 100125 199 100216 333
rect 98001 17 98070 111
rect 98114 56 98166 145
rect 98210 17 98262 111
rect 98306 56 98357 145
rect 98401 17 98461 111
rect 98641 17 98699 162
rect 98739 139 99982 173
rect 98943 17 99009 105
rect 99053 56 99091 139
rect 99135 17 99201 105
rect 99245 56 99283 139
rect 99327 17 99403 105
rect 99437 56 99475 139
rect 99519 17 99605 105
rect 99649 56 99687 139
rect 99731 17 99817 105
rect 100021 17 100079 162
rect 100253 150 100343 491
rect 100377 291 100429 525
rect 100481 294 100539 527
rect 100575 299 100640 527
rect 100155 17 100219 149
rect 100253 63 100405 150
rect 100481 17 100539 162
rect 100573 149 100641 265
rect 100677 259 100745 493
rect 100793 293 100848 527
rect 100887 259 100953 493
rect 101001 293 101057 527
rect 101125 294 101183 527
rect 101255 382 101321 527
rect 100677 203 100953 259
rect 100677 136 100747 203
rect 100575 17 100641 115
rect 100677 51 100789 136
rect 100891 17 100956 155
rect 101125 17 101183 162
rect 101217 51 101321 348
rect 101355 183 101459 493
rect 101493 294 101551 527
rect 101586 393 101637 493
rect 101671 427 101747 527
rect 101586 359 101746 393
rect 101586 195 101656 325
rect 101355 17 101423 149
rect 101493 17 101551 162
rect 101700 161 101746 359
rect 101586 127 101746 161
rect 101586 69 101637 127
rect 101671 17 101747 93
rect 101791 69 101825 493
rect 101922 435 101956 527
rect 102002 427 102052 493
rect 102105 427 102241 493
rect 102002 401 102036 427
rect 101859 333 101922 401
rect 101983 367 102036 401
rect 101859 123 101949 333
rect 101983 95 102017 367
rect 102070 315 102173 393
rect 102053 153 102105 277
rect 102139 197 102173 315
rect 102207 271 102241 427
rect 102275 407 102309 475
rect 102366 441 102432 527
rect 102476 407 102510 475
rect 102569 435 102653 527
rect 102275 373 102510 407
rect 102697 401 102731 493
rect 102778 425 102969 493
rect 103036 435 103086 527
rect 102599 367 102731 401
rect 102599 339 102633 367
rect 102313 305 102633 339
rect 102797 333 102900 391
rect 102207 237 102565 271
rect 102139 153 102210 197
rect 102254 95 102288 237
rect 102329 153 102497 203
rect 102531 201 102565 237
rect 102599 167 102633 305
rect 101883 17 101949 89
rect 101983 61 102067 95
rect 102107 61 102288 95
rect 102473 17 102539 109
rect 102581 89 102633 167
rect 102689 331 102900 333
rect 102935 349 102969 425
rect 103130 417 103164 475
rect 103200 451 103276 527
rect 103130 383 103290 417
rect 102689 299 102831 331
rect 102935 315 103222 349
rect 102689 141 102723 299
rect 102935 297 102979 315
rect 102757 141 102831 265
rect 102865 263 102979 297
rect 102865 107 102899 263
rect 102959 173 103013 229
rect 102959 139 103035 173
rect 102581 55 102661 89
rect 102715 51 102899 107
rect 102933 17 102967 105
rect 103001 93 103035 139
rect 103069 127 103149 281
rect 103256 259 103290 383
rect 103330 315 103364 527
rect 103226 257 103290 259
rect 103226 215 103382 257
rect 103226 93 103295 215
rect 103001 59 103295 93
rect 103330 17 103364 179
rect 103416 51 103483 493
rect 103517 294 103575 527
rect 103610 393 103661 493
rect 103695 427 103771 527
rect 103610 359 103770 393
rect 103610 195 103680 325
rect 103517 17 103575 162
rect 103724 161 103770 359
rect 103610 127 103770 161
rect 103610 69 103661 127
rect 103695 17 103771 93
rect 103815 69 103849 493
rect 103946 435 103980 527
rect 104026 427 104076 493
rect 104129 427 104265 493
rect 104026 401 104060 427
rect 103883 333 103946 401
rect 104007 367 104060 401
rect 103883 123 103973 333
rect 104007 95 104041 367
rect 104094 315 104197 393
rect 104077 153 104129 277
rect 104163 197 104197 315
rect 104231 271 104265 427
rect 104299 407 104333 475
rect 104390 441 104456 527
rect 104500 407 104534 475
rect 104593 435 104677 527
rect 104299 373 104534 407
rect 104721 401 104755 493
rect 104802 425 104993 493
rect 105060 435 105110 527
rect 104623 367 104755 401
rect 104623 339 104657 367
rect 104337 305 104657 339
rect 104821 333 104924 391
rect 104231 237 104589 271
rect 104163 153 104234 197
rect 104278 95 104312 237
rect 104353 153 104521 203
rect 104555 201 104589 237
rect 104623 167 104657 305
rect 103907 17 103973 89
rect 104007 61 104091 95
rect 104131 61 104312 95
rect 104497 17 104563 109
rect 104605 89 104657 167
rect 104713 331 104924 333
rect 104959 349 104993 425
rect 105154 417 105188 475
rect 105224 451 105300 527
rect 105154 383 105314 417
rect 104713 299 104855 331
rect 104959 315 105246 349
rect 104713 141 104747 299
rect 104959 297 105003 315
rect 104781 141 104855 265
rect 104889 263 105003 297
rect 104889 107 104923 263
rect 104983 173 105037 229
rect 104983 139 105059 173
rect 104605 55 104685 89
rect 104739 51 104923 107
rect 104957 17 104991 105
rect 105025 93 105059 139
rect 105093 127 105173 281
rect 105280 259 105314 383
rect 105354 315 105388 527
rect 105440 325 105498 493
rect 105542 359 105576 527
rect 105440 291 105594 325
rect 105633 294 105691 527
rect 105726 393 105777 493
rect 105811 427 105887 527
rect 105726 359 105886 393
rect 105250 257 105314 259
rect 105250 215 105459 257
rect 105250 93 105319 215
rect 105517 181 105594 291
rect 105726 195 105796 325
rect 105025 59 105319 93
rect 105354 17 105388 179
rect 105422 147 105594 181
rect 105422 51 105498 147
rect 105542 17 105576 111
rect 105633 17 105691 162
rect 105840 161 105886 359
rect 105726 127 105886 161
rect 105726 69 105777 127
rect 105811 17 105887 93
rect 105931 69 105965 493
rect 105999 333 106064 490
rect 106098 435 106148 527
rect 106192 427 106242 493
rect 106295 427 106441 493
rect 106192 401 106226 427
rect 106137 367 106226 401
rect 105999 123 106103 333
rect 106137 95 106171 367
rect 106260 315 106363 393
rect 106215 153 106295 277
rect 106329 197 106363 315
rect 106407 271 106441 427
rect 106475 407 106509 475
rect 106566 441 106632 527
rect 106676 407 106710 475
rect 106769 435 106853 527
rect 106475 373 106710 407
rect 106897 401 106931 493
rect 106978 425 107202 493
rect 107236 435 107286 527
rect 106809 367 106931 401
rect 106809 339 106843 367
rect 106513 305 106843 339
rect 107002 333 107114 391
rect 106407 237 106765 271
rect 106329 153 106410 197
rect 106444 95 106478 237
rect 106543 153 106697 203
rect 106731 201 106765 237
rect 106809 167 106843 305
rect 106037 17 106103 89
rect 106137 61 106246 95
rect 106297 61 106478 95
rect 106673 17 106739 109
rect 106781 89 106843 167
rect 106891 331 107114 333
rect 107158 349 107202 425
rect 107330 417 107364 475
rect 107400 451 107476 527
rect 107330 383 107500 417
rect 106891 299 107046 331
rect 107158 315 107432 349
rect 106891 141 106933 299
rect 107158 297 107202 315
rect 106967 141 107057 265
rect 107101 263 107202 297
rect 107101 107 107135 263
rect 107179 173 107233 229
rect 107269 207 107387 281
rect 107466 259 107500 383
rect 107535 315 107569 527
rect 107621 325 107679 493
rect 107723 359 107757 527
rect 107809 325 107859 493
rect 107911 359 107945 527
rect 107621 291 107989 325
rect 108025 294 108083 527
rect 108135 393 108169 493
rect 108203 427 108279 527
rect 108135 359 108278 393
rect 107179 139 107295 173
rect 106781 55 106861 89
rect 106915 51 107135 107
rect 107179 17 107227 105
rect 107261 93 107295 139
rect 107339 127 107387 207
rect 107431 257 107500 259
rect 107431 215 107867 257
rect 107431 164 107496 215
rect 107907 181 107989 291
rect 108118 195 108188 325
rect 107431 93 107495 164
rect 107261 59 107495 93
rect 107535 17 107569 179
rect 107603 147 107989 181
rect 107603 51 107679 147
rect 107723 17 107757 111
rect 107791 51 107867 147
rect 107911 17 107945 111
rect 108025 17 108083 162
rect 108232 161 108278 359
rect 108135 127 108278 161
rect 108135 69 108169 127
rect 108203 17 108279 93
rect 108323 69 108368 493
rect 108411 427 108477 527
rect 108521 393 108555 493
rect 108602 450 108788 484
rect 108846 451 108922 527
rect 108406 359 108555 393
rect 108406 165 108440 359
rect 108474 201 108566 325
rect 108600 315 108720 391
rect 108406 127 108555 165
rect 108600 141 108654 315
rect 108754 281 108788 450
rect 108968 417 109002 475
rect 109036 451 109112 527
rect 109212 433 109358 483
rect 109394 451 109488 527
rect 109314 417 109358 433
rect 109528 417 109576 475
rect 108822 367 109122 417
rect 108822 315 108882 367
rect 108994 281 109054 313
rect 108754 247 109054 281
rect 108754 246 108848 247
rect 108690 129 108770 203
rect 108411 17 108477 93
rect 108521 61 108555 127
rect 108804 93 108848 246
rect 109088 213 109122 367
rect 108882 147 109002 213
rect 109058 145 109122 213
rect 109166 331 109280 393
rect 109314 383 109576 417
rect 109642 389 109708 527
rect 109166 179 109200 331
rect 109244 213 109280 295
rect 109314 281 109358 383
rect 109742 353 109776 475
rect 109830 383 109896 485
rect 109742 349 109810 353
rect 109392 315 109810 349
rect 109314 247 109734 281
rect 109374 179 109450 203
rect 109166 145 109450 179
rect 108625 53 108848 93
rect 108882 17 108974 105
rect 109058 59 109092 145
rect 109128 17 109206 109
rect 109484 95 109518 247
rect 109658 235 109734 247
rect 109552 201 109628 213
rect 109552 147 109656 201
rect 109768 136 109810 315
rect 109338 61 109518 95
rect 109564 17 109706 113
rect 109742 70 109810 136
rect 109846 265 109896 383
rect 109930 367 110014 527
rect 110048 331 110105 465
rect 109846 199 110016 265
rect 109846 69 109896 199
rect 110060 159 110105 331
rect 110141 294 110199 527
rect 110251 393 110285 493
rect 110319 427 110395 527
rect 110251 359 110394 393
rect 110234 195 110304 325
rect 109930 17 110017 109
rect 110051 53 110105 159
rect 110141 17 110199 162
rect 110348 161 110394 359
rect 110251 127 110394 161
rect 110251 69 110285 127
rect 110319 17 110395 93
rect 110439 69 110484 493
rect 110527 427 110593 527
rect 110637 393 110671 493
rect 110718 450 110904 484
rect 110962 451 111038 527
rect 110522 359 110671 393
rect 110522 165 110556 359
rect 110590 201 110682 325
rect 110716 315 110836 391
rect 110522 127 110671 165
rect 110716 141 110770 315
rect 110870 281 110904 450
rect 111084 417 111118 475
rect 111152 451 111228 527
rect 111328 433 111474 483
rect 111510 451 111604 527
rect 111430 417 111474 433
rect 111644 417 111692 475
rect 110938 367 111238 417
rect 110938 315 110998 367
rect 111110 281 111170 313
rect 110870 247 111170 281
rect 110870 246 110964 247
rect 110806 129 110886 203
rect 110527 17 110593 93
rect 110637 61 110671 127
rect 110920 93 110964 246
rect 111204 213 111238 367
rect 110998 147 111118 213
rect 111174 145 111238 213
rect 111282 331 111396 393
rect 111430 383 111692 417
rect 111758 389 111824 527
rect 111282 179 111316 331
rect 111360 213 111396 295
rect 111430 281 111474 383
rect 111858 353 111892 475
rect 111946 383 112012 485
rect 111858 349 111926 353
rect 111508 315 111926 349
rect 111430 247 111850 281
rect 111490 179 111566 203
rect 111282 145 111566 179
rect 110741 53 110964 93
rect 110998 17 111090 105
rect 111174 59 111208 145
rect 111244 17 111322 109
rect 111600 95 111634 247
rect 111774 235 111850 247
rect 111668 201 111744 213
rect 111668 147 111772 201
rect 111884 136 111926 315
rect 111454 61 111634 95
rect 111680 17 111822 113
rect 111858 70 111926 136
rect 111962 265 112012 383
rect 112056 299 112090 527
rect 112124 323 112219 492
rect 112253 357 112306 527
rect 112124 299 112313 323
rect 111962 199 112132 265
rect 111962 69 111996 199
rect 112166 165 112313 299
rect 112349 294 112407 527
rect 112459 393 112493 493
rect 112527 427 112603 527
rect 112459 359 112602 393
rect 112442 195 112512 325
rect 112030 17 112106 165
rect 112153 149 112313 165
rect 112153 53 112219 149
rect 112253 17 112306 115
rect 112349 17 112407 162
rect 112556 161 112602 359
rect 112459 127 112602 161
rect 112459 69 112493 127
rect 112527 17 112603 93
rect 112647 69 112692 493
rect 112735 427 112801 527
rect 112845 393 112879 493
rect 112926 450 113112 484
rect 113170 451 113246 527
rect 112730 359 112879 393
rect 112730 165 112764 359
rect 112798 201 112890 325
rect 112924 315 113044 391
rect 112730 127 112879 165
rect 112924 141 112978 315
rect 113078 281 113112 450
rect 113292 417 113326 475
rect 113360 451 113436 527
rect 113536 433 113682 483
rect 113718 451 113812 527
rect 113638 417 113682 433
rect 113852 417 113900 475
rect 113146 367 113446 417
rect 113146 315 113206 367
rect 113318 281 113378 313
rect 113078 247 113378 281
rect 113078 246 113172 247
rect 113014 129 113094 203
rect 112735 17 112801 93
rect 112845 61 112879 127
rect 113128 93 113172 246
rect 113412 213 113446 367
rect 113206 147 113326 213
rect 113382 145 113446 213
rect 113490 331 113604 393
rect 113638 383 113900 417
rect 113966 389 114032 527
rect 113490 179 113524 331
rect 113568 213 113604 295
rect 113638 281 113682 383
rect 114066 353 114100 475
rect 114154 383 114220 485
rect 114066 349 114134 353
rect 113716 315 114134 349
rect 113638 247 114058 281
rect 113698 179 113774 203
rect 113490 145 113774 179
rect 112949 53 113172 93
rect 113206 17 113298 105
rect 113382 59 113416 145
rect 113452 17 113530 109
rect 113808 95 113842 247
rect 113982 235 114058 247
rect 113876 201 113952 213
rect 113876 147 113980 201
rect 114092 136 114134 315
rect 113662 61 113842 95
rect 113888 17 114030 113
rect 114066 70 114134 136
rect 114170 255 114220 383
rect 114262 367 114333 527
rect 114369 328 114423 493
rect 114457 362 114508 527
rect 114557 328 114591 493
rect 114635 362 114711 527
rect 114745 328 114796 493
rect 114369 294 114796 328
rect 114833 294 114891 527
rect 114943 393 114977 493
rect 115011 427 115087 527
rect 114943 359 115074 393
rect 114170 211 114712 255
rect 114170 69 114220 211
rect 114746 177 114796 294
rect 114925 197 114974 325
rect 115040 280 115074 359
rect 115131 337 115176 493
rect 115040 214 115086 280
rect 114369 143 114796 177
rect 114262 17 114319 109
rect 114369 53 114429 143
rect 114463 17 114523 109
rect 114557 53 114591 143
rect 114635 17 114711 109
rect 114745 53 114796 143
rect 114833 17 114891 162
rect 115040 161 115074 214
rect 114943 127 115074 161
rect 114943 69 114977 127
rect 115011 17 115087 93
rect 115131 69 115165 337
rect 115219 333 115285 483
rect 115329 367 115392 527
rect 115512 451 115678 485
rect 115219 299 115366 333
rect 115201 191 115286 265
rect 115332 219 115366 299
rect 115442 271 115499 401
rect 115542 283 115610 399
rect 115332 157 115416 219
rect 115542 207 115576 283
rect 115235 153 115416 157
rect 115235 123 115366 153
rect 115485 141 115576 207
rect 115644 265 115678 451
rect 115718 427 115778 527
rect 115822 373 115866 487
rect 115722 307 115866 373
rect 115832 265 115866 307
rect 115912 299 115966 527
rect 115644 199 115794 265
rect 115832 199 115992 265
rect 115235 69 115269 123
rect 115644 107 115678 199
rect 115832 165 115866 199
rect 115303 17 115379 89
rect 115509 73 115678 107
rect 115712 17 115768 165
rect 115822 83 115866 165
rect 115912 17 115966 165
rect 116026 83 116083 491
rect 116121 294 116179 527
rect 116231 393 116265 493
rect 116299 427 116375 527
rect 116231 359 116362 393
rect 116213 197 116262 325
rect 116328 280 116362 359
rect 116419 337 116464 493
rect 116328 214 116374 280
rect 116121 17 116179 162
rect 116328 161 116362 214
rect 116231 127 116362 161
rect 116231 69 116265 127
rect 116299 17 116375 93
rect 116419 69 116453 337
rect 116507 333 116573 483
rect 116617 367 116680 527
rect 116825 451 116985 485
rect 116507 299 116654 333
rect 116489 191 116574 265
rect 116620 219 116654 299
rect 116730 271 116787 401
rect 116830 283 116898 399
rect 116620 157 116704 219
rect 116830 207 116864 283
rect 116951 265 116985 451
rect 117029 427 117089 527
rect 117133 373 117177 487
rect 117033 307 117177 373
rect 117143 265 117177 307
rect 117223 299 117277 527
rect 117321 299 117378 491
rect 117415 351 117465 527
rect 117344 265 117378 299
rect 117501 294 117559 527
rect 117611 393 117645 493
rect 117679 427 117755 527
rect 117611 359 117754 393
rect 116951 233 117105 265
rect 116523 153 116704 157
rect 116523 123 116654 153
rect 116779 141 116864 207
rect 116921 199 117105 233
rect 117143 199 117303 265
rect 117344 199 117465 265
rect 116523 69 116557 123
rect 116921 107 116955 199
rect 117143 165 117177 199
rect 117344 165 117378 199
rect 117593 197 117642 325
rect 116591 17 116667 89
rect 116813 73 116955 107
rect 117003 17 117079 165
rect 117133 83 117177 165
rect 117223 17 117277 165
rect 117321 83 117378 165
rect 117415 17 117467 110
rect 117501 17 117559 162
rect 117708 161 117754 359
rect 117611 127 117754 161
rect 117611 69 117645 127
rect 117679 17 117755 93
rect 117799 69 117833 493
rect 117887 333 117953 483
rect 117997 367 118060 527
rect 118181 451 118366 485
rect 117887 299 118034 333
rect 117871 191 117954 265
rect 118000 219 118034 299
rect 118110 271 118167 401
rect 118211 283 118289 399
rect 118000 157 118084 219
rect 118211 207 118245 283
rect 117903 153 118084 157
rect 117903 123 118034 153
rect 118159 141 118245 207
rect 118332 265 118366 451
rect 118400 427 118434 527
rect 118504 373 118548 487
rect 118404 307 118548 373
rect 118510 265 118548 307
rect 118594 299 118651 527
rect 118695 299 118755 491
rect 118789 299 118839 527
rect 118718 265 118755 299
rect 118883 265 118937 491
rect 118977 299 119011 527
rect 119065 294 119123 527
rect 119157 401 119216 493
rect 119260 435 119303 527
rect 119337 435 119424 493
rect 119157 357 119329 401
rect 118332 199 118476 265
rect 118510 199 118674 265
rect 118718 199 119023 265
rect 119157 211 119261 323
rect 119295 265 119329 357
rect 119295 199 119356 265
rect 119390 255 119424 435
rect 119463 349 119508 486
rect 119569 383 119643 527
rect 119463 315 119662 349
rect 119620 265 119662 315
rect 119712 299 119764 493
rect 119390 215 119540 255
rect 117903 69 117937 123
rect 118332 107 118366 199
rect 117971 17 118047 89
rect 118194 73 118366 107
rect 118400 17 118434 122
rect 118510 83 118548 199
rect 118718 149 118755 199
rect 118594 17 118651 143
rect 118695 83 118755 149
rect 118789 17 118839 165
rect 118883 77 118937 199
rect 119295 177 119329 199
rect 118977 17 119011 143
rect 119065 17 119123 162
rect 119159 143 119329 177
rect 119159 51 119216 143
rect 119390 109 119424 215
rect 119620 199 119686 265
rect 119620 181 119662 199
rect 119260 17 119303 109
rect 119337 51 119424 109
rect 119463 147 119662 181
rect 119730 165 119764 299
rect 119801 294 119859 527
rect 119893 401 119952 493
rect 119996 435 120039 527
rect 120073 435 120160 493
rect 119893 357 120065 401
rect 119893 211 119997 323
rect 120031 265 120065 357
rect 120031 199 120092 265
rect 120126 255 120160 435
rect 120199 349 120244 416
rect 120305 383 120379 527
rect 120199 315 120398 349
rect 120356 265 120398 315
rect 120432 299 120498 493
rect 120126 215 120295 255
rect 120031 177 120065 199
rect 119463 51 119508 147
rect 119569 17 119651 113
rect 119706 51 119764 165
rect 119801 17 119859 162
rect 119895 143 120065 177
rect 119895 51 119952 143
rect 120126 109 120160 215
rect 120356 199 120414 265
rect 120356 181 120398 199
rect 119996 17 120039 109
rect 120073 51 120160 109
rect 120199 147 120398 181
rect 120448 165 120498 299
rect 120537 294 120595 527
rect 120629 401 120688 493
rect 120733 435 120783 527
rect 120873 435 120960 493
rect 120629 357 120801 401
rect 120629 211 120733 323
rect 120767 265 120801 357
rect 120767 199 120892 265
rect 120926 255 120960 435
rect 120994 349 121038 416
rect 121150 383 121216 527
rect 120994 315 121216 349
rect 121174 265 121216 315
rect 121250 299 121331 493
rect 120926 215 121107 255
rect 120767 177 120801 199
rect 120199 102 120244 147
rect 120305 17 120387 113
rect 120432 51 120498 165
rect 120537 17 120595 162
rect 120631 143 120801 177
rect 120631 51 120688 143
rect 120926 109 120960 215
rect 121174 199 121243 265
rect 121174 181 121216 199
rect 120732 17 120775 109
rect 120873 51 120960 109
rect 120994 147 121216 181
rect 121277 165 121331 299
rect 121365 294 121423 527
rect 121457 401 121509 493
rect 121543 435 121618 527
rect 121663 401 121714 492
rect 121748 435 121820 527
rect 121457 357 121598 401
rect 121663 360 121821 401
rect 121457 199 121511 323
rect 121545 165 121598 357
rect 121632 215 121698 326
rect 121732 265 121821 360
rect 121865 299 122157 493
rect 121732 215 121989 265
rect 120994 102 121040 147
rect 121150 17 121216 113
rect 121250 51 121331 165
rect 121365 17 121423 162
rect 121457 123 121687 165
rect 121732 127 121798 215
rect 122023 199 122069 265
rect 122023 181 122057 199
rect 121832 147 122057 181
rect 122103 165 122157 299
rect 122193 294 122251 527
rect 121457 56 121509 123
rect 121653 93 121687 123
rect 121832 93 121875 147
rect 121543 17 121619 89
rect 121653 51 121875 93
rect 121909 17 122057 113
rect 122091 51 122157 165
rect 122193 17 122251 162
rect 122285 56 122337 493
rect 122371 369 122468 527
rect 122512 353 122570 493
rect 122608 421 122650 493
rect 122684 455 122760 527
rect 122804 459 123153 493
rect 122804 421 122943 459
rect 122608 387 122943 421
rect 122987 353 123067 425
rect 123101 359 123153 459
rect 122371 153 122423 335
rect 122512 289 122631 353
rect 122665 325 123067 353
rect 122665 289 123160 325
rect 123205 294 123263 527
rect 123297 353 123349 493
rect 123383 369 123476 527
rect 123520 353 123571 493
rect 123613 421 123662 493
rect 123696 455 123772 527
rect 123816 421 123850 493
rect 123894 455 123960 527
rect 124004 421 124537 493
rect 123613 387 124537 421
rect 123679 379 124537 387
rect 122578 255 122631 289
rect 122457 153 122528 255
rect 122578 205 122911 255
rect 122967 205 123059 255
rect 122578 119 122634 205
rect 123114 171 123160 289
rect 122371 17 122448 119
rect 122482 51 122634 119
rect 122668 131 122943 171
rect 122668 51 122732 131
rect 122766 17 122842 97
rect 122886 93 122943 131
rect 122977 127 123160 171
rect 122886 55 123148 93
rect 123205 17 123263 162
rect 123297 133 123344 353
rect 123378 153 123446 335
rect 123520 319 123645 353
rect 123480 153 123556 285
rect 123590 255 123645 319
rect 123679 289 124547 345
rect 124585 294 124643 527
rect 124677 357 124749 527
rect 124793 323 124830 493
rect 124864 373 124941 527
rect 123590 205 124112 255
rect 124146 205 124467 255
rect 123297 56 123349 133
rect 123590 119 123645 205
rect 124501 171 124547 289
rect 124677 199 124746 323
rect 123383 17 123476 119
rect 123520 51 123645 119
rect 123679 131 124145 171
rect 123679 51 123745 131
rect 123779 17 123855 97
rect 123899 55 123933 131
rect 123967 17 124043 97
rect 124087 89 124145 131
rect 124179 123 124547 171
rect 124087 51 124537 89
rect 124585 17 124643 162
rect 124677 17 124749 165
rect 124790 56 124830 323
rect 124864 265 124941 339
rect 124975 299 125055 493
rect 125089 413 125139 493
rect 125173 447 125259 527
rect 125303 413 125337 493
rect 125381 447 125467 527
rect 125511 413 125545 493
rect 125589 447 125675 527
rect 125719 413 125753 493
rect 125797 447 125883 527
rect 125927 413 126845 493
rect 125089 379 126845 413
rect 124864 199 124966 265
rect 125010 255 125055 299
rect 125089 289 126845 345
rect 126885 294 126943 527
rect 126977 413 127034 493
rect 127068 447 127144 527
rect 126977 379 127144 413
rect 125010 205 126035 255
rect 126085 205 126751 255
rect 124864 124 124941 199
rect 125010 165 125087 205
rect 126795 171 126845 289
rect 126977 191 127062 345
rect 127107 323 127144 379
rect 127240 357 127495 493
rect 127107 288 127280 323
rect 124864 17 124941 89
rect 124975 51 125087 165
rect 125121 131 126071 171
rect 125121 51 125197 131
rect 125231 17 125317 97
rect 125361 55 125405 131
rect 125439 17 125525 97
rect 125569 51 125613 131
rect 125647 17 125733 97
rect 125777 55 125821 131
rect 125855 17 125941 97
rect 125985 89 126071 131
rect 126105 123 126845 171
rect 125985 51 126845 89
rect 126885 17 126943 162
rect 127184 161 127280 288
rect 127107 157 127280 161
rect 126977 123 127280 157
rect 126977 51 127034 123
rect 127354 119 127402 357
rect 127446 153 127495 323
rect 127529 294 127587 527
rect 127621 345 127673 493
rect 127707 379 127793 527
rect 127838 417 127872 493
rect 127906 451 128099 527
rect 128143 417 128177 493
rect 127838 373 128177 417
rect 127621 311 127793 345
rect 127621 199 127669 277
rect 127703 255 127793 311
rect 127838 289 127989 373
rect 128211 339 128311 493
rect 128033 289 128311 339
rect 128357 294 128415 527
rect 128449 333 128501 493
rect 128535 367 128611 527
rect 128645 333 128700 493
rect 128734 367 128810 527
rect 128854 333 128888 493
rect 128922 367 129010 527
rect 129054 459 129472 493
rect 129054 333 129096 459
rect 128449 299 128611 333
rect 128645 299 129096 333
rect 127703 199 128040 255
rect 127703 165 127782 199
rect 127068 17 127278 89
rect 127354 51 127495 119
rect 127529 17 127587 162
rect 127621 131 127782 165
rect 127817 131 128058 165
rect 127621 51 127673 131
rect 127707 17 127783 97
rect 127817 51 127880 131
rect 127924 17 127990 97
rect 128024 85 128058 131
rect 128093 119 128167 289
rect 128535 265 128611 299
rect 129130 296 129206 415
rect 129250 330 129284 459
rect 129318 296 129394 415
rect 129438 330 129472 459
rect 128201 215 128311 255
rect 128449 199 128501 265
rect 128535 199 129096 265
rect 128535 165 128611 199
rect 128237 85 128291 155
rect 128024 51 128291 85
rect 128357 17 128415 162
rect 128449 131 128611 165
rect 128645 131 129091 165
rect 128449 51 128501 131
rect 128535 17 128611 97
rect 128645 51 128709 131
rect 128753 17 128819 97
rect 128863 51 128897 131
rect 128941 17 129007 97
rect 129057 90 129091 131
rect 129130 124 129394 296
rect 129553 294 129611 527
rect 129646 333 129697 493
rect 129731 367 129807 527
rect 129841 333 129896 493
rect 129930 367 130006 527
rect 130050 333 130084 493
rect 130118 367 130194 527
rect 130238 333 130272 493
rect 130306 367 130382 527
rect 130426 333 130460 493
rect 130494 367 130574 527
rect 130618 459 131447 493
rect 130618 333 130668 459
rect 129646 299 129807 333
rect 129841 299 130668 333
rect 130702 325 130778 425
rect 130822 359 130856 459
rect 130890 325 130966 425
rect 131010 359 131044 459
rect 131078 325 131154 425
rect 131198 359 131232 459
rect 131266 325 131342 425
rect 131386 359 131447 459
rect 129731 265 129807 299
rect 130702 291 131447 325
rect 131485 294 131543 527
rect 131577 413 131629 493
rect 131663 447 131908 527
rect 131956 425 132085 493
rect 131577 379 131898 413
rect 129428 124 129515 265
rect 129646 199 129697 265
rect 129731 199 130623 265
rect 130657 199 131358 257
rect 129731 165 129807 199
rect 131402 165 131447 291
rect 131577 199 131679 345
rect 131713 165 131898 379
rect 129057 51 129519 90
rect 129553 17 129611 162
rect 129646 131 129807 165
rect 129841 131 130668 165
rect 129646 51 129697 131
rect 129731 17 129807 97
rect 129841 51 129905 131
rect 129949 17 130015 97
rect 130059 51 130093 131
rect 130137 17 130203 97
rect 130247 51 130281 131
rect 130325 17 130391 97
rect 130435 51 130469 131
rect 130513 17 130581 97
rect 130625 90 130668 131
rect 130702 124 131447 165
rect 130625 51 131447 90
rect 131485 17 131543 162
rect 131577 131 131898 165
rect 131956 161 131991 425
rect 132037 195 132085 391
rect 132129 294 132187 527
rect 132221 391 132273 493
rect 132307 425 132389 527
rect 132221 357 132389 391
rect 132221 199 132270 323
rect 132304 265 132389 357
rect 132433 345 132481 493
rect 132525 379 132591 527
rect 132641 459 132910 493
rect 132641 345 132675 459
rect 132433 311 132675 345
rect 132304 199 132625 265
rect 132304 165 132389 199
rect 131577 51 131629 131
rect 131663 17 131860 97
rect 131956 51 132085 161
rect 132129 17 132187 162
rect 132221 131 132389 165
rect 132433 131 132699 165
rect 132221 51 132273 131
rect 132307 17 132389 97
rect 132433 51 132472 131
rect 132506 17 132580 97
rect 132632 85 132699 131
rect 132733 119 132819 425
rect 132853 357 132910 459
rect 132853 153 132911 323
rect 132957 294 133015 527
rect 133049 391 133101 493
rect 133135 425 133217 527
rect 133049 357 133217 391
rect 133049 199 133098 323
rect 133132 265 133217 357
rect 133267 345 133309 493
rect 133353 379 133419 527
rect 133463 345 133497 493
rect 133541 379 133613 527
rect 133657 459 134114 493
rect 133657 345 133691 459
rect 133267 311 133691 345
rect 133730 323 133806 425
rect 133850 357 133884 459
rect 133918 323 133994 425
rect 133730 289 133994 323
rect 134038 289 134114 459
rect 134153 294 134211 527
rect 134245 391 134297 493
rect 134331 425 134413 527
rect 134245 357 134413 391
rect 133132 199 133696 265
rect 133132 165 133181 199
rect 133730 170 133838 289
rect 133874 204 134114 255
rect 134245 199 134294 323
rect 134328 265 134413 357
rect 134463 345 134505 493
rect 134549 379 134615 527
rect 134659 345 134693 493
rect 134737 379 134803 527
rect 134847 345 134881 493
rect 134925 379 134991 527
rect 135035 345 135069 493
rect 135113 379 135179 527
rect 135223 459 136047 493
rect 135223 345 135268 459
rect 134463 311 135268 345
rect 135302 323 135378 425
rect 135422 357 135456 459
rect 135490 323 135566 425
rect 135610 357 135644 459
rect 135678 323 135754 425
rect 135798 357 135832 459
rect 135866 323 135942 425
rect 135302 289 135942 323
rect 135986 289 136047 459
rect 136085 294 136143 527
rect 136228 299 136270 527
rect 136314 297 136417 493
rect 134328 199 135268 265
rect 132853 85 132910 119
rect 132632 51 132910 85
rect 132957 17 133015 162
rect 133049 131 133181 165
rect 133259 131 133696 165
rect 133049 51 133101 131
rect 133135 17 133211 97
rect 133259 51 133293 131
rect 133327 17 133403 97
rect 133447 51 133481 131
rect 133515 17 133593 97
rect 133629 93 133696 131
rect 133730 127 134114 170
rect 134328 165 134377 199
rect 135302 170 135388 289
rect 135432 204 136038 255
rect 136179 215 136290 263
rect 133629 51 134114 93
rect 134153 17 134211 162
rect 134245 131 134377 165
rect 134455 131 135268 165
rect 134245 51 134297 131
rect 134331 17 134407 97
rect 134455 51 134489 131
rect 134523 17 134599 97
rect 134643 51 134677 131
rect 134711 17 134787 97
rect 134831 51 134865 131
rect 134899 17 134975 97
rect 135019 51 135053 131
rect 135087 17 135165 97
rect 135199 93 135268 131
rect 135302 127 136047 170
rect 135199 51 136047 93
rect 136085 17 136143 162
rect 136224 17 136270 181
rect 136359 177 136417 297
rect 136453 294 136511 527
rect 136579 367 136630 527
rect 136664 333 136740 493
rect 136784 367 136818 527
rect 136852 333 136928 493
rect 136972 367 137006 527
rect 137040 333 137116 493
rect 137160 367 137194 527
rect 137228 333 137304 493
rect 137348 367 137382 527
rect 137416 333 137492 493
rect 137536 367 137570 527
rect 137604 333 137680 493
rect 137723 367 137774 527
rect 136545 299 137792 333
rect 136314 51 136417 177
rect 136545 181 136630 299
rect 136664 215 137688 265
rect 137722 181 137792 299
rect 137833 294 137891 527
rect 137948 297 137990 527
rect 138024 333 138100 493
rect 138144 367 138178 527
rect 138212 333 138288 493
rect 138332 367 138366 527
rect 138400 333 138476 493
rect 138520 367 138554 527
rect 138588 333 138664 493
rect 138708 367 138742 527
rect 138776 333 138852 493
rect 138896 367 138930 527
rect 138964 333 139040 493
rect 139084 367 139118 527
rect 139152 333 139228 493
rect 139272 367 139306 527
rect 139340 333 139416 493
rect 139460 367 139502 527
rect 138024 299 139416 333
rect 137925 215 139133 263
rect 139311 181 139416 299
rect 139581 294 139639 527
rect 139681 299 139727 527
rect 139761 297 139837 493
rect 139881 299 139923 527
rect 139677 215 139743 265
rect 136453 17 136511 162
rect 136545 143 137792 181
rect 136579 17 136630 109
rect 136664 51 136740 143
rect 136784 17 136818 109
rect 136852 51 136928 143
rect 136972 17 137006 109
rect 137040 51 137116 143
rect 137160 17 137194 109
rect 137228 51 137304 143
rect 137348 17 137382 109
rect 137416 51 137492 143
rect 137536 17 137570 109
rect 137604 51 137680 143
rect 137720 17 137774 109
rect 137833 17 137891 162
rect 137944 17 137990 177
rect 138024 143 139416 181
rect 138024 51 138100 143
rect 138144 17 138178 109
rect 138212 51 138288 143
rect 138332 17 138366 109
rect 138400 51 138476 143
rect 138520 17 138554 109
rect 138588 51 138664 143
rect 138708 17 138742 109
rect 138776 51 138852 143
rect 138896 17 138930 109
rect 138964 51 139040 143
rect 139084 17 139118 109
rect 139152 51 139228 143
rect 139272 17 139306 109
rect 139340 51 139416 143
rect 139460 17 139502 177
rect 139581 17 139639 162
rect 139681 17 139727 181
rect 139777 177 139837 297
rect 140041 294 140099 527
rect 140142 299 140195 527
rect 140229 333 140305 493
rect 140349 367 140383 527
rect 140417 337 140493 493
rect 140537 435 140579 527
rect 140417 333 140649 337
rect 140229 299 140649 333
rect 140137 215 140493 265
rect 140595 181 140649 299
rect 140685 294 140743 527
rect 140795 299 140829 527
rect 140863 333 140939 493
rect 140983 367 141017 527
rect 141051 333 141127 493
rect 141171 367 141205 527
rect 141239 337 141315 493
rect 141359 435 141393 527
rect 141239 333 141413 337
rect 140863 299 141413 333
rect 140817 215 141299 265
rect 141333 181 141413 299
rect 141513 294 141571 527
rect 141639 367 141690 527
rect 141724 333 141800 493
rect 141844 367 141878 527
rect 141912 333 141988 493
rect 142032 367 142066 527
rect 142100 333 142176 493
rect 142220 367 142254 527
rect 142288 333 142364 493
rect 142408 367 142468 527
rect 141605 299 142489 333
rect 139761 51 139837 177
rect 139881 17 139923 181
rect 140041 17 140099 162
rect 140229 145 140649 181
rect 140142 17 140195 109
rect 140229 51 140305 145
rect 140349 17 140383 109
rect 140417 51 140493 145
rect 140537 17 140587 110
rect 140685 17 140743 162
rect 140889 145 141413 181
rect 141605 181 141674 299
rect 141724 215 142365 265
rect 142425 181 142489 299
rect 142525 294 142583 527
rect 142618 299 142685 493
rect 142729 299 142763 527
rect 142814 459 143283 493
rect 140786 17 140839 109
rect 140889 51 140923 145
rect 140983 17 141017 109
rect 141077 51 141111 145
rect 141171 17 141205 109
rect 141265 51 141299 145
rect 141333 17 141393 110
rect 141513 17 141571 162
rect 141605 143 142489 181
rect 141639 17 141690 109
rect 141724 51 141800 143
rect 141844 17 141878 109
rect 141912 51 141988 143
rect 142032 17 142066 109
rect 142100 51 142176 143
rect 142220 17 142254 109
rect 142288 51 142364 143
rect 142408 17 142469 109
rect 142525 17 142583 162
rect 142618 51 142669 299
rect 142814 265 142854 459
rect 142703 165 142737 265
rect 142799 199 142854 265
rect 142888 391 143150 425
rect 142888 165 142922 391
rect 142703 131 142922 165
rect 142956 323 143215 357
rect 142956 163 142990 323
rect 142887 124 142922 131
rect 142703 17 142779 97
rect 142887 51 142991 124
rect 143058 51 143123 283
rect 143171 51 143215 323
rect 143249 326 143283 459
rect 143317 375 143351 527
rect 143408 375 143500 457
rect 143249 288 143409 326
rect 143443 213 143500 375
rect 143537 294 143595 527
rect 143630 299 143681 527
rect 143715 319 143787 493
rect 143835 435 143869 527
rect 143903 451 144184 485
rect 143903 401 143937 451
rect 144304 435 144348 527
rect 144382 401 144459 493
rect 143831 367 143937 401
rect 143971 367 144459 401
rect 143257 179 143500 213
rect 143250 17 143353 124
rect 143407 58 143456 179
rect 143537 17 143595 162
rect 143630 17 143681 177
rect 143715 51 143772 319
rect 143831 265 143865 367
rect 143971 333 144005 367
rect 143806 199 143865 265
rect 143899 299 144005 333
rect 143899 199 143943 299
rect 144039 282 144227 325
rect 144037 265 144227 282
rect 143996 256 144227 265
rect 143831 161 143865 199
rect 143831 127 143953 161
rect 143996 153 144071 256
rect 144118 155 144227 221
rect 143919 119 143953 127
rect 143809 17 143885 93
rect 143919 53 144062 119
rect 144186 84 144227 155
rect 144283 151 144321 325
rect 144309 17 144349 117
rect 144409 51 144459 367
rect 144549 294 144607 527
rect 144642 333 144693 493
rect 144727 367 144798 527
rect 144832 455 145218 489
rect 144832 387 144912 455
rect 145279 421 145313 493
rect 145347 451 145423 527
rect 144950 387 145313 421
rect 144642 299 144860 333
rect 144549 17 144607 162
rect 144642 125 144676 299
rect 144710 199 144782 265
rect 144816 199 144860 299
rect 144914 199 144983 323
rect 145050 319 145421 353
rect 145017 199 145141 265
rect 145200 199 145343 265
rect 145387 249 145421 319
rect 145467 349 145501 493
rect 145535 383 145611 527
rect 145655 349 145689 493
rect 145723 383 145799 527
rect 145467 315 145800 349
rect 145387 215 145710 249
rect 144748 161 144782 199
rect 145200 161 145234 199
rect 145387 165 145421 215
rect 144748 127 145234 161
rect 145276 131 145421 165
rect 145754 161 145800 315
rect 145837 294 145895 527
rect 145930 383 145997 527
rect 146033 349 146075 493
rect 146109 383 146185 527
rect 146229 349 146263 493
rect 146297 383 146373 527
rect 146417 349 146451 493
rect 146485 383 146561 527
rect 146605 349 146639 493
rect 146673 451 146749 527
rect 146838 451 147193 485
rect 147247 435 147281 527
rect 147318 451 147801 485
rect 147845 451 147921 527
rect 147955 417 147989 493
rect 146033 315 146639 349
rect 146673 367 147707 401
rect 147795 383 147989 417
rect 144642 59 144693 125
rect 145276 93 145310 131
rect 145467 127 145800 161
rect 144727 17 144803 93
rect 145039 59 145310 93
rect 145347 17 145423 93
rect 145467 51 145501 127
rect 145535 17 145611 93
rect 145655 51 145689 127
rect 145723 17 145799 93
rect 145837 17 145895 162
rect 146033 161 146085 315
rect 146673 249 146707 367
rect 147795 333 147839 383
rect 147955 359 147989 383
rect 146129 215 146707 249
rect 146673 161 146707 215
rect 146741 299 147229 333
rect 146741 199 146785 299
rect 146853 255 146897 265
rect 146850 221 146897 255
rect 146853 199 146897 221
rect 146946 161 146980 187
rect 146033 127 146639 161
rect 146673 127 146980 161
rect 147028 163 147072 265
rect 147146 199 147229 299
rect 147291 299 147839 333
rect 147291 199 147335 299
rect 147437 233 147481 265
rect 147377 199 147481 233
rect 147689 199 147746 265
rect 147377 163 147411 199
rect 147028 129 147411 163
rect 147542 161 147586 187
rect 145930 17 145997 93
rect 146033 51 146075 127
rect 146109 17 146185 93
rect 146229 59 146263 127
rect 146297 17 146373 93
rect 146417 51 146451 127
rect 146485 17 146561 93
rect 146605 59 146639 127
rect 146673 17 146749 93
rect 146783 59 147017 93
rect 147063 85 147190 129
rect 147455 127 147586 161
rect 147795 163 147839 299
rect 147873 199 147959 323
rect 148045 294 148103 527
rect 148144 459 148465 493
rect 148144 291 148204 459
rect 148241 291 148298 425
rect 148137 212 148204 257
rect 147795 129 147989 163
rect 147244 17 147310 93
rect 147347 59 147625 93
rect 147845 17 147921 93
rect 147955 59 147989 129
rect 148045 17 148103 162
rect 148137 93 148189 177
rect 148241 119 148287 291
rect 148333 265 148373 422
rect 148421 330 148465 459
rect 148499 367 148555 527
rect 148593 330 148669 493
rect 148421 296 148669 330
rect 148321 199 148373 265
rect 148714 262 148759 493
rect 148815 367 148874 527
rect 148417 215 148759 262
rect 148435 165 148660 177
rect 148321 143 148660 165
rect 148321 131 148470 143
rect 148137 85 148208 93
rect 148333 85 148491 93
rect 148137 51 148491 85
rect 148525 17 148559 105
rect 148613 51 148660 143
rect 148706 51 148759 215
rect 148793 152 148870 324
rect 148965 294 149023 527
rect 149057 427 149109 493
rect 149143 451 149219 527
rect 149331 451 149407 527
rect 149451 427 149496 493
rect 149545 435 149595 527
rect 149633 451 150125 485
rect 149057 333 149092 427
rect 149462 401 149496 427
rect 149633 401 149990 417
rect 149237 367 149417 401
rect 149462 383 149990 401
rect 149462 367 149667 383
rect 149383 333 149417 367
rect 150080 357 150125 451
rect 149717 333 149793 343
rect 149057 299 149349 333
rect 149383 299 149793 333
rect 148823 17 148867 109
rect 148965 17 149023 162
rect 149057 135 149092 299
rect 149305 265 149349 299
rect 149126 199 149206 265
rect 149305 231 149477 265
rect 149401 215 149477 231
rect 149584 215 149845 255
rect 149982 199 150057 323
rect 149166 145 149206 199
rect 149057 69 149109 135
rect 149263 115 149311 187
rect 149143 17 149217 109
rect 149357 17 149407 177
rect 149451 147 149793 181
rect 149451 59 149485 147
rect 149717 131 149793 147
rect 149880 165 149941 187
rect 149880 131 149989 165
rect 149545 17 149579 109
rect 150091 93 150125 357
rect 150161 294 150219 527
rect 150255 451 151073 485
rect 151111 451 151177 527
rect 151289 451 151365 527
rect 151477 451 151553 527
rect 149633 59 150125 93
rect 150161 17 150219 162
rect 150255 97 150300 451
rect 151597 417 151631 493
rect 151665 451 151741 527
rect 151785 417 151819 493
rect 151883 451 151949 527
rect 150715 383 151819 417
rect 151597 359 151631 383
rect 151785 359 151819 383
rect 151993 359 152045 493
rect 150339 315 151462 349
rect 151508 285 151966 319
rect 150354 199 150483 265
rect 150707 199 151046 265
rect 151508 258 151542 285
rect 151085 215 151542 258
rect 151722 215 151898 249
rect 150527 165 150606 187
rect 151596 181 151656 187
rect 150339 131 150606 165
rect 150715 131 151443 165
rect 150255 63 151073 97
rect 151111 17 151177 93
rect 151221 51 151255 131
rect 151289 17 151365 93
rect 151409 51 151443 131
rect 151596 143 151819 181
rect 151477 17 151552 118
rect 151596 51 151631 143
rect 151685 17 151735 109
rect 151785 102 151819 143
rect 151854 165 151898 215
rect 151932 199 151966 285
rect 152010 165 152045 359
rect 152093 294 152151 527
rect 152185 299 152241 527
rect 152275 297 152351 493
rect 152395 299 152447 527
rect 152187 211 152254 265
rect 152298 177 152332 297
rect 152553 294 152611 527
rect 152645 299 152697 527
rect 152731 333 152807 493
rect 152851 367 152885 527
rect 152919 333 152995 493
rect 153039 367 153090 527
rect 152731 299 153074 333
rect 152366 215 152443 265
rect 152645 215 152807 265
rect 152841 215 152984 265
rect 153018 181 153074 299
rect 153197 294 153255 527
rect 153290 299 153341 527
rect 153375 333 153451 493
rect 153495 367 153529 527
rect 153563 333 153639 493
rect 153683 367 153717 527
rect 153751 333 153827 493
rect 153871 367 153905 527
rect 153939 333 154015 493
rect 154059 367 154109 527
rect 153375 299 154015 333
rect 153294 215 153648 265
rect 151854 131 152045 165
rect 151883 17 151949 93
rect 151993 51 152045 131
rect 152093 17 152151 162
rect 152185 17 152247 177
rect 152298 51 152447 177
rect 152553 17 152611 162
rect 152645 143 152885 177
rect 152645 51 152713 143
rect 152757 17 152791 109
rect 152825 97 152885 143
rect 152919 131 153074 181
rect 152825 51 153089 97
rect 153197 17 153255 162
rect 153290 143 153717 181
rect 153290 51 153357 143
rect 153401 17 153435 109
rect 153469 51 153545 143
rect 153589 17 153623 109
rect 153657 93 153717 143
rect 153751 161 153811 299
rect 154209 294 154267 527
rect 154302 299 154353 527
rect 154387 333 154463 493
rect 154507 367 154541 527
rect 154575 333 154651 493
rect 154695 367 154729 527
rect 154763 333 154839 493
rect 154883 367 154917 527
rect 154951 333 155027 493
rect 155071 367 155105 527
rect 155139 333 155215 493
rect 155259 367 155293 527
rect 155327 333 155403 493
rect 155447 367 155481 527
rect 155515 333 155591 493
rect 155635 367 155669 527
rect 155703 333 155779 493
rect 154387 293 155779 333
rect 155827 299 155898 527
rect 155957 294 156015 527
rect 156158 367 156208 527
rect 156242 401 156318 493
rect 156362 435 156405 527
rect 156242 367 156470 401
rect 156050 333 156106 365
rect 156050 299 156356 333
rect 153845 215 154095 265
rect 154386 215 155027 259
rect 155092 215 155198 293
rect 155232 215 155685 255
rect 155139 181 155198 215
rect 155729 181 155779 293
rect 156050 215 156116 263
rect 156150 215 156269 263
rect 156322 181 156356 299
rect 153751 127 154015 161
rect 154059 93 154109 177
rect 153657 51 154109 93
rect 154209 17 154267 162
rect 154302 147 155105 181
rect 154302 51 154369 147
rect 154413 17 154447 113
rect 154481 51 154557 147
rect 154601 17 154635 113
rect 154669 51 154745 147
rect 154789 17 154823 113
rect 154857 51 154933 147
rect 154977 17 155011 113
rect 155045 97 155105 147
rect 155139 131 155779 181
rect 155823 97 155898 181
rect 155045 51 155898 97
rect 155957 17 156015 162
rect 156050 147 156356 181
rect 156050 105 156104 147
rect 156396 109 156470 367
rect 156509 294 156567 527
rect 156606 333 156666 372
rect 156710 367 156761 527
rect 156811 401 156877 493
rect 156929 435 157004 527
rect 157041 401 157107 493
rect 156811 367 157107 401
rect 157153 367 157187 527
rect 156606 299 156822 333
rect 156606 168 156640 299
rect 156675 199 156754 265
rect 156788 199 156822 299
rect 156158 17 156224 109
rect 156304 51 156470 109
rect 156509 17 156567 162
rect 156606 102 156653 168
rect 156703 17 156737 155
rect 156875 127 156941 367
rect 157052 299 157107 367
rect 157165 255 157203 331
rect 157245 294 157303 527
rect 157338 333 157405 493
rect 157449 367 157587 527
rect 157338 289 157486 333
rect 157524 289 157587 367
rect 157621 333 157697 493
rect 157741 367 157775 527
rect 157809 333 157888 493
rect 157932 367 157966 527
rect 158000 333 158076 493
rect 158120 367 158154 527
rect 158188 333 158264 493
rect 157621 289 158264 333
rect 158314 299 158380 527
rect 158441 294 158499 527
rect 158534 299 158585 527
rect 158619 333 158695 493
rect 158739 367 158785 527
rect 158819 333 158895 493
rect 158619 299 158895 333
rect 157452 255 157486 289
rect 157006 215 157203 255
rect 157342 215 157408 255
rect 157452 215 157791 255
rect 157452 181 157486 215
rect 157835 181 157888 289
rect 158001 215 158398 255
rect 156975 139 157203 181
rect 156975 93 157025 139
rect 156791 51 157025 93
rect 157069 17 157103 105
rect 157137 51 157203 139
rect 157245 17 157303 162
rect 157338 143 157486 181
rect 157338 51 157405 143
rect 157449 17 157488 109
rect 157537 93 157587 181
rect 157621 127 157888 181
rect 157932 143 158380 181
rect 157932 93 157982 143
rect 157537 51 157982 93
rect 158026 17 158060 109
rect 158094 51 158170 143
rect 158214 17 158262 109
rect 158314 51 158380 143
rect 158441 17 158499 162
rect 158538 149 158582 265
rect 158619 119 158665 299
rect 158993 294 159051 527
rect 159086 299 159137 527
rect 159171 333 159247 493
rect 159291 367 159325 527
rect 159359 333 159435 493
rect 159479 367 159617 527
rect 159651 333 159727 493
rect 159171 289 159727 333
rect 159771 289 159847 527
rect 159913 294 159971 527
rect 160006 289 160057 527
rect 160091 333 160167 493
rect 160211 367 160245 527
rect 160279 333 160355 493
rect 160399 367 160433 527
rect 160467 333 160543 493
rect 160587 367 160621 527
rect 160655 333 160731 493
rect 160775 367 160913 527
rect 160947 333 161023 493
rect 161067 367 161101 527
rect 161135 333 161211 493
rect 161255 367 161308 527
rect 160091 289 161345 333
rect 161385 294 161443 527
rect 161477 319 161562 385
rect 158699 153 158773 265
rect 158811 199 158897 265
rect 159086 199 159134 265
rect 158819 119 158895 165
rect 158534 17 158585 115
rect 158619 51 158895 119
rect 158993 17 159051 162
rect 159086 93 159137 157
rect 159171 127 159247 289
rect 159302 215 159591 255
rect 159625 215 159868 255
rect 160010 215 160358 255
rect 160443 215 160793 255
rect 160838 215 161262 255
rect 161299 181 161345 289
rect 159359 127 159727 181
rect 159086 59 159529 93
rect 159567 17 159633 93
rect 159771 17 159847 177
rect 159913 17 159971 162
rect 160006 147 160825 181
rect 160006 51 160073 147
rect 160117 17 160151 113
rect 160185 51 160261 147
rect 160373 131 160449 147
rect 160561 131 160637 147
rect 160749 131 160825 147
rect 160947 131 161345 181
rect 161477 165 161511 319
rect 161612 299 161662 527
rect 161696 333 161772 493
rect 161818 367 161852 527
rect 161886 333 161995 493
rect 161696 299 161995 333
rect 161545 199 161625 265
rect 161663 199 161727 265
rect 161764 199 161819 265
rect 161860 165 161904 265
rect 160305 17 160339 113
rect 160467 51 161308 97
rect 161385 17 161443 162
rect 161477 131 161904 165
rect 161477 89 161562 131
rect 161942 97 161995 299
rect 162029 294 162087 527
rect 162122 413 162186 493
rect 162122 323 162156 413
rect 162230 367 162292 527
rect 162326 401 162402 493
rect 162446 435 162480 527
rect 162514 401 162590 493
rect 162634 435 162684 527
rect 162722 435 162782 527
rect 162326 391 162590 401
rect 162816 401 162876 493
rect 162936 435 162994 527
rect 162816 391 163002 401
rect 162326 357 163002 391
rect 162122 289 162904 323
rect 161612 17 161678 97
rect 161886 51 161995 97
rect 162029 17 162087 162
rect 162122 131 162156 289
rect 162190 215 162270 255
rect 162317 215 162482 255
rect 162534 215 162792 255
rect 162838 215 162904 289
rect 162954 181 163002 357
rect 163041 294 163099 527
rect 162122 51 162186 131
rect 162230 17 162292 181
rect 162326 143 162704 181
rect 162326 51 162402 143
rect 162544 127 162704 143
rect 162446 17 162496 109
rect 162748 93 162782 181
rect 162816 127 163002 181
rect 163133 289 163201 493
rect 163245 289 163383 527
rect 163417 333 163493 493
rect 163537 367 163571 527
rect 163605 401 163681 493
rect 163725 435 163759 527
rect 163793 401 163869 493
rect 163605 333 163869 401
rect 163913 367 163947 527
rect 163981 333 164057 493
rect 164101 367 164239 527
rect 164273 333 164349 493
rect 164393 367 164427 527
rect 164461 333 164537 493
rect 163417 289 164537 333
rect 164581 289 164647 527
rect 164697 294 164755 527
rect 164789 299 164841 527
rect 164875 333 164951 493
rect 164995 367 165029 527
rect 165079 333 165145 493
rect 165195 367 165251 527
rect 164875 299 165161 333
rect 163133 181 163168 289
rect 163202 215 163282 255
rect 163327 215 163681 255
rect 163725 215 163827 289
rect 163861 215 164102 255
rect 164153 215 164536 255
rect 163327 181 163383 215
rect 163725 181 163759 215
rect 164794 199 164851 265
rect 164891 199 164987 265
rect 165021 199 165093 265
rect 162544 51 162994 93
rect 163041 17 163099 162
rect 163133 143 163383 181
rect 163133 51 163201 143
rect 163417 127 163759 181
rect 163793 143 164537 181
rect 163793 127 164151 143
rect 163245 17 163295 109
rect 163333 51 164151 93
rect 164189 17 164239 109
rect 164273 51 164349 143
rect 164393 17 164427 109
rect 164461 51 164537 143
rect 164581 17 164647 181
rect 164697 17 164755 162
rect 164790 17 164857 165
rect 164891 60 164944 199
rect 165021 165 165055 199
rect 165127 165 165161 299
rect 165207 199 165300 333
rect 165341 294 165399 527
rect 165434 299 165485 527
rect 165519 333 165595 493
rect 165639 367 165673 527
rect 165707 333 165783 493
rect 165827 367 165893 527
rect 165927 333 166003 493
rect 166075 367 166151 527
rect 166205 333 166281 493
rect 165519 289 166281 333
rect 166325 289 166391 527
rect 166445 294 166503 527
rect 166538 289 166589 527
rect 166623 333 166699 493
rect 166743 367 166777 527
rect 166811 333 166887 493
rect 166931 367 166965 527
rect 166999 333 167075 493
rect 167119 367 167153 527
rect 167187 333 167263 493
rect 167307 367 167445 527
rect 167479 333 167555 493
rect 167599 367 167633 527
rect 167667 333 167743 493
rect 167794 367 167828 527
rect 167867 333 167943 493
rect 167987 367 168021 527
rect 168055 333 168131 493
rect 166623 289 168131 333
rect 168175 289 168227 527
rect 168285 294 168343 527
rect 168377 319 168461 385
rect 165438 215 165595 255
rect 165629 215 165786 255
rect 165903 215 166092 255
rect 166160 211 166281 289
rect 166339 215 166405 255
rect 166541 215 166887 255
rect 166958 215 167325 255
rect 167370 215 167743 255
rect 164978 60 165055 165
rect 165106 51 165255 165
rect 165341 17 165399 162
rect 165434 147 165673 181
rect 165434 51 165501 147
rect 165545 17 165579 109
rect 165613 93 165673 147
rect 165707 127 166093 181
rect 166137 93 166171 177
rect 166205 127 166281 211
rect 167829 181 167885 289
rect 167943 215 168222 255
rect 166325 93 166391 181
rect 165613 51 165881 93
rect 165919 51 166391 93
rect 166445 17 166503 162
rect 166538 131 166965 181
rect 166999 131 167743 181
rect 167829 131 168131 181
rect 166538 51 166589 131
rect 166623 17 166699 97
rect 166743 51 166777 131
rect 166931 97 166965 131
rect 168175 97 168226 181
rect 168377 165 168411 319
rect 168511 299 168561 527
rect 168595 333 168671 493
rect 168705 367 168760 527
rect 168795 333 168861 493
rect 168935 367 168978 527
rect 168595 299 168987 333
rect 168445 199 168524 265
rect 168562 199 168626 265
rect 168660 192 168712 265
rect 166811 17 166887 97
rect 166931 51 167357 97
rect 167395 51 168226 97
rect 168285 17 168343 162
rect 168377 131 168634 165
rect 168668 153 168712 192
rect 168746 153 168805 265
rect 168839 199 168901 265
rect 168377 89 168454 131
rect 168600 119 168634 131
rect 168839 119 168880 199
rect 168935 167 168987 299
rect 169021 294 169079 527
rect 169114 417 169165 493
rect 169199 451 169363 527
rect 169114 383 169240 417
rect 169114 199 169162 323
rect 169196 249 169240 383
rect 169313 289 169363 451
rect 169397 333 169473 493
rect 169517 367 169551 527
rect 169585 333 169661 493
rect 169705 367 169833 527
rect 169867 333 169943 493
rect 169987 367 170039 527
rect 170073 333 170149 493
rect 169397 289 170149 333
rect 170193 299 170272 527
rect 170309 294 170367 527
rect 170402 333 170469 493
rect 170513 367 170651 527
rect 170402 299 170555 333
rect 170593 299 170651 367
rect 170685 333 170761 493
rect 170805 367 170839 527
rect 170873 333 170949 493
rect 170993 367 171027 527
rect 171061 333 171137 493
rect 171181 367 171215 527
rect 171249 333 171325 493
rect 171369 367 171507 527
rect 171541 333 171617 493
rect 171661 367 171695 527
rect 171729 333 171805 493
rect 171849 367 171883 527
rect 171917 333 171993 493
rect 172037 367 172071 527
rect 172105 333 172181 493
rect 169196 215 169363 249
rect 168493 17 168566 97
rect 168600 85 168880 119
rect 168915 51 168987 167
rect 169021 17 169079 162
rect 169196 161 169240 215
rect 169114 127 169240 161
rect 169114 51 169165 127
rect 169313 93 169363 181
rect 169397 127 169473 289
rect 170516 255 170555 299
rect 170685 289 172181 333
rect 172225 289 172276 527
rect 172333 294 172391 527
rect 172425 413 172493 493
rect 169528 215 169766 255
rect 169818 215 170033 255
rect 170100 215 170273 255
rect 170406 215 170472 255
rect 170516 215 170779 255
rect 170516 181 170555 215
rect 170866 181 170952 289
rect 171020 215 171392 255
rect 171432 215 171806 255
rect 171917 215 172285 255
rect 172425 181 172460 413
rect 172537 367 172603 527
rect 172639 333 172705 493
rect 172747 367 172811 527
rect 172846 401 172924 493
rect 172958 435 173112 527
rect 173156 401 173219 493
rect 172846 333 172944 401
rect 172494 215 172573 331
rect 172639 299 172944 333
rect 172607 215 172673 265
rect 169517 127 169755 181
rect 169793 143 170254 181
rect 169793 127 170057 143
rect 169517 93 169551 127
rect 169997 123 170057 127
rect 169199 17 169275 93
rect 169313 51 169551 93
rect 169585 51 169953 93
rect 169997 51 170049 123
rect 170109 17 170143 109
rect 170187 51 170254 143
rect 170309 17 170367 162
rect 170402 147 170555 181
rect 170402 51 170469 147
rect 170513 17 170563 109
rect 170601 93 170651 181
rect 170685 127 170952 181
rect 171061 127 171805 181
rect 171849 147 172276 181
rect 171849 93 171899 147
rect 170601 51 171419 93
rect 171457 51 171899 93
rect 171943 17 171977 109
rect 172011 51 172087 147
rect 172131 17 172165 109
rect 172199 51 172276 147
rect 172333 17 172391 162
rect 172425 143 172652 181
rect 172707 147 172760 265
rect 172425 97 172493 143
rect 172618 111 172652 143
rect 172806 111 172856 265
rect 172537 17 172584 109
rect 172618 73 172856 111
rect 172890 165 172944 299
rect 172978 367 173219 401
rect 172978 199 173033 367
rect 172890 51 173008 165
rect 173068 145 173150 323
rect 173185 109 173219 367
rect 173253 294 173311 527
rect 173345 396 173402 488
rect 173436 439 173491 527
rect 173525 430 173663 493
rect 173345 357 173594 396
rect 173345 214 173394 323
rect 173440 214 173516 323
rect 173560 180 173594 357
rect 173046 17 173116 109
rect 173150 51 173219 109
rect 173253 17 173311 162
rect 173345 146 173594 180
rect 173345 51 173397 146
rect 173628 112 173663 430
rect 173697 299 173731 527
rect 173765 333 173825 493
rect 173859 367 173919 527
rect 173953 333 174029 493
rect 174073 367 174205 527
rect 174239 333 174315 493
rect 174359 367 174393 527
rect 174427 333 174503 493
rect 173765 289 174503 333
rect 174547 289 174597 527
rect 174633 294 174691 527
rect 174725 396 174782 488
rect 174816 439 174871 527
rect 174905 430 175077 493
rect 174725 357 175009 396
rect 173765 131 173854 289
rect 173917 215 173993 255
rect 174027 215 174137 289
rect 174176 215 174318 255
rect 174391 215 174587 255
rect 174728 199 174774 323
rect 174825 199 174913 323
rect 173953 131 174315 181
rect 174359 147 174597 181
rect 173431 17 173491 109
rect 173525 51 173663 112
rect 173697 97 173731 117
rect 174359 97 174409 147
rect 173697 51 174123 97
rect 174161 51 174409 97
rect 174453 17 174487 113
rect 174521 51 174597 147
rect 174633 17 174691 162
rect 174947 161 175009 357
rect 174725 127 175009 161
rect 175043 261 175077 430
rect 175111 299 175145 527
rect 175179 333 175239 493
rect 175273 367 175333 527
rect 175367 333 175443 493
rect 175487 367 175521 527
rect 175555 333 175631 493
rect 175675 367 175709 527
rect 175743 333 175819 493
rect 175873 367 176001 527
rect 176041 333 176117 493
rect 176161 367 176195 527
rect 176229 333 176305 493
rect 176349 367 176383 527
rect 176417 333 176493 493
rect 176537 367 176571 527
rect 176605 333 176681 493
rect 175179 289 176681 333
rect 176725 289 176780 527
rect 176841 294 176899 527
rect 176935 333 177001 490
rect 176935 299 177071 333
rect 177139 299 177241 527
rect 175043 215 175113 261
rect 175179 215 175348 249
rect 174725 51 174777 127
rect 175043 93 175077 215
rect 175441 181 175511 289
rect 175545 215 175819 255
rect 175917 215 176305 255
rect 176387 215 176776 255
rect 176933 215 177003 265
rect 174811 17 174887 93
rect 174931 51 175077 93
rect 175111 97 175145 181
rect 175179 131 175511 181
rect 175555 131 176310 181
rect 177037 179 177071 299
rect 177301 294 177359 527
rect 177394 333 177449 493
rect 177483 367 177559 527
rect 177603 459 177851 493
rect 177603 333 177637 459
rect 177394 291 177637 333
rect 177671 333 177747 425
rect 177791 367 177851 459
rect 177671 289 177838 333
rect 177945 294 178003 527
rect 178038 333 178093 493
rect 178127 367 178203 527
rect 178247 333 178281 493
rect 178315 367 178375 527
rect 178409 459 178878 493
rect 178409 333 178485 459
rect 178038 291 178485 333
rect 178529 349 178563 425
rect 178597 387 178673 459
rect 178717 349 178751 425
rect 178785 383 178878 459
rect 178529 289 178918 349
rect 178957 294 179015 527
rect 179050 333 179113 493
rect 179157 367 179207 527
rect 179251 333 179301 493
rect 179345 367 179395 527
rect 179439 333 179489 493
rect 179533 367 179583 527
rect 179627 333 179677 493
rect 179721 367 179771 527
rect 179815 459 180617 493
rect 179815 333 179865 459
rect 179050 291 179865 333
rect 179909 323 179959 425
rect 180003 357 180053 459
rect 180097 323 180147 425
rect 180191 357 180241 459
rect 180285 323 180335 425
rect 180379 357 180429 459
rect 180473 323 180523 425
rect 180567 357 180617 459
rect 179909 289 180637 323
rect 180705 294 180763 527
rect 180935 451 181001 527
rect 180799 383 181077 417
rect 177125 215 177195 265
rect 177394 215 177548 255
rect 177582 215 177756 255
rect 177795 181 177838 289
rect 178048 215 178410 255
rect 178484 215 178787 255
rect 178839 181 178918 289
rect 179104 215 179818 255
rect 179872 215 180490 255
rect 180524 181 180637 289
rect 176349 131 176765 165
rect 176349 97 176383 131
rect 175111 51 175913 97
rect 175961 51 176383 97
rect 176427 17 176493 97
rect 176615 17 176681 97
rect 176841 17 176899 162
rect 176937 17 176985 179
rect 177019 51 177095 179
rect 177129 17 177231 179
rect 177301 17 177359 162
rect 177394 17 177449 181
rect 177483 147 177838 181
rect 177483 145 177747 147
rect 177483 51 177559 145
rect 177603 17 177637 111
rect 177671 51 177747 145
rect 177804 17 177872 111
rect 177945 17 178003 162
rect 178038 17 178093 181
rect 178127 145 178918 181
rect 178127 51 178203 145
rect 178247 17 178281 111
rect 178315 51 178391 145
rect 178435 17 178469 111
rect 178503 51 178579 145
rect 178623 17 178657 111
rect 178691 51 178767 145
rect 178811 17 178868 111
rect 178957 17 179015 162
rect 179050 17 179105 181
rect 179139 145 180637 181
rect 179139 51 179215 145
rect 179259 17 179293 111
rect 179327 51 179403 145
rect 179447 17 179481 111
rect 179515 51 179591 145
rect 179635 17 179669 111
rect 179703 51 179779 145
rect 179823 17 179857 111
rect 179891 51 179967 145
rect 180011 17 180045 111
rect 180079 51 180155 145
rect 180199 17 180233 111
rect 180267 51 180343 145
rect 180387 17 180421 111
rect 180455 51 180531 145
rect 180575 17 180633 111
rect 180705 17 180763 162
rect 180799 58 180849 383
rect 180883 195 180937 349
rect 181043 333 181077 383
rect 181111 370 181223 493
rect 181043 299 181111 333
rect 181077 265 181111 299
rect 180971 213 181037 265
rect 181077 215 181153 265
rect 181187 179 181223 370
rect 181257 294 181315 527
rect 181349 331 181413 493
rect 181457 365 181507 527
rect 181551 459 181797 493
rect 181551 331 181601 459
rect 181349 289 181601 331
rect 181428 213 181584 255
rect 181645 179 181695 425
rect 181739 289 181797 459
rect 181851 249 181885 492
rect 181969 429 182019 527
rect 181986 255 182039 393
rect 182085 294 182143 527
rect 182177 333 182233 493
rect 182267 367 182343 527
rect 182387 333 182421 493
rect 182455 367 182515 527
rect 182549 459 183005 493
rect 182549 333 182625 459
rect 182177 291 182625 333
rect 182669 349 182703 425
rect 182737 387 182813 459
rect 182857 349 182891 425
rect 182669 283 182891 349
rect 182925 315 183005 459
rect 181747 215 181885 249
rect 181007 145 181223 179
rect 180915 17 180973 125
rect 181007 51 181083 145
rect 181127 17 181204 111
rect 181257 17 181315 162
rect 181349 17 181405 179
rect 181439 145 181703 179
rect 181439 51 181519 145
rect 181559 17 181593 111
rect 181627 51 181703 145
rect 181747 17 181781 179
rect 181851 89 181885 215
rect 181924 213 182039 255
rect 182232 215 182550 255
rect 182669 181 182735 283
rect 183039 249 183111 493
rect 183155 299 183236 527
rect 183281 294 183339 527
rect 183374 456 183639 490
rect 183374 299 183441 456
rect 183475 265 183532 401
rect 182773 215 183111 249
rect 183145 215 183245 264
rect 181969 17 182020 169
rect 182085 17 182143 162
rect 182177 17 182233 181
rect 182267 145 182907 181
rect 182267 51 182343 145
rect 182387 17 182421 111
rect 182455 51 182531 145
rect 182575 17 182609 111
rect 182643 51 182719 145
rect 182763 17 182797 111
rect 182831 51 182907 145
rect 182951 17 182985 181
rect 183039 51 183111 215
rect 183374 199 183441 265
rect 183475 199 183571 265
rect 183155 17 183213 181
rect 183605 165 183639 456
rect 183673 367 183791 527
rect 183281 17 183339 162
rect 183374 131 183639 165
rect 183704 131 183797 333
rect 183833 294 183891 527
rect 183938 325 183989 493
rect 184033 359 184083 527
rect 184127 325 184177 493
rect 184221 459 184680 493
rect 184221 359 184271 459
rect 184315 325 184363 425
rect 184450 359 184492 459
rect 184544 325 184586 425
rect 184630 359 184680 459
rect 183938 291 184363 325
rect 184397 257 184495 325
rect 184544 291 184707 325
rect 184753 294 184811 527
rect 184858 325 184909 493
rect 184953 359 185003 527
rect 185047 325 185097 493
rect 185141 359 185191 527
rect 185235 417 185473 493
rect 185235 325 185285 417
rect 184858 291 185285 325
rect 185329 325 185379 383
rect 185423 359 185473 417
rect 185517 459 185943 493
rect 185517 325 185567 459
rect 185705 427 185755 459
rect 185893 427 185943 459
rect 185987 425 186037 493
rect 185611 393 185661 425
rect 185799 393 185849 425
rect 185611 391 185849 393
rect 185611 357 186097 391
rect 185329 291 185567 325
rect 183935 215 184111 257
rect 184155 215 184363 257
rect 184397 215 184570 257
rect 184604 181 184707 291
rect 185611 289 185971 323
rect 185611 257 185645 289
rect 184846 215 185233 257
rect 185287 215 185645 257
rect 185937 257 185971 289
rect 185679 215 185891 255
rect 185937 215 186005 257
rect 186039 181 186097 357
rect 186133 294 186191 527
rect 183374 77 183425 131
rect 183459 17 183535 97
rect 183579 77 183613 131
rect 183647 17 183791 97
rect 183833 17 183891 162
rect 183926 17 183981 181
rect 184015 145 184707 181
rect 184015 51 184091 145
rect 184135 17 184169 111
rect 184203 51 184279 145
rect 184323 17 184484 111
rect 184518 51 184594 145
rect 184638 17 184696 111
rect 184753 17 184811 162
rect 184846 17 184901 181
rect 184935 145 186097 181
rect 186225 289 186317 491
rect 186551 425 186627 527
rect 186351 357 186743 391
rect 186225 165 186259 289
rect 186351 249 186385 357
rect 186293 215 186385 249
rect 186419 199 186469 323
rect 186503 199 186571 323
rect 186605 199 186675 323
rect 186709 165 186743 357
rect 186777 294 186835 527
rect 186870 325 186933 493
rect 186977 359 187027 527
rect 187071 325 187121 493
rect 187165 455 187608 493
rect 187165 359 187215 455
rect 187251 325 187317 407
rect 186870 291 187317 325
rect 186874 215 187055 257
rect 187099 215 187292 257
rect 187426 181 187523 409
rect 187559 291 187608 455
rect 187650 291 187721 374
rect 187765 308 187815 527
rect 187881 294 187939 527
rect 187978 325 188037 493
rect 188081 359 188131 527
rect 188175 393 188225 493
rect 188269 427 188319 527
rect 188363 393 188413 493
rect 188457 427 188507 527
rect 188561 459 189363 493
rect 188561 427 188611 459
rect 188749 427 188799 459
rect 188655 393 188705 425
rect 188843 393 188893 425
rect 188175 359 188893 393
rect 188937 359 188987 459
rect 189031 325 189081 425
rect 189125 359 189175 459
rect 189219 325 189269 425
rect 189313 359 189363 459
rect 187978 291 188987 325
rect 189031 291 189405 325
rect 189445 294 189503 527
rect 189538 333 189605 490
rect 189538 299 189675 333
rect 187650 257 187684 291
rect 187559 215 187684 257
rect 187718 215 187835 257
rect 187978 215 188045 257
rect 184935 51 185011 145
rect 185055 17 185089 111
rect 185123 51 185199 145
rect 185243 17 185277 111
rect 185311 51 185387 145
rect 185431 17 185465 111
rect 185499 51 185575 145
rect 185619 17 185653 111
rect 185687 51 185763 145
rect 185807 17 185841 111
rect 185875 51 185951 145
rect 185995 17 186029 111
rect 186133 17 186191 162
rect 186225 131 186517 165
rect 186225 51 186329 131
rect 186363 17 186439 97
rect 186483 62 186517 131
rect 186551 17 186627 165
rect 186684 131 186743 165
rect 186684 81 186718 131
rect 186777 17 186835 162
rect 186870 17 186925 181
rect 186959 145 187523 181
rect 187650 181 187684 215
rect 188089 181 188123 291
rect 188953 257 188987 291
rect 188198 215 188510 257
rect 188613 215 188896 257
rect 188953 215 189300 257
rect 189337 181 189405 291
rect 186959 51 187035 145
rect 187079 17 187113 111
rect 187147 51 187223 145
rect 187267 17 187405 111
rect 187439 51 187523 145
rect 187567 17 187608 179
rect 187650 76 187721 181
rect 187765 17 187823 165
rect 187881 17 187939 162
rect 187978 147 188123 181
rect 187978 51 188045 147
rect 188157 145 189405 181
rect 188089 17 188123 111
rect 188157 51 188233 145
rect 188277 17 188311 111
rect 188345 51 188421 145
rect 188465 17 188603 111
rect 188637 51 188713 145
rect 188757 17 188791 111
rect 188825 51 188901 145
rect 188945 17 188979 111
rect 189013 51 189089 145
rect 189133 17 189167 111
rect 189201 51 189277 145
rect 189321 17 189355 111
rect 189445 17 189503 162
rect 189537 149 189587 265
rect 189623 165 189675 299
rect 189713 199 189777 490
rect 189811 199 189869 490
rect 189947 367 190027 527
rect 189623 131 189873 165
rect 189907 131 189961 333
rect 190089 294 190147 527
rect 190194 325 190245 493
rect 190289 359 190339 527
rect 190383 325 190433 493
rect 190477 459 190827 493
rect 190477 359 190527 459
rect 190571 325 190621 425
rect 190194 291 190621 325
rect 190683 325 190733 425
rect 190777 359 190827 459
rect 190871 459 191109 493
rect 190871 325 190921 459
rect 190683 291 190921 325
rect 190972 325 191022 425
rect 191059 359 191109 459
rect 190972 291 191154 325
rect 191193 294 191251 527
rect 191286 325 191349 493
rect 191393 359 191443 527
rect 191487 325 191537 493
rect 191581 359 191631 527
rect 191675 459 192112 493
rect 191675 325 191725 459
rect 191286 291 191725 325
rect 191769 325 191819 425
rect 191863 359 191913 459
rect 191957 325 192007 425
rect 192051 359 192112 459
rect 192149 459 192957 493
rect 192149 359 192205 459
rect 192249 325 192299 425
rect 192343 359 192393 459
rect 192437 325 192487 425
rect 192531 359 192581 459
rect 191769 291 192487 325
rect 192625 325 192675 425
rect 192719 359 192769 459
rect 192813 325 192863 425
rect 192907 359 192957 459
rect 192625 291 192994 325
rect 193033 294 193091 527
rect 190204 215 190367 257
rect 190411 215 190592 257
rect 190646 215 190835 257
rect 190892 215 191019 257
rect 191087 181 191154 291
rect 191304 215 191673 257
rect 191727 215 192162 257
rect 192207 215 192529 257
rect 192563 215 192877 257
rect 192940 181 192994 291
rect 189537 17 189589 115
rect 189623 77 189683 131
rect 189727 17 189793 97
rect 189839 77 189873 131
rect 189921 17 190024 97
rect 190089 17 190147 162
rect 190182 17 190237 181
rect 190278 145 191154 181
rect 190278 51 190354 145
rect 190391 17 190425 111
rect 190466 51 190542 145
rect 190579 17 190725 111
rect 190766 51 190842 145
rect 190879 17 190913 111
rect 190954 51 191030 145
rect 191067 17 191125 111
rect 191193 17 191251 162
rect 191286 17 191341 181
rect 191375 145 192994 181
rect 193125 165 193177 490
rect 193573 437 193649 527
rect 193213 359 193821 401
rect 193213 199 193257 359
rect 193295 199 193365 323
rect 193403 199 193495 323
rect 193543 199 193639 323
rect 193673 199 193753 323
rect 193787 165 193821 359
rect 193861 294 193919 527
rect 193953 325 194021 493
rect 194065 359 194107 527
rect 194151 325 194201 493
rect 194245 459 194594 493
rect 194245 359 194287 459
rect 194321 325 194397 425
rect 193953 291 194397 325
rect 194431 325 194508 425
rect 194552 359 194594 459
rect 194638 459 194875 493
rect 194638 325 194688 459
rect 194431 291 194688 325
rect 194732 325 194782 425
rect 194826 359 194875 459
rect 194909 407 194980 490
rect 195024 427 195074 527
rect 194732 291 194834 325
rect 193956 215 194204 257
rect 194241 215 194466 257
rect 194508 215 194668 257
rect 194749 215 194834 291
rect 194909 249 194943 407
rect 195059 257 195113 391
rect 195149 294 195207 527
rect 195243 325 195309 493
rect 195353 359 195395 527
rect 195439 325 195489 493
rect 195533 359 195583 527
rect 195627 459 196053 493
rect 195627 325 195677 459
rect 195243 291 195677 325
rect 195721 325 195771 425
rect 195815 359 195865 459
rect 195909 325 195959 425
rect 196003 359 196053 459
rect 196107 459 196909 493
rect 196107 359 196157 459
rect 196201 325 196251 425
rect 196295 359 196345 459
rect 196389 325 196439 425
rect 195721 291 196439 325
rect 196483 291 196533 459
rect 196577 325 196627 425
rect 196671 359 196721 459
rect 196765 325 196815 425
rect 196859 359 196909 459
rect 196954 325 197021 493
rect 196577 291 196815 325
rect 196878 291 197021 325
rect 197065 291 197111 527
rect 197173 294 197231 527
rect 197265 414 197317 491
rect 197351 448 197427 527
rect 197475 459 197771 493
rect 197475 414 197509 459
rect 197265 377 197509 414
rect 197563 391 197690 425
rect 194880 215 194943 249
rect 194977 215 195113 257
rect 195303 215 195625 257
rect 195679 215 196054 257
rect 196101 215 196481 257
rect 194749 181 194790 215
rect 191375 51 191451 145
rect 191495 17 191529 111
rect 191563 51 191639 145
rect 191683 17 191717 111
rect 191751 51 191827 145
rect 191871 17 191905 111
rect 191939 51 192015 145
rect 192059 17 192197 111
rect 192231 51 192307 145
rect 192351 17 192385 111
rect 192419 51 192495 145
rect 192539 17 192573 111
rect 192607 51 192683 145
rect 192727 17 192761 111
rect 192795 51 192871 145
rect 192915 17 192949 111
rect 193033 17 193091 162
rect 193125 131 193523 165
rect 193179 17 193245 96
rect 193289 60 193329 131
rect 193373 17 193439 97
rect 193483 62 193523 131
rect 193557 17 193655 165
rect 193726 131 193821 165
rect 193726 81 193760 131
rect 193861 17 193919 162
rect 193953 17 194005 181
rect 194039 145 194790 181
rect 194909 181 194943 215
rect 196577 181 196674 291
rect 196878 257 196912 291
rect 196708 215 196912 257
rect 196995 215 197134 257
rect 196878 181 196912 215
rect 194039 51 194115 145
rect 194159 17 194193 111
rect 194227 51 194303 145
rect 194347 17 194492 111
rect 194526 51 194602 145
rect 194646 17 194680 111
rect 194714 51 194790 145
rect 194834 17 194875 179
rect 194909 76 194980 181
rect 195024 17 195074 165
rect 195149 17 195207 162
rect 195259 17 195293 179
rect 195327 145 196823 181
rect 196878 147 197021 181
rect 195327 51 195403 145
rect 195447 17 195481 111
rect 195515 51 195591 145
rect 195635 17 195669 111
rect 195703 51 195779 145
rect 195823 17 195857 111
rect 195891 51 195967 145
rect 196011 17 196149 111
rect 196183 51 196259 145
rect 196303 17 196337 111
rect 196371 51 196447 145
rect 196491 17 196525 111
rect 196559 51 196635 145
rect 196679 17 196713 111
rect 196747 51 196823 145
rect 196867 17 196901 111
rect 196946 51 197021 147
rect 197065 17 197111 181
rect 197265 165 197300 377
rect 197334 199 197414 339
rect 197468 305 197606 343
rect 197448 199 197516 265
rect 197572 165 197606 305
rect 197173 17 197231 162
rect 197265 90 197329 165
rect 197389 17 197423 165
rect 197483 131 197606 165
rect 197640 165 197690 391
rect 197724 199 197771 459
rect 197812 199 197874 482
rect 197950 375 198046 527
rect 197920 199 197981 341
rect 198093 294 198151 527
rect 198185 411 198237 491
rect 198271 448 198347 527
rect 198503 445 198945 493
rect 198987 443 199233 493
rect 198185 377 198558 411
rect 198185 165 198219 377
rect 198253 199 198334 339
rect 198377 305 198490 343
rect 198368 199 198422 265
rect 198456 249 198490 305
rect 198524 317 198558 377
rect 198597 375 199147 409
rect 198524 283 198741 317
rect 198775 289 199014 341
rect 199089 291 199147 375
rect 199191 325 199233 443
rect 199277 359 199319 527
rect 199353 325 199429 493
rect 199191 291 199429 325
rect 199473 294 199531 527
rect 199565 409 199621 493
rect 199655 443 199731 527
rect 199871 459 200687 493
rect 199871 443 200313 459
rect 199565 375 200313 409
rect 199565 307 199715 375
rect 199749 307 199895 341
rect 198707 255 198741 283
rect 198456 215 198663 249
rect 198707 215 198896 255
rect 198456 165 198490 215
rect 198930 181 199014 289
rect 199048 215 199227 255
rect 199261 215 199434 255
rect 199570 215 199637 273
rect 197640 131 197916 165
rect 197483 90 197517 131
rect 197572 17 197638 96
rect 197682 60 197722 131
rect 197766 17 197832 97
rect 197876 62 197916 131
rect 197950 17 198046 165
rect 198093 17 198151 162
rect 198185 90 198261 165
rect 198305 17 198339 165
rect 198399 131 198490 165
rect 198587 145 199335 181
rect 198399 90 198438 131
rect 198487 17 198553 96
rect 198587 51 198663 145
rect 198707 17 198741 111
rect 198775 51 198851 145
rect 198895 17 199037 111
rect 199071 51 199147 145
rect 199191 17 199225 111
rect 199259 51 199335 145
rect 199379 17 199434 181
rect 199681 179 199715 307
rect 199749 215 199827 265
rect 199861 249 199895 307
rect 199936 283 200235 341
rect 199861 215 200167 249
rect 199861 181 199895 215
rect 200201 181 200235 283
rect 200279 257 200313 375
rect 200357 325 200399 425
rect 200443 359 200493 459
rect 200537 325 200587 425
rect 200631 359 200687 459
rect 200724 459 201161 493
rect 200724 359 200785 459
rect 200829 325 200879 425
rect 200923 359 200973 459
rect 201017 325 201067 425
rect 200357 291 201067 325
rect 201111 325 201161 459
rect 201205 359 201255 527
rect 201299 325 201349 493
rect 201393 359 201443 527
rect 201487 325 201550 493
rect 201111 291 201550 325
rect 201589 294 201647 527
rect 201681 299 201749 493
rect 201793 299 201827 527
rect 201881 367 201931 527
rect 202081 333 202157 493
rect 202216 367 202282 527
rect 202358 333 202424 493
rect 201865 299 202424 333
rect 200279 215 200629 257
rect 200678 215 201109 257
rect 201163 215 201550 257
rect 199473 17 199531 162
rect 199565 145 199715 179
rect 199749 147 199895 181
rect 199565 51 199637 145
rect 199681 17 199715 111
rect 199749 51 199825 147
rect 199955 145 201451 181
rect 199887 17 199921 111
rect 199955 51 200031 145
rect 200075 17 200109 111
rect 200143 51 200219 145
rect 200263 17 200297 111
rect 200331 51 200407 145
rect 200451 17 200485 111
rect 200519 51 200595 145
rect 200639 17 200777 111
rect 200811 51 200887 145
rect 200931 17 200965 111
rect 200999 51 201075 145
rect 201119 17 201153 111
rect 201187 51 201263 145
rect 201307 17 201341 111
rect 201375 51 201451 145
rect 201495 17 201550 181
rect 201681 177 201716 299
rect 201865 249 201899 299
rect 201750 215 201899 249
rect 201934 215 202027 255
rect 202061 215 202138 255
rect 202172 215 202280 255
rect 201589 17 201647 162
rect 201681 51 201749 177
rect 201793 17 201843 177
rect 201881 147 202146 181
rect 201881 51 201947 147
rect 201991 17 202036 109
rect 202070 51 202146 147
rect 202227 87 202280 215
rect 202314 173 202358 299
rect 202509 294 202567 527
rect 202602 353 202655 493
rect 202689 387 202765 527
rect 202809 353 202948 493
rect 203059 387 203155 527
rect 203201 415 203239 493
rect 203273 451 203349 527
rect 203201 381 203391 415
rect 202602 347 202948 353
rect 202602 302 203189 347
rect 202392 215 202465 265
rect 202601 199 202656 265
rect 202314 51 202424 173
rect 202690 165 202736 302
rect 203155 265 203189 302
rect 202770 199 202846 265
rect 202885 199 202973 265
rect 203017 199 203119 265
rect 203155 199 203297 265
rect 202509 17 202567 162
rect 202603 85 202736 165
rect 202770 127 203059 165
rect 203337 157 203391 381
rect 203429 294 203487 527
rect 203600 374 203676 527
rect 203720 340 203756 493
rect 203792 374 203868 527
rect 203912 340 203950 493
rect 203984 440 204060 527
rect 204104 405 204176 493
rect 204211 439 204287 527
rect 204321 405 204387 493
rect 204423 439 204476 527
rect 204597 405 204673 493
rect 203521 287 203950 340
rect 203984 371 204673 405
rect 204789 383 204865 527
rect 203173 123 203391 157
rect 202603 51 202670 85
rect 202891 17 202958 93
rect 203092 17 203139 105
rect 203173 51 203249 123
rect 203293 17 203359 89
rect 203429 17 203487 162
rect 203521 161 203577 287
rect 203984 253 204028 371
rect 203611 213 204028 253
rect 203984 163 204028 213
rect 204062 289 204424 337
rect 204062 199 204121 289
rect 204155 207 204322 255
rect 204358 207 204424 289
rect 204469 299 204867 337
rect 204469 207 204535 299
rect 204572 207 204727 265
rect 204764 207 204867 299
rect 204901 294 204959 527
rect 204995 299 205055 527
rect 205089 265 205141 450
rect 205175 409 205241 489
rect 205284 455 205350 527
rect 205391 409 205511 493
rect 205175 363 205511 409
rect 205175 319 205241 363
rect 205275 269 205325 323
rect 204993 199 205055 265
rect 205089 199 205192 265
rect 205260 199 205325 269
rect 205359 204 205430 323
rect 203521 127 203855 161
rect 203984 127 204268 163
rect 204399 139 204865 173
rect 205464 165 205511 363
rect 205545 294 205603 527
rect 205643 435 205695 527
rect 205637 199 205695 394
rect 205729 342 205791 493
rect 205825 383 205901 527
rect 205945 342 205983 493
rect 206017 383 206093 527
rect 206139 459 206383 493
rect 206139 420 206191 459
rect 206225 342 206301 425
rect 205729 308 206301 342
rect 206345 339 206383 459
rect 206417 373 206493 527
rect 206537 339 206589 493
rect 203633 123 203855 127
rect 203523 17 203589 93
rect 203633 51 203667 123
rect 203711 17 203777 89
rect 203821 51 203855 123
rect 204399 93 204465 139
rect 203889 17 203972 93
rect 204020 51 204465 93
rect 204500 17 204563 105
rect 204597 51 204673 139
rect 204717 17 204755 105
rect 204789 51 204865 139
rect 204901 17 204959 162
rect 204995 123 205266 165
rect 204995 51 205056 123
rect 205090 17 205156 89
rect 205190 51 205266 123
rect 205321 51 205511 165
rect 205545 17 205603 162
rect 205729 134 205805 308
rect 206345 305 206589 339
rect 206649 294 206707 527
rect 206742 333 206801 527
rect 206925 455 207001 527
rect 207045 455 207481 493
rect 206845 421 206889 438
rect 207045 421 207081 455
rect 207527 439 207581 527
rect 207701 455 207777 527
rect 207890 455 207966 527
rect 208078 455 208155 527
rect 208355 455 208421 527
rect 206845 387 207081 421
rect 207115 405 207488 421
rect 207623 405 208420 421
rect 206845 372 206889 387
rect 207115 371 208420 405
rect 206927 303 207530 337
rect 205863 215 206062 273
rect 206154 215 206347 271
rect 206927 266 207036 303
rect 206381 215 206603 259
rect 206804 215 207036 266
rect 207095 215 207430 269
rect 205849 93 205887 178
rect 205921 127 206479 169
rect 206513 153 206603 215
rect 207464 199 207530 303
rect 207666 303 208284 337
rect 207666 282 207829 303
rect 207564 199 207829 282
rect 207918 215 208152 269
rect 208240 199 208284 303
rect 208320 268 208420 371
rect 208489 294 208547 527
rect 206441 103 206479 127
rect 205849 89 206093 93
rect 205639 51 206093 89
rect 206139 17 206205 89
rect 206325 17 206401 89
rect 206513 17 206594 89
rect 206649 17 206707 162
rect 206755 159 207420 181
rect 208320 165 208356 268
rect 206755 125 207571 159
rect 207605 127 208098 163
rect 208177 131 208356 165
rect 208581 206 208637 493
rect 208671 372 208817 527
rect 208860 338 208926 493
rect 208684 295 208926 338
rect 206755 107 206795 125
rect 206829 17 206905 89
rect 206949 85 206992 125
rect 207525 91 207571 125
rect 207031 17 207097 91
rect 207213 17 207289 89
rect 207405 17 207481 89
rect 207525 51 207818 91
rect 208177 90 208221 131
rect 208388 96 208422 119
rect 207890 54 208221 90
rect 208270 62 208422 96
rect 208489 17 208547 162
rect 208581 51 208649 206
rect 208684 181 208741 295
rect 208775 215 208875 261
rect 208961 255 208995 478
rect 209040 383 209184 527
rect 208909 215 208995 255
rect 209029 215 209099 323
rect 209225 294 209283 527
rect 209318 327 209369 527
rect 208684 143 208841 181
rect 208687 17 208721 109
rect 208769 51 208841 143
rect 208875 143 209106 181
rect 208875 111 208917 143
rect 208960 17 208994 109
rect 209040 51 209106 143
rect 209225 17 209283 162
rect 209321 17 209369 177
rect 209406 51 209465 493
rect 209499 437 209679 527
rect 209723 401 209775 493
rect 209537 357 209775 401
rect 209537 266 209571 357
rect 209499 168 209571 266
rect 209605 202 209691 323
rect 209860 280 209915 397
rect 209949 330 210006 527
rect 210053 294 210111 527
rect 210211 374 210287 527
rect 210331 340 210369 493
rect 210403 374 210479 527
rect 210523 340 210559 493
rect 210595 451 210675 527
rect 210719 421 210767 493
rect 210831 455 210897 527
rect 211027 421 211103 489
rect 210719 417 211103 421
rect 210146 306 210559 340
rect 210593 375 211103 417
rect 211219 387 211301 527
rect 210593 366 210767 375
rect 209764 205 209915 280
rect 209955 199 210007 290
rect 209499 127 209679 168
rect 209499 17 209575 93
rect 209613 51 209679 127
rect 209723 127 210006 165
rect 209723 93 209765 127
rect 209951 99 210006 127
rect 209799 17 209907 93
rect 210053 17 210111 162
rect 210146 161 210198 306
rect 210593 267 210641 366
rect 210232 199 210641 267
rect 210675 215 210825 323
rect 210880 299 211304 341
rect 210591 174 210641 199
rect 210880 198 210951 299
rect 211012 199 211142 265
rect 211210 199 211304 299
rect 211341 294 211399 527
rect 211434 299 211498 527
rect 211532 265 211583 475
rect 211617 301 211699 493
rect 211745 367 211838 527
rect 211445 199 211498 265
rect 211532 199 211631 265
rect 211665 225 211699 301
rect 211747 259 211859 331
rect 211893 294 211951 527
rect 211989 357 212055 527
rect 212099 459 212341 493
rect 212099 357 212143 459
rect 212303 427 212341 459
rect 212380 435 212456 527
rect 212187 393 212247 425
rect 212507 393 212590 493
rect 212187 357 212590 393
rect 211992 289 212427 323
rect 211665 191 211838 225
rect 211992 211 212058 289
rect 212102 215 212282 255
rect 212318 215 212427 289
rect 210146 127 210501 161
rect 210591 131 210805 174
rect 210257 123 210501 127
rect 210839 123 211295 157
rect 210839 97 210905 123
rect 210147 17 210213 93
rect 210339 17 210405 89
rect 210531 17 210597 93
rect 210645 51 210905 97
rect 210939 17 211007 89
rect 211123 17 211199 89
rect 211341 17 211399 162
rect 211434 123 211697 157
rect 211434 53 211492 123
rect 211541 17 211617 89
rect 211651 62 211697 123
rect 211745 55 211838 191
rect 211893 17 211951 162
rect 211989 143 212461 177
rect 211989 51 212055 143
rect 212101 17 212135 109
rect 212171 51 212247 143
rect 212303 17 212337 109
rect 212395 85 212461 143
rect 212507 119 212590 357
rect 212624 314 212674 527
rect 212721 294 212779 527
rect 212820 364 212877 527
rect 212921 417 212968 493
rect 213002 451 213078 527
rect 213122 455 213558 493
rect 213122 417 213160 455
rect 213602 439 213658 527
rect 212921 383 213160 417
rect 213702 417 213744 493
rect 213778 451 213854 527
rect 213898 417 213936 493
rect 213702 405 213936 417
rect 213194 371 213936 405
rect 213970 376 214046 527
rect 213663 340 213936 371
rect 212921 303 213615 337
rect 212624 153 212682 280
rect 212921 264 213121 303
rect 212821 203 213121 264
rect 213233 214 213521 269
rect 213555 198 213615 303
rect 213663 289 214062 340
rect 214101 294 214159 527
rect 214193 296 214261 493
rect 214295 441 214377 527
rect 214530 443 214596 527
rect 214632 407 214693 493
rect 214305 373 214693 407
rect 213657 203 213916 255
rect 213980 169 214062 289
rect 212624 85 212674 119
rect 212395 51 212674 85
rect 212721 17 212779 162
rect 212820 123 213648 164
rect 213682 123 214062 169
rect 214193 165 214244 296
rect 214305 265 214348 373
rect 214391 305 214520 339
rect 214278 199 214348 265
rect 214382 199 214452 265
rect 214486 165 214520 305
rect 213602 89 213648 123
rect 212906 17 212982 89
rect 213098 17 213174 89
rect 213290 17 213366 89
rect 213482 17 213558 89
rect 213602 51 214046 89
rect 214101 17 214159 162
rect 214193 90 214265 165
rect 214311 17 214345 165
rect 214418 131 214520 165
rect 214554 291 214693 373
rect 214810 307 214886 527
rect 214929 294 214987 527
rect 215108 441 215196 527
rect 215308 441 215480 527
rect 215524 407 215589 493
rect 215021 373 215421 407
rect 215021 299 215083 373
rect 214418 90 214452 131
rect 214554 51 214588 291
rect 214622 215 214746 257
rect 214780 215 214890 257
rect 214632 147 214889 181
rect 215021 165 215055 299
rect 215125 265 215169 339
rect 215089 199 215169 265
rect 215203 299 215295 339
rect 214632 51 214698 147
rect 214742 17 214776 111
rect 214823 54 214889 147
rect 214929 17 214987 162
rect 215021 86 215073 165
rect 215133 17 215169 165
rect 215203 93 215251 299
rect 215285 165 215319 265
rect 215387 199 215421 373
rect 215455 291 215589 407
rect 215694 375 215770 527
rect 215455 165 215498 291
rect 215533 215 215640 257
rect 215674 215 215783 325
rect 215849 294 215907 527
rect 215941 409 216011 493
rect 216051 443 216127 527
rect 216239 443 216315 527
rect 216427 443 216503 527
rect 215941 375 216487 409
rect 215941 291 216011 375
rect 215285 131 215498 165
rect 215203 59 215280 93
rect 215316 17 215389 93
rect 215432 51 215498 131
rect 215543 147 215782 181
rect 215941 171 215975 291
rect 216045 257 216111 341
rect 216009 215 216111 257
rect 216155 289 216409 341
rect 216453 323 216487 375
rect 216547 393 216581 493
rect 216634 427 216684 527
rect 216731 459 216977 493
rect 216731 427 216789 459
rect 216841 393 216890 425
rect 216547 359 216890 393
rect 216453 289 216565 323
rect 216155 182 216265 289
rect 216299 216 216487 250
rect 215543 73 215593 147
rect 215637 17 215671 111
rect 215715 54 215782 147
rect 215849 17 215907 162
rect 215941 53 216033 171
rect 216077 17 216111 181
rect 216155 145 216399 182
rect 216155 51 216221 145
rect 216265 17 216299 111
rect 216333 51 216399 145
rect 216453 179 216487 216
rect 216521 249 216565 289
rect 216521 215 216611 249
rect 216673 179 216711 359
rect 216841 289 216890 359
rect 216943 333 216977 459
rect 217011 367 217087 527
rect 217131 333 217186 493
rect 216943 291 217186 333
rect 217229 294 217287 527
rect 217321 269 217375 489
rect 217409 341 217474 442
rect 217518 375 217584 527
rect 217409 307 217517 341
rect 217631 325 217735 493
rect 216760 215 216988 255
rect 217032 215 217195 255
rect 217321 199 217411 269
rect 217458 199 217517 307
rect 217551 289 217735 325
rect 217798 307 217916 527
rect 217965 294 218023 527
rect 218076 333 218110 383
rect 218167 375 218233 527
rect 218076 299 218223 333
rect 216453 129 216711 179
rect 216755 145 217186 181
rect 217458 165 217492 199
rect 216755 95 216805 145
rect 216437 17 216503 95
rect 216545 51 216805 95
rect 216849 17 216883 111
rect 216917 51 216993 145
rect 217037 17 217071 111
rect 217105 53 217186 145
rect 217229 17 217287 162
rect 217321 17 217376 165
rect 217439 99 217492 165
rect 217551 51 217595 289
rect 217639 215 217743 255
rect 217777 215 217889 257
rect 218057 199 218136 265
rect 218170 249 218223 299
rect 218277 323 218311 493
rect 218364 359 218414 527
rect 218461 459 218707 493
rect 218461 359 218527 459
rect 218571 323 218620 425
rect 218277 289 218620 323
rect 218673 333 218707 459
rect 218741 367 218817 527
rect 218861 333 218916 493
rect 218673 291 218916 333
rect 218977 294 219035 527
rect 219081 325 219147 487
rect 219191 359 219225 527
rect 219259 325 219327 493
rect 219371 359 219421 527
rect 219465 325 219515 493
rect 219559 359 219609 527
rect 219657 459 220099 493
rect 219657 359 219723 459
rect 219767 325 219817 425
rect 219861 359 219911 459
rect 219955 325 220005 425
rect 219081 291 219222 325
rect 219259 291 220005 325
rect 220049 325 220099 459
rect 220143 359 220193 527
rect 220237 325 220287 493
rect 220331 359 220381 527
rect 220425 325 220475 493
rect 220049 291 220475 325
rect 220541 294 220599 527
rect 220633 344 220689 493
rect 220728 417 220788 527
rect 220916 409 221087 493
rect 220822 375 221165 409
rect 220822 344 220863 375
rect 220633 299 220863 344
rect 220633 291 220767 299
rect 218170 215 218308 249
rect 217632 147 217887 181
rect 217632 51 217698 147
rect 217743 17 217777 111
rect 217811 54 217887 147
rect 217965 17 218023 162
rect 218076 17 218110 165
rect 218170 89 218204 215
rect 218252 95 218308 181
rect 218342 129 218441 289
rect 219188 257 219222 291
rect 219591 289 220005 291
rect 218475 215 218718 255
rect 218762 215 218931 255
rect 219069 215 219154 257
rect 219188 215 219557 257
rect 219591 215 219691 289
rect 219725 215 220047 255
rect 220081 215 220502 257
rect 218485 145 218916 181
rect 219188 179 219241 215
rect 218485 95 218535 145
rect 218252 51 218535 95
rect 218579 17 218613 111
rect 218647 51 218723 145
rect 218767 17 218801 111
rect 218835 53 218916 145
rect 218977 17 219035 162
rect 219097 17 219131 179
rect 219165 58 219241 179
rect 219591 163 219637 215
rect 220633 199 220699 257
rect 219356 129 219637 163
rect 219681 145 220483 181
rect 220733 165 220767 291
rect 220801 197 220863 265
rect 220897 197 220974 341
rect 221012 251 221079 341
rect 221131 325 221165 375
rect 221199 359 221275 527
rect 221309 375 221422 493
rect 221131 291 221325 325
rect 221012 197 221139 251
rect 221179 215 221245 257
rect 221291 199 221325 291
rect 221359 165 221422 375
rect 221461 294 221519 527
rect 221586 334 221652 493
rect 221696 370 221738 527
rect 221876 409 222027 493
rect 221772 375 222129 409
rect 221772 334 221806 375
rect 221586 299 221806 334
rect 221645 289 221806 299
rect 221553 195 221605 265
rect 219681 95 219731 145
rect 219288 61 219731 95
rect 219775 17 219809 111
rect 219843 51 219919 145
rect 219963 17 219997 111
rect 220031 51 220107 145
rect 220151 17 220185 111
rect 220219 51 220295 145
rect 220339 17 220373 111
rect 220407 51 220483 145
rect 220541 17 220599 162
rect 220650 129 220767 165
rect 220823 129 221203 163
rect 220650 51 220716 129
rect 220756 61 220997 95
rect 221033 17 221101 95
rect 221137 54 221203 129
rect 221237 17 221271 128
rect 221305 53 221422 165
rect 221461 17 221519 162
rect 221645 161 221689 289
rect 221723 215 221802 255
rect 221840 215 221917 341
rect 221983 215 222059 341
rect 222095 325 222129 375
rect 222165 359 222211 527
rect 222245 409 222305 493
rect 222339 443 222417 527
rect 222245 375 222434 409
rect 222095 291 222279 325
rect 222235 257 222279 291
rect 222103 215 222201 257
rect 222235 215 222311 257
rect 222372 181 222434 375
rect 222473 294 222531 527
rect 222577 291 222627 527
rect 222671 391 222721 493
rect 222765 425 222815 527
rect 222859 459 223097 493
rect 222859 425 222909 459
rect 223047 425 223097 459
rect 223141 425 223293 527
rect 223337 459 223575 493
rect 223337 425 223387 459
rect 223525 425 223575 459
rect 223619 425 223669 527
rect 223721 391 223763 493
rect 223807 425 223857 527
rect 222671 357 223677 391
rect 223721 357 223848 391
rect 222566 215 222636 255
rect 221570 127 221689 161
rect 221763 147 222133 181
rect 221763 129 221850 147
rect 221570 51 221636 127
rect 221670 59 221937 93
rect 221989 17 222023 111
rect 222057 54 222133 147
rect 222177 17 222211 181
rect 222245 147 222434 181
rect 222245 53 222321 147
rect 222365 17 222399 113
rect 222473 17 222531 162
rect 222565 95 222617 179
rect 222671 173 222727 357
rect 223643 323 223677 357
rect 223814 323 223848 357
rect 223901 323 223951 493
rect 223995 359 224045 527
rect 222761 289 223157 323
rect 222761 215 222894 289
rect 222938 215 223047 255
rect 223081 215 223157 289
rect 223209 289 223593 323
rect 223643 289 223733 323
rect 223814 289 224090 323
rect 224129 294 224187 527
rect 224221 341 224277 493
rect 224324 375 224520 527
rect 224584 436 224705 493
rect 224584 341 224697 436
rect 224221 299 224697 341
rect 224775 323 224829 481
rect 223209 215 223339 289
rect 223543 255 223593 289
rect 223689 255 223733 289
rect 223373 215 223499 255
rect 223543 215 223655 255
rect 223689 215 223959 255
rect 224021 181 224090 289
rect 224221 199 224297 265
rect 222651 129 222727 173
rect 222771 95 222805 181
rect 222839 145 223583 181
rect 222839 129 223395 145
rect 222565 51 223199 95
rect 223235 17 223301 93
rect 223345 51 223395 129
rect 223439 17 223473 111
rect 223507 51 223583 145
rect 223627 17 223661 181
rect 223695 147 224090 181
rect 224339 165 224373 299
rect 224731 289 224829 323
rect 224867 291 224919 527
rect 224957 294 225015 527
rect 225060 291 225110 527
rect 225154 391 225204 493
rect 225248 425 225402 527
rect 225446 459 225684 493
rect 225446 425 225496 459
rect 225634 425 225684 459
rect 225728 425 225794 527
rect 225838 459 226076 493
rect 225838 425 225888 459
rect 225540 391 225590 425
rect 225932 391 225982 425
rect 225154 357 225982 391
rect 226026 357 226076 459
rect 225154 289 225212 357
rect 224407 199 224523 265
rect 224567 199 224669 265
rect 224731 249 224783 289
rect 224705 215 224783 249
rect 224817 215 224919 255
rect 225049 215 225119 255
rect 224693 165 224919 173
rect 223695 145 223959 147
rect 223695 51 223771 145
rect 223815 17 223849 111
rect 223883 51 223959 145
rect 224003 17 224054 113
rect 224129 17 224187 162
rect 224221 129 224373 165
rect 224454 139 224919 165
rect 224454 129 224716 139
rect 224221 73 224273 129
rect 224307 61 224617 95
rect 224661 56 224716 129
rect 224773 17 224807 105
rect 224841 56 224919 139
rect 224957 17 225015 162
rect 225052 95 225102 179
rect 225163 173 225212 289
rect 225256 289 225744 323
rect 225256 215 225469 289
rect 225503 215 225634 255
rect 225668 215 225744 289
rect 225778 289 226085 323
rect 226129 291 226170 527
rect 226245 294 226303 527
rect 226351 297 226401 527
rect 226445 323 226495 493
rect 226539 365 226589 527
rect 226633 391 226683 493
rect 226727 425 226881 527
rect 226925 391 226975 493
rect 227019 425 227069 527
rect 227113 453 227547 493
rect 227113 391 227155 453
rect 227591 435 227641 527
rect 227675 453 228119 493
rect 226633 323 226785 391
rect 226925 357 227155 391
rect 227189 357 228033 401
rect 228077 391 228119 453
rect 228163 425 228213 527
rect 228257 391 228307 493
rect 228077 357 228307 391
rect 227189 323 227233 357
rect 226445 289 227233 323
rect 227267 289 227599 323
rect 225778 215 225854 289
rect 226051 255 226085 289
rect 225888 215 226007 255
rect 226051 215 226199 255
rect 226338 215 226700 255
rect 225136 129 225212 173
rect 225256 129 225692 181
rect 225736 147 226178 181
rect 225256 95 225306 129
rect 225736 95 225802 147
rect 225914 145 226178 147
rect 225052 51 225306 95
rect 225344 51 225802 95
rect 225846 17 225880 111
rect 225914 51 225990 145
rect 226034 17 226068 111
rect 226102 51 226178 145
rect 226245 17 226303 162
rect 226343 95 226393 179
rect 226744 173 226785 289
rect 227267 255 227305 289
rect 226832 215 227305 255
rect 227339 199 227487 255
rect 227523 215 227599 289
rect 227633 289 228184 323
rect 228257 289 228307 357
rect 228351 289 228401 527
rect 228453 294 228511 527
rect 227633 215 227709 289
rect 228121 255 228184 289
rect 227745 215 228067 255
rect 228121 215 228347 255
rect 226427 129 226785 173
rect 227523 164 228409 181
rect 226823 147 228409 164
rect 226823 129 227657 147
rect 226343 51 227547 95
rect 227591 51 227657 129
rect 227769 145 228033 147
rect 227701 17 227735 111
rect 227769 51 227845 145
rect 227889 17 227923 111
rect 227957 51 228033 145
rect 228145 145 228409 147
rect 228077 17 228111 111
rect 228145 51 228221 145
rect 228265 17 228299 111
rect 228333 51 228409 145
rect 228453 17 228511 162
rect 228545 73 228601 493
rect 228649 375 228800 527
rect 228889 341 228983 493
rect 228635 299 228983 341
rect 228635 179 228700 299
rect 229017 265 229061 481
rect 229125 291 229236 527
rect 229281 294 229339 527
rect 229379 289 229429 527
rect 228741 215 228835 265
rect 228874 215 228959 265
rect 228995 215 229061 265
rect 229095 215 229190 255
rect 228635 143 228889 179
rect 228816 129 228889 143
rect 228941 139 229199 173
rect 228651 17 228685 109
rect 228941 95 229007 139
rect 228739 59 229007 95
rect 229053 17 229087 105
rect 229121 56 229199 139
rect 229281 17 229339 162
rect 229393 17 229427 177
rect 229477 73 229527 493
rect 229575 375 229735 527
rect 229824 341 229895 493
rect 229571 291 229895 341
rect 229571 179 229627 291
rect 229937 255 229991 481
rect 230070 359 230134 527
rect 229661 215 229734 255
rect 229778 215 229881 255
rect 229915 215 229991 255
rect 230025 215 230097 323
rect 230201 294 230259 527
rect 230320 365 230370 527
rect 230414 323 230464 493
rect 230508 359 230558 527
rect 230602 323 230652 493
rect 230696 425 230850 527
rect 230894 459 231132 493
rect 230894 425 230944 459
rect 231082 425 231132 459
rect 231176 425 231242 527
rect 231286 459 231524 493
rect 231286 425 231336 459
rect 230988 391 231038 425
rect 231380 391 231430 425
rect 230293 289 230652 323
rect 230696 357 231430 391
rect 231474 357 231524 459
rect 230293 181 230350 289
rect 230696 255 230762 357
rect 230384 215 230762 255
rect 230800 289 231184 323
rect 230800 215 230912 289
rect 230946 215 231082 255
rect 231116 215 231184 289
rect 231218 289 231533 323
rect 231577 291 231618 527
rect 231673 294 231731 527
rect 231775 435 231817 527
rect 231974 409 232084 493
rect 231218 215 231302 289
rect 231491 255 231533 289
rect 231346 215 231457 255
rect 231491 215 231639 255
rect 230704 181 230762 215
rect 229571 143 229829 179
rect 229746 129 229829 143
rect 229874 139 230134 173
rect 229581 17 229617 109
rect 229874 95 229942 139
rect 229669 59 229942 95
rect 229995 17 230029 105
rect 230067 56 230134 139
rect 230201 17 230259 162
rect 230293 145 230660 181
rect 230704 147 231140 181
rect 230328 17 230362 111
rect 230396 53 230472 145
rect 230516 17 230550 111
rect 230584 51 230660 145
rect 230799 129 231140 147
rect 231184 147 231626 181
rect 230704 17 230738 111
rect 231184 95 231250 147
rect 231362 145 231626 147
rect 230792 51 231250 95
rect 231294 17 231328 111
rect 231362 51 231438 145
rect 231482 17 231516 111
rect 231550 51 231626 145
rect 231673 17 231731 162
rect 231765 133 231813 398
rect 231847 367 232084 409
rect 231847 165 231906 367
rect 231958 199 232018 333
rect 232132 323 232182 481
rect 232098 289 232182 323
rect 232216 291 232280 527
rect 232317 294 232375 527
rect 232422 325 232473 493
rect 232517 359 232567 527
rect 232611 459 232849 493
rect 232611 325 232661 459
rect 232422 291 232661 325
rect 232705 325 232755 425
rect 232799 359 232849 459
rect 232911 459 233149 493
rect 232911 359 232961 459
rect 233005 325 233055 425
rect 232705 289 233055 325
rect 233099 325 233149 459
rect 233193 359 233243 527
rect 233287 325 233338 493
rect 233099 291 233338 325
rect 233421 294 233479 527
rect 233529 289 233579 527
rect 233623 391 233673 493
rect 233717 425 233767 527
rect 233811 459 234245 493
rect 233811 391 233853 459
rect 233999 425 234049 459
rect 234187 425 234245 459
rect 234289 425 234333 527
rect 234367 425 234438 493
rect 234481 425 234529 527
rect 234573 459 234999 493
rect 233623 357 233853 391
rect 233887 391 233955 425
rect 234093 391 234143 425
rect 234404 391 234438 425
rect 234573 391 234623 459
rect 234761 425 234811 459
rect 234949 427 234999 459
rect 235043 425 235099 527
rect 233887 357 234370 391
rect 234404 357 234623 391
rect 234667 391 234717 425
rect 234855 391 234905 425
rect 234667 357 235130 391
rect 233623 289 233673 357
rect 234336 323 234370 357
rect 233746 289 234302 323
rect 234336 289 234411 323
rect 232098 249 232144 289
rect 232061 215 232144 249
rect 232178 215 232280 255
rect 232432 215 232615 257
rect 232657 215 232817 255
rect 232873 181 232921 289
rect 232959 215 233103 255
rect 233145 215 233305 257
rect 233746 255 233809 289
rect 233513 215 233809 255
rect 233863 215 234185 255
rect 234221 215 234302 289
rect 232040 165 232280 173
rect 231847 129 231927 165
rect 232006 139 232280 165
rect 232006 95 232072 139
rect 231765 59 232072 95
rect 232126 17 232160 105
rect 232202 56 232280 139
rect 232317 17 232375 162
rect 232410 95 232465 181
rect 232499 129 232921 181
rect 232955 145 233345 181
rect 232955 95 232989 145
rect 232410 61 232989 95
rect 233023 17 233057 111
rect 233091 51 233157 145
rect 233201 17 233235 111
rect 233269 51 233345 145
rect 233421 17 233479 162
rect 233521 147 234333 181
rect 233521 145 233775 147
rect 233521 51 233587 145
rect 233631 17 233665 111
rect 233699 51 233775 145
rect 233887 145 234151 147
rect 233819 17 233853 111
rect 233887 51 233963 145
rect 234007 17 234041 111
rect 234075 51 234151 145
rect 234195 17 234229 111
rect 234263 95 234333 147
rect 234367 164 234411 289
rect 234445 289 235043 323
rect 234445 199 234594 289
rect 234628 215 234928 255
rect 234989 199 235043 289
rect 235077 164 235130 357
rect 235169 294 235227 527
rect 235261 359 235313 493
rect 235347 447 235423 527
rect 235617 447 235697 527
rect 235755 411 235831 458
rect 235385 377 235831 411
rect 234367 129 235130 164
rect 235261 165 235296 359
rect 235385 323 235419 377
rect 235330 289 235419 323
rect 235453 299 235676 343
rect 235330 199 235374 289
rect 235621 271 235676 299
rect 235710 299 235831 377
rect 235408 215 235508 255
rect 235542 181 235587 220
rect 234263 51 235105 95
rect 235169 17 235227 162
rect 235261 51 235329 165
rect 235378 17 235412 150
rect 235447 147 235587 181
rect 235447 76 235504 147
rect 235621 113 235655 271
rect 235710 249 235744 299
rect 235911 265 235951 485
rect 235985 363 236055 527
rect 235705 215 235744 249
rect 235788 215 235951 265
rect 235985 215 236055 329
rect 236089 294 236147 527
rect 236186 282 236237 527
rect 236271 359 236332 493
rect 236366 447 236442 527
rect 236636 447 236717 527
rect 236771 411 236851 485
rect 236404 377 236851 411
rect 235705 138 235739 215
rect 235556 79 235655 113
rect 235689 64 235739 138
rect 235783 145 236055 181
rect 235783 64 235833 145
rect 235871 17 235941 111
rect 235977 64 236055 145
rect 236089 17 236147 162
rect 236186 17 236237 182
rect 236271 165 236315 359
rect 236404 323 236438 377
rect 236349 289 236438 323
rect 236472 299 236696 343
rect 236349 199 236393 289
rect 236643 271 236696 299
rect 236730 299 236851 377
rect 236895 383 236963 485
rect 236427 215 236531 255
rect 236565 181 236609 220
rect 236271 51 236348 165
rect 236391 17 236425 150
rect 236468 147 236609 181
rect 236468 76 236541 147
rect 236643 113 236677 271
rect 236730 249 236764 299
rect 236895 265 236929 383
rect 236997 363 237060 527
rect 236726 215 236764 249
rect 236808 215 236929 265
rect 236964 215 237057 329
rect 237101 294 237159 527
rect 237204 359 237245 527
rect 237297 459 237535 493
rect 237297 357 237347 459
rect 237485 425 237535 459
rect 237579 425 237629 527
rect 237391 391 237441 425
rect 237673 393 237731 493
rect 237775 427 237921 527
rect 238059 427 238109 527
rect 237965 393 238015 425
rect 238153 393 238203 493
rect 237673 391 237749 393
rect 237391 357 237749 391
rect 237193 289 237595 323
rect 237193 215 237301 289
rect 237347 215 237465 255
rect 237519 215 237595 289
rect 237629 283 237749 357
rect 237827 357 238203 393
rect 238247 359 238297 527
rect 238341 391 238391 493
rect 238435 433 238485 527
rect 238529 391 238579 493
rect 238341 357 238579 391
rect 238623 365 238673 527
rect 237629 215 237715 283
rect 237827 249 237865 357
rect 238529 331 238579 357
rect 237749 215 237865 249
rect 237899 289 238269 323
rect 237899 215 237975 289
rect 238009 215 238153 255
rect 238187 215 238269 289
rect 238309 249 238377 323
rect 238529 283 238718 331
rect 238757 294 238815 527
rect 238862 291 238912 527
rect 238956 333 239006 493
rect 239050 367 239188 527
rect 239222 333 239287 493
rect 238956 299 239120 333
rect 238309 215 238593 249
rect 236726 138 236760 215
rect 236575 79 236677 113
rect 236711 64 236760 138
rect 236805 145 237045 181
rect 236805 64 236851 145
rect 236899 17 236933 111
rect 236967 64 237045 145
rect 237101 17 237159 162
rect 237195 147 237621 181
rect 237195 145 237449 147
rect 237195 51 237261 145
rect 237305 17 237339 111
rect 237373 51 237449 145
rect 237493 17 237527 111
rect 237561 95 237621 147
rect 237655 163 237715 215
rect 237827 181 237865 215
rect 238657 181 238718 283
rect 239086 265 239120 299
rect 239184 289 239287 333
rect 238849 197 238919 257
rect 238953 199 239052 265
rect 239086 199 239148 265
rect 237655 129 237731 163
rect 237827 145 238117 181
rect 238041 129 238117 145
rect 237561 51 237825 95
rect 237879 17 237913 111
rect 238161 95 238211 179
rect 237947 61 238211 95
rect 238255 17 238289 179
rect 238323 145 238718 181
rect 238323 55 238399 145
rect 238443 17 238477 111
rect 238511 55 238587 145
rect 238631 17 238665 111
rect 238757 17 238815 162
rect 238850 17 238917 163
rect 238953 56 238997 199
rect 239086 165 239120 199
rect 239032 56 239120 165
rect 239184 158 239218 289
rect 239321 255 239355 485
rect 239422 291 239472 527
rect 239585 294 239643 527
rect 239690 359 239740 527
rect 239785 393 239835 493
rect 239879 427 239929 527
rect 240067 427 240205 527
rect 239785 357 240157 393
rect 239678 289 240089 323
rect 239262 215 239355 255
rect 239405 215 239481 257
rect 239678 215 239795 289
rect 239829 215 239960 255
rect 240013 215 240089 289
rect 240123 265 240157 357
rect 240239 391 240307 493
rect 240351 425 240408 527
rect 240452 459 240690 493
rect 240452 425 240502 459
rect 240546 391 240596 425
rect 240239 357 240596 391
rect 240640 357 240690 459
rect 240743 359 240784 527
rect 240123 199 240205 265
rect 240239 215 240353 357
rect 240390 289 240752 323
rect 240873 294 240931 527
rect 240979 359 241029 527
rect 241073 325 241123 493
rect 241167 359 241217 527
rect 241261 325 241311 493
rect 241355 359 241405 527
rect 241449 325 241499 493
rect 241543 359 241593 527
rect 241637 325 241687 493
rect 241731 359 241879 527
rect 241923 325 241973 493
rect 242017 359 242067 527
rect 242111 325 242161 493
rect 242205 359 242255 527
rect 242303 459 242735 493
rect 242303 359 242359 459
rect 242403 325 242453 425
rect 242497 359 242547 459
rect 242591 325 242641 425
rect 240390 215 240468 289
rect 240512 215 240640 255
rect 240686 215 240752 289
rect 240965 291 241811 325
rect 241923 291 242641 325
rect 242685 325 242735 459
rect 242779 359 242829 527
rect 242873 325 242923 493
rect 242967 359 243017 527
rect 243061 325 243123 493
rect 242685 291 243123 325
rect 243173 294 243231 527
rect 243265 299 243332 527
rect 240123 181 240157 199
rect 239154 86 239218 158
rect 239252 145 239480 181
rect 239252 85 239302 145
rect 239336 17 239370 111
rect 239404 55 239480 145
rect 239585 17 239643 162
rect 239699 17 239733 179
rect 239767 95 239827 179
rect 239861 145 240157 181
rect 239861 129 239937 145
rect 240239 129 240315 215
rect 240965 181 240999 291
rect 241777 257 241811 291
rect 241033 215 241353 257
rect 241407 215 241729 257
rect 241777 215 242209 257
rect 242243 181 242309 291
rect 242361 215 242683 257
rect 242717 215 243136 257
rect 243266 215 243335 265
rect 243369 215 243469 493
rect 243539 265 243587 481
rect 243511 215 243587 265
rect 240359 147 240792 181
rect 239767 61 240031 95
rect 240067 17 240101 111
rect 240155 95 240205 111
rect 240359 95 240416 147
rect 240528 145 240792 147
rect 240155 51 240416 95
rect 240460 17 240494 111
rect 240528 51 240604 145
rect 240648 17 240682 111
rect 240716 51 240792 145
rect 240873 17 240931 162
rect 240965 129 241319 181
rect 241363 145 241789 181
rect 241363 95 241413 145
rect 240968 51 241413 95
rect 241457 17 241491 111
rect 241525 51 241601 145
rect 241645 17 241679 111
rect 241713 51 241789 145
rect 241840 95 241877 167
rect 241921 129 242309 181
rect 242343 147 243119 181
rect 242343 95 242377 147
rect 242479 145 243119 147
rect 241840 51 242377 95
rect 242411 17 242445 111
rect 242479 51 242555 145
rect 242599 17 242633 111
rect 242667 51 242743 145
rect 242787 17 242821 111
rect 242855 51 242931 145
rect 242975 17 243009 111
rect 243043 51 243119 145
rect 243173 17 243231 162
rect 243283 17 243317 181
rect 243351 147 243591 181
rect 243351 51 243427 147
rect 243473 17 243507 113
rect 243541 92 243591 147
rect 243625 165 243679 493
rect 243719 299 243753 527
rect 243817 294 243875 527
rect 243910 333 243981 493
rect 244025 367 244059 527
rect 244093 333 244169 493
rect 244213 459 244553 493
rect 244213 367 244247 459
rect 244281 333 244357 425
rect 243910 299 244357 333
rect 244409 333 244475 425
rect 244519 367 244553 459
rect 244587 333 244663 493
rect 244707 367 244773 527
rect 244817 333 244885 493
rect 244409 299 244885 333
rect 243713 199 243778 265
rect 243910 211 244154 265
rect 244192 211 244376 265
rect 244432 211 244603 265
rect 243625 52 243747 165
rect 243817 17 243875 162
rect 243910 143 244663 177
rect 243910 51 243981 143
rect 244025 17 244059 109
rect 244093 51 244169 143
rect 244213 17 244325 109
rect 244377 51 244443 143
rect 244477 17 244553 109
rect 244587 85 244663 143
rect 244707 119 244783 299
rect 244921 294 244979 527
rect 245014 379 245085 493
rect 245129 413 245163 527
rect 245197 379 245273 493
rect 245317 413 245351 527
rect 245385 441 245853 493
rect 245385 379 245461 441
rect 245014 319 245461 379
rect 245505 353 245539 407
rect 245573 387 245649 441
rect 245902 407 246236 493
rect 245693 373 246236 407
rect 245693 353 245797 373
rect 245505 319 245797 353
rect 246280 339 246314 493
rect 246348 378 246424 527
rect 246468 339 246502 493
rect 246536 378 246612 527
rect 246656 339 246721 493
rect 245831 289 246721 339
rect 246761 294 246819 527
rect 246854 299 246908 527
rect 246942 357 247142 493
rect 244818 151 244886 265
rect 245014 211 245382 285
rect 245426 211 245797 285
rect 245831 211 246314 255
rect 246348 177 246395 289
rect 246429 211 246713 255
rect 244818 85 244885 117
rect 244587 51 244885 85
rect 244921 17 244979 162
rect 245014 143 246314 177
rect 245014 51 245085 143
rect 245129 17 245163 109
rect 245197 51 245273 143
rect 245317 17 245351 109
rect 245385 51 245461 143
rect 245505 17 245539 109
rect 245573 51 245649 143
rect 245693 17 245727 109
rect 245761 51 245837 143
rect 245885 17 246024 109
rect 246068 79 246102 143
rect 246154 17 246228 109
rect 246280 95 246314 143
rect 246348 129 246612 177
rect 246656 95 246713 177
rect 246280 51 246713 95
rect 246761 17 246819 162
rect 246854 137 246908 265
rect 246942 165 246986 357
rect 247020 199 247097 323
rect 247131 199 247185 323
rect 247219 199 247277 493
rect 247393 299 247463 527
rect 247497 294 247555 527
rect 247590 459 247845 493
rect 247590 299 247641 459
rect 247675 333 247751 419
rect 247795 401 247845 459
rect 247889 435 247923 527
rect 247957 401 248033 491
rect 247795 367 248033 401
rect 248089 451 248539 489
rect 248089 367 248139 451
rect 248177 333 248253 417
rect 247675 299 248253 333
rect 248297 299 248331 451
rect 248375 333 248441 417
rect 248489 367 248539 451
rect 248586 367 248627 527
rect 248671 333 248737 492
rect 248375 299 248737 333
rect 248781 299 248825 527
rect 247315 199 247434 265
rect 247590 215 247751 265
rect 247785 215 247935 265
rect 247969 221 248046 299
rect 248877 294 248935 527
rect 248970 451 249400 493
rect 248970 299 249021 451
rect 249055 333 249131 417
rect 249175 367 249209 451
rect 249243 333 249322 417
rect 249366 401 249400 451
rect 249434 435 249510 527
rect 249554 401 249588 485
rect 249622 435 249698 527
rect 249742 401 249792 493
rect 249366 367 249792 401
rect 249830 451 250648 493
rect 249830 367 249880 451
rect 249924 333 249990 417
rect 250034 367 250068 451
rect 250102 333 250178 417
rect 250222 367 250256 451
rect 249055 299 250178 333
rect 250290 333 250366 417
rect 250410 367 250444 451
rect 250478 333 250554 417
rect 250598 367 250648 451
rect 250686 367 250736 527
rect 250770 333 250846 493
rect 250890 367 250924 527
rect 250958 333 251034 493
rect 250290 299 251034 333
rect 251087 299 251137 527
rect 247969 181 248021 221
rect 248103 215 248245 265
rect 248316 215 248558 265
rect 248612 215 248831 265
rect 248974 215 249319 255
rect 249363 181 249399 299
rect 251177 294 251235 527
rect 251276 333 251354 368
rect 251471 367 251537 527
rect 251581 369 251695 493
rect 251276 299 251601 333
rect 249433 215 249740 255
rect 249786 215 250148 255
rect 250256 215 250554 255
rect 250770 215 251137 255
rect 246942 131 247015 165
rect 247049 131 247347 165
rect 247049 97 247124 131
rect 246853 51 247124 97
rect 247165 17 247231 97
rect 247313 75 247347 131
rect 247381 17 247455 165
rect 247497 17 247555 162
rect 247590 97 247641 181
rect 247675 131 248021 181
rect 248069 143 248833 181
rect 248069 97 248103 143
rect 247590 51 248103 97
rect 248146 17 248222 109
rect 248259 51 248335 143
rect 248379 17 248413 109
rect 248473 51 248607 143
rect 248643 17 248719 109
rect 248767 51 248833 143
rect 248877 17 248935 162
rect 248970 93 249021 181
rect 249055 131 249698 181
rect 249742 147 251137 181
rect 249742 93 249792 147
rect 248970 51 249792 93
rect 249836 17 249870 109
rect 249904 51 249980 147
rect 250024 17 250090 109
rect 250134 51 250268 147
rect 250316 17 250350 109
rect 250384 51 250460 147
rect 250504 17 250538 109
rect 250572 51 250720 147
rect 250796 17 250830 109
rect 250864 51 250940 147
rect 250984 17 251027 109
rect 251061 51 251137 147
rect 251177 17 251235 162
rect 251269 153 251340 265
rect 251374 119 251408 299
rect 251442 153 251509 265
rect 251557 199 251601 299
rect 251635 165 251695 369
rect 251729 294 251787 527
rect 251835 333 251907 368
rect 252044 367 252078 527
rect 252112 401 252188 493
rect 252232 435 252266 527
rect 252112 367 252287 401
rect 251835 299 252157 333
rect 251274 17 251322 119
rect 251374 53 251422 119
rect 251478 17 251521 119
rect 251555 51 251695 165
rect 251729 17 251787 162
rect 251829 153 251873 265
rect 251907 119 251953 299
rect 251987 153 252079 265
rect 252113 199 252157 299
rect 252191 165 252287 367
rect 252373 294 252431 527
rect 252479 333 252551 493
rect 252680 367 252714 527
rect 252766 401 252842 493
rect 252876 435 252910 527
rect 252954 401 253030 493
rect 252766 367 253030 401
rect 253064 367 253098 527
rect 252954 333 253030 367
rect 252479 299 252801 333
rect 252954 299 253082 333
rect 252138 131 252287 165
rect 251825 17 251873 119
rect 251907 51 251975 119
rect 252031 17 252094 119
rect 252138 77 252172 131
rect 252206 17 252282 97
rect 252373 17 252431 162
rect 252466 153 252517 265
rect 252551 165 252597 299
rect 252631 199 252716 265
rect 252750 249 252801 299
rect 252750 215 252972 249
rect 253013 181 253082 299
rect 253201 294 253259 527
rect 253294 299 253345 527
rect 253384 417 253643 483
rect 253405 265 253439 377
rect 253484 333 253568 383
rect 253689 367 253745 527
rect 253484 299 253753 333
rect 253797 299 253894 493
rect 253719 265 253753 299
rect 253294 215 253361 265
rect 253405 199 253553 265
rect 253719 199 253765 265
rect 253405 181 253455 199
rect 252469 17 252517 119
rect 252551 58 252627 165
rect 252680 17 252714 165
rect 252766 147 253082 181
rect 252766 53 252842 147
rect 252876 17 252910 113
rect 252954 53 253030 147
rect 253064 17 253098 113
rect 253201 17 253259 162
rect 253298 147 253455 181
rect 253719 165 253753 199
rect 253298 53 253360 147
rect 253595 131 253753 165
rect 253817 152 253894 299
rect 253937 294 253995 527
rect 254029 299 254081 527
rect 254120 417 254378 483
rect 254141 265 254175 377
rect 254219 333 254303 383
rect 254424 367 254480 527
rect 254219 299 254500 333
rect 254029 215 254097 265
rect 254141 199 254288 265
rect 254141 181 254190 199
rect 253404 17 253551 113
rect 253595 61 253629 131
rect 253663 17 253749 97
rect 253797 83 253894 152
rect 253937 17 253995 162
rect 254033 147 254190 181
rect 254466 165 254500 299
rect 254033 53 254096 147
rect 254330 131 254500 165
rect 254140 17 254286 113
rect 254330 61 254364 131
rect 254418 17 254484 97
rect 254570 83 254634 493
rect 254669 292 254716 527
rect 254765 294 254823 527
rect 254858 425 254909 527
rect 254858 215 254925 391
rect 254969 265 255003 493
rect 255048 323 255152 493
rect 255253 367 255309 527
rect 255353 391 255403 493
rect 255447 427 255497 527
rect 255541 391 255591 493
rect 255353 357 255591 391
rect 255635 359 255685 527
rect 255456 323 255591 357
rect 255048 299 255412 323
rect 255108 289 255412 299
rect 255456 289 255738 323
rect 255777 294 255835 527
rect 255869 425 256127 483
rect 255873 357 256127 391
rect 256171 367 256227 527
rect 255873 299 255938 357
rect 256093 333 256127 357
rect 254969 199 255074 265
rect 254669 17 254716 185
rect 254969 181 255019 199
rect 254765 17 254823 162
rect 254862 147 255019 181
rect 255108 181 255152 289
rect 255186 215 255334 255
rect 255378 249 255412 289
rect 255378 215 255600 249
rect 255661 181 255738 289
rect 255973 265 256021 323
rect 256093 299 256247 333
rect 256320 299 256375 493
rect 255869 199 255938 265
rect 255973 199 256150 265
rect 255108 147 255209 181
rect 254862 53 254924 147
rect 254968 17 255099 113
rect 255133 61 255209 147
rect 255266 17 255301 181
rect 255335 147 255738 181
rect 256213 165 256247 299
rect 255335 58 255411 147
rect 255455 17 255489 110
rect 255523 58 255599 147
rect 255643 17 255677 110
rect 255777 17 255835 162
rect 255872 131 256247 165
rect 256341 152 256375 299
rect 256421 294 256479 527
rect 256513 425 256772 483
rect 256517 357 256770 391
rect 256816 367 256910 527
rect 256517 299 256573 357
rect 256736 333 256770 357
rect 256607 265 256672 323
rect 256736 299 256918 333
rect 256962 299 257027 493
rect 256874 265 256918 299
rect 256513 199 256573 265
rect 256607 199 256812 265
rect 256874 199 256956 265
rect 256874 165 256918 199
rect 255872 61 255923 131
rect 255957 17 256033 97
rect 256077 61 256111 131
rect 256145 17 256231 97
rect 256320 83 256375 152
rect 256421 17 256479 162
rect 256517 131 256918 165
rect 256990 152 257027 299
rect 257061 286 257119 527
rect 257157 294 257215 527
rect 257249 459 257505 493
rect 257249 299 257317 459
rect 257351 265 257398 410
rect 257452 333 257505 459
rect 257549 367 257689 527
rect 257452 299 257680 333
rect 257249 215 257317 265
rect 257351 215 257463 265
rect 257497 215 257602 265
rect 257636 249 257680 299
rect 257741 323 257791 493
rect 257835 359 257885 527
rect 257929 323 257979 493
rect 258023 359 258073 527
rect 257741 289 258123 323
rect 258169 294 258227 527
rect 258261 299 258313 527
rect 258371 425 258714 491
rect 257636 215 258021 249
rect 256517 61 256568 131
rect 256602 17 256678 97
rect 256722 61 256756 131
rect 256790 17 256914 97
rect 256962 83 257027 152
rect 257061 17 257119 183
rect 257636 181 257680 215
rect 258055 181 258123 289
rect 258373 265 258407 377
rect 258459 357 258714 391
rect 258758 367 258814 527
rect 258459 299 258511 357
rect 258680 333 258714 357
rect 258549 265 258598 323
rect 258680 299 258822 333
rect 258866 299 258951 493
rect 258788 265 258822 299
rect 258262 215 258329 265
rect 258373 199 258498 265
rect 258549 199 258737 265
rect 258788 199 258843 265
rect 258373 181 258423 199
rect 257157 17 257215 162
rect 257249 145 257680 181
rect 257723 147 258123 181
rect 257249 51 257317 145
rect 257361 17 257395 111
rect 257429 51 257505 145
rect 257549 17 257689 111
rect 257723 53 257799 147
rect 257843 17 257877 111
rect 257911 53 257987 147
rect 258031 17 258065 111
rect 258169 17 258227 162
rect 258261 17 258313 181
rect 258347 97 258423 181
rect 258788 165 258822 199
rect 258459 131 258822 165
rect 258887 152 258951 299
rect 258997 294 259055 527
rect 259089 408 259141 444
rect 259192 442 259264 527
rect 259409 442 259475 527
rect 259511 425 259781 473
rect 259089 391 259468 408
rect 259089 374 259676 391
rect 259089 362 259235 374
rect 259089 215 259157 328
rect 259201 181 259235 362
rect 259434 357 259676 374
rect 258459 51 258511 131
rect 258545 17 258621 97
rect 258665 61 258699 131
rect 258733 17 258818 97
rect 258866 83 258951 152
rect 258997 17 259055 162
rect 259089 147 259235 181
rect 259269 299 259358 340
rect 259089 58 259141 147
rect 259269 119 259319 299
rect 259369 181 259403 265
rect 259463 215 259580 323
rect 259642 265 259676 357
rect 259720 299 259781 385
rect 259642 199 259712 265
rect 259369 165 259579 181
rect 259747 165 259781 299
rect 259825 294 259883 527
rect 259917 408 259969 444
rect 260020 442 260092 527
rect 260204 442 260280 527
rect 260391 442 260469 527
rect 260674 442 260791 485
rect 259917 374 260706 408
rect 259917 362 260063 374
rect 259917 215 259985 328
rect 260029 181 260063 362
rect 259369 147 259781 165
rect 259545 131 259781 147
rect 259201 17 259235 113
rect 259269 53 259349 119
rect 259445 17 259479 113
rect 259545 61 259579 131
rect 259620 17 259686 97
rect 259720 61 259781 131
rect 259825 17 259883 162
rect 259917 147 260063 181
rect 260102 283 260384 340
rect 260102 181 260154 283
rect 260188 215 260423 249
rect 260102 147 260348 181
rect 259917 58 259969 147
rect 260034 17 260068 113
rect 260102 57 260186 147
rect 260230 17 260264 113
rect 260301 51 260348 147
rect 260389 165 260423 215
rect 260460 199 260522 340
rect 260566 199 260614 340
rect 260672 199 260706 374
rect 260750 165 260791 442
rect 260837 294 260895 527
rect 260930 425 261291 483
rect 260930 357 261278 391
rect 261335 367 261391 527
rect 260930 299 260994 357
rect 261244 333 261278 357
rect 260389 131 260791 165
rect 260392 17 260468 97
rect 260580 17 260668 97
rect 260837 17 260895 162
rect 260930 151 261000 265
rect 261044 199 261183 323
rect 261244 299 261399 333
rect 261473 299 261527 493
rect 261365 265 261399 299
rect 261217 199 261331 265
rect 261365 199 261423 265
rect 261365 165 261399 199
rect 261047 131 261399 165
rect 261493 152 261527 299
rect 261573 294 261631 527
rect 261665 425 262027 483
rect 261665 357 262014 391
rect 262071 367 262127 527
rect 261665 299 261730 357
rect 261980 333 262014 357
rect 260931 17 260997 117
rect 261047 61 261081 131
rect 261121 17 261197 97
rect 261241 61 261275 131
rect 261309 17 261395 97
rect 261473 83 261527 152
rect 261573 17 261631 162
rect 261665 151 261735 265
rect 261769 199 261909 323
rect 261980 299 262135 333
rect 262212 299 262273 493
rect 262101 265 262135 299
rect 261943 199 262067 265
rect 262101 199 262188 265
rect 262101 165 262135 199
rect 261783 131 262135 165
rect 262226 152 262273 299
rect 262311 291 262355 527
rect 262401 294 262459 527
rect 262499 333 262566 490
rect 262499 299 262628 333
rect 261666 17 261733 117
rect 261783 61 261817 131
rect 261857 17 261933 97
rect 261977 61 262011 131
rect 262045 17 262131 97
rect 262212 83 262273 152
rect 262311 17 262355 200
rect 262401 17 262459 162
rect 262493 151 262550 265
rect 262584 165 262628 299
rect 262662 324 262742 475
rect 262776 357 262850 475
rect 262917 359 262967 527
rect 262662 199 262696 324
rect 262776 290 262828 357
rect 263022 325 263072 493
rect 263116 359 263166 527
rect 263210 325 263260 493
rect 263304 359 263354 527
rect 262752 199 262828 290
rect 262864 289 262971 323
rect 263022 291 263373 325
rect 263413 294 263471 527
rect 263505 312 263573 527
rect 263620 425 264060 483
rect 262864 199 262918 289
rect 262952 215 263274 249
rect 262952 165 262986 215
rect 263318 181 263373 291
rect 263617 265 263665 384
rect 263704 357 264060 391
rect 264104 367 264160 527
rect 263704 299 263768 357
rect 264026 333 264060 357
rect 262584 131 262986 165
rect 263030 145 263373 181
rect 262500 17 262550 117
rect 262626 61 262660 131
rect 262700 17 262776 97
rect 262820 61 262854 131
rect 262908 17 262984 97
rect 263030 51 263080 145
rect 263124 17 263158 111
rect 263192 51 263268 145
rect 263312 17 263346 111
rect 263413 17 263471 162
rect 263505 151 263573 265
rect 263617 199 263748 265
rect 263812 199 263970 323
rect 264026 299 264171 333
rect 264212 299 264287 493
rect 264137 265 264171 299
rect 264014 199 264103 265
rect 264137 199 264189 265
rect 263505 17 263573 117
rect 263617 61 263666 199
rect 264137 165 264171 199
rect 263821 131 264171 165
rect 264233 152 264287 299
rect 264333 294 264391 527
rect 264511 467 264587 527
rect 264734 467 264801 527
rect 264510 399 264781 433
rect 264845 425 264992 483
rect 265040 443 265147 477
rect 264510 378 264571 399
rect 264425 321 264571 378
rect 264716 391 264781 399
rect 265040 391 265074 443
rect 264425 215 264493 287
rect 264537 181 264571 321
rect 263705 17 263771 117
rect 263821 61 263855 131
rect 263890 17 263966 97
rect 264010 61 264044 131
rect 264078 17 264164 97
rect 264212 83 264287 152
rect 264333 17 264391 162
rect 264425 147 264571 181
rect 264612 299 264678 365
rect 264716 357 265074 391
rect 265113 323 265190 356
rect 264612 158 264655 299
rect 264712 289 265190 323
rect 265253 294 265311 527
rect 265345 427 265401 527
rect 264712 265 264755 289
rect 264689 192 264755 265
rect 264789 215 264912 255
rect 264968 215 265188 255
rect 265349 199 265417 391
rect 265457 265 265495 491
rect 265545 349 265611 490
rect 265545 315 265673 349
rect 265457 199 265581 265
rect 264721 174 264755 192
rect 264425 65 264478 147
rect 264544 17 264578 113
rect 264612 52 264678 158
rect 264721 140 265069 174
rect 264715 17 264801 97
rect 264845 54 264879 140
rect 264925 17 264991 97
rect 265035 54 265069 140
rect 265113 17 265189 117
rect 265253 17 265311 162
rect 265345 17 265397 165
rect 265457 87 265495 199
rect 265629 165 265673 315
rect 265707 199 265765 475
rect 265803 199 265869 475
rect 265962 359 266012 527
rect 266067 325 266117 493
rect 266161 359 266211 527
rect 266255 325 266305 493
rect 266349 359 266399 527
rect 265903 289 266016 323
rect 266067 291 266411 325
rect 266449 294 266507 527
rect 266541 407 266593 491
rect 266627 441 266703 527
rect 266846 441 267005 475
rect 266541 373 266927 407
rect 265903 199 265963 289
rect 265997 215 266319 249
rect 265997 165 266031 215
rect 266363 181 266411 291
rect 265629 131 266031 165
rect 266075 145 266411 181
rect 266541 165 266575 373
rect 266609 199 266686 339
rect 266732 305 266859 339
rect 266720 199 266791 265
rect 266825 249 266859 305
rect 266893 317 266927 373
rect 266971 391 267005 441
rect 267060 425 267198 491
rect 266971 357 267198 391
rect 267242 367 267298 527
rect 267164 333 267198 357
rect 266893 283 267033 317
rect 267164 299 267306 333
rect 267350 299 267415 493
rect 266825 215 266955 249
rect 266825 165 266859 215
rect 266999 199 267033 283
rect 267272 265 267306 299
rect 267087 199 267238 265
rect 267272 199 267330 265
rect 267272 165 267306 199
rect 265545 17 265595 117
rect 265671 61 265705 131
rect 265745 17 265821 97
rect 265865 61 265899 131
rect 265953 17 266029 97
rect 266075 51 266125 145
rect 266169 17 266203 111
rect 266237 51 266313 145
rect 266357 17 266391 111
rect 266449 17 266507 162
rect 266541 90 266604 165
rect 266665 17 266699 165
rect 266759 131 266859 165
rect 266957 131 267306 165
rect 267371 152 267415 299
rect 267461 294 267519 527
rect 267553 407 267605 491
rect 267639 441 267715 527
rect 267863 441 268022 475
rect 267553 373 267944 407
rect 267553 165 267588 373
rect 267622 199 267702 339
rect 267745 305 267876 339
rect 267736 199 267804 265
rect 267838 249 267876 305
rect 267910 317 267944 373
rect 267988 391 268022 441
rect 268077 425 268215 491
rect 267988 357 268215 391
rect 268259 367 268315 527
rect 268181 333 268215 357
rect 267910 283 268050 317
rect 268181 299 268323 333
rect 268367 299 268427 493
rect 267838 215 267927 249
rect 267838 165 267876 215
rect 268016 199 268050 283
rect 268289 265 268323 299
rect 268104 199 268255 265
rect 268289 199 268344 265
rect 268289 165 268323 199
rect 266759 90 266793 131
rect 266838 17 266913 97
rect 266957 61 266991 131
rect 267028 17 267104 97
rect 267148 61 267182 131
rect 267216 17 267302 97
rect 267350 83 267415 152
rect 267461 17 267519 162
rect 267553 90 267617 165
rect 267678 17 267712 165
rect 267772 131 267876 165
rect 267974 131 268323 165
rect 268388 152 268427 299
rect 268466 288 268500 527
rect 268565 294 268623 527
rect 268659 414 268709 491
rect 268743 448 268819 527
rect 268885 459 269153 493
rect 268885 414 268919 459
rect 268659 380 268919 414
rect 268962 391 269085 425
rect 267772 90 267806 131
rect 267855 17 267930 97
rect 267974 61 268008 131
rect 268045 17 268121 97
rect 268165 61 268199 131
rect 268233 17 268319 97
rect 268367 83 268427 152
rect 268466 17 268500 183
rect 268659 165 268693 380
rect 268727 199 268805 339
rect 268848 312 268979 346
rect 268941 265 268979 312
rect 268839 199 268907 265
rect 268941 199 268999 265
rect 268941 165 268979 199
rect 268565 17 268623 162
rect 268659 90 268720 165
rect 268781 17 268815 165
rect 268875 131 268979 165
rect 269047 165 269085 391
rect 269119 199 269153 459
rect 269209 199 269269 475
rect 269372 359 269422 527
rect 269477 325 269527 493
rect 269571 359 269621 527
rect 269665 325 269715 493
rect 269759 359 269809 527
rect 269303 280 269375 323
rect 269477 291 269811 325
rect 269853 294 269911 527
rect 269962 393 269997 493
rect 270031 427 270107 527
rect 269962 359 270105 393
rect 269331 199 269375 280
rect 269409 215 269729 249
rect 269409 165 269443 215
rect 269765 181 269811 291
rect 269945 195 270015 325
rect 269047 131 269443 165
rect 269485 145 269811 181
rect 268875 90 268909 131
rect 268963 17 269029 96
rect 269089 61 269123 131
rect 269157 17 269233 97
rect 269277 61 269311 131
rect 269363 17 269439 97
rect 269485 51 269535 145
rect 269579 17 269613 111
rect 269647 51 269723 145
rect 269767 17 269801 111
rect 269853 17 269911 162
rect 270059 161 270105 359
rect 269962 127 270105 161
rect 269962 69 269997 127
rect 270031 17 270107 93
rect 270151 69 270192 493
rect 270239 377 270305 527
rect 270405 375 270481 477
rect 270547 381 270581 493
rect 270630 443 270706 527
rect 270226 205 270281 337
rect 270315 203 270379 339
rect 270438 273 270481 375
rect 270517 349 270581 381
rect 270517 315 270707 349
rect 270438 237 270583 273
rect 270485 215 270583 237
rect 270673 219 270707 315
rect 270759 265 270823 475
rect 270315 153 270449 203
rect 270315 152 270379 153
rect 270239 17 270289 127
rect 270323 69 270379 152
rect 270485 119 270519 215
rect 270673 159 270742 219
rect 270438 53 270519 119
rect 270553 153 270742 159
rect 270553 125 270707 153
rect 270553 61 270593 125
rect 270652 17 270718 89
rect 270857 61 270891 493
rect 270935 450 271111 484
rect 270925 315 271043 391
rect 270925 141 270977 315
rect 271077 281 271111 450
rect 271169 441 271245 527
rect 271315 407 271349 475
rect 271145 357 271445 407
rect 271493 383 271559 527
rect 271788 450 271974 484
rect 272032 451 272108 527
rect 271145 315 271205 357
rect 271317 281 271367 297
rect 271077 247 271367 281
rect 271077 239 271171 247
rect 271013 129 271093 203
rect 271127 93 271171 239
rect 271323 231 271367 247
rect 271411 213 271445 357
rect 271489 283 271710 331
rect 271750 315 271797 397
rect 271489 247 271555 283
rect 271855 261 271906 381
rect 271617 213 271703 247
rect 271205 147 271287 213
rect 271411 179 271703 213
rect 271762 225 271906 261
rect 271940 281 271974 450
rect 272166 417 272200 475
rect 272316 451 272614 527
rect 272008 383 272614 417
rect 272008 315 272068 383
rect 271940 247 272230 281
rect 271411 153 271459 179
rect 271383 119 271459 153
rect 270948 53 271171 93
rect 271205 17 271239 105
rect 271283 85 271349 93
rect 271498 85 271537 143
rect 271762 141 271830 225
rect 271940 93 271974 247
rect 272186 215 272230 247
rect 272059 147 272144 213
rect 272274 163 272311 383
rect 272235 129 272311 163
rect 272354 315 272509 349
rect 272354 185 272397 315
rect 272580 265 272614 383
rect 272671 326 272747 493
rect 272781 345 272832 483
rect 272877 353 272936 527
rect 272692 304 272747 326
rect 272431 219 272546 265
rect 272580 199 272633 265
rect 272354 151 272491 185
rect 271283 51 271537 85
rect 271586 17 271663 93
rect 271811 53 271974 93
rect 272010 17 272072 105
rect 272124 85 272204 93
rect 272353 85 272388 117
rect 272124 51 272388 85
rect 272451 53 272491 151
rect 272548 17 272614 161
rect 272692 143 272751 304
rect 272671 51 272751 143
rect 272791 265 272832 345
rect 272980 321 273037 493
rect 272791 199 272946 265
rect 272791 51 272832 199
rect 272990 165 273037 321
rect 273073 294 273131 527
rect 273166 393 273217 493
rect 273254 427 273330 527
rect 273166 359 273331 393
rect 273176 195 273246 325
rect 273290 265 273331 359
rect 273375 346 273421 493
rect 273570 417 273624 480
rect 273668 451 273734 527
rect 273570 383 273694 417
rect 273290 199 273353 265
rect 272878 17 272936 109
rect 272980 51 273037 165
rect 273073 17 273131 162
rect 273290 161 273325 199
rect 273167 127 273325 161
rect 273387 135 273421 346
rect 273465 267 273592 349
rect 273465 214 273546 267
rect 273643 237 273694 383
rect 273772 271 273879 493
rect 273922 421 273956 493
rect 274119 455 274189 527
rect 274244 437 274318 487
rect 274244 421 274278 437
rect 274367 427 274440 493
rect 273922 387 274278 421
rect 273643 233 273837 237
rect 273601 199 273837 233
rect 273922 215 273957 387
rect 273601 180 273635 199
rect 273167 69 273217 127
rect 273251 17 273327 93
rect 273371 69 273421 135
rect 273487 146 273635 180
rect 273487 79 273521 146
rect 273555 17 273631 112
rect 273679 17 273755 165
rect 273803 85 273837 199
rect 273881 135 273957 215
rect 274001 85 274035 337
rect 274070 142 274139 340
rect 274176 179 274210 387
rect 274312 315 274372 391
rect 274244 213 274278 279
rect 274328 207 274372 315
rect 274406 277 274440 427
rect 274484 421 274518 475
rect 274575 471 274641 527
rect 274702 421 274736 475
rect 274778 435 274862 527
rect 274484 387 274736 421
rect 274911 401 274945 493
rect 274987 425 275191 493
rect 275231 439 275281 527
rect 274794 367 274945 401
rect 274794 353 274856 367
rect 274540 319 274856 353
rect 274985 333 275117 391
rect 274406 243 274778 277
rect 274176 143 274292 179
rect 273803 51 274035 85
rect 274149 17 274218 108
rect 274258 101 274292 143
rect 274328 141 274478 207
rect 274258 67 274326 101
rect 274516 95 274550 243
rect 274594 153 274710 209
rect 274744 201 274778 243
rect 274822 167 274856 319
rect 274370 61 274550 95
rect 274686 17 274752 109
rect 274794 89 274856 167
rect 274890 332 275117 333
rect 275156 349 275191 425
rect 275330 417 275364 475
rect 275399 451 275475 527
rect 275330 383 275494 417
rect 274890 299 275037 332
rect 275156 315 275422 349
rect 274890 141 274942 299
rect 275156 297 275205 315
rect 274995 184 275029 265
rect 275082 263 275205 297
rect 275460 265 275494 383
rect 275529 299 275586 527
rect 275082 107 275126 263
rect 275178 173 275222 229
rect 275268 213 275422 255
rect 275178 139 275294 173
rect 274794 55 274870 89
rect 274904 51 275126 107
rect 275170 17 275214 105
rect 275260 93 275294 139
rect 275361 127 275422 213
rect 275460 199 275589 265
rect 275460 93 275495 199
rect 275260 59 275495 93
rect 275529 17 275586 142
rect 275632 53 275702 479
rect 275736 341 275770 493
rect 275805 375 275887 527
rect 275736 307 275869 341
rect 275835 265 275869 307
rect 275925 295 275981 493
rect 275835 199 275901 265
rect 275835 161 275869 199
rect 275935 174 275981 295
rect 276017 294 276075 527
rect 276110 393 276161 493
rect 276198 427 276274 527
rect 276110 359 276275 393
rect 276120 195 276190 325
rect 276234 265 276275 359
rect 276319 346 276365 493
rect 276514 417 276568 480
rect 276612 451 276678 527
rect 276514 383 276638 417
rect 276234 199 276297 265
rect 275736 127 275869 161
rect 275736 51 275770 127
rect 275805 17 275887 93
rect 275925 51 275981 174
rect 276017 17 276075 162
rect 276234 161 276269 199
rect 276111 127 276269 161
rect 276331 135 276365 346
rect 276409 267 276536 349
rect 276409 214 276490 267
rect 276587 237 276638 383
rect 276716 271 276823 493
rect 276866 421 276900 493
rect 277063 455 277133 527
rect 277188 437 277262 487
rect 277188 421 277222 437
rect 277311 427 277384 493
rect 276866 387 277222 421
rect 276587 233 276781 237
rect 276545 199 276781 233
rect 276866 215 276901 387
rect 276545 180 276579 199
rect 276111 69 276161 127
rect 276195 17 276271 93
rect 276315 69 276365 135
rect 276431 146 276579 180
rect 276431 79 276465 146
rect 276499 17 276575 112
rect 276623 17 276699 165
rect 276747 85 276781 199
rect 276825 135 276901 215
rect 276945 85 276979 337
rect 277014 142 277083 340
rect 277120 179 277154 387
rect 277256 315 277316 391
rect 277188 213 277222 279
rect 277272 207 277316 315
rect 277350 277 277384 427
rect 277428 421 277462 475
rect 277519 471 277585 527
rect 277646 421 277680 475
rect 277722 435 277806 527
rect 277428 387 277680 421
rect 277855 401 277889 493
rect 277931 425 278135 493
rect 278175 439 278225 527
rect 277738 367 277889 401
rect 277738 353 277800 367
rect 277484 319 277800 353
rect 277929 333 278061 391
rect 277350 243 277722 277
rect 277120 143 277236 179
rect 276747 51 276979 85
rect 277093 17 277162 108
rect 277202 101 277236 143
rect 277272 141 277422 207
rect 277202 67 277270 101
rect 277460 95 277494 243
rect 277538 153 277654 209
rect 277688 201 277722 243
rect 277766 167 277800 319
rect 277314 61 277494 95
rect 277630 17 277696 109
rect 277738 89 277800 167
rect 277834 332 278061 333
rect 278100 349 278135 425
rect 278274 417 278308 475
rect 278343 451 278419 527
rect 278274 383 278438 417
rect 277834 299 277981 332
rect 278100 315 278366 349
rect 277834 141 277886 299
rect 278100 297 278149 315
rect 277939 184 277973 265
rect 278026 263 278149 297
rect 278404 265 278438 383
rect 278472 407 278507 493
rect 278543 441 278635 527
rect 278746 451 278837 527
rect 278472 373 278812 407
rect 278472 359 278620 373
rect 278026 107 278070 263
rect 278122 173 278166 229
rect 278212 213 278366 255
rect 278122 139 278238 173
rect 277738 55 277814 89
rect 277848 51 278070 107
rect 278114 17 278158 105
rect 278204 93 278238 139
rect 278305 127 278366 213
rect 278404 199 278533 265
rect 278404 93 278438 199
rect 278585 165 278620 359
rect 278204 59 278438 93
rect 278472 131 278620 165
rect 278472 69 278506 131
rect 278557 17 278623 97
rect 278664 53 278744 339
rect 278778 265 278812 373
rect 278846 307 278933 416
rect 278778 199 278865 265
rect 278899 165 278933 307
rect 278967 299 279017 527
rect 279053 294 279111 527
rect 279146 393 279197 493
rect 279234 427 279310 527
rect 279146 359 279311 393
rect 279156 195 279226 325
rect 279270 265 279311 359
rect 279355 346 279401 493
rect 279550 417 279604 480
rect 279648 451 279714 527
rect 279550 383 279674 417
rect 279270 199 279333 265
rect 278780 17 278814 165
rect 278848 62 278933 165
rect 278967 17 279001 186
rect 279053 17 279111 162
rect 279270 161 279305 199
rect 279147 127 279305 161
rect 279367 135 279401 346
rect 279445 267 279572 349
rect 279445 214 279526 267
rect 279623 237 279674 383
rect 279752 271 279859 493
rect 279902 421 279936 493
rect 280099 455 280169 527
rect 280224 437 280298 487
rect 280224 421 280258 437
rect 280347 427 280420 493
rect 279902 387 280258 421
rect 279623 233 279817 237
rect 279581 199 279817 233
rect 279902 215 279937 387
rect 279581 180 279615 199
rect 279147 69 279197 127
rect 279231 17 279307 93
rect 279351 69 279401 135
rect 279467 146 279615 180
rect 279467 79 279501 146
rect 279535 17 279611 112
rect 279659 17 279735 165
rect 279783 85 279817 199
rect 279861 135 279937 215
rect 279981 85 280015 337
rect 280050 142 280119 340
rect 280156 179 280190 387
rect 280292 315 280352 391
rect 280224 213 280258 279
rect 280308 207 280352 315
rect 280386 277 280420 427
rect 280464 421 280498 475
rect 280555 471 280621 527
rect 280682 421 280716 475
rect 280758 435 280842 527
rect 280464 387 280716 421
rect 280891 401 280925 493
rect 280967 425 281171 493
rect 281211 439 281261 527
rect 280774 367 280925 401
rect 280774 353 280836 367
rect 280520 319 280836 353
rect 280965 333 281097 391
rect 280386 243 280758 277
rect 280156 143 280272 179
rect 279783 51 280015 85
rect 280129 17 280198 108
rect 280238 101 280272 143
rect 280308 141 280458 207
rect 280238 67 280306 101
rect 280496 95 280530 243
rect 280574 153 280690 209
rect 280724 201 280758 243
rect 280802 167 280836 319
rect 280350 61 280530 95
rect 280666 17 280732 109
rect 280774 89 280836 167
rect 280870 332 281097 333
rect 281136 349 281171 425
rect 281310 417 281344 475
rect 281379 451 281455 527
rect 281310 383 281474 417
rect 280870 299 281017 332
rect 281136 315 281402 349
rect 280870 141 280922 299
rect 281136 297 281185 315
rect 280975 184 281009 265
rect 281062 263 281185 297
rect 281440 265 281474 383
rect 281509 299 281566 527
rect 281062 107 281106 263
rect 281158 173 281202 229
rect 281248 213 281402 255
rect 281158 139 281274 173
rect 280774 55 280850 89
rect 280884 51 281106 107
rect 281150 17 281194 105
rect 281240 93 281274 139
rect 281341 127 281402 213
rect 281440 199 281569 265
rect 281440 93 281475 199
rect 281240 59 281475 93
rect 281509 17 281566 142
rect 281612 53 281685 465
rect 281721 294 281779 527
rect 281814 393 281865 493
rect 281902 427 281978 527
rect 281814 359 281979 393
rect 281824 195 281894 325
rect 281938 265 281979 359
rect 282023 346 282069 493
rect 282218 417 282272 480
rect 282316 451 282382 527
rect 282218 383 282342 417
rect 281938 199 282001 265
rect 281721 17 281779 162
rect 281938 161 281973 199
rect 281815 127 281973 161
rect 282035 135 282069 346
rect 282113 267 282240 349
rect 282113 214 282194 267
rect 282291 237 282342 383
rect 282420 271 282527 493
rect 282570 421 282604 493
rect 282767 455 282837 527
rect 282892 437 282966 487
rect 282892 421 282926 437
rect 283015 427 283088 493
rect 282570 387 282926 421
rect 282291 233 282485 237
rect 282249 199 282485 233
rect 282570 215 282605 387
rect 282249 180 282283 199
rect 281815 69 281865 127
rect 281899 17 281975 93
rect 282019 69 282069 135
rect 282135 146 282283 180
rect 282135 79 282169 146
rect 282203 17 282279 112
rect 282327 17 282403 165
rect 282451 85 282485 199
rect 282529 135 282605 215
rect 282649 85 282683 337
rect 282718 142 282787 340
rect 282824 179 282858 387
rect 282960 315 283020 391
rect 282892 213 282926 279
rect 282976 207 283020 315
rect 283054 277 283088 427
rect 283132 421 283166 475
rect 283223 471 283289 527
rect 283350 421 283384 475
rect 283426 435 283510 527
rect 283132 387 283384 421
rect 283559 401 283593 493
rect 283635 425 283839 493
rect 283879 439 283929 527
rect 283442 367 283593 401
rect 283442 353 283504 367
rect 283188 319 283504 353
rect 283633 333 283765 391
rect 283054 243 283426 277
rect 282824 143 282940 179
rect 282451 51 282683 85
rect 282797 17 282866 108
rect 282906 101 282940 143
rect 282976 141 283126 207
rect 282906 67 282974 101
rect 283164 95 283198 243
rect 283242 153 283358 209
rect 283392 201 283426 243
rect 283470 167 283504 319
rect 283018 61 283198 95
rect 283334 17 283400 109
rect 283442 89 283504 167
rect 283538 332 283765 333
rect 283804 349 283839 425
rect 283978 417 284012 475
rect 284047 451 284123 527
rect 283978 383 284142 417
rect 283538 299 283685 332
rect 283804 315 284070 349
rect 283538 141 283590 299
rect 283804 297 283853 315
rect 283643 184 283677 265
rect 283730 263 283853 297
rect 284108 265 284142 383
rect 284177 299 284234 527
rect 283730 107 283774 263
rect 283826 173 283870 229
rect 283916 213 284070 255
rect 283826 139 283942 173
rect 283442 55 283518 89
rect 283552 51 283774 107
rect 283818 17 283862 105
rect 283908 93 283942 139
rect 284009 127 284070 213
rect 284108 199 284237 265
rect 284108 93 284143 199
rect 283908 59 284143 93
rect 284177 17 284234 142
rect 284280 53 284353 465
rect 284389 294 284447 527
rect 284482 393 284533 493
rect 284570 427 284646 527
rect 284482 359 284647 393
rect 284492 195 284562 325
rect 284606 265 284647 359
rect 284691 346 284737 493
rect 284886 417 284940 480
rect 284984 451 285050 527
rect 284886 383 285010 417
rect 284606 199 284669 265
rect 284389 17 284447 162
rect 284606 161 284641 199
rect 284483 127 284641 161
rect 284703 135 284737 346
rect 284781 267 284908 349
rect 284781 214 284862 267
rect 284959 237 285010 383
rect 285088 271 285195 493
rect 285238 421 285272 493
rect 285435 455 285505 527
rect 285560 437 285634 487
rect 285560 421 285594 437
rect 285683 427 285756 493
rect 285238 387 285594 421
rect 284959 233 285153 237
rect 284917 199 285153 233
rect 285238 215 285273 387
rect 284917 180 284951 199
rect 284483 69 284533 127
rect 284567 17 284643 93
rect 284687 69 284737 135
rect 284803 146 284951 180
rect 284803 79 284837 146
rect 284871 17 284947 112
rect 284995 17 285071 165
rect 285119 85 285153 199
rect 285197 135 285273 215
rect 285317 85 285351 337
rect 285386 142 285455 340
rect 285492 179 285526 387
rect 285628 315 285688 391
rect 285560 213 285594 279
rect 285644 207 285688 315
rect 285722 277 285756 427
rect 285800 421 285834 475
rect 285891 471 285957 527
rect 286018 421 286052 475
rect 286094 435 286178 527
rect 285800 387 286052 421
rect 286227 401 286261 493
rect 286303 425 286507 493
rect 286547 439 286597 527
rect 286110 367 286261 401
rect 286110 353 286172 367
rect 285856 319 286172 353
rect 286301 333 286433 391
rect 285722 243 286094 277
rect 285492 143 285608 179
rect 285119 51 285351 85
rect 285465 17 285534 108
rect 285574 101 285608 143
rect 285644 141 285794 207
rect 285574 67 285642 101
rect 285832 95 285866 243
rect 285910 153 286026 209
rect 286060 201 286094 243
rect 286138 167 286172 319
rect 285686 61 285866 95
rect 286002 17 286068 109
rect 286110 89 286172 167
rect 286206 332 286433 333
rect 286472 349 286507 425
rect 286646 417 286680 475
rect 286715 451 286791 527
rect 286646 383 286810 417
rect 286206 299 286353 332
rect 286472 315 286738 349
rect 286206 141 286258 299
rect 286472 297 286521 315
rect 286311 184 286345 265
rect 286398 263 286521 297
rect 286776 265 286810 383
rect 286845 299 286930 527
rect 286398 107 286442 263
rect 286494 173 286538 229
rect 286584 213 286738 255
rect 286494 139 286610 173
rect 286110 55 286186 89
rect 286220 51 286442 107
rect 286486 17 286530 105
rect 286576 93 286610 139
rect 286677 127 286738 213
rect 286776 199 286911 265
rect 286776 93 286811 199
rect 286576 59 286811 93
rect 286845 17 286929 134
rect 286964 53 287021 465
rect 287063 299 287113 527
rect 287149 294 287207 527
rect 287241 405 287293 493
rect 287327 439 287387 527
rect 287431 451 287673 493
rect 287431 405 287465 451
rect 287718 417 287761 493
rect 287812 428 287880 527
rect 287241 369 287465 405
rect 287503 374 287593 415
rect 287063 17 287097 109
rect 287149 17 287207 162
rect 287241 153 287297 335
rect 287334 153 287396 335
rect 287430 153 287509 335
rect 287241 17 287310 119
rect 287555 112 287593 374
rect 287637 354 287761 417
rect 287637 181 287704 354
rect 287795 344 287891 394
rect 287925 391 287959 465
rect 287993 455 288069 527
rect 288113 427 288182 493
rect 287925 355 288083 391
rect 287855 318 287891 344
rect 287738 215 287814 310
rect 287855 211 287987 318
rect 287637 143 287767 181
rect 288031 177 288083 355
rect 287419 56 287593 112
rect 287629 17 287665 109
rect 287716 51 287767 143
rect 287928 143 288083 177
rect 288127 284 288182 427
rect 288216 318 288260 493
rect 288310 427 288465 493
rect 288513 455 288579 527
rect 288127 218 288192 284
rect 287812 17 287880 111
rect 287928 51 287965 143
rect 288127 117 288161 218
rect 288226 184 288260 318
rect 288345 315 288397 391
rect 288431 279 288465 427
rect 288644 421 288697 490
rect 288755 425 288966 527
rect 289000 425 289171 492
rect 289233 447 289309 527
rect 288509 387 288697 421
rect 289137 413 289171 425
rect 289353 413 289396 490
rect 289451 447 289517 527
rect 288509 315 288543 387
rect 288662 289 288769 353
rect 288806 299 288975 391
rect 288321 255 288611 279
rect 288814 255 288896 265
rect 288010 17 288072 109
rect 288116 51 288161 117
rect 288195 51 288260 184
rect 288304 245 288896 255
rect 288304 51 288402 245
rect 288436 161 288519 203
rect 288574 195 288896 245
rect 288931 179 288975 299
rect 289047 215 289103 381
rect 289137 379 289517 413
rect 289161 305 289439 345
rect 289473 305 289517 379
rect 289161 283 289216 305
rect 289561 271 289613 493
rect 289658 297 289700 527
rect 289146 179 289202 249
rect 288436 127 288641 161
rect 288931 139 289202 179
rect 289252 237 289613 271
rect 289252 171 289297 237
rect 289345 169 289533 203
rect 288436 17 288543 93
rect 288579 51 288641 127
rect 288732 17 288879 138
rect 289345 89 289379 169
rect 289056 55 289379 89
rect 289468 17 289502 109
rect 289577 108 289613 237
rect 289536 51 289613 108
rect 289658 17 289700 177
rect 289734 51 289810 493
rect 289856 265 289898 493
rect 289969 315 290003 527
rect 290037 299 290149 490
rect 289856 199 290034 265
rect 289856 51 289898 199
rect 290078 165 290149 299
rect 290185 294 290243 527
rect 290277 405 290329 493
rect 290363 439 290423 527
rect 290467 451 290709 493
rect 290467 405 290501 451
rect 290754 417 290797 493
rect 290848 428 290916 527
rect 290277 369 290501 405
rect 290539 374 290629 415
rect 289962 17 290003 165
rect 290037 55 290149 165
rect 290185 17 290243 162
rect 290277 153 290333 335
rect 290370 153 290432 335
rect 290466 153 290545 335
rect 290277 17 290346 119
rect 290591 112 290629 374
rect 290673 354 290797 417
rect 290673 181 290740 354
rect 290831 344 290927 394
rect 290961 391 290995 465
rect 291029 455 291105 527
rect 291149 427 291218 493
rect 290961 355 291119 391
rect 290891 318 290927 344
rect 290774 215 290850 310
rect 290891 211 291023 318
rect 290673 143 290803 181
rect 291067 177 291119 355
rect 290455 56 290629 112
rect 290665 17 290701 109
rect 290752 51 290803 143
rect 290964 143 291119 177
rect 291163 284 291218 427
rect 291252 318 291296 493
rect 291346 427 291501 493
rect 291549 455 291615 527
rect 291163 218 291228 284
rect 290848 17 290916 111
rect 290964 51 291001 143
rect 291163 117 291197 218
rect 291262 184 291296 318
rect 291381 315 291433 391
rect 291467 279 291501 427
rect 291680 421 291733 490
rect 291791 425 292002 527
rect 292036 425 292207 492
rect 292269 447 292345 527
rect 291545 387 291733 421
rect 292173 413 292207 425
rect 292389 413 292432 490
rect 292487 447 292553 527
rect 291545 315 291579 387
rect 291698 289 291805 353
rect 291842 299 292011 391
rect 291357 255 291647 279
rect 291850 255 291932 265
rect 291046 17 291108 109
rect 291152 51 291197 117
rect 291231 51 291296 184
rect 291340 245 291932 255
rect 291340 51 291438 245
rect 291472 161 291555 203
rect 291610 195 291932 245
rect 291967 179 292011 299
rect 292083 215 292139 381
rect 292173 379 292553 413
rect 292197 305 292475 345
rect 292509 305 292553 379
rect 292197 283 292252 305
rect 292597 271 292649 493
rect 292694 297 292736 527
rect 292182 179 292238 249
rect 291472 127 291677 161
rect 291967 139 292238 179
rect 292288 237 292649 271
rect 292288 171 292333 237
rect 292381 169 292569 203
rect 291472 17 291579 93
rect 291615 51 291677 127
rect 291768 17 291915 138
rect 292381 89 292415 169
rect 292092 55 292415 89
rect 292504 17 292538 109
rect 292613 108 292649 237
rect 292572 51 292649 108
rect 292694 17 292736 177
rect 292771 51 292860 493
rect 292903 297 292961 527
rect 293004 265 293041 493
rect 293075 327 293156 527
rect 293200 299 293276 490
rect 293004 199 293177 265
rect 292903 17 292961 177
rect 293004 51 293041 199
rect 293221 165 293276 299
rect 293310 297 293363 527
rect 293405 294 293463 527
rect 293497 405 293549 493
rect 293583 439 293647 527
rect 293691 451 293929 493
rect 293691 405 293725 451
rect 293974 417 294024 493
rect 294068 428 294127 527
rect 293497 369 293725 405
rect 293759 369 293849 417
rect 293075 17 293156 165
rect 293200 55 293276 165
rect 293310 17 293363 177
rect 293405 17 293463 162
rect 293497 153 293548 335
rect 293588 153 293654 335
rect 293688 153 293777 335
rect 293811 119 293849 369
rect 293893 354 294024 417
rect 294181 400 294215 465
rect 294249 455 294325 527
rect 294369 427 294438 493
rect 294181 366 294339 400
rect 293893 181 293960 354
rect 293994 215 294070 320
rect 294111 211 294243 330
rect 293893 143 294024 181
rect 294287 177 294339 366
rect 293497 17 293630 119
rect 293664 51 293849 119
rect 293885 17 293938 109
rect 293972 51 294024 143
rect 294184 143 294339 177
rect 294375 284 294438 427
rect 294473 318 294516 493
rect 294567 427 294721 493
rect 294769 455 294846 527
rect 294375 217 294448 284
rect 294068 17 294150 111
rect 294184 51 294221 143
rect 294265 17 294331 109
rect 294375 51 294417 217
rect 294482 156 294516 318
rect 294601 315 294653 391
rect 294687 279 294721 427
rect 294911 421 294964 490
rect 295022 425 295205 527
rect 295239 425 295418 492
rect 295452 447 295518 527
rect 294765 387 294964 421
rect 295384 413 295418 425
rect 295559 413 295599 490
rect 295655 447 295731 527
rect 294765 315 294799 387
rect 294918 289 295023 353
rect 295057 334 295237 391
rect 294451 51 294516 156
rect 294573 255 294875 279
rect 295061 255 295143 265
rect 294573 245 295143 255
rect 294573 51 294658 245
rect 294699 161 294775 203
rect 294841 195 295143 245
rect 295177 181 295237 334
rect 295271 215 295338 381
rect 295384 379 295731 413
rect 295396 309 295619 345
rect 295655 321 295731 379
rect 295396 285 295452 309
rect 295765 273 295817 493
rect 295384 181 295450 251
rect 294699 127 294887 161
rect 294692 17 294799 93
rect 294837 51 294887 127
rect 294931 17 295143 161
rect 295177 144 295450 181
rect 295487 239 295817 273
rect 295487 171 295536 239
rect 295570 157 295737 203
rect 295570 109 295610 157
rect 295771 117 295817 239
rect 295285 55 295610 109
rect 295647 17 295697 109
rect 295749 51 295817 117
rect 295851 265 295919 493
rect 295967 369 296018 527
rect 295851 199 296029 265
rect 295851 51 295903 199
rect 295937 17 296018 110
rect 296063 55 296128 490
rect 296165 294 296223 527
rect 296257 405 296309 493
rect 296343 439 296407 527
rect 296451 451 296689 493
rect 296451 405 296485 451
rect 296734 417 296784 493
rect 296828 428 296887 527
rect 296257 369 296485 405
rect 296519 369 296609 417
rect 296165 17 296223 162
rect 296257 153 296308 335
rect 296348 153 296414 335
rect 296448 153 296537 335
rect 296571 119 296609 369
rect 296653 354 296784 417
rect 296941 400 296975 465
rect 297009 455 297085 527
rect 297129 427 297198 493
rect 296941 366 297099 400
rect 296653 181 296720 354
rect 296754 215 296830 320
rect 296871 211 297003 330
rect 296653 143 296784 181
rect 297047 177 297099 366
rect 296257 17 296390 119
rect 296424 51 296609 119
rect 296645 17 296698 109
rect 296732 51 296784 143
rect 296944 143 297099 177
rect 297135 284 297198 427
rect 297233 318 297276 493
rect 297327 427 297481 493
rect 297529 455 297606 527
rect 297135 217 297208 284
rect 296828 17 296910 111
rect 296944 51 296981 143
rect 297025 17 297091 109
rect 297135 51 297177 217
rect 297242 156 297276 318
rect 297361 315 297413 391
rect 297447 279 297481 427
rect 297671 421 297724 490
rect 297782 425 297993 527
rect 298027 425 298208 492
rect 298252 447 298328 527
rect 297525 387 297724 421
rect 298174 413 298208 425
rect 298362 413 298443 490
rect 298481 447 298557 527
rect 297525 315 297559 387
rect 297678 289 297783 353
rect 297817 334 298017 391
rect 297211 51 297276 156
rect 297333 255 297635 279
rect 297841 255 297923 265
rect 297333 245 297923 255
rect 297333 51 297418 245
rect 297459 161 297535 203
rect 297601 195 297923 245
rect 297957 181 298017 334
rect 298075 215 298140 381
rect 298174 379 298557 413
rect 298186 309 298439 345
rect 298481 321 298557 379
rect 298186 285 298247 309
rect 298591 273 298643 493
rect 298174 181 298241 251
rect 297459 127 297647 161
rect 297452 17 297559 93
rect 297597 51 297647 127
rect 297691 17 297923 161
rect 297957 144 298241 181
rect 298284 239 298643 273
rect 298284 171 298336 239
rect 298382 157 298563 203
rect 298382 109 298422 157
rect 298597 117 298643 239
rect 298093 55 298422 109
rect 298473 17 298523 109
rect 298575 51 298643 117
rect 298677 265 298745 493
rect 298793 369 298844 527
rect 298889 299 298971 490
rect 299005 299 299039 527
rect 298677 199 298865 265
rect 298677 51 298729 199
rect 298910 165 298971 299
rect 299109 294 299167 527
rect 299201 405 299253 493
rect 299287 439 299351 527
rect 299395 451 299633 493
rect 299395 405 299429 451
rect 299678 417 299728 493
rect 299772 428 299831 527
rect 299201 369 299429 405
rect 299463 369 299553 417
rect 298763 17 298844 110
rect 298889 55 298971 165
rect 299005 17 299039 177
rect 299109 17 299167 162
rect 299201 153 299252 335
rect 299292 153 299358 335
rect 299392 153 299481 335
rect 299515 119 299553 369
rect 299597 354 299728 417
rect 299885 400 299919 465
rect 299953 455 300029 527
rect 300073 427 300142 493
rect 299885 366 300043 400
rect 299597 181 299664 354
rect 299698 215 299774 320
rect 299815 211 299947 330
rect 299597 143 299728 181
rect 299991 177 300043 366
rect 299201 17 299334 119
rect 299368 51 299553 119
rect 299589 17 299642 109
rect 299676 51 299728 143
rect 299888 143 300043 177
rect 300079 284 300142 427
rect 300177 318 300220 493
rect 300271 427 300425 493
rect 300473 455 300550 527
rect 300079 217 300152 284
rect 299772 17 299854 111
rect 299888 51 299925 143
rect 299969 17 300035 109
rect 300079 51 300121 217
rect 300186 156 300220 318
rect 300305 315 300357 391
rect 300391 279 300425 427
rect 300615 421 300668 490
rect 300726 425 300937 527
rect 300971 425 301152 492
rect 301196 447 301272 527
rect 300469 387 300668 421
rect 301118 413 301152 425
rect 301306 413 301387 490
rect 301425 447 301501 527
rect 300469 315 300503 387
rect 300622 289 300727 353
rect 300761 334 300961 391
rect 300155 51 300220 156
rect 300277 255 300579 279
rect 300785 255 300867 265
rect 300277 245 300867 255
rect 300277 51 300362 245
rect 300403 161 300479 203
rect 300545 195 300867 245
rect 300901 181 300961 334
rect 301019 215 301084 381
rect 301118 379 301501 413
rect 301130 309 301383 345
rect 301425 321 301501 379
rect 301130 285 301191 309
rect 301535 273 301587 493
rect 301118 181 301185 251
rect 300403 127 300591 161
rect 300396 17 300503 93
rect 300541 51 300591 127
rect 300635 17 300867 161
rect 300901 144 301185 181
rect 301228 239 301587 273
rect 301228 171 301280 239
rect 301326 157 301507 203
rect 301326 109 301366 157
rect 301541 117 301587 239
rect 301037 55 301366 109
rect 301417 17 301467 109
rect 301519 51 301587 117
rect 301621 265 301673 493
rect 301707 299 301788 527
rect 301832 299 301898 490
rect 301942 299 301976 527
rect 301853 265 301898 299
rect 302010 265 302106 493
rect 302140 299 302197 527
rect 302237 294 302295 527
rect 302347 393 302381 493
rect 302415 427 302491 527
rect 302347 359 302491 393
rect 301621 199 301809 265
rect 301853 211 302106 265
rect 301621 51 301673 199
rect 301853 165 301898 211
rect 301707 17 301788 165
rect 301832 55 301898 165
rect 301942 17 301976 177
rect 302010 51 302106 211
rect 302331 195 302401 325
rect 302445 194 302491 359
rect 302140 17 302197 177
rect 302237 17 302295 162
rect 302445 161 302484 194
rect 302347 127 302484 161
rect 302347 69 302381 127
rect 302415 17 302491 93
rect 302535 69 302569 493
rect 302616 415 302673 489
rect 302707 449 302783 527
rect 302887 449 303086 483
rect 302616 372 303018 415
rect 302616 89 302650 372
rect 302684 157 302718 337
rect 302762 225 302796 372
rect 302979 337 303018 372
rect 303052 399 303086 449
rect 303130 433 303164 527
rect 303215 414 303272 488
rect 303311 438 303555 472
rect 303215 399 303249 414
rect 303052 365 303249 399
rect 302863 271 302937 337
rect 302979 271 303023 337
rect 302762 191 302851 225
rect 302975 157 303019 223
rect 303075 211 303181 331
rect 303215 177 303249 365
rect 302684 123 303019 157
rect 303053 143 303249 177
rect 303053 89 303087 143
rect 302616 51 302693 89
rect 302741 17 302807 89
rect 302922 55 303087 89
rect 303131 17 303171 109
rect 303215 107 303249 143
rect 303283 207 303341 381
rect 303379 331 303477 402
rect 303511 315 303555 438
rect 303589 367 303623 527
rect 303657 427 303717 493
rect 303762 433 303969 467
rect 303511 297 303623 315
rect 303453 263 303623 297
rect 303283 141 303409 207
rect 303453 107 303487 263
rect 303589 249 303623 263
rect 303531 213 303565 219
rect 303657 213 303701 427
rect 303735 249 303783 393
rect 303817 315 303891 381
rect 303531 153 303701 213
rect 303817 207 303855 315
rect 303935 281 303969 433
rect 304015 427 304076 527
rect 304134 381 304192 491
rect 304009 315 304192 381
rect 304236 325 304270 527
rect 303215 73 303285 107
rect 303329 73 303487 107
rect 303547 17 303621 117
rect 303657 107 303701 153
rect 303735 141 303855 207
rect 303899 265 303969 281
rect 304155 265 304192 315
rect 304308 301 304400 493
rect 303899 199 304121 265
rect 304155 199 304322 265
rect 303899 107 303943 199
rect 304155 165 304192 199
rect 304356 165 304400 301
rect 303657 73 303759 107
rect 303815 73 303943 107
rect 303988 17 304072 123
rect 304126 60 304192 165
rect 304236 17 304270 139
rect 304304 61 304400 165
rect 304434 265 304484 485
rect 304530 299 304591 527
rect 304434 199 304600 265
rect 304434 69 304484 199
rect 304525 17 304591 161
rect 304635 53 304686 465
rect 304721 294 304779 527
rect 304831 393 304865 493
rect 304899 427 304975 527
rect 304831 359 304975 393
rect 304815 195 304885 325
rect 304929 194 304975 359
rect 304721 17 304779 162
rect 304929 161 304968 194
rect 304831 127 304968 161
rect 304831 69 304865 127
rect 304899 17 304975 93
rect 305019 69 305053 493
rect 305100 415 305157 489
rect 305191 449 305267 527
rect 305371 449 305570 483
rect 305100 372 305502 415
rect 305100 89 305134 372
rect 305168 157 305202 337
rect 305246 225 305280 372
rect 305463 337 305502 372
rect 305536 399 305570 449
rect 305614 433 305648 527
rect 305699 414 305756 488
rect 305795 438 306039 472
rect 305699 399 305733 414
rect 305536 365 305733 399
rect 305347 271 305421 337
rect 305463 271 305507 337
rect 305246 191 305335 225
rect 305459 157 305503 223
rect 305559 211 305665 331
rect 305699 177 305733 365
rect 305168 123 305503 157
rect 305537 143 305733 177
rect 305537 89 305571 143
rect 305100 51 305177 89
rect 305225 17 305291 89
rect 305406 55 305571 89
rect 305615 17 305655 109
rect 305699 107 305733 143
rect 305767 207 305825 381
rect 305863 331 305961 402
rect 305995 315 306039 438
rect 306073 367 306107 527
rect 306141 427 306201 493
rect 306246 433 306453 467
rect 305995 297 306107 315
rect 305937 263 306107 297
rect 305767 141 305893 207
rect 305937 107 305971 263
rect 306073 249 306107 263
rect 306015 213 306049 219
rect 306141 213 306185 427
rect 306219 249 306267 393
rect 306301 315 306375 381
rect 306015 153 306185 213
rect 306301 207 306339 315
rect 306419 281 306453 433
rect 306499 427 306560 527
rect 306610 381 306676 491
rect 306493 315 306676 381
rect 306710 325 306794 527
rect 305699 73 305769 107
rect 305813 73 305971 107
rect 306031 17 306105 117
rect 306141 107 306185 153
rect 306219 141 306339 207
rect 306383 265 306453 281
rect 306639 265 306676 315
rect 306383 199 306605 265
rect 306639 199 306796 265
rect 306383 107 306427 199
rect 306639 165 306676 199
rect 306141 73 306243 107
rect 306299 73 306427 107
rect 306472 17 306556 123
rect 306603 60 306676 165
rect 306710 17 306794 139
rect 306838 51 306894 491
rect 306934 323 306968 527
rect 307022 265 307088 485
rect 307134 299 307255 527
rect 307022 199 307264 265
rect 306932 17 306978 138
rect 307022 69 307072 199
rect 307129 17 307255 161
rect 307299 53 307353 465
rect 307393 279 307427 527
rect 307481 294 307539 527
rect 307592 393 307626 493
rect 307660 427 307736 527
rect 307592 359 307735 393
rect 307575 195 307645 325
rect 307393 17 307427 191
rect 307481 17 307539 162
rect 307689 161 307735 359
rect 307591 127 307735 161
rect 307591 69 307625 127
rect 307659 17 307735 93
rect 307779 69 307825 493
rect 307863 415 307918 489
rect 307952 449 308028 527
rect 308135 449 308334 483
rect 307863 372 308264 415
rect 307863 89 307897 372
rect 307932 157 307999 337
rect 308033 225 308067 372
rect 308105 271 308186 337
rect 308222 271 308264 372
rect 308300 399 308334 449
rect 308378 433 308412 527
rect 308469 413 308516 488
rect 308565 438 308802 472
rect 308469 399 308503 413
rect 308300 365 308503 399
rect 308033 191 308099 225
rect 308223 157 308257 223
rect 308301 207 308375 331
rect 308469 173 308503 365
rect 307932 123 308257 157
rect 308301 139 308503 173
rect 308537 207 308595 381
rect 308633 331 308731 402
rect 308765 315 308802 438
rect 308836 367 308870 527
rect 308765 297 308893 315
rect 308697 263 308893 297
rect 308537 141 308663 207
rect 308301 89 308335 139
rect 308469 107 308503 139
rect 308697 107 308731 263
rect 308927 219 308968 493
rect 309006 433 309213 467
rect 309002 249 309050 393
rect 308765 153 308968 219
rect 309103 207 309145 381
rect 307863 55 307937 89
rect 307971 17 308037 89
rect 308170 55 308335 89
rect 308379 17 308419 105
rect 308469 73 308539 107
rect 308583 73 308731 107
rect 308801 17 308875 117
rect 308911 107 308968 153
rect 309006 141 309145 207
rect 309179 265 309213 433
rect 309249 427 309310 527
rect 309380 381 309437 491
rect 309247 315 309437 381
rect 309474 325 309508 527
rect 309400 265 309437 315
rect 309542 309 309650 479
rect 309179 199 309366 265
rect 309400 199 309562 265
rect 309179 107 309213 199
rect 309400 165 309436 199
rect 308911 73 309008 107
rect 309047 73 309213 107
rect 309247 17 309310 123
rect 309364 60 309436 165
rect 309602 164 309650 309
rect 309689 294 309747 527
rect 309800 393 309834 493
rect 309868 427 309944 527
rect 309800 359 309943 393
rect 309783 195 309853 325
rect 309474 17 309508 139
rect 309542 61 309650 164
rect 309689 17 309747 162
rect 309897 161 309943 359
rect 309799 127 309943 161
rect 309799 69 309833 127
rect 309867 17 309943 93
rect 309987 69 310033 493
rect 310071 415 310126 489
rect 310160 449 310236 527
rect 310343 449 310542 483
rect 310071 372 310469 415
rect 310071 89 310105 372
rect 310140 157 310207 337
rect 310241 225 310275 372
rect 310313 271 310394 337
rect 310430 271 310469 372
rect 310508 399 310542 449
rect 310586 433 310620 527
rect 310677 413 310724 488
rect 310773 438 311017 472
rect 310677 399 310711 413
rect 310508 365 310711 399
rect 310241 191 310307 225
rect 310431 157 310465 223
rect 310509 207 310583 331
rect 310677 173 310711 365
rect 310140 123 310465 157
rect 310509 139 310711 173
rect 310745 207 310803 381
rect 310841 331 310939 402
rect 310973 315 311017 438
rect 311051 367 311085 527
rect 311119 427 311179 493
rect 311224 433 311431 467
rect 310973 297 311085 315
rect 310909 249 311085 297
rect 310745 141 310871 207
rect 310509 89 310543 139
rect 310677 107 310711 139
rect 310909 107 310943 249
rect 311119 213 311163 427
rect 311197 249 311245 393
rect 311279 315 311353 381
rect 310977 153 311163 213
rect 311279 207 311317 315
rect 311397 281 311431 433
rect 311477 427 311538 527
rect 311608 381 311665 491
rect 311475 315 311665 381
rect 311702 325 311736 527
rect 310071 55 310145 89
rect 310189 17 310255 89
rect 310378 55 310543 89
rect 310587 17 310627 105
rect 310677 73 310747 107
rect 310791 73 310943 107
rect 311009 17 311083 117
rect 311119 107 311163 153
rect 311197 141 311317 207
rect 311361 265 311431 281
rect 311628 265 311665 315
rect 311770 309 311864 479
rect 311898 369 311932 527
rect 311361 199 311594 265
rect 311628 199 311790 265
rect 311361 107 311405 199
rect 311628 165 311664 199
rect 311119 73 311221 107
rect 311277 73 311405 107
rect 311454 17 311538 123
rect 311592 60 311664 165
rect 311830 164 311864 309
rect 311989 294 312047 527
rect 312100 393 312134 493
rect 312168 427 312244 527
rect 312100 359 312243 393
rect 312083 195 312153 325
rect 311702 17 311736 139
rect 311770 61 311864 164
rect 311898 17 311932 113
rect 311989 17 312047 162
rect 312197 161 312243 359
rect 312099 127 312243 161
rect 312099 69 312133 127
rect 312167 17 312243 93
rect 312287 69 312333 493
rect 312371 415 312426 489
rect 312460 449 312536 527
rect 312643 449 312842 483
rect 312371 372 312769 415
rect 312371 89 312405 372
rect 312440 157 312507 337
rect 312541 225 312575 372
rect 312613 271 312694 337
rect 312730 271 312769 372
rect 312808 399 312842 449
rect 312886 433 312920 527
rect 312977 413 313024 488
rect 313073 438 313317 472
rect 312977 399 313011 413
rect 312808 365 313011 399
rect 312541 191 312607 225
rect 312731 157 312765 223
rect 312809 207 312883 331
rect 312977 173 313011 365
rect 312440 123 312765 157
rect 312809 139 313011 173
rect 313045 207 313103 381
rect 313141 331 313239 402
rect 313273 315 313317 438
rect 313351 367 313385 527
rect 313419 427 313479 493
rect 313524 433 313731 467
rect 313273 297 313385 315
rect 313209 249 313385 297
rect 313045 141 313171 207
rect 312809 89 312843 139
rect 312977 107 313011 139
rect 313209 107 313243 249
rect 313419 213 313463 427
rect 313497 249 313545 393
rect 313579 315 313653 381
rect 313277 153 313463 213
rect 313579 207 313617 315
rect 313697 281 313731 433
rect 313777 427 313838 527
rect 313908 381 313965 491
rect 313775 315 313965 381
rect 314002 325 314036 527
rect 314070 335 314146 479
rect 314192 369 314226 527
rect 314260 335 314336 479
rect 314380 369 314414 527
rect 312371 55 312445 89
rect 312489 17 312555 89
rect 312678 55 312843 89
rect 312887 17 312927 105
rect 312977 73 313047 107
rect 313091 73 313243 107
rect 313309 17 313383 117
rect 313419 107 313463 153
rect 313497 141 313617 207
rect 313661 265 313731 281
rect 313928 265 313965 315
rect 314070 301 314434 335
rect 313661 199 313894 265
rect 313928 215 314340 265
rect 313661 107 313705 199
rect 313928 165 313964 215
rect 314374 181 314434 301
rect 314473 294 314531 527
rect 314565 367 314617 527
rect 314651 425 314804 493
rect 314870 425 315008 493
rect 314565 191 314614 333
rect 313419 73 313521 107
rect 313577 73 313705 107
rect 313754 17 313838 123
rect 313892 60 313964 165
rect 314070 147 314434 181
rect 314002 17 314036 139
rect 314070 61 314146 147
rect 314192 17 314226 113
rect 314260 61 314336 147
rect 314380 17 314414 113
rect 314473 17 314531 162
rect 314651 157 314685 425
rect 314719 191 314795 391
rect 314841 241 314940 391
rect 314974 275 315008 425
rect 315052 415 315169 527
rect 315213 417 315257 493
rect 315325 451 315695 527
rect 315739 417 315773 493
rect 315825 451 315891 527
rect 315213 383 315695 417
rect 315213 381 315257 383
rect 315042 327 315257 381
rect 315042 315 315081 327
rect 314974 241 315189 275
rect 314565 123 314807 157
rect 314841 141 314908 241
rect 314942 141 315009 207
rect 315043 199 315189 241
rect 314565 51 314617 123
rect 314651 17 314727 89
rect 314771 51 314807 123
rect 315043 107 315077 199
rect 314841 51 315077 107
rect 315130 17 315164 165
rect 315223 51 315257 327
rect 315295 315 315377 349
rect 315295 187 315329 315
rect 315421 299 315591 349
rect 315421 255 315458 299
rect 315363 221 315458 255
rect 315295 51 315361 187
rect 315424 157 315458 221
rect 315497 199 315560 265
rect 315625 199 315695 383
rect 315739 299 315911 417
rect 315739 199 315827 265
rect 315877 157 315911 299
rect 315424 123 315591 157
rect 315405 17 315471 89
rect 315541 51 315591 123
rect 315655 123 315911 157
rect 315655 51 315689 123
rect 315813 17 315885 89
rect 315945 51 315995 493
rect 316037 294 316095 527
rect 316129 367 316181 527
rect 316215 425 316368 493
rect 316434 425 316572 493
rect 316129 191 316178 333
rect 316037 17 316095 162
rect 316215 157 316256 425
rect 316290 191 316371 391
rect 316405 241 316504 391
rect 316538 275 316572 425
rect 316616 415 316733 527
rect 316777 417 316821 493
rect 316889 451 317263 527
rect 317307 417 317341 493
rect 317391 451 317457 527
rect 316777 383 317263 417
rect 316777 381 316821 383
rect 316606 327 316821 381
rect 316606 315 316645 327
rect 316538 241 316753 275
rect 316129 123 316371 157
rect 316405 141 316472 241
rect 316506 141 316573 207
rect 316607 199 316753 241
rect 316129 51 316181 123
rect 316215 17 316291 89
rect 316335 51 316371 123
rect 316607 107 316641 199
rect 316405 51 316641 107
rect 316694 17 316728 165
rect 316787 51 316821 327
rect 316859 315 316941 349
rect 316859 187 316893 315
rect 316985 299 317155 349
rect 316985 255 317046 299
rect 316927 221 317046 255
rect 316859 153 316944 187
rect 316988 157 317046 221
rect 317105 199 317149 265
rect 317193 199 317263 383
rect 317307 299 317462 417
rect 317307 199 317393 265
rect 317428 263 317462 299
rect 317506 331 317556 493
rect 317600 365 317650 527
rect 317506 297 317647 331
rect 317428 211 317566 263
rect 317428 157 317462 211
rect 317610 177 317647 297
rect 317693 294 317751 527
rect 317785 367 317837 527
rect 317871 425 318040 493
rect 318074 425 318249 493
rect 317785 191 317837 333
rect 316859 51 316925 153
rect 316988 123 317129 157
rect 316969 17 317035 89
rect 317079 51 317129 123
rect 317213 123 317462 157
rect 317506 143 317647 177
rect 317213 51 317247 123
rect 317506 89 317546 143
rect 317379 17 317446 89
rect 317480 51 317546 89
rect 317590 17 317624 109
rect 317693 17 317751 162
rect 317871 157 317915 425
rect 317949 289 318036 391
rect 317949 191 318027 289
rect 318070 265 318171 391
rect 318061 241 318171 265
rect 318215 275 318249 425
rect 318283 415 318421 527
rect 318465 417 318509 493
rect 318547 451 318951 527
rect 318995 417 319029 493
rect 319079 451 319145 527
rect 318465 383 318951 417
rect 318465 381 318509 383
rect 318283 327 318509 381
rect 318283 315 318327 327
rect 318215 241 318421 275
rect 317785 123 318027 157
rect 318061 141 318139 241
rect 318173 141 318240 207
rect 318274 199 318421 241
rect 317785 51 317837 123
rect 317871 17 317947 89
rect 317991 51 318027 123
rect 318274 107 318308 199
rect 318061 51 318308 107
rect 318352 17 318421 165
rect 318465 51 318509 327
rect 318547 315 318629 349
rect 318547 187 318581 315
rect 318673 299 318843 349
rect 318673 255 318734 299
rect 318615 221 318734 255
rect 318547 153 318632 187
rect 318676 157 318734 221
rect 318779 199 318837 265
rect 318881 199 318951 383
rect 318995 299 319150 417
rect 318995 199 319081 265
rect 319116 263 319150 299
rect 319194 331 319244 493
rect 319288 365 319338 527
rect 319194 297 319332 331
rect 319298 263 319332 297
rect 319409 263 319487 493
rect 319521 297 319575 527
rect 319625 294 319683 527
rect 319735 393 319769 493
rect 319803 427 319879 527
rect 319735 359 319879 393
rect 319116 211 319254 263
rect 319298 211 319579 263
rect 319116 157 319150 211
rect 319298 177 319332 211
rect 318547 51 318613 153
rect 318676 123 318817 157
rect 318647 17 318723 89
rect 318767 51 318817 123
rect 318851 123 319150 157
rect 319194 143 319332 177
rect 318851 51 318935 123
rect 319194 89 319244 143
rect 318969 17 319134 89
rect 319168 51 319244 89
rect 319288 17 319338 109
rect 319409 51 319487 211
rect 319719 195 319789 325
rect 319521 17 319575 177
rect 319625 17 319683 162
rect 319833 161 319879 359
rect 319735 127 319879 161
rect 319735 69 319769 127
rect 319803 17 319879 93
rect 319923 69 319957 493
rect 319991 378 320077 493
rect 320177 378 320253 527
rect 319991 103 320025 378
rect 320291 344 320357 485
rect 320403 365 320442 527
rect 320585 404 320661 493
rect 320707 442 320773 493
rect 320585 364 320673 404
rect 320059 153 320131 344
rect 320165 237 320205 274
rect 320239 271 320357 344
rect 320165 153 320253 237
rect 320296 235 320357 271
rect 320521 264 320605 330
rect 320296 169 320477 235
rect 319991 51 320077 103
rect 320177 17 320253 103
rect 320296 51 320341 169
rect 320521 137 320555 264
rect 320639 230 320673 364
rect 320589 196 320673 230
rect 320717 357 320773 442
rect 320858 401 320926 493
rect 320970 435 321039 527
rect 321192 430 321258 493
rect 321300 435 321538 475
rect 320858 367 321174 401
rect 320377 17 320453 122
rect 320589 51 320653 196
rect 320717 165 320751 357
rect 320821 221 320877 323
rect 320911 187 320945 367
rect 320989 221 321090 333
rect 321124 271 321174 367
rect 321208 373 321258 430
rect 321208 237 321242 373
rect 320699 129 320751 165
rect 320699 51 320739 129
rect 320879 103 320945 187
rect 320773 51 320945 103
rect 320989 17 321039 181
rect 321160 113 321242 237
rect 321276 225 321323 344
rect 321357 331 321460 401
rect 321357 191 321391 331
rect 321494 315 321538 435
rect 321572 367 321619 527
rect 321494 297 321619 315
rect 321280 147 321391 191
rect 321439 263 321619 297
rect 321439 113 321473 263
rect 321585 249 321619 263
rect 321653 275 321729 493
rect 321771 421 321829 527
rect 321952 433 322175 471
rect 321511 213 321561 219
rect 321653 213 321846 275
rect 321925 249 321973 393
rect 321511 209 321846 213
rect 321511 153 321744 209
rect 322007 207 322081 399
rect 321160 51 321284 113
rect 321328 51 321473 113
rect 321536 17 321615 112
rect 321653 51 321744 153
rect 321975 141 322081 207
rect 321790 17 321845 123
rect 322125 107 322175 433
rect 322219 299 322253 527
rect 321982 66 322175 107
rect 322209 17 322258 180
rect 322292 51 322363 493
rect 322421 244 322489 493
rect 322533 293 322580 527
rect 322397 178 322489 244
rect 322523 214 322589 259
rect 322421 51 322489 178
rect 322533 17 322580 180
rect 322631 51 322714 484
rect 322753 294 322811 527
rect 322863 393 322897 493
rect 322931 427 323007 527
rect 322863 359 323007 393
rect 322847 195 322917 325
rect 322753 17 322811 162
rect 322961 161 323007 359
rect 322863 127 323007 161
rect 322863 69 322897 127
rect 322931 17 323007 93
rect 323051 69 323085 493
rect 323119 378 323205 493
rect 323305 378 323381 527
rect 323119 103 323153 378
rect 323419 344 323485 485
rect 323531 365 323570 527
rect 323713 404 323789 493
rect 323835 442 323901 493
rect 323713 364 323801 404
rect 323187 153 323259 344
rect 323293 237 323333 274
rect 323367 271 323485 344
rect 323293 153 323381 237
rect 323424 235 323485 271
rect 323649 264 323733 330
rect 323424 169 323605 235
rect 323119 51 323205 103
rect 323305 17 323381 103
rect 323424 51 323469 169
rect 323649 137 323683 264
rect 323767 230 323801 364
rect 323717 196 323801 230
rect 323845 357 323901 442
rect 323986 401 324054 493
rect 324098 435 324167 527
rect 324320 430 324386 493
rect 324428 435 324666 475
rect 323986 367 324302 401
rect 323505 17 323581 122
rect 323717 51 323781 196
rect 323845 165 323879 357
rect 323949 221 324005 323
rect 324039 187 324073 367
rect 324117 221 324218 333
rect 324252 271 324302 367
rect 324336 373 324386 430
rect 324336 237 324370 373
rect 323827 129 323879 165
rect 323827 51 323867 129
rect 324007 103 324073 187
rect 323901 51 324073 103
rect 324117 17 324167 181
rect 324288 113 324370 237
rect 324404 225 324451 344
rect 324485 331 324588 401
rect 324485 191 324519 331
rect 324622 315 324666 435
rect 324700 367 324747 527
rect 324622 297 324747 315
rect 324408 147 324519 191
rect 324567 263 324747 297
rect 324567 113 324601 263
rect 324713 249 324747 263
rect 324781 275 324857 493
rect 324899 421 324957 527
rect 325080 433 325303 471
rect 324639 213 324689 219
rect 324781 213 324974 275
rect 325053 249 325101 393
rect 324639 209 324974 213
rect 324639 153 324872 209
rect 325135 207 325209 399
rect 324288 51 324412 113
rect 324456 51 324601 113
rect 324664 17 324743 112
rect 324781 51 324872 153
rect 325106 141 325209 207
rect 324918 17 324973 123
rect 325253 107 325303 433
rect 325347 299 325381 527
rect 325415 260 325491 493
rect 325535 293 325585 527
rect 325619 315 325665 402
rect 325415 213 325514 260
rect 325699 244 325767 493
rect 325811 293 325858 527
rect 325110 66 325303 107
rect 325354 17 325404 180
rect 325448 51 325514 213
rect 325558 17 325608 180
rect 325642 178 325767 244
rect 325699 51 325767 178
rect 325811 17 325858 180
rect 325892 51 325968 484
rect 326012 293 326064 527
rect 326157 294 326215 527
rect 326249 425 326309 527
rect 326343 391 326419 493
rect 326463 425 326599 527
rect 326735 425 326811 459
rect 326855 425 326915 527
rect 326777 391 326811 425
rect 326249 357 326743 391
rect 326012 17 326064 180
rect 326249 165 326283 357
rect 326317 289 326665 323
rect 326317 199 326394 289
rect 326428 215 326587 255
rect 326621 249 326665 289
rect 326699 317 326743 357
rect 326777 351 326951 391
rect 326699 283 326851 317
rect 326621 215 326761 249
rect 326807 199 326851 283
rect 326157 17 326215 162
rect 326249 56 326342 165
rect 326463 17 326497 181
rect 326903 165 326951 351
rect 326985 294 327043 527
rect 327077 393 327140 493
rect 327184 427 327234 527
rect 327278 393 327328 493
rect 327372 427 327422 527
rect 327466 393 327516 493
rect 327578 425 327628 493
rect 327672 427 327722 527
rect 327766 459 328011 493
rect 327766 425 327831 459
rect 327961 427 328011 459
rect 328065 427 328115 527
rect 327077 391 327516 393
rect 327875 393 327917 425
rect 328159 393 328209 425
rect 327077 357 327816 391
rect 327875 359 328209 393
rect 328253 359 328328 527
rect 326531 131 326811 165
rect 326531 51 326607 131
rect 326651 17 326731 95
rect 326765 51 326811 131
rect 326867 69 326951 165
rect 327077 179 327123 357
rect 327782 325 327816 357
rect 328159 325 328209 359
rect 327228 289 327730 323
rect 327782 291 328101 325
rect 327228 257 327262 289
rect 327157 215 327262 257
rect 327696 257 327730 289
rect 327331 215 327641 255
rect 327696 215 327921 257
rect 328067 249 328101 291
rect 328159 283 328328 325
rect 328365 294 328423 527
rect 328457 323 328532 493
rect 328576 367 328626 527
rect 328670 401 328720 493
rect 328764 435 328814 527
rect 328858 401 328908 493
rect 328952 435 329002 527
rect 329046 401 329096 493
rect 329140 435 329190 527
rect 329234 401 329284 493
rect 328670 357 329284 401
rect 329325 401 329388 493
rect 329432 435 329482 527
rect 329526 401 329576 493
rect 329620 435 329670 527
rect 329714 443 330148 493
rect 329714 401 329756 443
rect 330186 409 330252 493
rect 329325 357 329756 401
rect 329790 357 330252 409
rect 330288 367 330338 527
rect 328670 323 328720 357
rect 330186 333 330252 357
rect 330382 333 330432 493
rect 330476 367 330526 527
rect 330562 333 330628 493
rect 328067 215 328209 249
rect 326985 17 327043 162
rect 327077 129 327242 179
rect 327286 145 327524 181
rect 327286 95 327336 145
rect 327081 51 327336 95
rect 327380 17 327414 111
rect 327448 51 327524 145
rect 327586 17 327620 181
rect 327654 145 328211 181
rect 327654 51 327730 145
rect 327774 17 327808 111
rect 327842 51 327925 145
rect 328141 129 328211 145
rect 327969 17 328003 111
rect 328250 95 328328 283
rect 328457 289 328720 323
rect 328807 289 329694 323
rect 329738 289 330152 323
rect 330186 289 330628 333
rect 330665 294 330723 527
rect 328457 181 328504 289
rect 328807 255 328841 289
rect 329660 255 329694 289
rect 330118 255 330152 289
rect 328538 215 328841 255
rect 328915 215 329626 255
rect 329660 215 330074 255
rect 330118 215 330547 255
rect 330581 181 330628 289
rect 328057 61 328328 95
rect 328365 17 328423 162
rect 328457 129 328822 181
rect 328866 145 329292 181
rect 328866 95 328916 145
rect 328474 51 328916 95
rect 328960 17 328994 111
rect 329028 51 329104 145
rect 329148 17 329182 111
rect 329216 51 329292 145
rect 329326 17 329380 181
rect 329414 147 330236 181
rect 329414 145 330074 147
rect 329414 51 329490 145
rect 329534 17 329568 111
rect 329602 51 329678 145
rect 329722 17 329756 111
rect 329790 51 329866 145
rect 329910 17 329944 111
rect 329978 51 330054 145
rect 330098 17 330132 111
rect 330186 95 330236 147
rect 330270 131 330628 181
rect 330757 288 330813 493
rect 330847 443 330924 527
rect 330960 447 331274 481
rect 331425 447 331491 527
rect 331578 455 332237 489
rect 332323 455 332459 527
rect 330960 409 331004 447
rect 331578 413 331612 455
rect 330847 375 331004 409
rect 331072 379 331612 413
rect 330186 61 330628 95
rect 330665 17 330723 162
rect 330757 70 330809 288
rect 330847 266 330891 375
rect 330937 307 331274 341
rect 330843 173 330891 266
rect 330843 139 330981 173
rect 330843 17 330903 105
rect 330937 85 330981 139
rect 331015 119 331049 307
rect 331240 265 331274 307
rect 331318 305 331395 339
rect 331339 275 331395 305
rect 331083 215 331206 265
rect 331240 199 331305 265
rect 331109 159 331185 181
rect 331339 159 331373 275
rect 331429 241 331463 379
rect 331509 289 331613 343
rect 331109 125 331373 159
rect 331407 207 331463 241
rect 331407 91 331441 207
rect 331174 85 331271 91
rect 330937 51 331271 85
rect 331315 57 331441 91
rect 331475 17 331509 173
rect 331555 83 331613 289
rect 331649 119 331683 421
rect 331717 178 331751 455
rect 332503 421 332562 493
rect 331797 323 331880 409
rect 331997 387 332562 421
rect 331797 289 331963 323
rect 331800 199 331885 254
rect 331717 165 331769 178
rect 331717 144 331809 165
rect 331725 131 331809 144
rect 331649 97 331691 119
rect 331649 53 331731 97
rect 331775 64 331809 131
rect 331843 126 331885 199
rect 331929 85 331963 289
rect 331997 119 332031 387
rect 332455 375 332562 387
rect 332065 289 332191 323
rect 332235 299 332472 341
rect 332065 199 332109 289
rect 332438 265 332472 299
rect 332143 189 332205 255
rect 332239 215 332383 265
rect 332438 199 332494 265
rect 332143 146 332184 189
rect 332438 181 332472 199
rect 332251 150 332472 181
rect 332243 147 332472 150
rect 332065 85 332168 93
rect 331929 51 332168 85
rect 332243 59 332301 147
rect 332528 117 332562 375
rect 332597 294 332655 527
rect 332689 298 332747 527
rect 332350 17 332442 113
rect 332502 51 332562 117
rect 332597 17 332655 162
rect 332689 17 332747 147
rect 332781 70 332845 493
rect 332881 443 332958 527
rect 332994 447 333308 481
rect 333459 447 333525 527
rect 333612 455 334271 489
rect 334363 455 334430 527
rect 332994 409 333038 447
rect 333612 413 333646 455
rect 332881 375 333038 409
rect 333106 379 333646 413
rect 332881 173 332925 375
rect 332971 307 333308 341
rect 332881 139 333015 173
rect 332879 17 332937 105
rect 332971 85 333015 139
rect 333049 119 333083 307
rect 333274 265 333308 307
rect 333352 305 333429 339
rect 333373 275 333429 305
rect 333117 215 333240 265
rect 333274 199 333339 265
rect 333143 159 333219 181
rect 333373 159 333407 275
rect 333463 241 333497 379
rect 333543 289 333647 343
rect 333143 125 333407 159
rect 333441 207 333497 241
rect 333441 91 333475 207
rect 333208 85 333305 91
rect 332971 51 333305 85
rect 333349 57 333475 91
rect 333509 17 333543 173
rect 333589 83 333647 289
rect 333683 119 333717 421
rect 333751 178 333785 455
rect 334510 421 334569 493
rect 333831 323 333914 409
rect 334031 387 334569 421
rect 333831 289 333997 323
rect 333834 199 333919 254
rect 333751 165 333803 178
rect 333751 144 333843 165
rect 333759 131 333843 144
rect 333683 97 333725 119
rect 333683 53 333765 97
rect 333809 64 333843 131
rect 333877 126 333919 199
rect 333963 85 333997 289
rect 334031 119 334065 387
rect 334462 375 334569 387
rect 334099 289 334225 323
rect 334269 299 334479 341
rect 334099 199 334143 289
rect 334445 265 334479 299
rect 334177 189 334239 255
rect 334283 215 334411 265
rect 334445 199 334501 265
rect 334177 146 334218 189
rect 334445 181 334479 199
rect 334285 150 334479 181
rect 334277 147 334479 150
rect 334099 85 334202 93
rect 333963 51 334202 85
rect 334277 59 334335 147
rect 334535 117 334569 375
rect 334621 294 334679 527
rect 334753 298 334787 527
rect 334821 265 334897 485
rect 334941 299 334975 527
rect 335009 288 335075 493
rect 335109 443 335186 527
rect 335222 447 335536 481
rect 335687 447 335753 527
rect 335840 455 336499 489
rect 336581 455 336658 527
rect 335222 409 335266 447
rect 335840 413 335874 455
rect 335109 375 335266 409
rect 335334 379 335874 413
rect 335009 265 335068 288
rect 335109 265 335153 375
rect 335199 307 335536 341
rect 334821 199 335068 265
rect 335102 199 335153 265
rect 334379 17 334413 113
rect 334509 51 334569 117
rect 334621 17 334679 162
rect 334753 17 334787 147
rect 334821 75 334881 199
rect 335009 185 335068 199
rect 334941 17 334975 147
rect 335009 70 335071 185
rect 335108 173 335153 199
rect 335108 139 335243 173
rect 335105 17 335165 105
rect 335199 85 335243 139
rect 335277 119 335311 307
rect 335502 265 335536 307
rect 335580 305 335657 339
rect 335601 275 335657 305
rect 335345 215 335468 265
rect 335502 199 335567 265
rect 335371 159 335447 181
rect 335601 159 335635 275
rect 335691 241 335725 379
rect 335771 289 335875 343
rect 335371 125 335635 159
rect 335669 207 335725 241
rect 335669 91 335703 207
rect 335436 85 335533 91
rect 335199 51 335533 85
rect 335577 57 335703 91
rect 335737 17 335771 173
rect 335817 83 335875 289
rect 335911 97 335945 421
rect 335979 165 336013 455
rect 336702 421 336761 493
rect 336059 323 336142 409
rect 336259 387 336761 421
rect 336059 289 336225 323
rect 336062 199 336147 254
rect 335979 131 336071 165
rect 335911 53 336000 97
rect 336037 64 336071 131
rect 336105 126 336147 199
rect 336191 85 336225 289
rect 336259 119 336293 387
rect 336654 375 336761 387
rect 336327 289 336453 323
rect 336497 299 336671 341
rect 336327 199 336371 289
rect 336637 265 336671 299
rect 336405 189 336467 255
rect 336511 215 336603 265
rect 336637 199 336693 265
rect 336405 146 336446 189
rect 336637 181 336671 199
rect 336513 150 336671 181
rect 336505 147 336671 150
rect 336327 85 336430 93
rect 336191 51 336430 85
rect 336505 59 336563 147
rect 336727 117 336761 375
rect 336829 294 336887 527
rect 336921 357 336997 493
rect 337137 357 337171 527
rect 337205 391 337281 493
rect 337327 425 337361 527
rect 337395 391 337475 493
rect 337205 357 337475 391
rect 336921 165 336955 357
rect 336989 289 337282 323
rect 337549 307 337613 493
rect 336989 199 337059 289
rect 337095 215 337204 255
rect 337248 249 337282 289
rect 337487 273 337613 307
rect 337657 294 337715 527
rect 337756 427 337812 493
rect 337856 427 337906 527
rect 337950 459 338188 493
rect 337950 427 338000 459
rect 338138 427 338188 459
rect 337761 425 337795 427
rect 337965 425 337999 427
rect 338229 425 338292 493
rect 338336 427 338386 527
rect 338044 391 338094 425
rect 338250 391 338292 425
rect 338430 391 338480 493
rect 338524 427 338585 527
rect 338629 459 338971 493
rect 338629 391 338783 459
rect 337756 357 338216 391
rect 338250 357 338783 391
rect 337248 215 337335 249
rect 337407 165 337453 265
rect 336607 17 336641 113
rect 336701 51 336761 117
rect 336829 17 336887 162
rect 336921 131 337453 165
rect 336931 17 336997 95
rect 337041 67 337075 131
rect 337487 97 337521 273
rect 337111 17 337187 95
rect 337280 63 337521 97
rect 337555 17 337613 184
rect 337756 181 337790 357
rect 338182 323 338216 357
rect 338827 325 338877 425
rect 338921 359 338971 459
rect 337883 289 338148 323
rect 338182 289 338769 323
rect 337883 255 337917 289
rect 338104 255 338148 289
rect 337841 215 337917 255
rect 337961 215 338070 255
rect 338104 215 338438 255
rect 338476 215 338630 255
rect 338735 249 338769 289
rect 338827 283 339002 325
rect 339037 294 339095 527
rect 339129 401 339192 493
rect 339236 435 339286 527
rect 339330 401 339380 493
rect 339424 435 339474 527
rect 339518 459 339944 493
rect 339518 401 339568 459
rect 339706 425 339756 459
rect 339129 357 339568 401
rect 339612 391 339662 425
rect 339800 391 339850 425
rect 339612 357 339850 391
rect 339894 359 339944 459
rect 339998 401 340048 493
rect 340092 435 340142 527
rect 340186 401 340236 493
rect 340280 435 340330 527
rect 340374 401 340424 493
rect 340468 435 340518 527
rect 340562 401 340612 493
rect 340656 435 340706 527
rect 340750 459 341188 493
rect 340750 401 340800 459
rect 339998 357 340800 401
rect 339612 323 339646 357
rect 338735 215 338877 249
rect 338929 181 339002 283
rect 337657 17 337715 162
rect 337756 145 338102 181
rect 337770 17 337804 111
rect 337838 51 337914 145
rect 337958 17 337992 111
rect 338026 51 338102 145
rect 338234 145 338472 181
rect 338146 17 338180 111
rect 338234 51 338300 145
rect 338344 17 338378 111
rect 338412 95 338472 145
rect 338527 145 339002 181
rect 339129 289 339646 323
rect 339688 289 340475 323
rect 340562 291 340612 357
rect 340848 333 340906 425
rect 340950 367 341000 459
rect 341044 333 341094 425
rect 341138 359 341188 459
rect 340848 325 341094 333
rect 341222 325 341303 493
rect 340714 289 340814 323
rect 340848 289 341303 325
rect 341337 294 341395 527
rect 339129 181 339163 289
rect 339688 255 339732 289
rect 340431 255 340475 289
rect 340780 255 340814 289
rect 339197 215 339732 255
rect 339766 221 340380 255
rect 339766 215 340212 221
rect 340431 215 340736 255
rect 340780 215 341138 255
rect 340242 181 340338 187
rect 341239 181 341303 289
rect 338527 129 338593 145
rect 338809 129 338885 145
rect 338412 51 338688 95
rect 338741 17 338775 111
rect 338929 17 338963 111
rect 339037 17 339095 162
rect 339129 147 339858 181
rect 339218 145 339858 147
rect 339129 17 339184 113
rect 339218 51 339294 145
rect 339338 17 339372 111
rect 339406 51 339482 145
rect 339526 17 339560 111
rect 339594 51 339670 145
rect 339714 17 339748 111
rect 339782 51 339858 145
rect 339902 17 339956 179
rect 340025 129 340338 181
rect 340382 145 340808 181
rect 340842 147 341303 181
rect 341429 288 341534 493
rect 341578 443 341645 527
rect 341682 447 342021 481
rect 342074 447 342155 481
rect 342189 447 342255 527
rect 342342 455 343001 489
rect 343083 455 343222 527
rect 341682 409 341726 447
rect 342121 413 342155 447
rect 342342 413 342376 455
rect 341572 375 341726 409
rect 341806 379 342087 413
rect 342121 379 342376 413
rect 341429 185 341492 288
rect 340842 145 341008 147
rect 340382 95 340432 145
rect 339990 51 340432 95
rect 340476 17 340510 111
rect 340544 51 340620 145
rect 340664 17 340698 111
rect 340732 51 340808 145
rect 340864 17 340898 111
rect 340932 51 341008 145
rect 341052 17 341086 111
rect 341120 51 341196 147
rect 341240 17 341274 111
rect 341337 17 341395 162
rect 341429 70 341530 185
rect 341572 173 341612 375
rect 341659 307 342009 341
rect 341572 139 341702 173
rect 341574 17 341624 105
rect 341658 85 341702 139
rect 341736 119 341770 307
rect 341975 265 342009 307
rect 342053 339 342087 379
rect 342053 305 342159 339
rect 342102 275 342159 305
rect 341804 199 341941 265
rect 341975 199 342040 265
rect 341826 131 342068 165
rect 341910 85 341990 91
rect 341658 51 341990 85
rect 342024 85 342068 131
rect 342102 119 342136 275
rect 342193 241 342227 379
rect 342273 289 342376 343
rect 342170 207 342227 241
rect 342170 85 342204 207
rect 342024 51 342204 85
rect 342238 17 342272 173
rect 342318 83 342376 289
rect 342411 119 342445 421
rect 342479 178 342513 455
rect 343266 421 343325 493
rect 342561 323 342644 409
rect 342761 387 343325 421
rect 342561 289 342727 323
rect 342564 199 342649 254
rect 342479 165 342533 178
rect 342479 144 342572 165
rect 342489 131 342572 144
rect 342411 97 342455 119
rect 342411 53 342494 97
rect 342538 64 342572 131
rect 342606 126 342649 199
rect 342693 85 342727 289
rect 342761 119 342795 387
rect 343218 375 343325 387
rect 342829 289 342955 345
rect 342999 299 343235 341
rect 342829 199 342873 289
rect 343201 265 343235 299
rect 342907 189 342969 255
rect 343013 215 343151 265
rect 343201 199 343257 265
rect 342907 146 342948 189
rect 343201 181 343235 199
rect 343015 150 343235 181
rect 343007 147 343235 150
rect 342829 85 342932 93
rect 342693 51 342932 85
rect 343007 59 343065 147
rect 343291 117 343325 375
rect 343361 294 343419 527
rect 343457 443 343523 527
rect 343567 409 343617 493
rect 343661 443 343728 527
rect 343765 447 344104 481
rect 344157 447 344238 481
rect 344272 447 344338 527
rect 344425 455 345084 489
rect 345166 455 345243 527
rect 343765 409 343809 447
rect 344204 413 344238 447
rect 344425 413 344459 455
rect 343502 288 343617 409
rect 343661 375 343809 409
rect 343889 379 344170 413
rect 344204 379 344459 413
rect 343502 185 343575 288
rect 343661 265 343695 375
rect 343742 307 344092 341
rect 343655 199 343695 265
rect 343109 17 343199 113
rect 343265 51 343325 117
rect 343361 17 343419 162
rect 343502 132 343622 185
rect 343661 173 343695 199
rect 343661 139 343785 173
rect 343457 17 343523 93
rect 343572 70 343622 132
rect 343657 17 343707 105
rect 343741 85 343785 139
rect 343819 119 343853 307
rect 344058 265 344092 307
rect 344136 339 344170 379
rect 344136 305 344242 339
rect 344185 275 344242 305
rect 343887 199 344024 265
rect 344058 199 344123 265
rect 343909 131 344151 165
rect 343993 85 344074 91
rect 343741 51 344074 85
rect 344108 85 344151 131
rect 344185 119 344219 275
rect 344276 241 344310 379
rect 344356 289 344459 343
rect 344253 207 344310 241
rect 344253 85 344287 207
rect 344108 51 344287 85
rect 344321 17 344355 173
rect 344401 83 344459 289
rect 344494 119 344528 421
rect 344562 178 344596 455
rect 345287 421 345346 493
rect 344644 323 344727 409
rect 344844 387 345346 421
rect 344644 289 344810 323
rect 344647 199 344732 254
rect 344562 165 344616 178
rect 344562 144 344655 165
rect 344572 131 344655 144
rect 344494 97 344538 119
rect 344494 53 344577 97
rect 344621 64 344655 131
rect 344689 126 344732 199
rect 344776 85 344810 289
rect 344844 119 344878 387
rect 345239 375 345346 387
rect 344912 289 345038 333
rect 345082 299 345256 341
rect 344912 199 344956 289
rect 345222 265 345256 299
rect 344990 189 345054 255
rect 345096 215 345188 265
rect 345222 199 345278 265
rect 344990 146 345031 189
rect 345222 181 345256 199
rect 345098 150 345256 181
rect 345090 147 345256 150
rect 344912 85 345015 93
rect 344776 51 345015 85
rect 345090 59 345148 147
rect 345312 117 345346 375
rect 345385 294 345443 527
rect 345515 427 345549 527
rect 345609 409 345643 493
rect 345687 443 345753 527
rect 345797 409 345831 493
rect 345875 443 345941 527
rect 345975 447 346303 481
rect 346356 447 346437 481
rect 346471 447 346537 527
rect 346624 455 347283 489
rect 347383 455 347449 527
rect 345975 409 346019 447
rect 346403 413 346437 447
rect 346624 413 346658 455
rect 345609 291 345831 409
rect 345875 375 346019 409
rect 346088 379 346369 413
rect 346403 379 346658 413
rect 345609 288 345774 291
rect 345701 185 345774 288
rect 345875 265 345909 375
rect 345974 307 346291 341
rect 345864 193 345909 265
rect 345192 17 345226 113
rect 345286 51 345346 117
rect 345385 17 345443 162
rect 345589 132 345811 185
rect 345875 173 345909 193
rect 345875 139 345973 173
rect 345495 17 345529 109
rect 345589 70 345623 132
rect 345657 17 345733 93
rect 345777 70 345811 132
rect 345871 17 345905 105
rect 345939 85 345973 139
rect 346018 119 346052 307
rect 346257 265 346291 307
rect 346335 339 346369 379
rect 346335 305 346441 339
rect 346384 275 346441 305
rect 346086 199 346223 265
rect 346257 199 346341 265
rect 346108 131 346350 165
rect 346192 85 346272 91
rect 345939 51 346272 85
rect 346306 85 346350 131
rect 346384 119 346418 275
rect 346475 241 346509 379
rect 346555 289 346658 343
rect 346452 210 346509 241
rect 346452 209 346508 210
rect 346452 208 346506 209
rect 346452 207 346503 208
rect 346452 85 346486 207
rect 346306 51 346486 85
rect 346520 17 346554 177
rect 346600 83 346658 289
rect 346693 119 346727 421
rect 346765 178 346799 455
rect 347493 421 347545 493
rect 346843 323 346926 409
rect 347043 387 347545 421
rect 346843 289 347009 323
rect 346846 199 346931 254
rect 346765 165 346815 178
rect 346765 144 346854 165
rect 346771 131 346854 144
rect 346693 97 346737 119
rect 346693 53 346776 97
rect 346820 64 346854 131
rect 346888 126 346931 199
rect 346975 85 347009 289
rect 347043 119 347077 387
rect 347438 375 347545 387
rect 347111 289 347188 323
rect 347281 299 347455 341
rect 347111 199 347155 289
rect 347421 265 347455 299
rect 347189 189 347251 255
rect 347295 215 347387 265
rect 347421 199 347467 265
rect 347189 146 347230 189
rect 347421 181 347455 199
rect 347297 150 347455 181
rect 347289 147 347455 150
rect 347111 85 347214 93
rect 346975 51 347214 85
rect 347289 59 347347 147
rect 347511 117 347545 375
rect 347593 294 347651 527
rect 347686 393 347737 493
rect 347774 427 347850 527
rect 347686 359 347851 393
rect 347696 195 347766 325
rect 347810 265 347851 359
rect 347895 346 347941 493
rect 348090 417 348144 480
rect 348188 451 348254 527
rect 348090 383 348214 417
rect 347810 199 347873 265
rect 347399 17 347433 113
rect 347493 51 347545 117
rect 347593 17 347651 162
rect 347810 161 347845 199
rect 347687 127 347845 161
rect 347907 135 347941 346
rect 347985 267 348112 349
rect 347985 214 348066 267
rect 348163 237 348214 383
rect 348292 271 348399 493
rect 348442 421 348476 493
rect 348639 455 348709 527
rect 348764 437 348838 487
rect 348764 421 348798 437
rect 348887 427 348960 493
rect 348442 387 348798 421
rect 348163 233 348357 237
rect 348121 199 348357 233
rect 348442 215 348477 387
rect 348121 180 348155 199
rect 347687 69 347737 127
rect 347771 17 347847 93
rect 347891 69 347941 135
rect 348007 146 348155 180
rect 348007 79 348041 146
rect 348075 17 348151 112
rect 348199 17 348275 165
rect 348323 85 348357 199
rect 348401 135 348477 215
rect 348521 85 348555 337
rect 348590 142 348659 340
rect 348696 179 348730 387
rect 348832 315 348892 391
rect 348764 213 348798 279
rect 348848 207 348892 315
rect 348926 277 348960 427
rect 349004 421 349038 475
rect 349095 471 349161 527
rect 349222 421 349256 475
rect 349298 435 349382 527
rect 349004 387 349256 421
rect 349431 401 349465 493
rect 349507 425 349711 493
rect 349751 439 349801 527
rect 349314 367 349465 401
rect 349314 353 349376 367
rect 349060 319 349376 353
rect 349505 333 349637 391
rect 348926 243 349298 277
rect 348696 143 348812 179
rect 348323 51 348555 85
rect 348669 17 348738 108
rect 348778 101 348812 143
rect 348848 141 348998 207
rect 348778 67 348846 101
rect 349036 95 349070 243
rect 349114 153 349230 209
rect 349264 201 349298 243
rect 349342 167 349376 319
rect 348890 61 349070 95
rect 349206 17 349272 109
rect 349314 89 349376 167
rect 349410 332 349637 333
rect 349676 349 349711 425
rect 349850 417 349884 475
rect 349919 451 349995 527
rect 349850 383 350014 417
rect 349410 299 349557 332
rect 349676 315 349942 349
rect 349410 141 349462 299
rect 349676 297 349725 315
rect 349515 184 349549 265
rect 349602 263 349725 297
rect 349980 265 350014 383
rect 350049 299 350099 527
rect 350153 265 350219 465
rect 350263 299 350313 527
rect 350357 265 350407 465
rect 350451 299 350501 527
rect 350537 294 350595 527
rect 350637 393 350693 527
rect 350737 349 350797 459
rect 350847 383 350913 527
rect 350961 383 351053 493
rect 349602 107 349646 263
rect 349698 173 349742 229
rect 349788 213 349942 255
rect 349698 139 349814 173
rect 349314 55 349390 89
rect 349424 51 349646 107
rect 349690 17 349734 105
rect 349780 93 349814 139
rect 349881 127 349942 213
rect 349980 199 350109 265
rect 350153 199 350407 265
rect 350632 265 350685 337
rect 350737 315 350951 349
rect 350632 215 350730 265
rect 350783 215 350867 265
rect 349980 93 350015 199
rect 349780 59 350015 93
rect 350049 17 350083 109
rect 350153 53 350219 199
rect 350263 17 350297 109
rect 350357 53 350407 199
rect 350917 181 350951 315
rect 350451 17 350485 109
rect 350537 17 350595 162
rect 350637 143 350951 181
rect 350637 71 350703 143
rect 351003 109 351053 383
rect 351089 294 351147 527
rect 351199 403 351233 489
rect 351267 437 351343 527
rect 351199 357 351343 403
rect 350847 17 350897 109
rect 350931 51 351053 109
rect 351089 17 351147 162
rect 351193 153 351253 323
rect 351293 227 351343 357
rect 351377 295 351431 484
rect 351477 433 351629 527
rect 351465 329 351531 391
rect 351665 316 351780 473
rect 351377 265 351541 295
rect 351377 261 351659 265
rect 351293 161 351400 227
rect 351434 189 351659 261
rect 351182 17 351249 118
rect 351293 56 351341 161
rect 351434 122 351482 189
rect 351745 155 351780 316
rect 351825 294 351883 527
rect 351918 299 351969 527
rect 352008 417 352279 483
rect 352029 265 352063 377
rect 352108 333 352192 383
rect 352325 367 352381 527
rect 352108 299 352401 333
rect 352435 299 352516 493
rect 351918 215 351985 265
rect 352029 199 352177 265
rect 352029 181 352079 199
rect 351397 83 351482 122
rect 351397 54 351431 83
rect 351578 17 351644 116
rect 351688 51 351780 155
rect 351825 17 351883 162
rect 351922 147 352079 181
rect 352367 165 352401 299
rect 351922 53 351984 147
rect 352231 131 352401 165
rect 352482 152 352516 299
rect 352561 294 352619 527
rect 352666 333 352744 368
rect 352873 367 352939 527
rect 352995 369 353079 493
rect 352666 299 352977 333
rect 352028 17 352175 113
rect 352231 61 352265 131
rect 352299 17 352385 97
rect 352435 83 352516 152
rect 352561 17 352619 162
rect 352653 153 352724 265
rect 352758 119 352802 299
rect 352836 153 352899 265
rect 352943 199 352977 299
rect 353016 165 353079 369
rect 353113 294 353171 527
rect 353271 336 353323 381
rect 353373 371 353439 527
rect 353539 370 353629 493
rect 353271 302 353559 336
rect 352674 17 352722 119
rect 352758 53 352824 119
rect 352880 17 352923 119
rect 352969 51 353079 165
rect 353113 17 353171 162
rect 353208 145 353253 265
rect 353287 109 353323 302
rect 353390 213 353473 265
rect 353515 197 353559 302
rect 353254 74 353323 109
rect 353369 17 353411 179
rect 353593 163 353629 370
rect 353665 294 353723 527
rect 353757 331 353821 493
rect 353865 365 353915 527
rect 353959 459 354205 493
rect 353959 331 354009 459
rect 353757 289 354009 331
rect 353836 213 353934 255
rect 354045 179 354103 425
rect 354147 378 354205 459
rect 354147 289 354198 378
rect 354259 323 354293 492
rect 354345 429 354395 527
rect 354232 289 354293 323
rect 354232 249 354266 289
rect 354408 255 354451 393
rect 354493 294 354551 527
rect 354585 333 354641 493
rect 354675 367 354751 527
rect 354795 333 354829 493
rect 354863 367 354923 527
rect 354957 459 355419 493
rect 354957 333 355033 459
rect 354585 291 355033 333
rect 355077 349 355111 425
rect 355145 387 355221 459
rect 355265 349 355299 425
rect 355077 289 355299 349
rect 355333 315 355419 459
rect 355453 315 355519 493
rect 354155 215 354266 249
rect 354223 179 354266 215
rect 354300 213 354451 255
rect 354640 215 354958 255
rect 355077 181 355143 289
rect 355453 255 355503 315
rect 355563 299 355644 527
rect 355689 294 355747 527
rect 355789 291 355833 527
rect 355867 291 355953 493
rect 355997 291 356056 527
rect 356099 333 356163 493
rect 356207 367 356257 527
rect 356301 333 356351 493
rect 356395 367 356445 527
rect 356489 333 356539 493
rect 356583 367 356633 527
rect 356677 333 356727 493
rect 356771 367 356821 527
rect 356865 459 357667 493
rect 356865 333 356915 459
rect 356099 291 356915 333
rect 356959 323 357009 425
rect 357053 357 357103 459
rect 357147 323 357197 425
rect 357241 357 357291 459
rect 357335 323 357385 425
rect 357429 357 357479 459
rect 357523 323 357573 425
rect 357617 357 357667 459
rect 355187 215 355503 255
rect 355537 215 355653 264
rect 355909 257 355953 291
rect 356959 289 357677 323
rect 357713 294 357771 527
rect 357848 299 357891 527
rect 357925 299 358011 493
rect 353445 129 353629 163
rect 353445 51 353515 129
rect 353549 17 353615 95
rect 353665 17 353723 162
rect 353757 17 353813 179
rect 353847 145 354111 179
rect 353847 51 353923 145
rect 353967 17 354001 111
rect 354035 51 354111 145
rect 354155 17 354189 179
rect 354223 145 354293 179
rect 354259 89 354293 145
rect 354345 17 354396 169
rect 354493 17 354551 162
rect 354585 17 354641 181
rect 354675 145 355315 181
rect 354675 51 354751 145
rect 354795 17 354829 111
rect 354863 51 354939 145
rect 354983 17 355017 111
rect 355051 51 355127 145
rect 355171 17 355205 111
rect 355239 51 355315 145
rect 355359 17 355417 181
rect 355453 163 355503 215
rect 355781 213 355865 257
rect 355909 215 356868 257
rect 356922 215 357540 255
rect 355909 213 356011 215
rect 355453 51 355519 163
rect 355563 17 355621 181
rect 355689 17 355747 162
rect 355781 51 355827 213
rect 355861 17 355905 179
rect 355939 51 356011 213
rect 357574 181 357677 289
rect 356053 17 356155 181
rect 356189 145 357677 181
rect 357805 199 357921 265
rect 357965 257 358011 299
rect 358055 291 358099 527
rect 358133 257 358219 493
rect 358263 291 358322 527
rect 358363 333 358427 493
rect 358471 367 358521 527
rect 358565 333 358615 493
rect 358659 367 358709 527
rect 358753 333 358803 493
rect 358847 367 358897 527
rect 358941 333 358991 493
rect 359035 367 359085 527
rect 359129 333 359179 493
rect 359223 367 359273 527
rect 359317 333 359367 493
rect 359411 367 359461 527
rect 359505 333 359555 493
rect 359599 367 359649 527
rect 359693 333 359743 493
rect 359787 367 359837 527
rect 359881 459 361435 493
rect 359881 333 359931 459
rect 358363 291 359931 333
rect 359975 325 360025 425
rect 360069 359 360119 459
rect 360163 325 360213 425
rect 360257 359 360307 459
rect 360351 325 360401 425
rect 360445 359 360495 459
rect 360539 325 360589 425
rect 360633 359 360683 459
rect 360727 325 360777 425
rect 360821 359 360871 459
rect 360915 325 360965 425
rect 361009 359 361059 459
rect 361103 325 361153 425
rect 361197 359 361247 459
rect 361291 325 361341 425
rect 361385 359 361435 459
rect 359975 291 361449 325
rect 361485 294 361543 527
rect 361577 309 361819 527
rect 357965 215 359884 257
rect 359918 215 361308 257
rect 357965 213 358265 215
rect 356189 51 356265 145
rect 356309 17 356343 111
rect 356377 51 356453 145
rect 356497 17 356531 111
rect 356565 51 356641 145
rect 356685 17 356719 111
rect 356753 51 356829 145
rect 356873 17 356907 111
rect 356941 51 357017 145
rect 357061 17 357095 111
rect 357129 51 357205 145
rect 357249 17 357283 111
rect 357317 51 357393 145
rect 357437 17 357471 111
rect 357505 51 357581 145
rect 357625 17 357679 111
rect 357713 17 357771 162
rect 357805 51 357851 199
rect 357885 17 357961 165
rect 358005 51 358057 213
rect 358101 17 358161 179
rect 358205 51 358265 213
rect 361342 181 361449 291
rect 358309 17 358419 181
rect 358453 145 361449 181
rect 361577 167 361681 275
rect 361715 201 361819 309
rect 361853 294 361911 527
rect 361945 309 362279 527
rect 361945 171 362095 275
rect 362129 205 362279 309
rect 362313 294 362371 527
rect 362405 309 362923 527
rect 362405 171 362647 275
rect 362681 205 362923 309
rect 362957 294 363015 527
rect 363049 309 363751 527
rect 363049 171 363379 275
rect 363413 205 363751 309
rect 363785 294 363843 527
rect 363877 309 364946 527
rect 363877 171 364393 275
rect 364427 205 364946 309
rect 364981 294 365039 527
rect 366453 294 366511 527
rect 366545 294 366603 527
rect 366639 299 366705 527
rect 366838 397 366904 493
rect 366800 361 366904 397
rect 366800 351 366879 361
rect 366687 211 366766 265
rect 358453 51 358529 145
rect 358573 17 358607 111
rect 358641 51 358717 145
rect 358761 17 358795 111
rect 358829 51 358905 145
rect 358949 17 358983 111
rect 359017 51 359093 145
rect 359137 17 359171 111
rect 359205 51 359281 145
rect 359325 17 359359 111
rect 359393 51 359469 145
rect 359513 17 359547 111
rect 359581 51 359657 145
rect 359701 17 359735 111
rect 359769 51 359845 145
rect 359889 17 359923 111
rect 359957 51 360033 145
rect 360077 17 360111 111
rect 360145 51 360221 145
rect 360265 17 360299 111
rect 360333 51 360409 145
rect 360453 17 360487 111
rect 360521 51 360597 145
rect 360641 17 360675 111
rect 360709 51 360785 145
rect 360829 17 360863 111
rect 360897 51 360973 145
rect 361017 17 361051 111
rect 361085 51 361161 145
rect 361205 17 361239 111
rect 361273 51 361349 145
rect 361393 17 361447 111
rect 361485 17 361543 162
rect 361577 17 361819 167
rect 361853 17 361911 162
rect 361945 17 362279 171
rect 362313 17 362371 162
rect 362405 17 362923 171
rect 362957 17 363015 162
rect 363049 17 363751 171
rect 363785 17 363843 162
rect 363877 17 364946 171
rect 364981 17 365039 162
rect 366453 17 366511 162
rect 366545 17 366603 162
rect 366646 17 366698 177
rect 366732 125 366766 211
rect 366800 201 366834 351
rect 366942 327 367008 493
rect 366912 301 367008 327
rect 366868 293 367008 301
rect 367053 293 367113 527
rect 367152 327 367218 493
rect 367256 397 367322 493
rect 367256 361 367360 397
rect 367281 351 367360 361
rect 367152 301 367248 327
rect 367152 293 367292 301
rect 366868 235 366946 293
rect 366800 167 366878 201
rect 366732 79 366787 125
rect 366829 66 366878 167
rect 366912 151 366946 235
rect 366981 189 367051 259
rect 367109 189 367179 259
rect 367214 235 367292 293
rect 367214 151 367248 235
rect 367326 201 367360 351
rect 367455 299 367533 527
rect 367666 397 367732 493
rect 367628 361 367732 397
rect 367628 351 367707 361
rect 366912 117 367000 151
rect 366950 66 367000 117
rect 367047 17 367113 132
rect 367160 117 367248 151
rect 367282 167 367360 201
rect 367394 211 367473 265
rect 367515 211 367594 265
rect 367160 66 367210 117
rect 367282 66 367331 167
rect 367394 125 367428 211
rect 367373 79 367428 125
rect 367462 17 367526 177
rect 367560 125 367594 211
rect 367628 201 367662 351
rect 367770 327 367836 493
rect 367740 301 367836 327
rect 367696 293 367836 301
rect 367875 293 367935 527
rect 367980 327 368046 493
rect 368084 397 368150 493
rect 368084 361 368188 397
rect 368109 351 368188 361
rect 367980 301 368076 327
rect 367980 293 368120 301
rect 367696 235 367774 293
rect 367628 167 367706 201
rect 367560 79 367615 125
rect 367657 66 367706 167
rect 367740 151 367774 235
rect 367809 189 367879 259
rect 367937 189 368007 259
rect 368042 235 368120 293
rect 368042 151 368076 235
rect 368154 201 368188 351
rect 368283 299 368349 527
rect 368385 294 368443 527
rect 368479 442 368545 493
rect 368479 333 368539 442
rect 368579 421 368639 527
rect 368573 367 368639 421
rect 368683 459 368916 493
rect 368683 333 368717 459
rect 368753 351 368839 425
rect 368479 299 368717 333
rect 367740 117 367828 151
rect 367778 66 367828 117
rect 367875 17 367941 132
rect 367988 117 368076 151
rect 368110 167 368188 201
rect 368222 211 368301 265
rect 368479 211 368643 265
rect 367988 66 368038 117
rect 368110 66 368159 167
rect 368222 125 368256 211
rect 368666 177 368727 185
rect 368777 177 368811 351
rect 368882 329 368916 459
rect 368970 327 369036 493
rect 368950 295 369036 327
rect 368880 293 369036 295
rect 369071 293 369137 527
rect 369172 327 369238 493
rect 369292 459 369525 493
rect 369292 329 369326 459
rect 369369 351 369455 425
rect 369172 295 369258 327
rect 369172 293 369328 295
rect 368880 261 368984 293
rect 369224 261 369328 293
rect 368880 241 368963 261
rect 368201 79 368256 125
rect 368290 17 368342 177
rect 368385 17 368443 162
rect 368489 143 368727 177
rect 368489 51 368555 143
rect 368589 17 368632 109
rect 368666 85 368727 143
rect 368761 119 368827 177
rect 368861 85 368895 154
rect 368929 151 368963 241
rect 369018 205 369085 259
rect 369123 205 369190 259
rect 369245 241 369328 261
rect 369245 151 369279 241
rect 369397 177 369431 351
rect 369491 333 369525 459
rect 369569 421 369629 527
rect 369663 442 369729 493
rect 369569 367 369635 421
rect 369669 333 369729 442
rect 369491 299 369729 333
rect 369767 442 369833 493
rect 369767 333 369827 442
rect 369867 421 369927 527
rect 369861 367 369927 421
rect 369971 459 370204 493
rect 369971 333 370005 459
rect 370041 351 370127 425
rect 369767 299 370005 333
rect 369565 211 369729 265
rect 369767 211 369931 265
rect 369481 177 369542 185
rect 369954 177 370015 185
rect 370065 177 370099 351
rect 370170 329 370204 459
rect 370258 327 370324 493
rect 370238 295 370324 327
rect 370168 293 370324 295
rect 370359 293 370425 527
rect 370460 327 370526 493
rect 370580 459 370813 493
rect 370580 329 370614 459
rect 370657 351 370743 425
rect 370460 295 370546 327
rect 370460 293 370616 295
rect 370168 261 370272 293
rect 370512 261 370616 293
rect 370168 241 370251 261
rect 368929 117 369045 151
rect 368666 51 368895 85
rect 368995 66 369045 117
rect 369079 17 369129 132
rect 369163 117 369279 151
rect 369163 66 369213 117
rect 369313 85 369347 154
rect 369381 119 369447 177
rect 369481 143 369719 177
rect 369481 85 369542 143
rect 369313 51 369542 85
rect 369576 17 369619 109
rect 369653 51 369719 143
rect 369777 143 370015 177
rect 369777 51 369843 143
rect 369877 17 369920 109
rect 369954 85 370015 143
rect 370049 119 370115 177
rect 370149 85 370183 154
rect 370217 151 370251 241
rect 370306 205 370373 259
rect 370411 205 370478 259
rect 370533 241 370616 261
rect 370533 151 370567 241
rect 370685 177 370719 351
rect 370779 333 370813 459
rect 370857 421 370917 527
rect 370951 442 371017 493
rect 370857 367 370923 421
rect 370957 333 371017 442
rect 370779 299 371017 333
rect 371053 294 371111 527
rect 371153 299 371207 527
rect 371241 333 371307 493
rect 371341 367 371395 527
rect 371429 333 371495 493
rect 371529 367 371583 527
rect 371627 459 372069 493
rect 371627 333 371687 459
rect 371241 299 371687 333
rect 371721 273 371787 425
rect 371821 307 371875 459
rect 371909 273 371975 425
rect 372009 313 372069 459
rect 372118 321 372173 527
rect 372212 321 372278 493
rect 372312 321 372372 527
rect 372460 321 372520 527
rect 372554 321 372620 493
rect 372659 321 372714 527
rect 372763 459 373205 493
rect 372212 279 372246 321
rect 370853 211 371017 265
rect 371207 211 371485 265
rect 371721 213 371975 273
rect 372009 213 372246 279
rect 372586 279 372620 321
rect 372763 313 372823 459
rect 370769 177 370830 185
rect 371721 177 371767 213
rect 370217 117 370333 151
rect 369954 51 370183 85
rect 370283 66 370333 117
rect 370367 17 370417 132
rect 370451 117 370567 151
rect 370451 66 370501 117
rect 370601 85 370635 154
rect 370669 119 370735 177
rect 370769 143 371007 177
rect 370769 85 370830 143
rect 370601 51 370830 85
rect 370864 17 370907 109
rect 370941 51 371007 143
rect 371053 17 371111 162
rect 371157 17 371207 177
rect 371241 143 371667 177
rect 371241 51 371307 143
rect 371341 17 371395 109
rect 371429 51 371495 143
rect 371529 17 371579 109
rect 371613 85 371667 143
rect 371701 119 371767 177
rect 371801 85 371835 154
rect 371869 119 371935 213
rect 372212 165 372246 213
rect 372280 199 372399 265
rect 372433 199 372552 265
rect 372586 213 372823 279
rect 372857 273 372923 425
rect 372957 307 373011 459
rect 373045 273 373111 425
rect 373145 333 373205 459
rect 373249 367 373303 527
rect 373337 333 373403 493
rect 373437 367 373491 527
rect 373525 333 373591 493
rect 373145 299 373591 333
rect 373625 299 373679 527
rect 373729 299 373783 527
rect 373817 333 373883 493
rect 373917 367 373971 527
rect 374005 333 374071 493
rect 374105 367 374159 527
rect 374203 459 374645 493
rect 374203 333 374263 459
rect 373817 299 374263 333
rect 372857 213 373111 273
rect 374297 273 374363 425
rect 374397 307 374451 459
rect 374485 273 374551 425
rect 374585 313 374645 459
rect 374694 321 374749 527
rect 374788 321 374854 493
rect 374888 321 374948 527
rect 375036 321 375096 527
rect 375130 321 375196 493
rect 375235 321 375290 527
rect 375339 459 375781 493
rect 374788 279 374822 321
rect 372586 165 372620 213
rect 371969 85 372019 154
rect 371613 51 372019 85
rect 372120 17 372178 122
rect 372212 56 372262 165
rect 372304 17 372362 122
rect 372470 17 372528 122
rect 372570 56 372620 165
rect 372654 17 372712 122
rect 372813 85 372863 154
rect 372897 119 372963 213
rect 373065 177 373111 213
rect 373347 211 373625 265
rect 373783 211 374061 265
rect 374297 213 374551 273
rect 374585 213 374822 279
rect 375162 279 375196 321
rect 375339 313 375399 459
rect 374297 177 374343 213
rect 372997 85 373031 154
rect 373065 119 373131 177
rect 373165 143 373591 177
rect 373165 85 373219 143
rect 372813 51 373219 85
rect 373253 17 373303 109
rect 373337 51 373403 143
rect 373437 17 373491 109
rect 373525 51 373591 143
rect 373625 17 373675 177
rect 373733 17 373783 177
rect 373817 143 374243 177
rect 373817 51 373883 143
rect 373917 17 373971 109
rect 374005 51 374071 143
rect 374105 17 374155 109
rect 374189 85 374243 143
rect 374277 119 374343 177
rect 374377 85 374411 154
rect 374445 119 374511 213
rect 374788 165 374822 213
rect 374856 199 374975 265
rect 375009 199 375128 265
rect 375162 213 375399 279
rect 375433 273 375499 425
rect 375533 307 375587 459
rect 375621 273 375687 425
rect 375721 333 375781 459
rect 375825 367 375879 527
rect 375913 333 375979 493
rect 376013 367 376067 527
rect 376101 333 376167 493
rect 375721 299 376167 333
rect 376201 299 376255 527
rect 376297 294 376355 527
rect 376391 299 376457 527
rect 376590 397 376656 493
rect 376552 361 376656 397
rect 376552 351 376631 361
rect 375433 213 375687 273
rect 375162 165 375196 213
rect 374545 85 374595 154
rect 374189 51 374595 85
rect 374696 17 374754 122
rect 374788 56 374838 165
rect 374880 17 374938 122
rect 375046 17 375104 122
rect 375146 56 375196 165
rect 375230 17 375288 122
rect 375389 85 375439 154
rect 375473 119 375539 213
rect 375641 177 375687 213
rect 375923 211 376201 265
rect 376439 211 376518 265
rect 375573 85 375607 154
rect 375641 119 375707 177
rect 375741 143 376167 177
rect 375741 85 375795 143
rect 375389 51 375795 85
rect 375829 17 375879 109
rect 375913 51 375979 143
rect 376013 17 376067 109
rect 376101 51 376167 143
rect 376201 17 376251 177
rect 376297 17 376355 162
rect 376398 17 376450 177
rect 376484 125 376518 211
rect 376552 201 376586 351
rect 376694 327 376760 493
rect 376664 301 376760 327
rect 376620 293 376760 301
rect 376799 293 376865 527
rect 376904 327 376970 493
rect 377008 397 377074 493
rect 377008 361 377112 397
rect 377033 351 377112 361
rect 376904 301 377000 327
rect 376904 293 377044 301
rect 376620 235 376698 293
rect 376552 167 376630 201
rect 376484 79 376539 125
rect 376581 66 376630 167
rect 376664 151 376698 235
rect 376733 189 376813 259
rect 376851 189 376931 259
rect 376966 235 377044 293
rect 376966 151 377000 235
rect 377078 201 377112 351
rect 377207 299 377285 527
rect 377418 397 377484 493
rect 377380 361 377484 397
rect 377380 351 377459 361
rect 376664 117 376752 151
rect 376702 66 376752 117
rect 376799 17 376865 132
rect 376912 117 377000 151
rect 377034 167 377112 201
rect 377146 211 377225 265
rect 377267 211 377346 265
rect 376912 66 376962 117
rect 377034 66 377083 167
rect 377146 125 377180 211
rect 377125 79 377180 125
rect 377214 17 377278 177
rect 377312 125 377346 211
rect 377380 201 377414 351
rect 377522 327 377588 493
rect 377492 301 377588 327
rect 377448 293 377588 301
rect 377627 293 377693 527
rect 377732 327 377798 493
rect 377836 397 377902 493
rect 377836 361 377940 397
rect 377861 351 377940 361
rect 377732 301 377828 327
rect 377732 293 377872 301
rect 377448 235 377526 293
rect 377380 167 377458 201
rect 377312 79 377367 125
rect 377409 66 377458 167
rect 377492 151 377526 235
rect 377561 189 377641 259
rect 377679 189 377759 259
rect 377794 235 377872 293
rect 377794 151 377828 235
rect 377906 201 377940 351
rect 378035 299 378113 527
rect 378246 397 378312 493
rect 378208 361 378312 397
rect 378208 351 378287 361
rect 377492 117 377580 151
rect 377530 66 377580 117
rect 377627 17 377693 132
rect 377740 117 377828 151
rect 377862 167 377940 201
rect 377974 211 378053 265
rect 378095 211 378174 265
rect 377740 66 377790 117
rect 377862 66 377911 167
rect 377974 125 378008 211
rect 377953 79 378008 125
rect 378042 17 378106 177
rect 378140 125 378174 211
rect 378208 201 378242 351
rect 378350 327 378416 493
rect 378320 301 378416 327
rect 378276 293 378416 301
rect 378455 293 378521 527
rect 378560 327 378626 493
rect 378664 397 378730 493
rect 378664 361 378768 397
rect 378689 351 378768 361
rect 378560 301 378656 327
rect 378560 293 378700 301
rect 378276 235 378354 293
rect 378208 167 378286 201
rect 378140 79 378195 125
rect 378237 66 378286 167
rect 378320 151 378354 235
rect 378389 189 378469 259
rect 378507 189 378587 259
rect 378622 235 378700 293
rect 378622 151 378656 235
rect 378734 201 378768 351
rect 378863 299 378941 527
rect 379074 397 379140 493
rect 379036 361 379140 397
rect 379036 351 379115 361
rect 378320 117 378408 151
rect 378358 66 378408 117
rect 378455 17 378521 132
rect 378568 117 378656 151
rect 378690 167 378768 201
rect 378802 211 378881 265
rect 378923 211 379002 265
rect 378568 66 378618 117
rect 378690 66 378739 167
rect 378802 125 378836 211
rect 378781 79 378836 125
rect 378870 17 378934 177
rect 378968 125 379002 211
rect 379036 201 379070 351
rect 379178 327 379244 493
rect 379148 301 379244 327
rect 379104 293 379244 301
rect 379283 293 379349 527
rect 379388 327 379454 493
rect 379492 397 379558 493
rect 379492 361 379596 397
rect 379517 351 379596 361
rect 379388 301 379484 327
rect 379388 293 379528 301
rect 379104 235 379182 293
rect 379036 167 379114 201
rect 378968 79 379023 125
rect 379065 66 379114 167
rect 379148 151 379182 235
rect 379217 189 379297 259
rect 379335 189 379415 259
rect 379450 235 379528 293
rect 379450 151 379484 235
rect 379562 201 379596 351
rect 379691 299 379757 527
rect 379793 294 379851 527
rect 379887 442 379953 493
rect 379887 333 379947 442
rect 379987 421 380047 527
rect 379981 367 380047 421
rect 380091 459 380324 493
rect 380091 333 380125 459
rect 380161 351 380247 425
rect 379887 299 380125 333
rect 379148 117 379236 151
rect 379186 66 379236 117
rect 379283 17 379349 132
rect 379396 117 379484 151
rect 379518 167 379596 201
rect 379630 211 379709 265
rect 379887 211 380051 265
rect 379396 66 379446 117
rect 379518 66 379567 167
rect 379630 125 379664 211
rect 380074 177 380135 185
rect 380185 177 380219 351
rect 380290 329 380324 459
rect 380378 327 380444 493
rect 380358 295 380444 327
rect 380288 293 380444 295
rect 380479 293 380545 527
rect 380580 327 380646 493
rect 380700 459 380933 493
rect 380700 329 380734 459
rect 380777 351 380863 425
rect 380580 295 380666 327
rect 380580 293 380736 295
rect 380288 261 380392 293
rect 380632 261 380736 293
rect 380288 241 380371 261
rect 379609 79 379664 125
rect 379698 17 379750 177
rect 379793 17 379851 162
rect 379897 143 380135 177
rect 379897 51 379963 143
rect 379997 17 380040 109
rect 380074 85 380135 143
rect 380169 119 380235 177
rect 380269 85 380303 154
rect 380337 151 380371 241
rect 380426 205 380493 259
rect 380531 205 380598 259
rect 380653 241 380736 261
rect 380653 151 380687 241
rect 380805 177 380839 351
rect 380899 333 380933 459
rect 380977 421 381037 527
rect 381071 442 381137 493
rect 380977 367 381043 421
rect 381077 333 381137 442
rect 380899 299 381137 333
rect 381175 442 381241 493
rect 381175 333 381235 442
rect 381275 421 381335 527
rect 381269 367 381335 421
rect 381379 459 381612 493
rect 381379 333 381413 459
rect 381449 351 381535 425
rect 381175 299 381413 333
rect 380973 211 381137 265
rect 381175 211 381339 265
rect 380889 177 380950 185
rect 381362 177 381423 185
rect 381473 177 381507 351
rect 381578 329 381612 459
rect 381666 327 381732 493
rect 381646 295 381732 327
rect 381576 293 381732 295
rect 381767 293 381833 527
rect 381868 327 381934 493
rect 381988 459 382221 493
rect 381988 329 382022 459
rect 382065 351 382151 425
rect 381868 295 381954 327
rect 381868 293 382024 295
rect 381576 261 381680 293
rect 381920 261 382024 293
rect 381576 241 381659 261
rect 380337 117 380453 151
rect 380074 51 380303 85
rect 380403 66 380453 117
rect 380487 17 380537 132
rect 380571 117 380687 151
rect 380571 66 380621 117
rect 380721 85 380755 154
rect 380789 119 380855 177
rect 380889 143 381127 177
rect 380889 85 380950 143
rect 380721 51 380950 85
rect 380984 17 381027 109
rect 381061 51 381127 143
rect 381185 143 381423 177
rect 381185 51 381251 143
rect 381285 17 381328 109
rect 381362 85 381423 143
rect 381457 119 381523 177
rect 381557 85 381591 154
rect 381625 151 381659 241
rect 381714 205 381781 259
rect 381819 205 381886 259
rect 381941 241 382024 261
rect 381941 151 381975 241
rect 382093 177 382127 351
rect 382187 333 382221 459
rect 382265 421 382325 527
rect 382359 442 382425 493
rect 382265 367 382331 421
rect 382365 333 382425 442
rect 382187 299 382425 333
rect 382463 442 382529 493
rect 382463 333 382523 442
rect 382563 421 382623 527
rect 382557 367 382623 421
rect 382667 459 382900 493
rect 382667 333 382701 459
rect 382737 351 382823 425
rect 382463 299 382701 333
rect 382261 211 382425 265
rect 382463 211 382627 265
rect 382177 177 382238 185
rect 382650 177 382711 185
rect 382761 177 382795 351
rect 382866 329 382900 459
rect 382954 327 383020 493
rect 382934 295 383020 327
rect 382864 293 383020 295
rect 383055 293 383121 527
rect 383156 327 383222 493
rect 383276 459 383509 493
rect 383276 329 383310 459
rect 383353 351 383439 425
rect 383156 295 383242 327
rect 383156 293 383312 295
rect 382864 261 382968 293
rect 383208 261 383312 293
rect 382864 241 382947 261
rect 381625 117 381741 151
rect 381362 51 381591 85
rect 381691 66 381741 117
rect 381775 17 381825 132
rect 381859 117 381975 151
rect 381859 66 381909 117
rect 382009 85 382043 154
rect 382077 119 382143 177
rect 382177 143 382415 177
rect 382177 85 382238 143
rect 382009 51 382238 85
rect 382272 17 382315 109
rect 382349 51 382415 143
rect 382473 143 382711 177
rect 382473 51 382539 143
rect 382573 17 382616 109
rect 382650 85 382711 143
rect 382745 119 382811 177
rect 382845 85 382879 154
rect 382913 151 382947 241
rect 383002 205 383069 259
rect 383107 205 383174 259
rect 383229 241 383312 261
rect 383229 151 383263 241
rect 383381 177 383415 351
rect 383475 333 383509 459
rect 383553 421 383613 527
rect 383647 442 383713 493
rect 383553 367 383619 421
rect 383653 333 383713 442
rect 383475 299 383713 333
rect 383751 442 383817 493
rect 383751 333 383811 442
rect 383851 421 383911 527
rect 383845 367 383911 421
rect 383955 459 384188 493
rect 383955 333 383989 459
rect 384025 351 384111 425
rect 383751 299 383989 333
rect 383549 211 383713 265
rect 383751 211 383915 265
rect 383465 177 383526 185
rect 383938 177 383999 185
rect 384049 177 384083 351
rect 384154 329 384188 459
rect 384242 327 384308 493
rect 384222 295 384308 327
rect 384152 293 384308 295
rect 384343 293 384409 527
rect 384444 327 384510 493
rect 384564 459 384797 493
rect 384564 329 384598 459
rect 384641 351 384727 425
rect 384444 295 384530 327
rect 384444 293 384600 295
rect 384152 261 384256 293
rect 384496 261 384600 293
rect 384152 241 384235 261
rect 382913 117 383029 151
rect 382650 51 382879 85
rect 382979 66 383029 117
rect 383063 17 383113 132
rect 383147 117 383263 151
rect 383147 66 383197 117
rect 383297 85 383331 154
rect 383365 119 383431 177
rect 383465 143 383703 177
rect 383465 85 383526 143
rect 383297 51 383526 85
rect 383560 17 383603 109
rect 383637 51 383703 143
rect 383761 143 383999 177
rect 383761 51 383827 143
rect 383861 17 383904 109
rect 383938 85 383999 143
rect 384033 119 384099 177
rect 384133 85 384167 154
rect 384201 151 384235 241
rect 384290 205 384357 259
rect 384395 205 384462 259
rect 384517 241 384600 261
rect 384517 151 384551 241
rect 384669 177 384703 351
rect 384763 333 384797 459
rect 384841 421 384901 527
rect 384935 442 385001 493
rect 384841 367 384907 421
rect 384941 333 385001 442
rect 384763 299 385001 333
rect 385037 294 385095 527
rect 385130 299 385197 493
rect 385241 299 385275 527
rect 385326 459 385795 493
rect 384837 211 385001 265
rect 384753 177 384814 185
rect 384201 117 384317 151
rect 383938 51 384167 85
rect 384267 66 384317 117
rect 384351 17 384401 132
rect 384435 117 384551 151
rect 384435 66 384485 117
rect 384585 85 384619 154
rect 384653 119 384719 177
rect 384753 143 384991 177
rect 384753 85 384814 143
rect 384585 51 384814 85
rect 384848 17 384891 109
rect 384925 51 384991 143
rect 385037 17 385095 162
rect 385130 51 385181 299
rect 385326 265 385366 459
rect 385215 165 385249 265
rect 385311 199 385366 265
rect 385400 391 385689 425
rect 385400 165 385434 391
rect 385215 131 385434 165
rect 385468 323 385727 357
rect 385468 162 385502 323
rect 385399 124 385434 131
rect 385215 17 385291 97
rect 385399 51 385503 124
rect 385570 51 385635 283
rect 385669 51 385727 323
rect 385761 326 385795 459
rect 385829 367 385875 527
rect 385909 367 385989 493
rect 385761 288 385911 326
rect 385777 173 385811 237
rect 385873 211 385911 288
rect 385955 173 385989 367
rect 386049 294 386107 527
rect 386151 299 386200 527
rect 386235 299 386303 493
rect 386339 299 386389 527
rect 386430 459 386899 493
rect 385777 139 385989 173
rect 385762 17 385865 105
rect 385919 51 385968 139
rect 386049 17 386107 162
rect 386151 17 386201 131
rect 386235 51 386285 299
rect 386430 265 386470 459
rect 386319 165 386353 265
rect 386415 199 386470 265
rect 386504 391 386793 425
rect 386504 165 386538 391
rect 386319 131 386538 165
rect 386572 323 386831 357
rect 386572 162 386606 323
rect 386503 124 386538 131
rect 386319 17 386395 97
rect 386503 51 386640 124
rect 386674 51 386739 283
rect 386773 51 386831 323
rect 386865 326 386899 459
rect 386933 367 386979 527
rect 387013 367 387093 493
rect 386865 288 387015 326
rect 386881 173 386915 237
rect 386977 211 387015 288
rect 387059 173 387093 367
rect 387153 294 387211 527
rect 387255 299 387307 527
rect 387341 299 387407 493
rect 387441 299 387489 527
rect 387523 299 387595 493
rect 387629 299 387684 527
rect 387718 459 388187 493
rect 386881 139 387093 173
rect 387346 265 387398 299
rect 387523 265 387577 299
rect 387718 265 387758 459
rect 387346 213 387577 265
rect 386866 17 386969 105
rect 387023 51 387072 139
rect 387153 17 387211 162
rect 387263 17 387312 131
rect 387346 51 387398 213
rect 387439 17 387489 131
rect 387523 51 387577 213
rect 387611 165 387645 265
rect 387703 199 387758 265
rect 387792 391 388081 425
rect 387792 165 387826 391
rect 387611 131 387826 165
rect 387860 323 388119 357
rect 387860 162 387894 323
rect 387791 124 387826 131
rect 387611 17 387683 97
rect 387791 51 387928 124
rect 387962 51 388027 283
rect 388061 51 388119 323
rect 388153 326 388187 459
rect 388221 367 388267 527
rect 388301 367 388381 493
rect 388153 288 388303 326
rect 388169 173 388203 237
rect 388265 211 388303 288
rect 388347 173 388381 367
rect 388441 294 388499 527
rect 388560 321 388620 527
rect 388654 321 388720 493
rect 388759 321 388814 527
rect 388686 279 388720 321
rect 388863 313 388923 493
rect 388533 199 388652 265
rect 388686 213 388923 279
rect 388957 273 389023 815
rect 389057 595 389111 781
rect 389057 307 389111 493
rect 389145 273 389211 815
rect 390305 815 390559 875
rect 389245 755 389691 789
rect 389245 595 389305 755
rect 389349 561 389403 721
rect 389437 595 389503 755
rect 389537 561 389591 721
rect 389625 595 389691 755
rect 389725 561 389791 789
rect 389825 755 390271 789
rect 389825 595 389891 755
rect 389925 561 389979 721
rect 390013 595 390079 755
rect 390113 561 390167 721
rect 390211 595 390271 755
rect 389245 527 390271 561
rect 389245 333 389305 493
rect 389349 367 389403 527
rect 389437 333 389503 493
rect 389537 367 389591 527
rect 389625 333 389691 493
rect 389245 299 389691 333
rect 389725 299 389791 527
rect 389825 333 389891 493
rect 389925 367 389979 527
rect 390013 333 390079 493
rect 390113 367 390167 527
rect 390211 333 390271 493
rect 389825 299 390271 333
rect 388957 213 389211 273
rect 390305 273 390371 815
rect 390405 595 390459 781
rect 390405 307 390459 493
rect 390493 273 390559 815
rect 390593 809 390830 875
rect 390864 823 390983 889
rect 391017 823 391136 889
rect 391170 875 391204 923
rect 391481 875 391547 969
rect 391581 934 391615 1003
rect 391649 911 391715 969
rect 391749 945 391803 1003
rect 391837 979 391887 1071
rect 391921 945 391987 1037
rect 392021 979 392075 1071
rect 392109 945 392175 1037
rect 391749 911 392175 945
rect 392209 911 392275 1071
rect 392309 945 392375 1037
rect 392409 979 392463 1071
rect 392497 945 392563 1037
rect 392597 979 392647 1071
rect 392681 1003 393087 1037
rect 392681 945 392735 1003
rect 392309 911 392735 945
rect 392769 911 392835 969
rect 392869 934 392903 1003
rect 391649 875 391695 911
rect 390593 595 390653 775
rect 390796 767 390830 809
rect 391170 809 391407 875
rect 391441 815 391695 875
rect 391931 823 392209 877
rect 392275 823 392553 877
rect 392789 875 392835 911
rect 392937 875 393003 969
rect 393037 934 393087 1003
rect 393188 966 393246 1071
rect 393280 923 393330 1032
rect 393372 966 393430 1071
rect 393501 926 393559 1071
rect 393280 875 393314 923
rect 393602 911 393654 1071
rect 393688 963 393743 1009
rect 391170 767 391204 809
rect 390702 561 390757 767
rect 390796 595 390862 767
rect 390896 561 390956 767
rect 391044 561 391104 767
rect 391138 595 391204 767
rect 391243 561 391298 767
rect 391347 595 391407 775
rect 390593 527 391407 561
rect 390593 313 390653 493
rect 390702 321 390757 527
rect 390796 321 390862 493
rect 390896 321 390956 527
rect 391044 321 391104 527
rect 391138 321 391204 493
rect 391243 321 391298 527
rect 390796 279 390830 321
rect 388169 139 388381 173
rect 388686 165 388720 213
rect 388154 17 388257 105
rect 388311 51 388360 139
rect 388441 17 388499 162
rect 388570 17 388628 122
rect 388670 56 388720 165
rect 388754 17 388812 122
rect 388913 85 388963 154
rect 388997 119 389063 213
rect 389165 177 389211 213
rect 389447 211 389725 265
rect 389791 211 390069 265
rect 390305 213 390559 273
rect 390593 213 390830 279
rect 391170 279 391204 321
rect 391347 313 391407 493
rect 390305 177 390351 213
rect 389097 85 389131 154
rect 389165 119 389231 177
rect 389265 143 389691 177
rect 389265 85 389319 143
rect 388913 51 389319 85
rect 389353 17 389403 109
rect 389437 51 389503 143
rect 389537 17 389591 109
rect 389625 51 389691 143
rect 389725 17 389791 177
rect 389825 143 390251 177
rect 389825 51 389891 143
rect 389925 17 389979 109
rect 390013 51 390079 143
rect 390113 17 390163 109
rect 390197 85 390251 143
rect 390285 119 390351 177
rect 390385 85 390419 154
rect 390453 119 390519 213
rect 390796 165 390830 213
rect 390864 199 390983 265
rect 391017 199 391136 265
rect 391170 213 391407 279
rect 391441 273 391507 815
rect 391541 595 391595 781
rect 391541 307 391595 493
rect 391629 273 391695 815
rect 392789 815 393043 875
rect 391729 755 392175 789
rect 391729 595 391789 755
rect 391833 561 391887 721
rect 391921 595 391987 755
rect 392021 561 392075 721
rect 392109 595 392175 755
rect 392209 561 392275 789
rect 392309 755 392755 789
rect 392309 595 392375 755
rect 392409 561 392463 721
rect 392497 595 392563 755
rect 392597 561 392651 721
rect 392695 595 392755 755
rect 391729 527 392755 561
rect 391729 333 391789 493
rect 391833 367 391887 527
rect 391921 333 391987 493
rect 392021 367 392075 527
rect 392109 333 392175 493
rect 391729 299 392175 333
rect 392209 299 392275 527
rect 392309 333 392375 493
rect 392409 367 392463 527
rect 392497 333 392563 493
rect 392597 367 392651 527
rect 392695 333 392755 493
rect 392309 299 392755 333
rect 391441 213 391695 273
rect 392789 273 392855 815
rect 392889 595 392943 781
rect 392889 307 392943 493
rect 392977 273 393043 815
rect 393077 809 393314 875
rect 393348 823 393467 889
rect 393688 877 393722 963
rect 393785 921 393834 1022
rect 393906 971 393956 1022
rect 393643 823 393722 877
rect 393756 887 393834 921
rect 393868 937 393956 971
rect 394003 956 394069 1071
rect 394116 971 394166 1022
rect 394116 937 394204 971
rect 393077 595 393137 775
rect 393280 767 393314 809
rect 393186 561 393241 767
rect 393280 595 393346 767
rect 393380 561 393440 767
rect 393501 561 393559 794
rect 393595 561 393661 789
rect 393756 737 393790 887
rect 393868 853 393902 937
rect 393824 795 393902 853
rect 393937 829 394017 899
rect 394055 829 394135 899
rect 394170 853 394204 937
rect 394238 921 394287 1022
rect 394329 963 394384 1009
rect 394238 887 394316 921
rect 394170 795 394248 853
rect 393824 787 393964 795
rect 393868 761 393964 787
rect 393756 727 393835 737
rect 393756 691 393860 727
rect 393794 595 393860 691
rect 393898 595 393964 761
rect 393077 527 393760 561
rect 393077 313 393137 493
rect 393186 321 393241 527
rect 393280 321 393346 493
rect 393380 321 393440 527
rect 393280 279 393314 321
rect 393501 294 393559 527
rect 393595 299 393661 527
rect 393794 493 393835 595
rect 394003 561 394069 795
rect 394108 787 394248 795
rect 394108 761 394204 787
rect 394108 595 394174 761
rect 394282 737 394316 887
rect 394350 877 394384 963
rect 394418 911 394482 1071
rect 394516 963 394571 1009
rect 394516 877 394550 963
rect 394613 921 394662 1022
rect 394734 971 394784 1022
rect 394350 823 394429 877
rect 394471 823 394550 877
rect 394584 887 394662 921
rect 394696 937 394784 971
rect 394831 956 394897 1071
rect 394944 971 394994 1022
rect 394944 937 395032 971
rect 394237 727 394316 737
rect 394212 691 394316 727
rect 394212 595 394278 691
rect 393869 527 394203 561
rect 393794 397 393860 493
rect 393756 361 393860 397
rect 393756 351 393835 361
rect 391170 165 391204 213
rect 390553 85 390603 154
rect 390197 51 390603 85
rect 390704 17 390762 122
rect 390796 56 390846 165
rect 390888 17 390946 122
rect 391054 17 391112 122
rect 391154 56 391204 165
rect 391238 17 391296 122
rect 391397 85 391447 154
rect 391481 119 391547 213
rect 391649 177 391695 213
rect 391931 211 392209 265
rect 392275 211 392553 265
rect 392789 213 393043 273
rect 393077 213 393314 279
rect 392789 177 392835 213
rect 391581 85 391615 154
rect 391649 119 391715 177
rect 391749 143 392175 177
rect 391749 85 391803 143
rect 391397 51 391803 85
rect 391837 17 391887 109
rect 391921 51 391987 143
rect 392021 17 392075 109
rect 392109 51 392175 143
rect 392209 17 392275 177
rect 392309 143 392735 177
rect 392309 51 392375 143
rect 392409 17 392463 109
rect 392497 51 392563 143
rect 392597 17 392647 109
rect 392681 85 392735 143
rect 392769 119 392835 177
rect 392869 85 392903 154
rect 392937 119 393003 213
rect 393280 165 393314 213
rect 393348 199 393467 265
rect 393643 211 393722 265
rect 393037 85 393087 154
rect 392681 51 393087 85
rect 393188 17 393246 122
rect 393280 56 393330 165
rect 393372 17 393430 122
rect 393501 17 393559 162
rect 393602 17 393654 177
rect 393688 125 393722 211
rect 393756 201 393790 351
rect 393898 327 393964 493
rect 393868 301 393964 327
rect 393824 293 393964 301
rect 394003 293 394069 527
rect 394237 493 394278 595
rect 394411 561 394489 789
rect 394584 737 394618 887
rect 394696 853 394730 937
rect 394652 795 394730 853
rect 394765 829 394845 899
rect 394883 829 394963 899
rect 394998 853 395032 937
rect 395066 921 395115 1022
rect 395157 963 395212 1009
rect 395066 887 395144 921
rect 394998 795 395076 853
rect 394652 787 394792 795
rect 394696 761 394792 787
rect 394584 727 394663 737
rect 394584 691 394688 727
rect 394622 595 394688 691
rect 394726 595 394792 761
rect 394312 527 394588 561
rect 394108 327 394174 493
rect 394212 397 394278 493
rect 394212 361 394316 397
rect 394237 351 394316 361
rect 394108 301 394204 327
rect 394108 293 394248 301
rect 393824 235 393902 293
rect 393756 167 393834 201
rect 393688 79 393743 125
rect 393785 66 393834 167
rect 393868 151 393902 235
rect 393937 189 394017 259
rect 394055 189 394135 259
rect 394170 235 394248 293
rect 394170 151 394204 235
rect 394282 201 394316 351
rect 394411 299 394489 527
rect 394622 493 394663 595
rect 394831 561 394897 795
rect 394936 787 395076 795
rect 394936 761 395032 787
rect 394936 595 395002 761
rect 395110 737 395144 887
rect 395178 877 395212 963
rect 395246 911 395310 1071
rect 395344 963 395399 1009
rect 395344 877 395378 963
rect 395441 921 395490 1022
rect 395562 971 395612 1022
rect 395178 823 395257 877
rect 395299 823 395378 877
rect 395412 887 395490 921
rect 395524 937 395612 971
rect 395659 956 395725 1071
rect 395772 971 395822 1022
rect 395772 937 395860 971
rect 395065 727 395144 737
rect 395040 691 395144 727
rect 395040 595 395106 691
rect 394697 527 395031 561
rect 394622 397 394688 493
rect 394584 361 394688 397
rect 394584 351 394663 361
rect 393868 117 393956 151
rect 393906 66 393956 117
rect 394003 17 394069 132
rect 394116 117 394204 151
rect 394238 167 394316 201
rect 394350 211 394429 265
rect 394471 211 394550 265
rect 394116 66 394166 117
rect 394238 66 394287 167
rect 394350 125 394384 211
rect 394329 79 394384 125
rect 394418 17 394482 177
rect 394516 125 394550 211
rect 394584 201 394618 351
rect 394726 327 394792 493
rect 394696 301 394792 327
rect 394652 293 394792 301
rect 394831 293 394897 527
rect 395065 493 395106 595
rect 395239 561 395317 789
rect 395412 737 395446 887
rect 395524 853 395558 937
rect 395480 795 395558 853
rect 395593 829 395673 899
rect 395711 829 395791 899
rect 395826 853 395860 937
rect 395894 921 395943 1022
rect 395985 963 396040 1009
rect 395894 887 395972 921
rect 395826 795 395904 853
rect 395480 787 395620 795
rect 395524 761 395620 787
rect 395412 727 395491 737
rect 395412 691 395516 727
rect 395450 595 395516 691
rect 395554 595 395620 761
rect 395140 527 395416 561
rect 394936 327 395002 493
rect 395040 397 395106 493
rect 395040 361 395144 397
rect 395065 351 395144 361
rect 394936 301 395032 327
rect 394936 293 395076 301
rect 394652 235 394730 293
rect 394584 167 394662 201
rect 394516 79 394571 125
rect 394613 66 394662 167
rect 394696 151 394730 235
rect 394765 189 394845 259
rect 394883 189 394963 259
rect 394998 235 395076 293
rect 394998 151 395032 235
rect 395110 201 395144 351
rect 395239 299 395317 527
rect 395450 493 395491 595
rect 395659 561 395725 795
rect 395764 787 395904 795
rect 395764 761 395860 787
rect 395764 595 395830 761
rect 395938 737 395972 887
rect 396006 877 396040 963
rect 396074 911 396138 1071
rect 396172 963 396227 1009
rect 396172 877 396206 963
rect 396269 921 396318 1022
rect 396390 971 396440 1022
rect 396006 823 396085 877
rect 396127 823 396206 877
rect 396240 887 396318 921
rect 396352 937 396440 971
rect 396487 956 396553 1071
rect 396600 971 396650 1022
rect 396600 937 396688 971
rect 395893 727 395972 737
rect 395868 691 395972 727
rect 395868 595 395934 691
rect 395525 527 395859 561
rect 395450 397 395516 493
rect 395412 361 395516 397
rect 395412 351 395491 361
rect 394696 117 394784 151
rect 394734 66 394784 117
rect 394831 17 394897 132
rect 394944 117 395032 151
rect 395066 167 395144 201
rect 395178 211 395257 265
rect 395299 211 395378 265
rect 394944 66 394994 117
rect 395066 66 395115 167
rect 395178 125 395212 211
rect 395157 79 395212 125
rect 395246 17 395310 177
rect 395344 125 395378 211
rect 395412 201 395446 351
rect 395554 327 395620 493
rect 395524 301 395620 327
rect 395480 293 395620 301
rect 395659 293 395725 527
rect 395893 493 395934 595
rect 396067 561 396145 789
rect 396240 737 396274 887
rect 396352 853 396386 937
rect 396308 795 396386 853
rect 396421 829 396501 899
rect 396539 829 396619 899
rect 396654 853 396688 937
rect 396722 921 396771 1022
rect 396813 963 396868 1009
rect 396722 887 396800 921
rect 396654 795 396732 853
rect 396308 787 396448 795
rect 396352 761 396448 787
rect 396240 727 396319 737
rect 396240 691 396344 727
rect 396278 595 396344 691
rect 396382 595 396448 761
rect 395968 527 396244 561
rect 395764 327 395830 493
rect 395868 397 395934 493
rect 395868 361 395972 397
rect 395893 351 395972 361
rect 395764 301 395860 327
rect 395764 293 395904 301
rect 395480 235 395558 293
rect 395412 167 395490 201
rect 395344 79 395399 125
rect 395441 66 395490 167
rect 395524 151 395558 235
rect 395593 189 395673 259
rect 395711 189 395791 259
rect 395826 235 395904 293
rect 395826 151 395860 235
rect 395938 201 395972 351
rect 396067 299 396145 527
rect 396278 493 396319 595
rect 396487 561 396553 795
rect 396592 787 396732 795
rect 396592 761 396688 787
rect 396592 595 396658 761
rect 396766 737 396800 887
rect 396834 877 396868 963
rect 396902 911 396954 1071
rect 396997 926 397055 1071
rect 397101 945 397167 1037
rect 397201 979 397244 1071
rect 397278 1003 397507 1037
rect 397278 945 397339 1003
rect 397101 911 397339 945
rect 397373 911 397439 969
rect 397473 934 397507 1003
rect 397607 971 397657 1022
rect 397541 937 397657 971
rect 397691 956 397741 1071
rect 397775 971 397825 1022
rect 397925 1003 398154 1037
rect 397775 937 397891 971
rect 397278 903 397339 911
rect 396834 823 396913 877
rect 397091 823 397255 877
rect 396721 727 396800 737
rect 396696 691 396800 727
rect 396696 595 396762 691
rect 396353 527 396687 561
rect 396278 397 396344 493
rect 396240 361 396344 397
rect 396240 351 396319 361
rect 395524 117 395612 151
rect 395562 66 395612 117
rect 395659 17 395725 132
rect 395772 117 395860 151
rect 395894 167 395972 201
rect 396006 211 396085 265
rect 396127 211 396206 265
rect 395772 66 395822 117
rect 395894 66 395943 167
rect 396006 125 396040 211
rect 395985 79 396040 125
rect 396074 17 396138 177
rect 396172 125 396206 211
rect 396240 201 396274 351
rect 396382 327 396448 493
rect 396352 301 396448 327
rect 396308 293 396448 301
rect 396487 293 396553 527
rect 396721 493 396762 595
rect 396895 561 396961 789
rect 396997 561 397055 794
rect 397091 755 397329 789
rect 397091 646 397151 755
rect 397185 667 397251 721
rect 397091 595 397157 646
rect 397191 561 397251 667
rect 397295 629 397329 755
rect 397389 737 397423 911
rect 397541 847 397575 937
rect 397492 827 397575 847
rect 397630 829 397697 883
rect 397735 829 397802 883
rect 397857 847 397891 937
rect 397925 934 397959 1003
rect 397993 911 398059 969
rect 398093 945 398154 1003
rect 398188 979 398231 1071
rect 398265 945 398331 1037
rect 398093 911 398331 945
rect 398389 945 398455 1037
rect 398489 979 398532 1071
rect 398566 1003 398795 1037
rect 398566 945 398627 1003
rect 398389 911 398627 945
rect 398661 911 398727 969
rect 398761 934 398795 1003
rect 398895 971 398945 1022
rect 398829 937 398945 971
rect 398979 956 399029 1071
rect 399063 971 399113 1022
rect 399213 1003 399442 1037
rect 399063 937 399179 971
rect 397857 827 397940 847
rect 397492 795 397596 827
rect 397836 795 397940 827
rect 397492 793 397648 795
rect 397562 761 397648 793
rect 397365 663 397451 737
rect 397295 595 397355 629
rect 396796 527 397355 561
rect 396592 327 396658 493
rect 396696 397 396762 493
rect 396696 361 396800 397
rect 396721 351 396800 361
rect 396592 301 396688 327
rect 396592 293 396732 301
rect 396308 235 396386 293
rect 396240 167 396318 201
rect 396172 79 396227 125
rect 396269 66 396318 167
rect 396352 151 396386 235
rect 396421 189 396501 259
rect 396539 189 396619 259
rect 396654 235 396732 293
rect 396654 151 396688 235
rect 396766 201 396800 351
rect 396895 299 396961 527
rect 396997 294 397055 527
rect 397091 442 397157 493
rect 397091 333 397151 442
rect 397191 421 397251 527
rect 397185 367 397251 421
rect 397295 459 397355 493
rect 397295 333 397329 459
rect 397389 425 397423 663
rect 397494 629 397528 759
rect 397457 595 397528 629
rect 397582 595 397648 761
rect 397683 561 397749 795
rect 397784 793 397940 795
rect 397784 761 397870 793
rect 397784 595 397850 761
rect 397904 629 397938 759
rect 398009 737 398043 911
rect 398093 903 398154 911
rect 398566 903 398627 911
rect 398177 823 398341 877
rect 398379 823 398543 877
rect 398103 755 398341 789
rect 397981 663 398067 737
rect 397904 595 397975 629
rect 397457 527 397975 561
rect 397457 459 397528 493
rect 397365 351 397451 425
rect 397091 299 397329 333
rect 396352 117 396440 151
rect 396390 66 396440 117
rect 396487 17 396553 132
rect 396600 117 396688 151
rect 396722 167 396800 201
rect 396834 211 396913 265
rect 397091 211 397255 265
rect 396600 66 396650 117
rect 396722 66 396771 167
rect 396834 125 396868 211
rect 397278 177 397339 185
rect 397389 177 397423 351
rect 397494 329 397528 459
rect 397582 327 397648 493
rect 397562 295 397648 327
rect 397492 293 397648 295
rect 397683 293 397749 527
rect 397784 327 397850 493
rect 397904 459 397975 493
rect 397904 329 397938 459
rect 398009 425 398043 663
rect 398103 629 398137 755
rect 398077 595 398137 629
rect 398181 667 398247 721
rect 398181 561 398241 667
rect 398281 646 398341 755
rect 398275 595 398341 646
rect 398379 755 398617 789
rect 398379 646 398439 755
rect 398473 667 398539 721
rect 398379 595 398445 646
rect 398479 561 398539 667
rect 398583 629 398617 755
rect 398677 737 398711 911
rect 398829 847 398863 937
rect 398780 827 398863 847
rect 398918 829 398985 883
rect 399023 829 399090 883
rect 399145 847 399179 937
rect 399213 934 399247 1003
rect 399281 911 399347 969
rect 399381 945 399442 1003
rect 399476 979 399519 1071
rect 399553 945 399619 1037
rect 399381 911 399619 945
rect 399677 945 399743 1037
rect 399777 979 399820 1071
rect 399854 1003 400083 1037
rect 399854 945 399915 1003
rect 399677 911 399915 945
rect 399949 911 400015 969
rect 400049 934 400083 1003
rect 400183 971 400233 1022
rect 400117 937 400233 971
rect 400267 956 400317 1071
rect 400351 971 400401 1022
rect 400501 1003 400730 1037
rect 400351 937 400467 971
rect 399145 827 399228 847
rect 398780 795 398884 827
rect 399124 795 399228 827
rect 398780 793 398936 795
rect 398850 761 398936 793
rect 398653 663 398739 737
rect 398583 595 398643 629
rect 398077 527 398643 561
rect 398077 459 398137 493
rect 397981 351 398067 425
rect 397784 295 397870 327
rect 397784 293 397940 295
rect 397492 261 397596 293
rect 397836 261 397940 293
rect 397492 241 397575 261
rect 396813 79 396868 125
rect 396902 17 396954 177
rect 396997 17 397055 162
rect 397101 143 397339 177
rect 397101 51 397167 143
rect 397201 17 397244 109
rect 397278 85 397339 143
rect 397373 119 397439 177
rect 397473 85 397507 154
rect 397541 151 397575 241
rect 397630 205 397697 259
rect 397735 205 397802 259
rect 397857 241 397940 261
rect 397857 151 397891 241
rect 398009 177 398043 351
rect 398103 333 398137 459
rect 398181 421 398241 527
rect 398275 442 398341 493
rect 398181 367 398247 421
rect 398281 333 398341 442
rect 398103 299 398341 333
rect 398379 442 398445 493
rect 398379 333 398439 442
rect 398479 421 398539 527
rect 398473 367 398539 421
rect 398583 459 398643 493
rect 398583 333 398617 459
rect 398677 425 398711 663
rect 398782 629 398816 759
rect 398745 595 398816 629
rect 398870 595 398936 761
rect 398971 561 399037 795
rect 399072 793 399228 795
rect 399072 761 399158 793
rect 399072 595 399138 761
rect 399192 629 399226 759
rect 399297 737 399331 911
rect 399381 903 399442 911
rect 399854 903 399915 911
rect 399465 823 399629 877
rect 399667 823 399831 877
rect 399391 755 399629 789
rect 399269 663 399355 737
rect 399192 595 399263 629
rect 398745 527 399263 561
rect 398745 459 398816 493
rect 398653 351 398739 425
rect 398379 299 398617 333
rect 398177 211 398341 265
rect 398379 211 398543 265
rect 398093 177 398154 185
rect 398566 177 398627 185
rect 398677 177 398711 351
rect 398782 329 398816 459
rect 398870 327 398936 493
rect 398850 295 398936 327
rect 398780 293 398936 295
rect 398971 293 399037 527
rect 399072 327 399138 493
rect 399192 459 399263 493
rect 399192 329 399226 459
rect 399297 425 399331 663
rect 399391 629 399425 755
rect 399365 595 399425 629
rect 399469 667 399535 721
rect 399469 561 399529 667
rect 399569 646 399629 755
rect 399563 595 399629 646
rect 399667 755 399905 789
rect 399667 646 399727 755
rect 399761 667 399827 721
rect 399667 595 399733 646
rect 399767 561 399827 667
rect 399871 629 399905 755
rect 399965 737 399999 911
rect 400117 847 400151 937
rect 400068 827 400151 847
rect 400206 829 400273 883
rect 400311 829 400378 883
rect 400433 847 400467 937
rect 400501 934 400535 1003
rect 400569 911 400635 969
rect 400669 945 400730 1003
rect 400764 979 400807 1071
rect 400841 945 400907 1037
rect 400669 911 400907 945
rect 400965 945 401031 1037
rect 401065 979 401108 1071
rect 401142 1003 401371 1037
rect 401142 945 401203 1003
rect 400965 911 401203 945
rect 401237 911 401303 969
rect 401337 934 401371 1003
rect 401471 971 401521 1022
rect 401405 937 401521 971
rect 401555 956 401605 1071
rect 401639 971 401689 1022
rect 401789 1003 402018 1037
rect 401639 937 401755 971
rect 400433 827 400516 847
rect 400068 795 400172 827
rect 400412 795 400516 827
rect 400068 793 400224 795
rect 400138 761 400224 793
rect 399941 663 400027 737
rect 399871 595 399931 629
rect 399365 527 399931 561
rect 399365 459 399425 493
rect 399269 351 399355 425
rect 399072 295 399158 327
rect 399072 293 399228 295
rect 398780 261 398884 293
rect 399124 261 399228 293
rect 398780 241 398863 261
rect 397541 117 397657 151
rect 397278 51 397507 85
rect 397607 66 397657 117
rect 397691 17 397741 132
rect 397775 117 397891 151
rect 397775 66 397825 117
rect 397925 85 397959 154
rect 397993 119 398059 177
rect 398093 143 398331 177
rect 398093 85 398154 143
rect 397925 51 398154 85
rect 398188 17 398231 109
rect 398265 51 398331 143
rect 398389 143 398627 177
rect 398389 51 398455 143
rect 398489 17 398532 109
rect 398566 85 398627 143
rect 398661 119 398727 177
rect 398761 85 398795 154
rect 398829 151 398863 241
rect 398918 205 398985 259
rect 399023 205 399090 259
rect 399145 241 399228 261
rect 399145 151 399179 241
rect 399297 177 399331 351
rect 399391 333 399425 459
rect 399469 421 399529 527
rect 399563 442 399629 493
rect 399469 367 399535 421
rect 399569 333 399629 442
rect 399391 299 399629 333
rect 399667 442 399733 493
rect 399667 333 399727 442
rect 399767 421 399827 527
rect 399761 367 399827 421
rect 399871 459 399931 493
rect 399871 333 399905 459
rect 399965 425 399999 663
rect 400070 629 400104 759
rect 400033 595 400104 629
rect 400158 595 400224 761
rect 400259 561 400325 795
rect 400360 793 400516 795
rect 400360 761 400446 793
rect 400360 595 400426 761
rect 400480 629 400514 759
rect 400585 737 400619 911
rect 400669 903 400730 911
rect 401142 903 401203 911
rect 400753 823 400917 877
rect 400955 823 401119 877
rect 400679 755 400917 789
rect 400557 663 400643 737
rect 400480 595 400551 629
rect 400033 527 400551 561
rect 400033 459 400104 493
rect 399941 351 400027 425
rect 399667 299 399905 333
rect 399465 211 399629 265
rect 399667 211 399831 265
rect 399381 177 399442 185
rect 399854 177 399915 185
rect 399965 177 399999 351
rect 400070 329 400104 459
rect 400158 327 400224 493
rect 400138 295 400224 327
rect 400068 293 400224 295
rect 400259 293 400325 527
rect 400360 327 400426 493
rect 400480 459 400551 493
rect 400480 329 400514 459
rect 400585 425 400619 663
rect 400679 629 400713 755
rect 400653 595 400713 629
rect 400757 667 400823 721
rect 400757 561 400817 667
rect 400857 646 400917 755
rect 400851 595 400917 646
rect 400955 755 401193 789
rect 400955 646 401015 755
rect 401049 667 401115 721
rect 400955 595 401021 646
rect 401055 561 401115 667
rect 401159 629 401193 755
rect 401253 737 401287 911
rect 401405 847 401439 937
rect 401356 827 401439 847
rect 401494 829 401561 883
rect 401599 829 401666 883
rect 401721 847 401755 937
rect 401789 934 401823 1003
rect 401857 911 401923 969
rect 401957 945 402018 1003
rect 402052 979 402095 1071
rect 402129 945 402195 1037
rect 401957 911 402195 945
rect 402241 926 402299 1071
rect 402345 911 402395 1071
rect 402429 945 402495 1037
rect 402529 979 402583 1071
rect 402617 945 402683 1037
rect 402717 979 402767 1071
rect 402801 1003 403207 1037
rect 402801 945 402855 1003
rect 402429 911 402855 945
rect 402889 911 402955 969
rect 402989 934 403023 1003
rect 401721 827 401804 847
rect 401356 795 401460 827
rect 401700 795 401804 827
rect 401356 793 401512 795
rect 401426 761 401512 793
rect 401229 663 401315 737
rect 401159 595 401219 629
rect 400653 527 401219 561
rect 400653 459 400713 493
rect 400557 351 400643 425
rect 400360 295 400446 327
rect 400360 293 400516 295
rect 400068 261 400172 293
rect 400412 261 400516 293
rect 400068 241 400151 261
rect 398829 117 398945 151
rect 398566 51 398795 85
rect 398895 66 398945 117
rect 398979 17 399029 132
rect 399063 117 399179 151
rect 399063 66 399113 117
rect 399213 85 399247 154
rect 399281 119 399347 177
rect 399381 143 399619 177
rect 399381 85 399442 143
rect 399213 51 399442 85
rect 399476 17 399519 109
rect 399553 51 399619 143
rect 399677 143 399915 177
rect 399677 51 399743 143
rect 399777 17 399820 109
rect 399854 85 399915 143
rect 399949 119 400015 177
rect 400049 85 400083 154
rect 400117 151 400151 241
rect 400206 205 400273 259
rect 400311 205 400378 259
rect 400433 241 400516 261
rect 400433 151 400467 241
rect 400585 177 400619 351
rect 400679 333 400713 459
rect 400757 421 400817 527
rect 400851 442 400917 493
rect 400757 367 400823 421
rect 400857 333 400917 442
rect 400679 299 400917 333
rect 400955 442 401021 493
rect 400955 333 401015 442
rect 401055 421 401115 527
rect 401049 367 401115 421
rect 401159 459 401219 493
rect 401159 333 401193 459
rect 401253 425 401287 663
rect 401358 629 401392 759
rect 401321 595 401392 629
rect 401446 595 401512 761
rect 401547 561 401613 795
rect 401648 793 401804 795
rect 401648 761 401734 793
rect 401648 595 401714 761
rect 401768 629 401802 759
rect 401873 737 401907 911
rect 401957 903 402018 911
rect 402041 823 402205 877
rect 402395 823 402673 877
rect 402909 875 402955 911
rect 403057 875 403123 969
rect 403157 934 403207 1003
rect 403308 966 403366 1071
rect 403400 923 403450 1032
rect 403492 966 403550 1071
rect 403658 966 403716 1071
rect 403758 923 403808 1032
rect 403842 966 403900 1071
rect 404001 1003 404407 1037
rect 404001 934 404051 1003
rect 403400 875 403434 923
rect 402909 815 403163 875
rect 401967 755 402205 789
rect 401845 663 401931 737
rect 401768 595 401839 629
rect 401321 527 401839 561
rect 401321 459 401392 493
rect 401229 351 401315 425
rect 400955 299 401193 333
rect 400753 211 400917 265
rect 400955 211 401119 265
rect 400669 177 400730 185
rect 401142 177 401203 185
rect 401253 177 401287 351
rect 401358 329 401392 459
rect 401446 327 401512 493
rect 401426 295 401512 327
rect 401356 293 401512 295
rect 401547 293 401613 527
rect 401648 327 401714 493
rect 401768 459 401839 493
rect 401768 329 401802 459
rect 401873 425 401907 663
rect 401967 629 402001 755
rect 401941 595 402001 629
rect 402045 667 402111 721
rect 402045 561 402105 667
rect 402145 646 402205 755
rect 402139 595 402205 646
rect 402241 561 402299 794
rect 402341 561 402395 789
rect 402429 755 402875 789
rect 402429 595 402495 755
rect 402529 561 402583 721
rect 402617 595 402683 755
rect 402717 561 402771 721
rect 402815 595 402875 755
rect 401941 527 402875 561
rect 401941 459 402001 493
rect 401845 351 401931 425
rect 401648 295 401734 327
rect 401648 293 401804 295
rect 401356 261 401460 293
rect 401700 261 401804 293
rect 401356 241 401439 261
rect 400117 117 400233 151
rect 399854 51 400083 85
rect 400183 66 400233 117
rect 400267 17 400317 132
rect 400351 117 400467 151
rect 400351 66 400401 117
rect 400501 85 400535 154
rect 400569 119 400635 177
rect 400669 143 400907 177
rect 400669 85 400730 143
rect 400501 51 400730 85
rect 400764 17 400807 109
rect 400841 51 400907 143
rect 400965 143 401203 177
rect 400965 51 401031 143
rect 401065 17 401108 109
rect 401142 85 401203 143
rect 401237 119 401303 177
rect 401337 85 401371 154
rect 401405 151 401439 241
rect 401494 205 401561 259
rect 401599 205 401666 259
rect 401721 241 401804 261
rect 401721 151 401755 241
rect 401873 177 401907 351
rect 401967 333 402001 459
rect 402045 421 402105 527
rect 402139 442 402205 493
rect 402045 367 402111 421
rect 402145 333 402205 442
rect 401967 299 402205 333
rect 402241 294 402299 527
rect 402341 299 402395 527
rect 402429 333 402495 493
rect 402529 367 402583 527
rect 402617 333 402683 493
rect 402717 367 402771 527
rect 402815 333 402875 493
rect 402429 299 402875 333
rect 402909 273 402975 815
rect 403009 595 403063 781
rect 403009 307 403063 493
rect 403097 273 403163 815
rect 403197 809 403434 875
rect 403468 823 403587 889
rect 403621 823 403740 889
rect 403774 875 403808 923
rect 404085 875 404151 969
rect 404185 934 404219 1003
rect 404253 911 404319 969
rect 404353 945 404407 1003
rect 404441 979 404491 1071
rect 404525 945 404591 1037
rect 404625 979 404679 1071
rect 404713 945 404779 1037
rect 404353 911 404779 945
rect 404813 911 404863 1071
rect 404921 911 404971 1071
rect 405005 945 405071 1037
rect 405105 979 405159 1071
rect 405193 945 405259 1037
rect 405293 979 405343 1071
rect 405377 1003 405783 1037
rect 405377 945 405431 1003
rect 405005 911 405431 945
rect 405465 911 405531 969
rect 405565 934 405599 1003
rect 404253 875 404299 911
rect 403197 595 403257 775
rect 403400 767 403434 809
rect 403774 809 404011 875
rect 404045 815 404299 875
rect 404535 823 404813 877
rect 404971 823 405249 877
rect 405485 875 405531 911
rect 405633 875 405699 969
rect 405733 934 405783 1003
rect 405884 966 405942 1071
rect 405976 923 406026 1032
rect 406068 966 406126 1071
rect 406234 966 406292 1071
rect 406334 923 406384 1032
rect 406418 966 406476 1071
rect 406577 1003 406983 1037
rect 406577 934 406627 1003
rect 405976 875 406010 923
rect 403774 767 403808 809
rect 403306 561 403361 767
rect 403400 595 403466 767
rect 403500 561 403560 767
rect 403648 561 403708 767
rect 403742 595 403808 767
rect 403847 561 403902 767
rect 403951 595 404011 775
rect 403197 527 404011 561
rect 403197 313 403257 493
rect 403306 321 403361 527
rect 403400 321 403466 493
rect 403500 321 403560 527
rect 403648 321 403708 527
rect 403742 321 403808 493
rect 403847 321 403902 527
rect 403400 279 403434 321
rect 402041 211 402205 265
rect 402395 211 402673 265
rect 402909 213 403163 273
rect 403197 213 403434 279
rect 403774 279 403808 321
rect 403951 313 404011 493
rect 401957 177 402018 185
rect 402909 177 402955 213
rect 401405 117 401521 151
rect 401142 51 401371 85
rect 401471 66 401521 117
rect 401555 17 401605 132
rect 401639 117 401755 151
rect 401639 66 401689 117
rect 401789 85 401823 154
rect 401857 119 401923 177
rect 401957 143 402195 177
rect 401957 85 402018 143
rect 401789 51 402018 85
rect 402052 17 402095 109
rect 402129 51 402195 143
rect 402241 17 402299 162
rect 402345 17 402395 177
rect 402429 143 402855 177
rect 402429 51 402495 143
rect 402529 17 402583 109
rect 402617 51 402683 143
rect 402717 17 402767 109
rect 402801 85 402855 143
rect 402889 119 402955 177
rect 402989 85 403023 154
rect 403057 119 403123 213
rect 403400 165 403434 213
rect 403468 199 403587 265
rect 403621 199 403740 265
rect 403774 213 404011 279
rect 404045 273 404111 815
rect 404145 595 404199 781
rect 404145 307 404199 493
rect 404233 273 404299 815
rect 405485 815 405739 875
rect 404333 755 404779 789
rect 404333 595 404393 755
rect 404437 561 404491 721
rect 404525 595 404591 755
rect 404625 561 404679 721
rect 404713 595 404779 755
rect 404813 561 404867 789
rect 404917 561 404971 789
rect 405005 755 405451 789
rect 405005 595 405071 755
rect 405105 561 405159 721
rect 405193 595 405259 755
rect 405293 561 405347 721
rect 405391 595 405451 755
rect 404333 527 405451 561
rect 404333 333 404393 493
rect 404437 367 404491 527
rect 404525 333 404591 493
rect 404625 367 404679 527
rect 404713 333 404779 493
rect 404333 299 404779 333
rect 404813 299 404867 527
rect 404917 299 404971 527
rect 405005 333 405071 493
rect 405105 367 405159 527
rect 405193 333 405259 493
rect 405293 367 405347 527
rect 405391 333 405451 493
rect 405005 299 405451 333
rect 404045 213 404299 273
rect 405485 273 405551 815
rect 405585 595 405639 781
rect 405585 307 405639 493
rect 405673 273 405739 815
rect 405773 809 406010 875
rect 406044 823 406163 889
rect 406197 823 406316 889
rect 406350 875 406384 923
rect 406661 875 406727 969
rect 406761 934 406795 1003
rect 406829 911 406895 969
rect 406929 945 406983 1003
rect 407017 979 407067 1071
rect 407101 945 407167 1037
rect 407201 979 407255 1071
rect 407289 945 407355 1037
rect 406929 911 407355 945
rect 407389 911 407439 1071
rect 407485 926 407543 1071
rect 407589 911 407639 1071
rect 407673 945 407739 1037
rect 407773 979 407827 1071
rect 407861 945 407927 1037
rect 407961 979 408011 1071
rect 408045 1003 408451 1037
rect 408045 945 408099 1003
rect 407673 911 408099 945
rect 408133 911 408199 969
rect 408233 934 408267 1003
rect 406829 875 406875 911
rect 405773 595 405833 775
rect 405976 767 406010 809
rect 406350 809 406587 875
rect 406621 815 406875 875
rect 407111 823 407389 877
rect 407639 823 407917 877
rect 408153 875 408199 911
rect 408301 875 408367 969
rect 408401 934 408451 1003
rect 408552 966 408610 1071
rect 408644 923 408694 1032
rect 408736 966 408794 1071
rect 408902 966 408960 1071
rect 409002 923 409052 1032
rect 409086 966 409144 1071
rect 409245 1003 409651 1037
rect 409245 934 409295 1003
rect 408644 875 408678 923
rect 406350 767 406384 809
rect 405882 561 405937 767
rect 405976 595 406042 767
rect 406076 561 406136 767
rect 406224 561 406284 767
rect 406318 595 406384 767
rect 406423 561 406478 767
rect 406527 595 406587 775
rect 405773 527 406587 561
rect 405773 313 405833 493
rect 405882 321 405937 527
rect 405976 321 406042 493
rect 406076 321 406136 527
rect 406224 321 406284 527
rect 406318 321 406384 493
rect 406423 321 406478 527
rect 405976 279 406010 321
rect 403774 165 403808 213
rect 403157 85 403207 154
rect 402801 51 403207 85
rect 403308 17 403366 122
rect 403400 56 403450 165
rect 403492 17 403550 122
rect 403658 17 403716 122
rect 403758 56 403808 165
rect 403842 17 403900 122
rect 404001 85 404051 154
rect 404085 119 404151 213
rect 404253 177 404299 213
rect 404535 211 404813 265
rect 404971 211 405249 265
rect 405485 213 405739 273
rect 405773 213 406010 279
rect 406350 279 406384 321
rect 406527 313 406587 493
rect 405485 177 405531 213
rect 404185 85 404219 154
rect 404253 119 404319 177
rect 404353 143 404779 177
rect 404353 85 404407 143
rect 404001 51 404407 85
rect 404441 17 404491 109
rect 404525 51 404591 143
rect 404625 17 404679 109
rect 404713 51 404779 143
rect 404813 17 404863 177
rect 404921 17 404971 177
rect 405005 143 405431 177
rect 405005 51 405071 143
rect 405105 17 405159 109
rect 405193 51 405259 143
rect 405293 17 405343 109
rect 405377 85 405431 143
rect 405465 119 405531 177
rect 405565 85 405599 154
rect 405633 119 405699 213
rect 405976 165 406010 213
rect 406044 199 406163 265
rect 406197 199 406316 265
rect 406350 213 406587 279
rect 406621 273 406687 815
rect 406721 595 406775 781
rect 406721 307 406775 493
rect 406809 273 406875 815
rect 408153 815 408407 875
rect 406909 755 407355 789
rect 406909 595 406969 755
rect 407013 561 407067 721
rect 407101 595 407167 755
rect 407201 561 407255 721
rect 407289 595 407355 755
rect 407389 561 407443 789
rect 407485 561 407543 794
rect 407585 561 407639 789
rect 407673 755 408119 789
rect 407673 595 407739 755
rect 407773 561 407827 721
rect 407861 595 407927 755
rect 407961 561 408015 721
rect 408059 595 408119 755
rect 406909 527 408119 561
rect 406909 333 406969 493
rect 407013 367 407067 527
rect 407101 333 407167 493
rect 407201 367 407255 527
rect 407289 333 407355 493
rect 406909 299 407355 333
rect 407389 299 407443 527
rect 407485 294 407543 527
rect 407585 299 407639 527
rect 407673 333 407739 493
rect 407773 367 407827 527
rect 407861 333 407927 493
rect 407961 367 408015 527
rect 408059 333 408119 493
rect 407673 299 408119 333
rect 406621 213 406875 273
rect 408153 273 408219 815
rect 408253 595 408307 781
rect 408253 307 408307 493
rect 408341 273 408407 815
rect 408441 809 408678 875
rect 408712 823 408831 889
rect 408865 823 408984 889
rect 409018 875 409052 923
rect 409329 875 409395 969
rect 409429 934 409463 1003
rect 409497 911 409563 969
rect 409597 945 409651 1003
rect 409685 979 409735 1071
rect 409769 945 409835 1037
rect 409869 979 409923 1071
rect 409957 945 410023 1037
rect 409597 911 410023 945
rect 410057 911 410107 1071
rect 410165 911 410215 1071
rect 410249 945 410315 1037
rect 410349 979 410403 1071
rect 410437 945 410503 1037
rect 410537 979 410587 1071
rect 410621 1003 411027 1037
rect 410621 945 410675 1003
rect 410249 911 410675 945
rect 410709 911 410775 969
rect 410809 934 410843 1003
rect 409497 875 409543 911
rect 408441 595 408501 775
rect 408644 767 408678 809
rect 409018 809 409255 875
rect 409289 815 409543 875
rect 409779 823 410057 877
rect 410215 823 410493 877
rect 410729 875 410775 911
rect 410877 875 410943 969
rect 410977 934 411027 1003
rect 411128 966 411186 1071
rect 411220 923 411270 1032
rect 411312 966 411370 1071
rect 411478 966 411536 1071
rect 411578 923 411628 1032
rect 411662 966 411720 1071
rect 411821 1003 412227 1037
rect 411821 934 411871 1003
rect 411220 875 411254 923
rect 409018 767 409052 809
rect 408550 561 408605 767
rect 408644 595 408710 767
rect 408744 561 408804 767
rect 408892 561 408952 767
rect 408986 595 409052 767
rect 409091 561 409146 767
rect 409195 595 409255 775
rect 408441 527 409255 561
rect 408441 313 408501 493
rect 408550 321 408605 527
rect 408644 321 408710 493
rect 408744 321 408804 527
rect 408892 321 408952 527
rect 408986 321 409052 493
rect 409091 321 409146 527
rect 408644 279 408678 321
rect 406350 165 406384 213
rect 405733 85 405783 154
rect 405377 51 405783 85
rect 405884 17 405942 122
rect 405976 56 406026 165
rect 406068 17 406126 122
rect 406234 17 406292 122
rect 406334 56 406384 165
rect 406418 17 406476 122
rect 406577 85 406627 154
rect 406661 119 406727 213
rect 406829 177 406875 213
rect 407111 211 407389 265
rect 407639 211 407917 265
rect 408153 213 408407 273
rect 408441 213 408678 279
rect 409018 279 409052 321
rect 409195 313 409255 493
rect 408153 177 408199 213
rect 406761 85 406795 154
rect 406829 119 406895 177
rect 406929 143 407355 177
rect 406929 85 406983 143
rect 406577 51 406983 85
rect 407017 17 407067 109
rect 407101 51 407167 143
rect 407201 17 407255 109
rect 407289 51 407355 143
rect 407389 17 407439 177
rect 407485 17 407543 162
rect 407589 17 407639 177
rect 407673 143 408099 177
rect 407673 51 407739 143
rect 407773 17 407827 109
rect 407861 51 407927 143
rect 407961 17 408011 109
rect 408045 85 408099 143
rect 408133 119 408199 177
rect 408233 85 408267 154
rect 408301 119 408367 213
rect 408644 165 408678 213
rect 408712 199 408831 265
rect 408865 199 408984 265
rect 409018 213 409255 279
rect 409289 273 409355 815
rect 409389 595 409443 781
rect 409389 307 409443 493
rect 409477 273 409543 815
rect 410729 815 410983 875
rect 409577 755 410023 789
rect 409577 595 409637 755
rect 409681 561 409735 721
rect 409769 595 409835 755
rect 409869 561 409923 721
rect 409957 595 410023 755
rect 410057 561 410111 789
rect 410161 561 410215 789
rect 410249 755 410695 789
rect 410249 595 410315 755
rect 410349 561 410403 721
rect 410437 595 410503 755
rect 410537 561 410591 721
rect 410635 595 410695 755
rect 409577 527 410695 561
rect 409577 333 409637 493
rect 409681 367 409735 527
rect 409769 333 409835 493
rect 409869 367 409923 527
rect 409957 333 410023 493
rect 409577 299 410023 333
rect 410057 299 410111 527
rect 410161 299 410215 527
rect 410249 333 410315 493
rect 410349 367 410403 527
rect 410437 333 410503 493
rect 410537 367 410591 527
rect 410635 333 410695 493
rect 410249 299 410695 333
rect 409289 213 409543 273
rect 410729 273 410795 815
rect 410829 595 410883 781
rect 410829 307 410883 493
rect 410917 273 410983 815
rect 411017 809 411254 875
rect 411288 823 411407 889
rect 411441 823 411560 889
rect 411594 875 411628 923
rect 411905 875 411971 969
rect 412005 934 412039 1003
rect 412073 911 412139 969
rect 412173 945 412227 1003
rect 412261 979 412311 1071
rect 412345 945 412411 1037
rect 412445 979 412499 1071
rect 412533 945 412599 1037
rect 412173 911 412599 945
rect 412633 911 412683 1071
rect 412729 926 412787 1071
rect 412073 875 412119 911
rect 411017 595 411077 775
rect 411220 767 411254 809
rect 411594 809 411831 875
rect 411865 815 412119 875
rect 412355 823 412633 877
rect 411594 767 411628 809
rect 411126 561 411181 767
rect 411220 595 411286 767
rect 411320 561 411380 767
rect 411468 561 411528 767
rect 411562 595 411628 767
rect 411667 561 411722 767
rect 411771 595 411831 775
rect 411017 527 411831 561
rect 411017 313 411077 493
rect 411126 321 411181 527
rect 411220 321 411286 493
rect 411320 321 411380 527
rect 411468 321 411528 527
rect 411562 321 411628 493
rect 411667 321 411722 527
rect 411220 279 411254 321
rect 409018 165 409052 213
rect 408401 85 408451 154
rect 408045 51 408451 85
rect 408552 17 408610 122
rect 408644 56 408694 165
rect 408736 17 408794 122
rect 408902 17 408960 122
rect 409002 56 409052 165
rect 409086 17 409144 122
rect 409245 85 409295 154
rect 409329 119 409395 213
rect 409497 177 409543 213
rect 409779 211 410057 265
rect 410215 211 410493 265
rect 410729 213 410983 273
rect 411017 213 411254 279
rect 411594 279 411628 321
rect 411771 313 411831 493
rect 410729 177 410775 213
rect 409429 85 409463 154
rect 409497 119 409563 177
rect 409597 143 410023 177
rect 409597 85 409651 143
rect 409245 51 409651 85
rect 409685 17 409735 109
rect 409769 51 409835 143
rect 409869 17 409923 109
rect 409957 51 410023 143
rect 410057 17 410107 177
rect 410165 17 410215 177
rect 410249 143 410675 177
rect 410249 51 410315 143
rect 410349 17 410403 109
rect 410437 51 410503 143
rect 410537 17 410587 109
rect 410621 85 410675 143
rect 410709 119 410775 177
rect 410809 85 410843 154
rect 410877 119 410943 213
rect 411220 165 411254 213
rect 411288 199 411407 265
rect 411441 199 411560 265
rect 411594 213 411831 279
rect 411865 273 411931 815
rect 411965 595 412019 781
rect 411965 307 412019 493
rect 412053 273 412119 815
rect 412153 755 412599 789
rect 412153 595 412213 755
rect 412257 561 412311 721
rect 412345 595 412411 755
rect 412445 561 412499 721
rect 412533 595 412599 755
rect 412633 561 412687 789
rect 412729 561 412787 794
rect 412153 527 412804 561
rect 412153 333 412213 493
rect 412257 367 412311 527
rect 412345 333 412411 493
rect 412445 367 412499 527
rect 412533 333 412599 493
rect 412153 299 412599 333
rect 412633 299 412687 527
rect 412729 294 412787 527
rect 411865 213 412119 273
rect 411594 165 411628 213
rect 410977 85 411027 154
rect 410621 51 411027 85
rect 411128 17 411186 122
rect 411220 56 411270 165
rect 411312 17 411370 122
rect 411478 17 411536 122
rect 411578 56 411628 165
rect 411662 17 411720 122
rect 411821 85 411871 154
rect 411905 119 411971 213
rect 412073 177 412119 213
rect 412355 211 412633 265
rect 412005 85 412039 154
rect 412073 119 412139 177
rect 412173 143 412599 177
rect 412173 85 412227 143
rect 411821 51 412227 85
rect 412261 17 412311 109
rect 412345 51 412411 143
rect 412445 17 412499 109
rect 412533 51 412599 143
rect 412633 17 412683 177
rect 412729 17 412787 162
rect 0 -17 412804 17
<< via1 >>
rect 35730 1062 35782 1114
rect 35794 1062 35846 1114
rect 31243 824 31295 876
rect 31307 824 31359 876
rect 35094 824 35146 876
rect 35158 824 35210 876
rect 35730 518 35782 570
rect 35794 518 35846 570
<< obsm1 >>
rect 0 1114 46920 1136
rect 0 1102 35730 1114
rect -76 1074 35730 1102
rect -76 14 -48 1074
rect 0 1062 35730 1074
rect 35782 1062 35794 1114
rect 35846 1062 46920 1114
rect 0 1040 46920 1062
rect 388424 1102 412804 1136
rect 388424 1074 412880 1102
rect 388424 1040 412804 1074
rect 10419 1000 10477 1009
rect 12319 1000 12377 1009
rect 10419 972 12377 1000
rect 10419 963 10477 972
rect 12319 963 12377 972
rect 13823 1000 13881 1009
rect 15723 1000 15781 1009
rect 13823 972 15781 1000
rect 13823 963 13881 972
rect 15723 963 15781 972
rect 31237 824 31243 876
rect 31295 824 31307 876
rect 31359 873 31365 876
rect 31359 827 31574 873
rect 31359 824 31365 827
rect 35088 824 35094 876
rect 35146 824 35158 876
rect 35210 864 35216 876
rect 35533 864 35663 873
rect 35210 836 35663 864
rect 35210 824 35216 836
rect 35533 827 35663 836
rect 36179 796 36237 805
rect 36505 796 36563 805
rect 36179 768 36563 796
rect 36179 759 36237 768
rect 36505 759 36563 768
rect 37461 796 37519 805
rect 37885 796 37943 805
rect 37461 768 37943 796
rect 37461 759 37519 768
rect 37885 759 37943 768
rect 38939 796 38997 805
rect 39265 796 39323 805
rect 38939 768 39323 796
rect 38939 759 38997 768
rect 39265 759 39323 768
rect 40313 796 40371 805
rect 40737 796 40795 805
rect 40313 768 40795 796
rect 40313 759 40371 768
rect 40737 759 40795 768
rect 41883 796 41941 805
rect 42209 796 42267 805
rect 41883 768 42267 796
rect 41883 759 41941 768
rect 42209 759 42267 768
rect 43441 796 43499 805
rect 43865 796 43923 805
rect 43441 768 43923 796
rect 43441 759 43499 768
rect 43865 759 43923 768
rect 10513 728 10571 737
rect 10701 728 10759 737
rect 11557 728 11615 737
rect 11745 728 11803 737
rect 12037 728 12095 737
rect 12225 728 12283 737
rect 10513 700 11803 728
rect 10513 691 10571 700
rect 10701 691 10759 700
rect 11557 691 11615 700
rect 11745 691 11803 700
rect 11900 700 12283 728
rect 10993 660 11051 669
rect 11181 660 11239 669
rect 11900 660 11928 700
rect 12037 691 12095 700
rect 12225 691 12283 700
rect 13917 728 13975 737
rect 14105 728 14163 737
rect 14961 728 15019 737
rect 15149 728 15207 737
rect 15441 728 15499 737
rect 15629 728 15687 737
rect 13917 700 15207 728
rect 13917 691 13975 700
rect 14105 691 14163 700
rect 14961 691 15019 700
rect 15149 691 15207 700
rect 15304 700 15687 728
rect 10993 632 11928 660
rect 14397 660 14455 669
rect 14585 660 14643 669
rect 15304 660 15332 700
rect 15441 691 15499 700
rect 15629 691 15687 700
rect 33321 691 33379 737
rect 36087 728 36145 737
rect 36616 728 36674 737
rect 36087 700 36674 728
rect 36087 691 36145 700
rect 36616 691 36674 700
rect 37563 728 37621 737
rect 37996 728 38054 737
rect 37563 700 38054 728
rect 37563 691 37621 700
rect 37996 691 38054 700
rect 38847 728 38905 737
rect 39376 728 39434 737
rect 38847 700 39434 728
rect 38847 691 38905 700
rect 39376 691 39434 700
rect 40415 728 40473 737
rect 40848 728 40906 737
rect 40415 700 40906 728
rect 40415 691 40473 700
rect 40848 691 40906 700
rect 41791 728 41849 737
rect 42320 728 42378 737
rect 41791 700 42378 728
rect 41791 691 41849 700
rect 42320 691 42378 700
rect 43543 728 43601 737
rect 43976 728 44034 737
rect 43543 700 44034 728
rect 43543 691 43601 700
rect 43976 691 44034 700
rect 388961 728 389019 737
rect 389149 728 389207 737
rect 390309 728 390367 737
rect 390497 728 390555 737
rect 391445 728 391503 737
rect 391633 728 391691 737
rect 392793 728 392851 737
rect 392981 728 393039 737
rect 388961 700 393039 728
rect 388961 691 389019 700
rect 389149 691 389207 700
rect 390309 691 390367 700
rect 390497 691 390555 700
rect 391445 691 391503 700
rect 391633 691 391691 700
rect 392793 691 392851 700
rect 392981 691 393039 700
rect 393777 728 393835 737
rect 394237 728 394295 737
rect 394605 728 394663 737
rect 395065 728 395123 737
rect 395433 728 395491 737
rect 395893 728 395951 737
rect 396261 728 396319 737
rect 396721 728 396779 737
rect 393777 700 396779 728
rect 393777 691 393835 700
rect 394237 691 394295 700
rect 394605 691 394663 700
rect 395065 691 395123 700
rect 395433 691 395491 700
rect 395893 691 395951 700
rect 396261 691 396319 700
rect 396721 691 396779 700
rect 397365 728 397423 737
rect 398009 728 398067 737
rect 398653 728 398711 737
rect 399297 728 399355 737
rect 399941 728 399999 737
rect 400585 728 400643 737
rect 401229 728 401287 737
rect 401873 728 401931 737
rect 397365 700 401931 728
rect 397365 691 397423 700
rect 398009 691 398067 700
rect 398653 691 398711 700
rect 399297 691 399355 700
rect 399941 691 399999 700
rect 400585 691 400643 700
rect 401229 691 401287 700
rect 401873 691 401931 700
rect 402913 728 402971 737
rect 403101 728 403159 737
rect 404049 728 404107 737
rect 404237 728 404295 737
rect 405489 728 405547 737
rect 405677 728 405735 737
rect 406625 728 406683 737
rect 406813 728 406871 737
rect 408157 728 408215 737
rect 408345 728 408403 737
rect 409293 728 409351 737
rect 409481 728 409539 737
rect 410733 728 410791 737
rect 410921 728 410979 737
rect 411869 728 411927 737
rect 412057 728 412115 737
rect 402913 700 412115 728
rect 402913 691 402971 700
rect 403101 691 403159 700
rect 404049 691 404107 700
rect 404237 691 404295 700
rect 405489 691 405547 700
rect 405677 691 405735 700
rect 406625 691 406683 700
rect 406813 691 406871 700
rect 408157 691 408215 700
rect 408345 691 408403 700
rect 409293 691 409351 700
rect 409481 691 409539 700
rect 410733 691 410791 700
rect 410921 691 410979 700
rect 411869 691 411927 700
rect 412057 691 412115 700
rect 14397 632 15332 660
rect 10993 623 11051 632
rect 11181 623 11239 632
rect 14397 623 14455 632
rect 14585 623 14643 632
rect 33229 623 33287 669
rect 33244 592 33272 623
rect 33336 592 33364 691
rect 388865 657 388923 666
rect 389055 657 389113 666
rect 389245 657 389303 666
rect 389441 657 389499 666
rect 389629 657 389687 666
rect 388865 629 389687 657
rect 388865 620 388923 629
rect 389055 620 389113 629
rect 389245 620 389303 629
rect 389441 620 389499 629
rect 389629 620 389687 629
rect 389829 657 389887 666
rect 390017 657 390075 666
rect 390213 657 390271 666
rect 390403 657 390461 666
rect 390593 657 390651 666
rect 389829 629 390651 657
rect 389829 620 389887 629
rect 390017 620 390075 629
rect 390213 620 390271 629
rect 390403 620 390461 629
rect 390593 620 390651 629
rect 391349 657 391407 666
rect 391539 657 391597 666
rect 391729 657 391787 666
rect 391925 657 391983 666
rect 392113 657 392171 666
rect 391349 629 392171 657
rect 391349 620 391407 629
rect 391539 620 391597 629
rect 391729 620 391787 629
rect 391925 620 391983 629
rect 392113 620 392171 629
rect 392313 657 392371 666
rect 392501 657 392559 666
rect 392697 657 392755 666
rect 392887 657 392945 666
rect 393077 657 393135 666
rect 392313 629 393135 657
rect 392313 620 392371 629
rect 392501 620 392559 629
rect 392697 620 392755 629
rect 392887 620 392945 629
rect 393077 620 393135 629
rect 397095 657 397153 666
rect 397283 657 397341 666
rect 397482 657 397540 666
rect 397095 629 397540 657
rect 397095 620 397153 629
rect 397283 620 397341 629
rect 397482 620 397540 629
rect 397892 657 397950 666
rect 398091 657 398149 666
rect 398279 657 398337 666
rect 397892 629 398337 657
rect 397892 620 397950 629
rect 398091 620 398149 629
rect 398279 620 398337 629
rect 398383 657 398441 666
rect 398571 657 398629 666
rect 398770 657 398828 666
rect 398383 629 398828 657
rect 398383 620 398441 629
rect 398571 620 398629 629
rect 398770 620 398828 629
rect 399180 657 399238 666
rect 399379 657 399437 666
rect 399567 657 399625 666
rect 399180 629 399625 657
rect 399180 620 399238 629
rect 399379 620 399437 629
rect 399567 620 399625 629
rect 399671 657 399729 666
rect 399859 657 399917 666
rect 400058 657 400116 666
rect 399671 629 400116 657
rect 399671 620 399729 629
rect 399859 620 399917 629
rect 400058 620 400116 629
rect 400468 657 400526 666
rect 400667 657 400725 666
rect 400855 657 400913 666
rect 400468 629 400913 657
rect 400468 620 400526 629
rect 400667 620 400725 629
rect 400855 620 400913 629
rect 400959 657 401017 666
rect 401147 657 401205 666
rect 401346 657 401404 666
rect 400959 629 401404 657
rect 400959 620 401017 629
rect 401147 620 401205 629
rect 401346 620 401404 629
rect 401756 657 401814 666
rect 401955 657 402013 666
rect 402143 657 402201 666
rect 401756 629 402201 657
rect 401756 620 401814 629
rect 401955 620 402013 629
rect 402143 620 402201 629
rect 402433 657 402491 666
rect 402621 657 402679 666
rect 402817 657 402875 666
rect 403007 657 403065 666
rect 403197 657 403255 666
rect 402433 629 403255 657
rect 402433 620 402491 629
rect 402621 620 402679 629
rect 402817 620 402875 629
rect 403007 620 403065 629
rect 403197 620 403255 629
rect 403953 657 404011 666
rect 404143 657 404201 666
rect 404333 657 404391 666
rect 404529 657 404587 666
rect 404717 657 404775 666
rect 403953 629 404775 657
rect 403953 620 404011 629
rect 404143 620 404201 629
rect 404333 620 404391 629
rect 404529 620 404587 629
rect 404717 620 404775 629
rect 405009 657 405067 666
rect 405197 657 405255 666
rect 405393 657 405451 666
rect 405583 657 405641 666
rect 405773 657 405831 666
rect 405009 629 405831 657
rect 405009 620 405067 629
rect 405197 620 405255 629
rect 405393 620 405451 629
rect 405583 620 405641 629
rect 405773 620 405831 629
rect 406529 657 406587 666
rect 406719 657 406777 666
rect 406909 657 406967 666
rect 407105 657 407163 666
rect 407293 657 407351 666
rect 406529 629 407351 657
rect 406529 620 406587 629
rect 406719 620 406777 629
rect 406909 620 406967 629
rect 407105 620 407163 629
rect 407293 620 407351 629
rect 407677 657 407735 666
rect 407865 657 407923 666
rect 408061 657 408119 666
rect 408251 657 408309 666
rect 408441 657 408499 666
rect 407677 629 408499 657
rect 407677 620 407735 629
rect 407865 620 407923 629
rect 408061 620 408119 629
rect 408251 620 408309 629
rect 408441 620 408499 629
rect 409197 657 409255 666
rect 409387 657 409445 666
rect 409577 657 409635 666
rect 409773 657 409831 666
rect 409961 657 410019 666
rect 409197 629 410019 657
rect 409197 620 409255 629
rect 409387 620 409445 629
rect 409577 620 409635 629
rect 409773 620 409831 629
rect 409961 620 410019 629
rect 410253 657 410311 666
rect 410441 657 410499 666
rect 410637 657 410695 666
rect 410827 657 410885 666
rect 411017 657 411075 666
rect 410253 629 411075 657
rect 410253 620 410311 629
rect 410441 620 410499 629
rect 410637 620 410695 629
rect 410827 620 410885 629
rect 411017 620 411075 629
rect 411773 657 411831 666
rect 411963 657 412021 666
rect 412153 657 412211 666
rect 412349 657 412407 666
rect 412537 657 412595 666
rect 411773 629 412595 657
rect 411773 620 411831 629
rect 411963 620 412021 629
rect 412153 620 412211 629
rect 412349 620 412407 629
rect 412537 620 412595 629
rect 0 570 412804 592
rect 0 518 35730 570
rect 35782 518 35794 570
rect 35846 518 412804 570
rect 0 496 412804 518
rect 185355 456 185424 467
rect 185967 456 186036 467
rect 185355 428 186036 456
rect 185355 413 185424 428
rect 185967 413 186036 428
rect 327581 456 327639 465
rect 327785 456 327843 465
rect 327581 428 327843 456
rect 327581 419 327639 428
rect 327785 419 327843 428
rect 337749 456 337807 465
rect 337953 456 338011 465
rect 337749 428 338011 456
rect 337749 419 337807 428
rect 337953 419 338011 428
rect 388865 459 388923 468
rect 389055 459 389113 468
rect 389245 459 389303 468
rect 389441 459 389499 468
rect 389629 459 389687 468
rect 388865 431 389687 459
rect 388865 422 388923 431
rect 389055 422 389113 431
rect 389245 422 389303 431
rect 389441 422 389499 431
rect 389629 422 389687 431
rect 389829 459 389887 468
rect 390017 459 390075 468
rect 390213 459 390271 468
rect 390403 459 390461 468
rect 390593 459 390651 468
rect 389829 431 390651 459
rect 389829 422 389887 431
rect 390017 422 390075 431
rect 390213 422 390271 431
rect 390403 422 390461 431
rect 390593 422 390651 431
rect 391349 459 391407 468
rect 391539 459 391597 468
rect 391729 459 391787 468
rect 391925 459 391983 468
rect 392113 459 392171 468
rect 391349 431 392171 459
rect 391349 422 391407 431
rect 391539 422 391597 431
rect 391729 422 391787 431
rect 391925 422 391983 431
rect 392113 422 392171 431
rect 392313 459 392371 468
rect 392501 459 392559 468
rect 392697 459 392755 468
rect 392887 459 392945 468
rect 393077 459 393135 468
rect 392313 431 393135 459
rect 392313 422 392371 431
rect 392501 422 392559 431
rect 392697 422 392755 431
rect 392887 422 392945 431
rect 393077 422 393135 431
rect 397095 459 397153 468
rect 397283 459 397341 468
rect 397482 459 397540 468
rect 397095 431 397540 459
rect 397095 422 397153 431
rect 397283 422 397341 431
rect 397482 422 397540 431
rect 397892 459 397950 468
rect 398091 459 398149 468
rect 398279 459 398337 468
rect 397892 431 398337 459
rect 397892 422 397950 431
rect 398091 422 398149 431
rect 398279 422 398337 431
rect 398383 459 398441 468
rect 398571 459 398629 468
rect 398770 459 398828 468
rect 398383 431 398828 459
rect 398383 422 398441 431
rect 398571 422 398629 431
rect 398770 422 398828 431
rect 399180 459 399238 468
rect 399379 459 399437 468
rect 399567 459 399625 468
rect 399180 431 399625 459
rect 399180 422 399238 431
rect 399379 422 399437 431
rect 399567 422 399625 431
rect 399671 459 399729 468
rect 399859 459 399917 468
rect 400058 459 400116 468
rect 399671 431 400116 459
rect 399671 422 399729 431
rect 399859 422 399917 431
rect 400058 422 400116 431
rect 400468 459 400526 468
rect 400667 459 400725 468
rect 400855 459 400913 468
rect 400468 431 400913 459
rect 400468 422 400526 431
rect 400667 422 400725 431
rect 400855 422 400913 431
rect 400959 459 401017 468
rect 401147 459 401205 468
rect 401346 459 401404 468
rect 400959 431 401404 459
rect 400959 422 401017 431
rect 401147 422 401205 431
rect 401346 422 401404 431
rect 401756 459 401814 468
rect 401955 459 402013 468
rect 402143 459 402201 468
rect 401756 431 402201 459
rect 401756 422 401814 431
rect 401955 422 402013 431
rect 402143 422 402201 431
rect 402433 459 402491 468
rect 402621 459 402679 468
rect 402817 459 402875 468
rect 403007 459 403065 468
rect 403197 459 403255 468
rect 402433 431 403255 459
rect 402433 422 402491 431
rect 402621 422 402679 431
rect 402817 422 402875 431
rect 403007 422 403065 431
rect 403197 422 403255 431
rect 403953 459 404011 468
rect 404143 459 404201 468
rect 404333 459 404391 468
rect 404529 459 404587 468
rect 404717 459 404775 468
rect 403953 431 404775 459
rect 403953 422 404011 431
rect 404143 422 404201 431
rect 404333 422 404391 431
rect 404529 422 404587 431
rect 404717 422 404775 431
rect 405009 459 405067 468
rect 405197 459 405255 468
rect 405393 459 405451 468
rect 405583 459 405641 468
rect 405773 459 405831 468
rect 405009 431 405831 459
rect 405009 422 405067 431
rect 405197 422 405255 431
rect 405393 422 405451 431
rect 405583 422 405641 431
rect 405773 422 405831 431
rect 406529 459 406587 468
rect 406719 459 406777 468
rect 406909 459 406967 468
rect 407105 459 407163 468
rect 407293 459 407351 468
rect 406529 431 407351 459
rect 406529 422 406587 431
rect 406719 422 406777 431
rect 406909 422 406967 431
rect 407105 422 407163 431
rect 407293 422 407351 431
rect 407677 459 407735 468
rect 407865 459 407923 468
rect 408061 459 408119 468
rect 408251 459 408309 468
rect 408441 459 408499 468
rect 407677 431 408499 459
rect 407677 422 407735 431
rect 407865 422 407923 431
rect 408061 422 408119 431
rect 408251 422 408309 431
rect 408441 422 408499 431
rect 409197 459 409255 468
rect 409387 459 409445 468
rect 409577 459 409635 468
rect 409773 459 409831 468
rect 409961 459 410019 468
rect 409197 431 410019 459
rect 409197 422 409255 431
rect 409387 422 409445 431
rect 409577 422 409635 431
rect 409773 422 409831 431
rect 409961 422 410019 431
rect 410253 459 410311 468
rect 410441 459 410499 468
rect 410637 459 410695 468
rect 410827 459 410885 468
rect 411017 459 411075 468
rect 410253 431 411075 459
rect 410253 422 410311 431
rect 410441 422 410499 431
rect 410637 422 410695 431
rect 410827 422 410885 431
rect 411017 422 411075 431
rect 411773 459 411831 468
rect 411963 459 412021 468
rect 412153 459 412211 468
rect 412349 459 412407 468
rect 412537 459 412595 468
rect 411773 431 412595 459
rect 411773 422 411831 431
rect 411963 422 412021 431
rect 412153 422 412211 431
rect 412349 422 412407 431
rect 412537 422 412595 431
rect 101769 388 101837 397
rect 102101 388 102159 397
rect 102850 388 102908 397
rect 101769 360 102908 388
rect 101769 351 101837 360
rect 102101 351 102159 360
rect 102850 351 102908 360
rect 103793 388 103861 397
rect 104125 388 104183 397
rect 104874 388 104932 397
rect 103793 360 104932 388
rect 103793 351 103861 360
rect 104125 351 104183 360
rect 104874 351 104932 360
rect 105909 388 105977 397
rect 106317 388 106375 397
rect 107001 388 107069 397
rect 115130 388 115188 397
rect 115430 388 115488 397
rect 105909 360 107069 388
rect 105909 351 105977 360
rect 106317 351 106375 360
rect 107001 351 107069 360
rect 108221 360 109287 388
rect 108221 342 108279 360
rect 108617 342 108675 360
rect 109229 342 109287 360
rect 110337 360 111403 388
rect 110337 342 110395 360
rect 110733 342 110791 360
rect 111345 342 111403 360
rect 112545 360 113611 388
rect 112545 342 112603 360
rect 112941 342 112999 360
rect 113553 342 113611 360
rect 115130 360 115488 388
rect 115130 351 115188 360
rect 115430 351 115488 360
rect 116418 388 116476 397
rect 116718 388 116776 397
rect 116418 360 116776 388
rect 116418 351 116476 360
rect 116718 351 116776 360
rect 117787 388 117845 394
rect 118098 388 118156 394
rect 117787 360 118156 388
rect 117787 348 117845 360
rect 118098 348 118156 360
rect 270047 388 270105 397
rect 270945 388 271003 397
rect 271751 388 271809 397
rect 270047 360 271809 388
rect 270047 351 270105 360
rect 270945 351 271003 360
rect 271751 351 271809 360
rect 273362 388 273422 397
rect 274326 388 274384 397
rect 275048 388 275107 397
rect 273362 360 275107 388
rect 273362 351 273422 360
rect 274326 351 274384 360
rect 275048 351 275107 360
rect 276306 388 276366 397
rect 277270 388 277328 397
rect 277992 388 278051 397
rect 276306 360 278051 388
rect 276306 351 276366 360
rect 277270 351 277328 360
rect 277992 351 278051 360
rect 279260 388 279320 397
rect 280306 388 280364 397
rect 281028 388 281087 397
rect 279260 360 281087 388
rect 279260 351 279320 360
rect 280306 351 280364 360
rect 281028 351 281087 360
rect 282010 388 282070 397
rect 282974 388 283032 397
rect 283696 388 283755 397
rect 282010 360 283755 388
rect 282010 351 282070 360
rect 282974 351 283032 360
rect 283696 351 283755 360
rect 284678 388 284738 397
rect 285642 388 285700 397
rect 286364 388 286423 397
rect 284678 360 286423 388
rect 284678 351 284738 360
rect 285642 351 285700 360
rect 286364 351 286423 360
rect 288037 388 288105 397
rect 288333 388 288401 397
rect 288853 388 288911 397
rect 288037 360 288911 388
rect 288037 351 288105 360
rect 288333 351 288401 360
rect 288853 351 288911 360
rect 291073 388 291141 397
rect 291369 388 291437 397
rect 291889 388 291947 397
rect 291073 360 291947 388
rect 291073 351 291141 360
rect 291369 351 291437 360
rect 291889 351 291947 360
rect 294293 388 294361 397
rect 294589 388 294657 397
rect 295110 388 295178 397
rect 294293 360 295178 388
rect 294293 351 294361 360
rect 294589 351 294657 360
rect 295110 351 295178 360
rect 297053 388 297121 397
rect 297349 388 297417 397
rect 297870 388 297938 397
rect 297053 360 297938 388
rect 297053 351 297121 360
rect 297349 351 297417 360
rect 297870 351 297938 360
rect 299997 388 300065 397
rect 300293 388 300361 397
rect 300814 388 300882 397
rect 299997 360 300882 388
rect 299997 351 300065 360
rect 300293 351 300361 360
rect 300814 351 300882 360
rect 302439 388 302497 397
rect 303423 388 303481 397
rect 303735 388 303793 397
rect 302439 360 303793 388
rect 302439 351 302497 360
rect 303423 351 303481 360
rect 303735 351 303793 360
rect 304923 388 304981 397
rect 305907 388 305965 397
rect 306219 388 306277 397
rect 319825 388 319883 397
rect 321357 388 321425 397
rect 321915 388 321983 397
rect 304923 360 306277 388
rect 304923 351 304981 360
rect 305907 351 305965 360
rect 306219 351 306277 360
rect 307677 360 309050 388
rect 307677 342 307735 360
rect 308667 342 308735 360
rect 308982 342 309050 360
rect 309885 360 311255 388
rect 309885 342 309943 360
rect 310875 342 310943 360
rect 311187 342 311255 360
rect 312185 360 313555 388
rect 312185 342 312243 360
rect 313175 342 313243 360
rect 313487 342 313555 360
rect 319825 360 321983 388
rect 319825 351 319883 360
rect 321357 351 321425 360
rect 321915 351 321983 360
rect 322953 388 323011 397
rect 324485 388 324553 397
rect 325043 388 325111 397
rect 322953 360 325111 388
rect 322953 351 323011 360
rect 324485 351 324553 360
rect 325043 351 325111 360
rect 325249 388 325307 397
rect 325613 388 325671 397
rect 325249 360 325671 388
rect 325249 351 325307 360
rect 325613 351 325671 360
rect 347882 388 347942 397
rect 348846 388 348904 397
rect 349568 388 349627 397
rect 347882 360 349627 388
rect 347882 351 347942 360
rect 348846 351 348904 360
rect 349568 351 349627 360
rect 366821 388 366879 397
rect 367281 388 367339 397
rect 367649 388 367707 397
rect 368109 388 368167 397
rect 366821 360 368167 388
rect 366821 351 366879 360
rect 367281 351 367339 360
rect 367649 351 367707 360
rect 368109 351 368167 360
rect 368753 388 368811 397
rect 369397 388 369455 397
rect 370041 388 370099 397
rect 370685 388 370743 397
rect 368753 360 370743 388
rect 368753 351 368811 360
rect 369397 351 369455 360
rect 370041 351 370099 360
rect 370685 351 370743 360
rect 371725 388 371783 397
rect 371913 388 371971 397
rect 372861 388 372919 397
rect 373049 388 373107 397
rect 374301 388 374359 397
rect 374489 388 374547 397
rect 375437 388 375495 397
rect 375625 388 375683 397
rect 371725 360 375683 388
rect 371725 351 371783 360
rect 371913 351 371971 360
rect 372861 351 372919 360
rect 373049 351 373107 360
rect 374301 351 374359 360
rect 374489 351 374547 360
rect 375437 351 375495 360
rect 375625 351 375683 360
rect 376573 388 376631 397
rect 377033 388 377091 397
rect 377401 388 377459 397
rect 377861 388 377919 397
rect 378229 388 378287 397
rect 378689 388 378747 397
rect 379057 388 379115 397
rect 379517 388 379575 397
rect 376573 360 379575 388
rect 376573 351 376631 360
rect 377033 351 377091 360
rect 377401 351 377459 360
rect 377861 351 377919 360
rect 378229 351 378287 360
rect 378689 351 378747 360
rect 379057 351 379115 360
rect 379517 351 379575 360
rect 380161 388 380219 397
rect 380805 388 380863 397
rect 381449 388 381507 397
rect 382093 388 382151 397
rect 382737 388 382795 397
rect 383381 388 383439 397
rect 384025 388 384083 397
rect 384669 388 384727 397
rect 380161 360 384727 388
rect 380161 351 380219 360
rect 380805 351 380863 360
rect 381449 351 381507 360
rect 382093 351 382151 360
rect 382737 351 382795 360
rect 383381 351 383439 360
rect 384025 351 384083 360
rect 384669 351 384727 360
rect 388961 388 389019 397
rect 389149 388 389207 397
rect 390309 388 390367 397
rect 390497 388 390555 397
rect 391445 388 391503 397
rect 391633 388 391691 397
rect 392793 388 392851 397
rect 392981 388 393039 397
rect 388961 360 393039 388
rect 388961 351 389019 360
rect 389149 351 389207 360
rect 390309 351 390367 360
rect 390497 351 390555 360
rect 391445 351 391503 360
rect 391633 351 391691 360
rect 392793 351 392851 360
rect 392981 351 393039 360
rect 393777 388 393835 397
rect 394237 388 394295 397
rect 394605 388 394663 397
rect 395065 388 395123 397
rect 395433 388 395491 397
rect 395893 388 395951 397
rect 396261 388 396319 397
rect 396721 388 396779 397
rect 393777 360 396779 388
rect 393777 351 393835 360
rect 394237 351 394295 360
rect 394605 351 394663 360
rect 395065 351 395123 360
rect 395433 351 395491 360
rect 395893 351 395951 360
rect 396261 351 396319 360
rect 396721 351 396779 360
rect 397365 388 397423 397
rect 398009 388 398067 397
rect 398653 388 398711 397
rect 399297 388 399355 397
rect 399941 388 399999 397
rect 400585 388 400643 397
rect 401229 388 401287 397
rect 401873 388 401931 397
rect 397365 360 401931 388
rect 397365 351 397423 360
rect 398009 351 398067 360
rect 398653 351 398711 360
rect 399297 351 399355 360
rect 399941 351 399999 360
rect 400585 351 400643 360
rect 401229 351 401287 360
rect 401873 351 401931 360
rect 402913 388 402971 397
rect 403101 388 403159 397
rect 404049 388 404107 397
rect 404237 388 404295 397
rect 405489 388 405547 397
rect 405677 388 405735 397
rect 406625 388 406683 397
rect 406813 388 406871 397
rect 408157 388 408215 397
rect 408345 388 408403 397
rect 409293 388 409351 397
rect 409481 388 409539 397
rect 410733 388 410791 397
rect 410921 388 410979 397
rect 411869 388 411927 397
rect 412057 388 412115 397
rect 402913 360 412115 388
rect 402913 351 402971 360
rect 403101 351 403159 360
rect 404049 351 404107 360
rect 404237 351 404295 360
rect 405489 351 405547 360
rect 405677 351 405735 360
rect 406625 351 406683 360
rect 406813 351 406871 360
rect 408157 351 408215 360
rect 408345 351 408403 360
rect 409293 351 409351 360
rect 409481 351 409539 360
rect 410733 351 410791 360
rect 410921 351 410979 360
rect 411869 351 411927 360
rect 412057 351 412115 360
rect 5905 320 5963 329
rect 6516 320 6574 329
rect 5905 292 6574 320
rect 5905 283 5963 292
rect 6516 283 6574 292
rect 33556 320 33624 329
rect 34162 320 34220 329
rect 33556 292 34220 320
rect 33556 283 33624 292
rect 34162 283 34220 292
rect 115028 320 115086 329
rect 115531 320 115589 329
rect 115028 292 115589 320
rect 115028 283 115086 292
rect 115531 283 115589 292
rect 116316 320 116374 329
rect 116819 320 116877 329
rect 147134 320 147192 329
rect 147861 320 147919 329
rect 116316 292 116877 320
rect 116316 283 116374 292
rect 116819 283 116877 292
rect 117696 292 118258 320
rect 117696 274 117754 292
rect 118199 274 118258 292
rect 147134 292 147919 320
rect 147134 283 147192 292
rect 147861 283 147919 292
rect 237703 320 237771 327
rect 238309 320 238368 329
rect 237703 292 238368 320
rect 237703 277 237771 292
rect 238309 279 238368 292
rect 271659 320 271717 329
rect 272349 320 272407 329
rect 271659 292 272407 320
rect 271659 283 271717 292
rect 272349 283 272407 292
rect 287547 320 287615 329
rect 288214 320 288272 329
rect 287547 292 288272 320
rect 287547 283 287615 292
rect 288214 283 288272 292
rect 288701 320 288769 329
rect 289159 320 289217 329
rect 288701 292 289217 320
rect 288701 283 288769 292
rect 289159 283 289217 292
rect 290583 320 290651 329
rect 291250 320 291308 329
rect 290583 292 291308 320
rect 290583 283 290651 292
rect 291250 283 291308 292
rect 291737 320 291805 329
rect 292195 320 292253 329
rect 291737 292 292253 320
rect 291737 283 291805 292
rect 292195 283 292253 292
rect 293803 320 293871 329
rect 294470 320 294528 329
rect 293803 292 294528 320
rect 293803 283 293871 292
rect 294470 283 294528 292
rect 294955 320 295023 329
rect 295393 320 295461 329
rect 294955 292 295461 320
rect 294955 283 295023 292
rect 295393 283 295461 292
rect 296563 320 296631 329
rect 297230 320 297288 329
rect 296563 292 297288 320
rect 296563 283 296631 292
rect 297230 283 297288 292
rect 297715 320 297783 329
rect 298186 320 298254 329
rect 297715 292 298254 320
rect 297715 283 297783 292
rect 298186 283 298254 292
rect 299507 320 299575 329
rect 300174 320 300232 329
rect 299507 292 300232 320
rect 299507 283 299575 292
rect 300174 283 300232 292
rect 300659 320 300727 329
rect 301130 320 301198 329
rect 300659 292 301198 320
rect 300659 283 300727 292
rect 301130 283 301198 292
rect 314861 320 314919 329
rect 315409 320 315467 329
rect 314861 292 315467 320
rect 314861 283 314919 292
rect 315409 283 315467 292
rect 316425 320 316483 329
rect 317000 320 317058 329
rect 316425 292 317058 320
rect 316425 283 316483 292
rect 317000 283 317058 292
rect 318092 320 318150 329
rect 318688 320 318746 329
rect 318092 292 318746 320
rect 318092 283 318150 292
rect 318688 283 318746 292
rect 319901 320 319969 329
rect 321265 320 321333 329
rect 322009 320 322077 329
rect 319901 292 322077 320
rect 319901 283 319969 292
rect 321265 283 321333 292
rect 322009 283 322077 292
rect 323029 320 323097 329
rect 324393 320 324461 329
rect 325137 320 325205 329
rect 323029 292 325205 320
rect 323029 283 323097 292
rect 324393 283 324461 292
rect 325137 283 325205 292
rect 328651 320 328719 329
rect 329771 320 329841 329
rect 328651 292 329841 320
rect 328651 283 328719 292
rect 329771 283 329841 292
rect 331349 320 331407 329
rect 331839 320 331897 329
rect 331349 292 331897 320
rect 331349 283 331407 292
rect 331839 283 331897 292
rect 333383 320 333441 329
rect 333873 320 333931 329
rect 333383 292 333931 320
rect 333383 283 333441 292
rect 333873 283 333931 292
rect 335611 320 335669 329
rect 336101 320 336159 329
rect 335611 292 336159 320
rect 335611 283 335669 292
rect 336101 283 336159 292
rect 339537 320 339595 329
rect 340761 320 340819 329
rect 339537 292 340819 320
rect 339537 283 339595 292
rect 340761 283 340819 292
rect 342113 320 342171 329
rect 342603 320 342661 329
rect 342113 292 342661 320
rect 342113 283 342171 292
rect 342603 283 342661 292
rect 344196 320 344254 329
rect 344686 320 344744 329
rect 344196 292 344744 320
rect 344196 283 344254 292
rect 344686 283 344744 292
rect 346395 320 346453 329
rect 346885 320 346943 329
rect 346395 292 346943 320
rect 346395 283 346453 292
rect 346885 283 346943 292
rect 95083 252 95243 261
rect 96817 252 96987 261
rect 95083 224 96987 252
rect 95083 215 95243 224
rect 96817 215 96987 224
rect 101688 252 101746 261
rect 102052 252 102110 261
rect 102760 252 102818 261
rect 101688 224 102818 252
rect 101688 215 101746 224
rect 102052 215 102110 224
rect 102760 215 102818 224
rect 103712 252 103770 261
rect 104076 252 104134 261
rect 104784 252 104842 261
rect 103712 224 104842 252
rect 103712 215 103770 224
rect 104076 215 104134 224
rect 104784 215 104842 224
rect 105828 252 105886 261
rect 106215 252 106273 261
rect 107001 252 107069 261
rect 105828 224 107069 252
rect 105828 215 105886 224
rect 106215 215 106273 224
rect 107001 215 107069 224
rect 102367 184 102517 193
rect 103083 184 103141 193
rect 102367 156 103141 184
rect 102367 147 102517 156
rect 103083 147 103141 156
rect 104391 184 104541 193
rect 105107 184 105165 193
rect 104391 156 105165 184
rect 104391 147 104541 156
rect 105107 147 105165 156
rect 106543 184 106693 193
rect 107270 184 107387 256
rect 109233 252 109291 262
rect 111349 252 111407 262
rect 113557 252 113615 262
rect 108734 224 109291 252
rect 108734 184 108777 224
rect 109233 216 109291 224
rect 110850 224 111407 252
rect 106543 156 107387 184
rect 106543 147 106693 156
rect 107329 147 107387 156
rect 108321 156 108777 184
rect 108321 138 108379 156
rect 108719 138 108777 156
rect 108944 184 109002 193
rect 109589 184 109647 193
rect 110850 184 110893 224
rect 111349 216 111407 224
rect 113058 224 113615 252
rect 108944 156 109647 184
rect 108944 147 109002 156
rect 109589 147 109647 156
rect 110437 156 110893 184
rect 110437 138 110495 156
rect 110835 138 110893 156
rect 111060 184 111118 193
rect 111705 184 111763 193
rect 113058 184 113101 224
rect 113557 216 113615 224
rect 122285 224 123050 252
rect 122285 206 122344 224
rect 122982 206 123050 224
rect 123297 233 124268 261
rect 146836 252 146904 261
rect 147665 252 147735 261
rect 123297 215 123356 233
rect 124210 215 124268 233
rect 124769 224 126232 252
rect 124769 206 124837 224
rect 126164 206 126232 224
rect 146836 224 147735 252
rect 146836 215 146904 224
rect 147665 215 147735 224
rect 173548 215 174005 261
rect 175055 252 175113 261
rect 175555 252 175623 261
rect 175055 224 175623 252
rect 175055 215 175113 224
rect 175555 215 175623 224
rect 270537 252 270595 261
rect 270845 252 270903 261
rect 271751 252 271809 261
rect 270537 224 270903 252
rect 270537 215 270595 224
rect 270845 215 270903 224
rect 271062 224 271809 252
rect 271062 193 271105 224
rect 271751 215 271809 224
rect 273307 252 273365 261
rect 274232 252 274290 261
rect 274979 252 275041 261
rect 273307 224 275041 252
rect 273307 215 273365 224
rect 274232 215 274290 224
rect 274979 215 275041 224
rect 276251 252 276309 261
rect 277176 252 277234 261
rect 277923 252 277985 261
rect 276251 224 277985 252
rect 276251 215 276309 224
rect 277176 215 277234 224
rect 277923 215 277985 224
rect 279355 252 279413 261
rect 280212 252 280270 261
rect 280959 252 281021 261
rect 279355 224 281021 252
rect 279355 215 279413 224
rect 280212 215 280270 224
rect 280959 215 281021 224
rect 281955 252 282013 261
rect 282880 252 282938 261
rect 283627 252 283689 261
rect 281955 224 283689 252
rect 281955 215 282013 224
rect 282880 215 282938 224
rect 283627 215 283689 224
rect 284623 252 284681 261
rect 285548 252 285606 261
rect 286295 252 286357 261
rect 284623 224 286357 252
rect 284623 215 284681 224
rect 285548 215 285606 224
rect 286295 215 286357 224
rect 287338 252 287396 261
rect 287741 252 287799 261
rect 287338 224 287799 252
rect 287338 215 287396 224
rect 287741 215 287799 224
rect 288129 252 288187 261
rect 289047 252 289115 261
rect 288129 224 289115 252
rect 288129 215 288187 224
rect 289047 215 289115 224
rect 290374 252 290432 261
rect 290777 252 290835 261
rect 290374 224 290835 252
rect 290374 215 290432 224
rect 290777 215 290835 224
rect 291165 252 291223 261
rect 292083 252 292151 261
rect 291165 224 292151 252
rect 291165 215 291223 224
rect 292083 215 292151 224
rect 293596 252 293654 261
rect 293997 252 294055 261
rect 293596 224 294055 252
rect 293596 215 293654 224
rect 293997 215 294055 224
rect 294395 252 294453 260
rect 295268 252 295346 261
rect 294395 224 295346 252
rect 294395 214 294453 224
rect 295268 215 295346 224
rect 296356 252 296414 261
rect 296757 252 296815 261
rect 296356 224 296815 252
rect 296356 215 296414 224
rect 296757 215 296815 224
rect 297155 252 297213 260
rect 298074 252 298152 261
rect 297155 224 298152 252
rect 297155 214 297213 224
rect 298074 215 298152 224
rect 299300 252 299358 261
rect 299701 252 299759 261
rect 299300 224 299759 252
rect 299300 215 299358 224
rect 299701 215 299759 224
rect 300099 252 300157 260
rect 301018 252 301096 261
rect 300099 224 301096 252
rect 300099 214 300157 224
rect 301018 215 301096 224
rect 315497 252 315555 261
rect 315736 252 315794 261
rect 315497 224 315794 252
rect 315497 215 315555 224
rect 315736 215 315794 224
rect 317102 252 317160 261
rect 317300 252 317358 261
rect 317102 224 317358 252
rect 317102 215 317160 224
rect 317300 215 317358 224
rect 318779 252 318837 261
rect 318988 252 319046 261
rect 318779 224 319046 252
rect 318779 215 318837 224
rect 318988 215 319046 224
rect 322121 252 322179 261
rect 322527 252 322585 261
rect 322121 224 322585 252
rect 322121 215 322179 224
rect 322527 215 322585 224
rect 337953 252 338011 261
rect 338485 252 338543 261
rect 337953 224 338543 252
rect 337953 215 338011 224
rect 338485 215 338543 224
rect 347827 252 347885 261
rect 348752 252 348810 261
rect 349499 252 349561 261
rect 347827 224 349561 252
rect 347827 215 347885 224
rect 348752 215 348810 224
rect 349499 215 349561 224
rect 349823 193 349881 262
rect 111060 156 111763 184
rect 111060 147 111118 156
rect 111705 147 111763 156
rect 112645 156 113101 184
rect 112645 138 112703 156
rect 113043 138 113101 156
rect 113268 184 113326 193
rect 113913 184 113971 193
rect 113268 156 113971 184
rect 113268 147 113326 156
rect 113913 147 113971 156
rect 146934 184 146992 193
rect 147530 184 147598 193
rect 146934 156 147598 184
rect 146934 147 146992 156
rect 147530 147 147598 156
rect 149262 184 149320 193
rect 149868 184 149936 193
rect 149262 156 149936 184
rect 149262 147 149320 156
rect 149868 147 149936 156
rect 150560 184 150618 193
rect 151574 184 151642 193
rect 150560 156 151642 184
rect 150560 147 150618 156
rect 151574 147 151642 156
rect 270146 184 270204 193
rect 271047 184 271105 193
rect 270146 156 271105 184
rect 270146 147 270204 156
rect 271047 147 271105 156
rect 271233 184 271291 193
rect 272059 184 272117 193
rect 271233 156 272117 184
rect 271233 147 271291 156
rect 272059 147 272117 156
rect 274577 184 274728 193
rect 275371 184 275429 193
rect 274577 156 275429 184
rect 274577 147 274728 156
rect 275371 147 275429 156
rect 277521 184 277672 193
rect 278315 184 278373 193
rect 277521 156 278373 184
rect 277521 147 277672 156
rect 278315 147 278373 156
rect 280557 184 280708 193
rect 281351 184 281409 193
rect 280557 156 281409 184
rect 280557 147 280708 156
rect 281351 147 281409 156
rect 283225 184 283376 193
rect 284019 184 284077 193
rect 283225 156 284077 184
rect 283225 147 283376 156
rect 284019 147 284077 156
rect 285893 184 286044 193
rect 286680 184 286738 193
rect 285893 156 286738 184
rect 285893 147 286044 156
rect 286680 147 286738 156
rect 303341 184 303399 193
rect 303737 184 303795 193
rect 303341 156 303795 184
rect 303341 147 303399 156
rect 303737 147 303795 156
rect 305813 184 305871 193
rect 306221 184 306279 193
rect 314963 184 315021 193
rect 315296 184 315354 193
rect 305813 156 306279 184
rect 305813 147 305871 156
rect 306221 147 306279 156
rect 307775 156 309064 184
rect 206946 116 207004 125
rect 208376 116 208434 125
rect 206946 88 208434 116
rect 206946 79 207004 88
rect 208376 79 208434 88
rect 302513 116 302581 125
rect 303341 116 303369 147
rect 302513 88 303369 116
rect 304997 116 305065 125
rect 305813 116 305841 147
rect 307775 138 307833 156
rect 308565 138 308633 156
rect 309002 138 309064 156
rect 309983 156 311255 184
rect 309983 138 310041 156
rect 310773 138 310841 156
rect 311187 138 311255 156
rect 312283 156 313555 184
rect 312283 138 312341 156
rect 313073 138 313141 156
rect 313487 138 313555 156
rect 314963 156 315354 184
rect 314963 147 315021 156
rect 315296 147 315354 156
rect 316527 184 316585 193
rect 316898 184 316956 193
rect 316527 156 316956 184
rect 316527 147 316585 156
rect 316898 147 316956 156
rect 318194 184 318252 193
rect 318586 184 318644 193
rect 318194 156 318644 184
rect 318194 147 318252 156
rect 318586 147 318644 156
rect 320509 184 320567 193
rect 322428 184 322486 193
rect 320509 156 322486 184
rect 320509 147 320567 156
rect 322428 147 322486 156
rect 323637 184 323695 193
rect 325705 184 325763 193
rect 323637 156 325763 184
rect 323637 147 323695 156
rect 325705 147 325763 156
rect 331543 184 331601 193
rect 331839 184 331897 193
rect 332135 184 332193 193
rect 331543 156 332193 184
rect 331543 147 331601 156
rect 331839 147 331897 156
rect 332135 147 332193 156
rect 333577 184 333635 193
rect 333873 184 333931 193
rect 334169 184 334227 193
rect 333577 156 334227 184
rect 333577 147 333635 156
rect 333873 147 333931 156
rect 334169 147 334227 156
rect 335805 184 335863 193
rect 336101 184 336159 193
rect 336397 184 336455 193
rect 335805 156 336455 184
rect 335805 147 335863 156
rect 336101 147 336159 156
rect 336397 147 336455 156
rect 340241 156 340911 185
rect 340241 139 340299 156
rect 340853 139 340911 156
rect 342307 184 342365 193
rect 342603 184 342661 193
rect 342899 184 342957 193
rect 342307 156 342957 184
rect 342307 147 342365 156
rect 342603 147 342661 156
rect 342899 147 342957 156
rect 344390 184 344448 193
rect 344686 184 344744 193
rect 344982 184 345040 193
rect 344390 156 345040 184
rect 344390 147 344448 156
rect 344686 147 344744 156
rect 344982 147 345040 156
rect 346589 184 346657 193
rect 346885 184 346943 193
rect 347181 184 347239 193
rect 346589 156 347239 184
rect 346589 147 346657 156
rect 346885 147 346943 156
rect 347181 147 347239 156
rect 349097 184 349248 193
rect 349823 184 349949 193
rect 349097 156 349949 184
rect 349097 147 349248 156
rect 349891 147 349949 156
rect 304997 88 305841 116
rect 319979 116 320037 125
rect 320585 116 320653 125
rect 302513 79 302581 88
rect 304997 79 305065 88
rect 319979 79 320653 116
rect 320681 116 320749 125
rect 321141 116 321209 125
rect 320681 79 321209 116
rect 323107 116 323165 125
rect 323713 116 323781 125
rect 323107 79 323781 116
rect 323809 116 323877 125
rect 324269 116 324337 125
rect 323809 79 324337 116
rect 331645 116 331703 125
rect 332237 116 332295 125
rect 331645 88 332295 116
rect 331645 79 331703 88
rect 332237 79 332295 88
rect 333679 116 333737 125
rect 334271 116 334329 125
rect 333679 88 334329 116
rect 333679 79 333737 88
rect 334271 79 334329 88
rect 335899 116 335959 125
rect 336499 116 336557 125
rect 335899 88 336557 116
rect 335899 79 335959 88
rect 336499 79 336557 88
rect 342409 116 342467 125
rect 343001 116 343059 125
rect 342409 88 343059 116
rect 342409 79 342467 88
rect 343001 79 343059 88
rect 344492 116 344550 125
rect 345084 116 345142 125
rect 344492 88 345142 116
rect 344492 79 344550 88
rect 345084 79 345142 88
rect 346691 116 346749 125
rect 347283 116 347341 125
rect 346691 88 347341 116
rect 346691 79 346749 88
rect 347283 79 347341 88
rect 0 14 412804 48
rect 412852 14 412880 1074
rect -76 -14 412880 14
rect 0 -48 412804 -14
<< via2 >>
rect 35720 1114 35776 1116
rect 35800 1114 35856 1116
rect 35720 1062 35730 1114
rect 35730 1062 35776 1114
rect 35800 1062 35846 1114
rect 35846 1062 35856 1114
rect 35720 1060 35776 1062
rect 35800 1060 35856 1062
rect 31233 876 31289 878
rect 31313 876 31369 878
rect 31233 824 31243 876
rect 31243 824 31289 876
rect 31313 824 31359 876
rect 31359 824 31369 876
rect 31233 822 31289 824
rect 31313 822 31369 824
rect 35071 876 35127 878
rect 35151 876 35207 878
rect 35071 824 35094 876
rect 35094 824 35127 876
rect 35151 824 35158 876
rect 35158 824 35207 876
rect 35071 822 35127 824
rect 35151 822 35207 824
rect 35720 570 35776 572
rect 35800 570 35856 572
rect 35720 518 35730 570
rect 35730 518 35776 570
rect 35800 518 35846 570
rect 35846 518 35856 570
rect 35720 516 35776 518
rect 35800 516 35856 518
<< obsm2 >>
rect 35711 1060 35720 1116
rect 35776 1114 35800 1116
rect 35782 1062 35794 1114
rect 35776 1060 35800 1062
rect 35856 1060 35865 1116
rect 31233 878 31369 887
rect 31289 876 31313 878
rect 31295 824 31307 876
rect 31289 822 31313 824
rect 35062 822 35071 878
rect 35127 876 35151 878
rect 35207 876 35216 878
rect 35146 824 35151 876
rect 35210 824 35216 876
rect 35127 822 35151 824
rect 35207 822 35216 824
rect 31233 813 31369 822
rect 35711 516 35720 572
rect 35776 570 35800 572
rect 35782 518 35794 570
rect 35776 516 35800 518
rect 35856 516 35865 572
<< obsm3 >>
rect 35710 1120 35866 1121
rect 35710 1056 35716 1120
rect 35780 1056 35796 1120
rect 35860 1056 35866 1120
rect 35710 1055 35866 1056
rect 31223 882 31379 883
rect 35061 882 35217 883
rect 31223 818 31229 882
rect 31293 818 31309 882
rect 31373 818 31379 882
rect 34541 818 34547 882
rect 34611 818 34627 882
rect 34691 818 34697 882
rect 35061 818 35067 882
rect 35131 818 35147 882
rect 35211 818 35217 882
rect 31223 817 31379 818
rect 35061 817 35217 818
rect 35710 576 35866 577
rect 35710 512 35716 576
rect 35780 512 35796 576
rect 35860 512 35866 576
rect 35710 511 35866 512
<< via3 >>
rect 35716 1116 35780 1120
rect 35716 1060 35720 1116
rect 35720 1060 35776 1116
rect 35776 1060 35780 1116
rect 35716 1056 35780 1060
rect 35796 1116 35860 1120
rect 35796 1060 35800 1116
rect 35800 1060 35856 1116
rect 35856 1060 35860 1116
rect 35796 1056 35860 1060
rect 31229 878 31293 882
rect 31229 822 31233 878
rect 31233 822 31289 878
rect 31289 822 31293 878
rect 31229 818 31293 822
rect 31309 878 31373 882
rect 31309 822 31313 878
rect 31313 822 31369 878
rect 31369 822 31373 878
rect 31309 818 31373 822
rect 34547 818 34611 882
rect 34627 818 34691 882
rect 35067 878 35131 882
rect 35067 822 35071 878
rect 35071 822 35127 878
rect 35127 822 35131 878
rect 35067 818 35131 822
rect 35147 878 35211 882
rect 35147 822 35151 878
rect 35151 822 35207 878
rect 35207 822 35211 878
rect 35147 818 35211 822
rect 35716 572 35780 576
rect 35716 516 35720 572
rect 35720 516 35776 572
rect 35776 516 35780 572
rect 35716 512 35780 516
rect 35796 572 35860 576
rect 35796 516 35800 572
rect 35800 516 35856 572
rect 35856 516 35860 572
rect 35796 512 35860 516
<< obsm4 >>
rect 35670 1120 35906 1267
rect 35670 1056 35716 1120
rect 35780 1056 35796 1120
rect 35860 1056 35906 1120
rect 35670 1031 35906 1056
rect 30818 716 31138 952
rect 34456 882 34692 934
rect 34456 818 34547 882
rect 34611 818 34627 882
rect 34691 818 34692 882
rect 34456 698 34692 818
rect 34976 882 35212 934
rect 34976 818 35067 882
rect 35131 818 35147 882
rect 35211 818 35212 882
rect 34976 698 35212 818
rect 35670 576 35906 601
rect 35670 512 35716 576
rect 35780 512 35796 576
rect 35860 512 35906 576
rect 35670 365 35906 512
<< via4 >>
rect 31138 882 31374 952
rect 31138 818 31229 882
rect 31229 818 31293 882
rect 31293 818 31309 882
rect 31309 818 31373 882
rect 31373 818 31374 882
rect 31138 716 31374 818
<< metal5 >>
rect 35556 1179 36019 1322
rect 35596 1119 36019 1179
rect 35556 976 36019 1119
rect 35556 513 36019 656
rect 35596 453 36019 513
rect 35556 310 36019 453
<< obsm5 >>
rect 30794 952 31398 976
rect 30794 716 31138 952
rect 31374 716 31398 952
rect 30794 699 31398 716
rect 30794 656 31398 698
rect 34432 656 34896 976
rect 34916 323 35236 1309
rect 35556 1139 35576 1159
rect 35556 473 35576 493
<< labels >>
rlabel metal5 s 35596 1119 36019 1179 6 VGND
port 1 nsew ground default
rlabel metal5 s 35556 1179 36019 1322 6 VGND
port 1 nsew ground default
rlabel metal5 s 35556 976 36019 1119 6 VGND
port 1 nsew ground default
rlabel metal5 s 35596 453 36019 513 6 VPWR
port 2 nsew power default
rlabel metal5 s 35556 513 36019 656 6 VPWR
port 2 nsew power default
rlabel metal5 s 35556 310 36019 453 6 VPWR
port 2 nsew power default
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX -2976 -3165 415786 3725
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3646290
string GDS_START 3609774
<< end >>
