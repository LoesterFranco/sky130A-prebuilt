magic
tech sky130A
magscale 1 2
timestamp 1599588209
<< nwell >>
rect -38 335 806 704
rect -38 332 232 335
rect 638 332 806 335
<< pwell >>
rect 0 0 768 49
<< scpmos >>
rect 86 368 116 592
rect 368 392 398 592
rect 452 392 482 592
rect 542 392 572 592
rect 650 392 680 592
<< nmoslvt >>
rect 84 74 114 222
rect 356 139 386 267
rect 450 139 480 267
rect 536 139 566 267
rect 654 130 684 258
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 192 171 222
rect 306 199 356 267
rect 114 158 125 192
rect 159 158 171 192
rect 114 120 171 158
rect 299 186 356 199
rect 299 152 311 186
rect 345 152 356 186
rect 299 139 356 152
rect 386 255 450 267
rect 386 221 401 255
rect 435 221 450 255
rect 386 139 450 221
rect 480 186 536 267
rect 480 152 491 186
rect 525 152 536 186
rect 480 139 536 152
rect 566 258 616 267
rect 566 176 654 258
rect 566 142 594 176
rect 628 142 654 176
rect 566 139 654 142
rect 114 86 125 120
rect 159 86 171 120
rect 114 74 171 86
rect 581 130 654 139
rect 684 256 734 258
rect 684 244 741 256
rect 684 210 695 244
rect 729 210 741 244
rect 684 176 741 210
rect 684 142 695 176
rect 729 142 741 176
rect 684 130 741 142
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 497 86 546
rect 27 463 39 497
rect 73 463 86 497
rect 27 414 86 463
rect 27 380 39 414
rect 73 380 86 414
rect 27 368 86 380
rect 116 583 368 592
rect 116 549 130 583
rect 164 549 230 583
rect 264 549 320 583
rect 354 549 368 583
rect 116 515 368 549
rect 116 481 130 515
rect 164 481 230 515
rect 264 481 320 515
rect 354 481 368 515
rect 116 447 368 481
rect 116 413 130 447
rect 164 413 230 447
rect 264 413 320 447
rect 354 413 368 447
rect 116 392 368 413
rect 398 392 452 592
rect 482 580 542 592
rect 482 546 495 580
rect 529 546 542 580
rect 482 512 542 546
rect 482 478 495 512
rect 529 478 542 512
rect 482 444 542 478
rect 482 410 495 444
rect 529 410 542 444
rect 482 392 542 410
rect 572 392 650 592
rect 680 580 739 592
rect 680 546 693 580
rect 727 546 739 580
rect 680 512 739 546
rect 680 478 693 512
rect 727 478 739 512
rect 680 444 739 478
rect 680 410 693 444
rect 727 410 739 444
rect 680 392 739 410
rect 116 368 169 392
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 125 158 159 192
rect 311 152 345 186
rect 401 221 435 255
rect 491 152 525 186
rect 594 142 628 176
rect 125 86 159 120
rect 695 210 729 244
rect 695 142 729 176
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 130 549 164 583
rect 230 549 264 583
rect 320 549 354 583
rect 130 481 164 515
rect 230 481 264 515
rect 320 481 354 515
rect 130 413 164 447
rect 230 413 264 447
rect 320 413 354 447
rect 495 546 529 580
rect 495 478 529 512
rect 495 410 529 444
rect 693 546 727 580
rect 693 478 727 512
rect 693 410 727 444
<< poly >>
rect 86 592 116 618
rect 368 592 398 618
rect 452 592 482 618
rect 542 592 572 618
rect 650 592 680 618
rect 368 377 398 392
rect 452 377 482 392
rect 542 377 572 392
rect 650 377 680 392
rect 86 353 116 368
rect 365 360 401 377
rect 83 326 119 353
rect 267 344 401 360
rect 83 310 219 326
rect 83 276 101 310
rect 135 276 169 310
rect 203 276 219 310
rect 267 310 283 344
rect 317 310 351 344
rect 385 310 401 344
rect 267 294 401 310
rect 83 260 219 276
rect 356 267 386 294
rect 449 282 485 377
rect 539 360 575 377
rect 647 360 683 377
rect 533 344 599 360
rect 533 310 549 344
rect 583 310 599 344
rect 533 294 599 310
rect 647 344 713 360
rect 647 310 663 344
rect 697 310 713 344
rect 647 294 713 310
rect 450 267 480 282
rect 536 267 566 294
rect 84 222 114 260
rect 654 258 684 294
rect 356 113 386 139
rect 450 117 480 139
rect 428 101 494 117
rect 536 113 566 139
rect 654 104 684 130
rect 84 48 114 74
rect 428 67 444 101
rect 478 67 494 101
rect 428 51 494 67
<< polycont >>
rect 101 276 135 310
rect 169 276 203 310
rect 283 310 317 344
rect 351 310 385 344
rect 549 310 583 344
rect 663 310 697 344
rect 444 67 478 101
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 17 580 89 596
rect 17 546 39 580
rect 73 546 89 580
rect 17 497 89 546
rect 17 463 39 497
rect 73 463 89 497
rect 17 414 89 463
rect 17 380 39 414
rect 73 380 89 414
rect 123 583 370 649
rect 123 549 130 583
rect 164 549 230 583
rect 264 549 320 583
rect 354 549 370 583
rect 123 515 370 549
rect 123 481 130 515
rect 164 481 230 515
rect 264 481 320 515
rect 354 481 370 515
rect 123 447 370 481
rect 123 413 130 447
rect 164 413 230 447
rect 264 413 320 447
rect 354 413 370 447
rect 479 580 545 596
rect 479 546 495 580
rect 529 546 545 580
rect 479 512 545 546
rect 479 478 495 512
rect 529 478 545 512
rect 479 444 545 478
rect 479 428 495 444
rect 123 397 370 413
rect 435 410 495 428
rect 529 410 545 444
rect 17 364 89 380
rect 435 394 545 410
rect 677 580 743 649
rect 677 546 693 580
rect 727 546 743 580
rect 677 512 743 546
rect 677 478 693 512
rect 727 478 743 512
rect 677 444 743 478
rect 677 410 693 444
rect 727 410 743 444
rect 677 394 743 410
rect 17 226 51 364
rect 267 344 401 360
rect 85 310 219 326
rect 85 276 101 310
rect 135 276 169 310
rect 203 276 219 310
rect 267 310 283 344
rect 317 310 351 344
rect 385 310 401 344
rect 267 294 401 310
rect 85 260 219 276
rect 435 260 469 394
rect 505 344 599 360
rect 505 310 549 344
rect 583 310 599 344
rect 505 294 599 310
rect 647 344 743 360
rect 647 310 663 344
rect 697 310 743 344
rect 647 294 743 310
rect 185 255 469 260
rect 185 226 401 255
rect 17 210 73 226
rect 381 221 401 226
rect 435 221 469 255
rect 507 244 745 260
rect 507 226 695 244
rect 17 176 39 210
rect 17 120 73 176
rect 17 86 39 120
rect 17 70 73 86
rect 109 158 125 192
rect 159 158 175 192
rect 507 187 541 226
rect 679 210 695 226
rect 729 210 745 244
rect 109 120 175 158
rect 295 186 541 187
rect 295 152 311 186
rect 345 152 491 186
rect 525 152 541 186
rect 295 151 541 152
rect 577 176 645 192
rect 577 142 594 176
rect 628 142 645 176
rect 109 86 125 120
rect 159 86 175 120
rect 109 17 175 86
rect 217 117 261 134
rect 217 101 494 117
rect 217 67 444 101
rect 478 67 494 101
rect 217 51 494 67
rect 577 17 645 142
rect 679 176 745 210
rect 679 142 695 176
rect 729 142 745 176
rect 679 126 745 142
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o22a_1
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 223 94 257 128 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 768 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1210476
string GDS_START 1202926
<< end >>
