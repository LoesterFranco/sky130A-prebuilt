magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1748 561
rect 119 359 161 527
rect 279 359 329 527
rect 1223 325 1273 425
rect 1391 325 1441 425
rect 1223 291 1441 325
rect 1671 291 1717 527
rect 79 215 361 257
rect 415 215 750 257
rect 797 215 1137 257
rect 1223 181 1293 291
rect 1562 215 1731 257
rect 35 17 69 179
rect 103 145 1449 181
rect 103 51 169 145
rect 203 17 237 111
rect 271 51 337 145
rect 371 17 405 111
rect 439 51 505 145
rect 539 17 573 111
rect 607 51 673 145
rect 707 17 845 111
rect 879 51 945 145
rect 979 17 1013 111
rect 1047 51 1113 145
rect 1147 17 1181 111
rect 1215 51 1281 145
rect 1315 17 1349 111
rect 1383 51 1449 145
rect 1483 17 1517 111
rect 1671 17 1717 181
rect 0 -17 1748 17
<< obsli1 >>
rect 19 325 85 493
rect 195 325 245 493
rect 363 459 749 493
rect 363 325 413 459
rect 19 291 413 325
rect 447 325 497 425
rect 531 359 581 459
rect 615 325 665 425
rect 699 359 749 459
rect 803 459 1525 493
rect 803 359 853 459
rect 887 325 937 425
rect 971 359 1021 459
rect 1055 325 1105 425
rect 447 291 1105 325
rect 1139 291 1189 459
rect 1307 359 1357 459
rect 1475 359 1525 459
rect 1570 325 1637 493
rect 1494 291 1637 325
rect 1494 257 1528 291
rect 1327 215 1528 257
rect 1494 181 1528 215
rect 1494 147 1637 181
rect 1562 51 1637 147
<< metal1 >>
rect 0 496 1748 592
rect 0 -48 1748 48
<< labels >>
rlabel locali s 79 215 361 257 6 A
port 1 nsew signal input
rlabel locali s 415 215 750 257 6 B
port 2 nsew signal input
rlabel locali s 797 215 1137 257 6 C
port 3 nsew signal input
rlabel locali s 1562 215 1731 257 6 D_N
port 4 nsew signal input
rlabel locali s 1391 325 1441 425 6 Y
port 5 nsew signal output
rlabel locali s 1383 51 1449 145 6 Y
port 5 nsew signal output
rlabel locali s 1223 325 1273 425 6 Y
port 5 nsew signal output
rlabel locali s 1223 291 1441 325 6 Y
port 5 nsew signal output
rlabel locali s 1223 181 1293 291 6 Y
port 5 nsew signal output
rlabel locali s 1215 51 1281 145 6 Y
port 5 nsew signal output
rlabel locali s 1047 51 1113 145 6 Y
port 5 nsew signal output
rlabel locali s 879 51 945 145 6 Y
port 5 nsew signal output
rlabel locali s 607 51 673 145 6 Y
port 5 nsew signal output
rlabel locali s 439 51 505 145 6 Y
port 5 nsew signal output
rlabel locali s 271 51 337 145 6 Y
port 5 nsew signal output
rlabel locali s 103 145 1449 181 6 Y
port 5 nsew signal output
rlabel locali s 103 51 169 145 6 Y
port 5 nsew signal output
rlabel locali s 1671 17 1717 181 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1483 17 1517 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1315 17 1349 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1147 17 1181 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 979 17 1013 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 707 17 845 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 539 17 573 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 371 17 405 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 203 17 237 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 35 17 69 179 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 1748 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1748 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1671 291 1717 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 279 359 329 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 119 359 161 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 1748 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 1748 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1748 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1191072
string GDS_START 1177578
<< end >>
