magic
tech sky130A
magscale 1 2
timestamp 1599588209
<< nwell >>
rect -38 332 1574 704
rect 782 316 996 332
<< pwell >>
rect 0 0 1536 49
<< scpmos >>
rect 86 424 116 592
rect 164 424 194 592
rect 383 368 413 536
rect 585 379 615 547
rect 692 492 722 576
rect 770 492 800 576
rect 871 352 901 576
rect 1073 403 1103 571
rect 1212 403 1242 571
rect 1302 403 1332 571
rect 1403 368 1433 592
<< nmoslvt >>
rect 84 112 114 222
rect 170 112 200 222
rect 288 74 318 222
rect 536 74 566 184
rect 637 80 667 164
rect 709 80 739 164
rect 845 74 875 222
rect 1041 74 1071 222
rect 1136 94 1166 222
rect 1208 94 1238 222
rect 1423 74 1453 222
<< ndiff >>
rect 27 183 84 222
rect 27 149 39 183
rect 73 149 84 183
rect 27 112 84 149
rect 114 183 170 222
rect 114 149 125 183
rect 159 149 170 183
rect 114 112 170 149
rect 200 112 288 222
rect 215 74 288 112
rect 318 210 375 222
rect 318 176 329 210
rect 363 176 375 210
rect 318 74 375 176
rect 429 130 536 184
rect 429 96 441 130
rect 475 96 536 130
rect 429 74 536 96
rect 566 169 622 184
rect 566 135 577 169
rect 611 164 622 169
rect 795 164 845 222
rect 611 135 637 164
rect 566 80 637 135
rect 667 80 709 164
rect 739 126 845 164
rect 739 92 750 126
rect 784 92 845 126
rect 739 80 845 92
rect 566 74 616 80
rect 215 40 227 74
rect 261 40 273 74
rect 795 74 845 80
rect 875 181 931 222
rect 875 147 886 181
rect 920 147 931 181
rect 875 74 931 147
rect 985 210 1041 222
rect 985 176 996 210
rect 1030 176 1041 210
rect 985 120 1041 176
rect 985 86 996 120
rect 1030 86 1041 120
rect 985 74 1041 86
rect 1071 210 1136 222
rect 1071 176 1082 210
rect 1116 176 1136 210
rect 1071 140 1136 176
rect 1071 106 1082 140
rect 1116 106 1136 140
rect 1071 94 1136 106
rect 1166 94 1208 222
rect 1238 208 1295 222
rect 1238 174 1249 208
rect 1283 174 1295 208
rect 1238 140 1295 174
rect 1238 106 1249 140
rect 1283 106 1295 140
rect 1238 94 1295 106
rect 1351 210 1423 222
rect 1351 176 1363 210
rect 1397 176 1423 210
rect 1351 120 1423 176
rect 1071 74 1121 94
rect 1351 86 1363 120
rect 1397 86 1423 120
rect 1351 74 1423 86
rect 1453 210 1509 222
rect 1453 176 1464 210
rect 1498 176 1509 210
rect 1453 120 1509 176
rect 1453 86 1464 120
rect 1498 86 1509 120
rect 1453 74 1509 86
rect 215 28 273 40
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 476 86 546
rect 27 442 39 476
rect 73 442 86 476
rect 27 424 86 442
rect 116 424 164 592
rect 194 580 253 592
rect 194 546 207 580
rect 241 546 253 580
rect 194 498 253 546
rect 194 464 207 498
rect 241 464 253 498
rect 194 424 253 464
rect 307 582 365 594
rect 307 548 319 582
rect 353 548 365 582
rect 1121 617 1194 629
rect 307 536 365 548
rect 639 547 692 576
rect 307 368 383 536
rect 413 414 472 536
rect 413 380 426 414
rect 460 380 472 414
rect 413 368 472 380
rect 526 535 585 547
rect 526 501 538 535
rect 572 501 585 535
rect 526 427 585 501
rect 526 393 538 427
rect 572 393 585 427
rect 526 379 585 393
rect 615 535 692 547
rect 615 501 628 535
rect 662 501 692 535
rect 615 492 692 501
rect 722 492 770 576
rect 800 551 871 576
rect 800 517 813 551
rect 847 517 871 551
rect 800 492 871 517
rect 615 427 674 492
rect 615 393 628 427
rect 662 393 674 427
rect 615 379 674 393
rect 818 352 871 492
rect 901 564 960 576
rect 1121 583 1140 617
rect 1174 583 1194 617
rect 1121 571 1194 583
rect 1350 571 1403 592
rect 901 530 914 564
rect 948 530 960 564
rect 901 481 960 530
rect 901 447 914 481
rect 948 447 960 481
rect 901 398 960 447
rect 1014 449 1073 571
rect 1014 415 1026 449
rect 1060 415 1073 449
rect 1014 403 1073 415
rect 1103 403 1212 571
rect 1242 559 1302 571
rect 1242 525 1255 559
rect 1289 525 1302 559
rect 1242 449 1302 525
rect 1242 415 1255 449
rect 1289 415 1302 449
rect 1242 403 1302 415
rect 1332 559 1403 571
rect 1332 525 1355 559
rect 1389 525 1403 559
rect 1332 462 1403 525
rect 1332 428 1355 462
rect 1389 428 1403 462
rect 1332 403 1403 428
rect 901 364 914 398
rect 948 364 960 398
rect 901 352 960 364
rect 1350 368 1403 403
rect 1433 580 1509 592
rect 1433 546 1463 580
rect 1497 546 1509 580
rect 1433 497 1509 546
rect 1433 463 1463 497
rect 1497 463 1509 497
rect 1433 414 1509 463
rect 1433 380 1463 414
rect 1497 380 1509 414
rect 1433 368 1509 380
<< ndiffc >>
rect 39 149 73 183
rect 125 149 159 183
rect 329 176 363 210
rect 441 96 475 130
rect 577 135 611 169
rect 750 92 784 126
rect 227 40 261 74
rect 886 147 920 181
rect 996 176 1030 210
rect 996 86 1030 120
rect 1082 176 1116 210
rect 1082 106 1116 140
rect 1249 174 1283 208
rect 1249 106 1283 140
rect 1363 176 1397 210
rect 1363 86 1397 120
rect 1464 176 1498 210
rect 1464 86 1498 120
<< pdiffc >>
rect 39 546 73 580
rect 39 442 73 476
rect 207 546 241 580
rect 207 464 241 498
rect 319 548 353 582
rect 426 380 460 414
rect 538 501 572 535
rect 538 393 572 427
rect 628 501 662 535
rect 813 517 847 551
rect 628 393 662 427
rect 1140 583 1174 617
rect 914 530 948 564
rect 914 447 948 481
rect 1026 415 1060 449
rect 1255 525 1289 559
rect 1255 415 1289 449
rect 1355 525 1389 559
rect 1355 428 1389 462
rect 914 364 948 398
rect 1463 546 1497 580
rect 1463 463 1497 497
rect 1463 380 1497 414
<< poly >>
rect 86 592 116 618
rect 164 592 194 618
rect 380 615 725 645
rect 380 551 416 615
rect 689 591 725 615
rect 692 576 722 591
rect 770 576 800 602
rect 871 576 901 602
rect 383 536 413 551
rect 585 547 615 573
rect 86 409 116 424
rect 164 409 194 424
rect 83 392 119 409
rect 44 376 119 392
rect 44 342 60 376
rect 94 342 119 376
rect 44 308 119 342
rect 161 392 197 409
rect 161 376 227 392
rect 161 342 177 376
rect 211 342 227 376
rect 692 466 722 492
rect 770 477 800 492
rect 767 424 803 477
rect 709 408 803 424
rect 383 353 413 368
rect 585 364 615 379
rect 709 374 736 408
rect 770 374 803 408
rect 161 326 227 342
rect 44 274 60 308
rect 94 274 119 308
rect 44 258 119 274
rect 84 222 114 258
rect 170 222 200 326
rect 380 272 416 353
rect 582 343 618 364
rect 709 358 803 374
rect 525 327 667 343
rect 525 293 541 327
rect 575 293 667 327
rect 525 277 667 293
rect 288 256 483 272
rect 288 242 433 256
rect 288 222 318 242
rect 417 222 433 242
rect 467 229 483 256
rect 467 222 566 229
rect 84 86 114 112
rect 170 86 200 112
rect 417 199 566 222
rect 536 184 566 199
rect 637 164 667 277
rect 709 164 739 358
rect 1073 571 1103 597
rect 1212 571 1242 597
rect 1302 571 1332 597
rect 1403 592 1433 618
rect 1073 388 1103 403
rect 1212 388 1242 403
rect 1302 388 1332 403
rect 1070 358 1245 388
rect 871 337 901 352
rect 1070 337 1166 358
rect 868 310 904 337
rect 798 294 904 310
rect 798 260 814 294
rect 848 260 904 294
rect 798 244 904 260
rect 1041 321 1166 337
rect 1041 287 1082 321
rect 1116 287 1166 321
rect 1299 310 1335 388
rect 1403 353 1433 368
rect 1400 345 1436 353
rect 1041 271 1166 287
rect 845 222 875 244
rect 1041 222 1071 271
rect 1136 222 1166 271
rect 1208 294 1335 310
rect 1208 260 1224 294
rect 1258 280 1335 294
rect 1383 310 1453 345
rect 1258 260 1329 280
rect 1208 244 1329 260
rect 1383 276 1399 310
rect 1433 276 1453 310
rect 1208 222 1238 244
rect 1383 237 1453 276
rect 1423 222 1453 237
rect 288 48 318 74
rect 536 48 566 74
rect 637 54 667 80
rect 709 54 739 80
rect 845 48 875 74
rect 1041 48 1071 74
rect 1136 68 1166 94
rect 1208 68 1238 94
rect 1423 48 1453 74
<< polycont >>
rect 60 342 94 376
rect 177 342 211 376
rect 736 374 770 408
rect 60 274 94 308
rect 541 293 575 327
rect 433 222 467 256
rect 814 260 848 294
rect 1082 287 1116 321
rect 1224 260 1258 294
rect 1399 276 1433 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 23 580 89 649
rect 23 546 39 580
rect 73 546 89 580
rect 23 476 89 546
rect 23 442 39 476
rect 73 442 89 476
rect 191 580 257 596
rect 191 546 207 580
rect 241 546 257 580
rect 191 498 257 546
rect 303 582 369 649
rect 303 548 319 582
rect 353 548 369 582
rect 797 551 863 649
rect 1117 617 1198 649
rect 1117 583 1140 617
rect 1174 583 1198 617
rect 303 532 369 548
rect 522 535 572 551
rect 522 501 538 535
rect 522 498 572 501
rect 191 464 207 498
rect 241 464 572 498
rect 612 535 678 551
rect 612 501 628 535
rect 662 501 678 535
rect 612 485 678 501
rect 797 517 813 551
rect 847 517 863 551
rect 797 488 863 517
rect 898 564 964 580
rect 1117 567 1198 583
rect 898 530 914 564
rect 948 533 964 564
rect 1239 559 1305 575
rect 948 530 1200 533
rect 898 499 1200 530
rect 23 426 89 442
rect 25 376 109 392
rect 25 342 60 376
rect 94 342 109 376
rect 25 308 109 342
rect 161 376 257 430
rect 161 342 177 376
rect 211 342 257 376
rect 161 326 257 342
rect 25 274 60 308
rect 94 274 109 308
rect 291 292 325 464
rect 25 258 109 274
rect 143 258 325 292
rect 359 414 476 430
rect 359 380 426 414
rect 460 380 476 414
rect 359 343 476 380
rect 522 427 572 464
rect 522 393 538 427
rect 522 377 572 393
rect 614 427 678 485
rect 614 393 628 427
rect 662 393 678 427
rect 898 481 964 499
rect 898 447 914 481
rect 948 447 964 481
rect 898 424 964 447
rect 359 327 580 343
rect 359 309 541 327
rect 143 224 177 258
rect 359 224 393 309
rect 525 293 541 309
rect 575 293 580 327
rect 525 277 580 293
rect 614 310 678 393
rect 720 408 964 424
rect 720 374 736 408
rect 770 398 964 408
rect 770 374 914 398
rect 720 364 914 374
rect 948 364 964 398
rect 720 348 964 364
rect 998 449 1076 465
rect 998 415 1026 449
rect 1060 415 1076 449
rect 998 399 1076 415
rect 614 294 864 310
rect 23 183 73 224
rect 23 149 39 183
rect 23 17 73 149
rect 109 183 177 224
rect 109 149 125 183
rect 159 149 177 183
rect 313 210 393 224
rect 313 176 329 210
rect 363 190 393 210
rect 427 256 483 272
rect 427 222 433 256
rect 467 240 483 256
rect 614 260 814 294
rect 848 260 864 294
rect 614 244 864 260
rect 467 222 543 240
rect 427 206 543 222
rect 363 176 379 190
rect 109 142 177 149
rect 425 142 475 156
rect 109 130 475 142
rect 109 108 441 130
rect 425 96 441 108
rect 211 40 227 74
rect 261 40 277 74
rect 425 70 475 96
rect 509 85 543 206
rect 614 185 648 244
rect 898 210 936 348
rect 998 226 1032 399
rect 1066 321 1132 356
rect 1066 287 1082 321
rect 1116 287 1132 321
rect 1066 271 1132 287
rect 1166 310 1200 499
rect 1239 525 1255 559
rect 1289 525 1305 559
rect 1239 449 1305 525
rect 1239 415 1255 449
rect 1289 415 1305 449
rect 1239 378 1305 415
rect 1339 559 1405 649
rect 1339 525 1355 559
rect 1389 525 1405 559
rect 1339 462 1405 525
rect 1339 428 1355 462
rect 1389 428 1405 462
rect 1339 412 1405 428
rect 1447 580 1517 596
rect 1447 546 1463 580
rect 1497 546 1517 580
rect 1447 497 1517 546
rect 1447 463 1463 497
rect 1497 463 1517 497
rect 1447 414 1517 463
rect 1447 380 1463 414
rect 1497 380 1517 414
rect 1239 344 1329 378
rect 1447 364 1517 380
rect 1295 326 1329 344
rect 1295 310 1449 326
rect 1166 294 1261 310
rect 1166 260 1224 294
rect 1258 260 1261 294
rect 1166 244 1261 260
rect 1295 276 1399 310
rect 1433 276 1449 310
rect 1295 260 1449 276
rect 577 169 648 185
rect 611 135 648 169
rect 577 119 648 135
rect 682 176 852 210
rect 682 85 716 176
rect 509 51 716 85
rect 750 126 784 142
rect 211 17 277 40
rect 750 17 784 92
rect 818 85 852 176
rect 886 181 936 210
rect 920 147 936 181
rect 886 119 936 147
rect 980 210 1046 226
rect 980 176 996 210
rect 1030 176 1046 210
rect 980 120 1046 176
rect 980 86 996 120
rect 1030 86 1046 120
rect 980 85 1046 86
rect 818 51 1046 85
rect 1082 210 1132 226
rect 1295 210 1329 260
rect 1483 226 1517 364
rect 1116 176 1132 210
rect 1082 140 1132 176
rect 1116 106 1132 140
rect 1082 17 1132 106
rect 1233 208 1329 210
rect 1233 174 1249 208
rect 1283 174 1329 208
rect 1233 140 1329 174
rect 1233 106 1249 140
rect 1283 106 1329 140
rect 1233 90 1329 106
rect 1363 210 1413 226
rect 1397 176 1413 210
rect 1363 120 1413 176
rect 1397 86 1413 120
rect 1363 17 1413 86
rect 1448 210 1517 226
rect 1448 176 1464 210
rect 1498 176 1517 210
rect 1448 120 1517 176
rect 1448 86 1464 120
rect 1498 86 1517 120
rect 1448 70 1517 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
rlabel comment s 0 0 0 0 4 sdlclkp_1
flabel pwell s 0 0 1536 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 0 617 1536 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 1536 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 1536 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 1471 390 1505 424 0 FreeSans 340 0 0 0 GCLK
port 8 nsew
flabel corelocali s 1471 464 1505 498 0 FreeSans 340 0 0 0 GCLK
port 8 nsew
flabel corelocali s 1471 538 1505 572 0 FreeSans 340 0 0 0 GCLK
port 8 nsew
flabel corelocali s 1087 316 1121 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 223 390 257 424 0 FreeSans 340 0 0 0 GATE
port 2 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 SCE
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 1536 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 267868
string GDS_START 256092
<< end >>
