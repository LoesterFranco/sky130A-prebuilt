magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 1190 704
<< pwell >>
rect 0 0 1152 49
<< scnmos >>
rect 92 74 122 222
rect 178 74 208 222
rect 434 74 464 222
rect 520 74 550 222
rect 606 74 636 222
rect 692 74 722 222
rect 778 74 808 222
rect 864 74 894 222
rect 950 74 980 222
rect 1040 74 1070 222
<< pmoshvt >>
rect 86 368 116 592
rect 181 368 211 592
rect 407 368 437 592
rect 497 368 527 592
rect 587 368 617 592
rect 677 368 707 592
rect 767 368 797 592
rect 857 368 887 592
rect 947 368 977 592
rect 1037 368 1067 592
<< ndiff >>
rect 35 210 92 222
rect 35 176 47 210
rect 81 176 92 210
rect 35 120 92 176
rect 35 86 47 120
rect 81 86 92 120
rect 35 74 92 86
rect 122 196 178 222
rect 122 162 133 196
rect 167 162 178 196
rect 122 116 178 162
rect 122 82 133 116
rect 167 82 178 116
rect 122 74 178 82
rect 208 186 265 222
rect 208 152 219 186
rect 253 152 265 186
rect 208 118 265 152
rect 208 84 219 118
rect 253 84 265 118
rect 208 74 265 84
rect 378 210 434 222
rect 378 176 389 210
rect 423 176 434 210
rect 378 120 434 176
rect 378 86 389 120
rect 423 86 434 120
rect 378 74 434 86
rect 464 188 520 222
rect 464 154 475 188
rect 509 154 520 188
rect 464 120 520 154
rect 464 86 475 120
rect 509 86 520 120
rect 464 74 520 86
rect 550 210 606 222
rect 550 176 561 210
rect 595 176 606 210
rect 550 120 606 176
rect 550 86 561 120
rect 595 86 606 120
rect 550 74 606 86
rect 636 146 692 222
rect 636 112 647 146
rect 681 112 692 146
rect 636 74 692 112
rect 722 210 778 222
rect 722 176 733 210
rect 767 176 778 210
rect 722 120 778 176
rect 722 86 733 120
rect 767 86 778 120
rect 722 74 778 86
rect 808 181 864 222
rect 808 147 819 181
rect 853 147 864 181
rect 808 74 864 147
rect 894 133 950 222
rect 894 99 905 133
rect 939 99 950 133
rect 894 74 950 99
rect 980 189 1040 222
rect 980 155 991 189
rect 1025 155 1040 189
rect 980 74 1040 155
rect 1070 210 1125 222
rect 1070 176 1081 210
rect 1115 176 1125 210
rect 1070 120 1125 176
rect 1070 86 1081 120
rect 1115 86 1125 120
rect 1070 74 1125 86
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 510 86 546
rect 27 476 39 510
rect 73 476 86 510
rect 27 440 86 476
rect 27 406 39 440
rect 73 406 86 440
rect 27 368 86 406
rect 116 580 181 592
rect 116 546 131 580
rect 165 546 181 580
rect 116 368 181 546
rect 211 421 270 592
rect 211 387 224 421
rect 258 387 270 421
rect 211 368 270 387
rect 348 530 407 592
rect 348 496 360 530
rect 394 496 407 530
rect 348 368 407 496
rect 437 582 497 592
rect 437 548 450 582
rect 484 548 497 582
rect 437 368 497 548
rect 527 580 587 592
rect 527 546 540 580
rect 574 546 587 580
rect 527 497 587 546
rect 527 463 540 497
rect 574 463 587 497
rect 527 414 587 463
rect 527 380 540 414
rect 574 380 587 414
rect 527 368 587 380
rect 617 580 677 592
rect 617 546 630 580
rect 664 546 677 580
rect 617 482 677 546
rect 617 448 630 482
rect 664 448 677 482
rect 617 368 677 448
rect 707 580 767 592
rect 707 546 720 580
rect 754 546 767 580
rect 707 497 767 546
rect 707 463 720 497
rect 754 463 767 497
rect 707 414 767 463
rect 707 380 720 414
rect 754 380 767 414
rect 707 368 767 380
rect 797 547 857 592
rect 797 513 810 547
rect 844 513 857 547
rect 797 479 857 513
rect 797 445 810 479
rect 844 445 857 479
rect 797 411 857 445
rect 797 377 810 411
rect 844 377 857 411
rect 797 368 857 377
rect 887 580 947 592
rect 887 546 900 580
rect 934 546 947 580
rect 887 482 947 546
rect 887 448 900 482
rect 934 448 947 482
rect 887 368 947 448
rect 977 547 1037 592
rect 977 513 990 547
rect 1024 513 1037 547
rect 977 479 1037 513
rect 977 445 990 479
rect 1024 445 1037 479
rect 977 411 1037 445
rect 977 377 990 411
rect 1024 377 1037 411
rect 977 368 1037 377
rect 1067 580 1125 592
rect 1067 546 1080 580
rect 1114 546 1125 580
rect 1067 497 1125 546
rect 1067 463 1080 497
rect 1114 463 1125 497
rect 1067 414 1125 463
rect 1067 380 1080 414
rect 1114 380 1125 414
rect 1067 368 1125 380
<< ndiffc >>
rect 47 176 81 210
rect 47 86 81 120
rect 133 162 167 196
rect 133 82 167 116
rect 219 152 253 186
rect 219 84 253 118
rect 389 176 423 210
rect 389 86 423 120
rect 475 154 509 188
rect 475 86 509 120
rect 561 176 595 210
rect 561 86 595 120
rect 647 112 681 146
rect 733 176 767 210
rect 733 86 767 120
rect 819 147 853 181
rect 905 99 939 133
rect 991 155 1025 189
rect 1081 176 1115 210
rect 1081 86 1115 120
<< pdiffc >>
rect 39 546 73 580
rect 39 476 73 510
rect 39 406 73 440
rect 131 546 165 580
rect 224 387 258 421
rect 360 496 394 530
rect 450 548 484 582
rect 540 546 574 580
rect 540 463 574 497
rect 540 380 574 414
rect 630 546 664 580
rect 630 448 664 482
rect 720 546 754 580
rect 720 463 754 497
rect 720 380 754 414
rect 810 513 844 547
rect 810 445 844 479
rect 810 377 844 411
rect 900 546 934 580
rect 900 448 934 482
rect 990 513 1024 547
rect 990 445 1024 479
rect 990 377 1024 411
rect 1080 546 1114 580
rect 1080 463 1114 497
rect 1080 380 1114 414
<< poly >>
rect 86 592 116 618
rect 181 592 211 618
rect 407 592 437 618
rect 497 592 527 618
rect 587 592 617 618
rect 677 592 707 618
rect 767 592 797 618
rect 857 592 887 618
rect 947 592 977 618
rect 1037 592 1067 618
rect 86 353 116 368
rect 181 353 211 368
rect 407 353 437 368
rect 497 353 527 368
rect 587 353 617 368
rect 677 353 707 368
rect 767 353 797 368
rect 857 353 887 368
rect 947 353 977 368
rect 1037 353 1067 368
rect 83 326 119 353
rect 178 345 214 353
rect 404 345 440 353
rect 494 345 530 353
rect 584 345 620 353
rect 674 345 710 353
rect 70 310 136 326
rect 70 276 86 310
rect 120 276 136 310
rect 70 260 136 276
rect 178 315 710 345
rect 764 330 800 353
rect 854 330 890 353
rect 944 330 980 353
rect 1034 330 1070 353
rect 178 294 248 315
rect 178 260 198 294
rect 232 260 248 294
rect 764 314 1070 330
rect 764 280 780 314
rect 814 280 848 314
rect 882 280 916 314
rect 950 280 1070 314
rect 92 222 122 260
rect 178 244 248 260
rect 290 246 722 267
rect 764 264 1070 280
rect 178 222 208 244
rect 290 212 306 246
rect 340 237 722 246
rect 340 212 356 237
rect 434 222 464 237
rect 520 222 550 237
rect 606 222 636 237
rect 692 222 722 237
rect 778 222 808 264
rect 864 222 894 264
rect 950 222 980 264
rect 1040 222 1070 264
rect 290 178 356 212
rect 290 144 306 178
rect 340 144 356 178
rect 290 110 356 144
rect 290 76 306 110
rect 340 76 356 110
rect 92 48 122 74
rect 178 48 208 74
rect 290 60 356 76
rect 434 48 464 74
rect 520 48 550 74
rect 606 48 636 74
rect 692 48 722 74
rect 778 48 808 74
rect 864 48 894 74
rect 950 48 980 74
rect 1040 48 1070 74
<< polycont >>
rect 86 276 120 310
rect 198 260 232 294
rect 780 280 814 314
rect 848 280 882 314
rect 916 280 950 314
rect 306 212 340 246
rect 306 144 340 178
rect 306 76 340 110
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 17 580 73 596
rect 17 546 39 580
rect 113 580 184 649
rect 113 546 131 580
rect 165 546 184 580
rect 434 582 500 649
rect 17 512 73 546
rect 360 530 394 564
rect 434 548 450 582
rect 484 548 500 582
rect 540 580 574 596
rect 17 510 326 512
rect 17 476 39 510
rect 73 478 326 510
rect 540 514 574 546
rect 394 497 574 514
rect 394 496 540 497
rect 360 480 540 496
rect 17 440 73 476
rect 292 446 326 478
rect 17 406 39 440
rect 17 390 73 406
rect 208 421 258 444
rect 17 226 51 390
rect 208 387 224 421
rect 292 412 506 446
rect 208 378 258 387
rect 85 310 161 356
rect 208 344 355 378
rect 85 276 86 310
rect 120 276 161 310
rect 85 260 161 276
rect 195 294 257 310
rect 195 260 198 294
rect 232 260 257 294
rect 195 236 257 260
rect 291 246 355 344
rect 472 330 506 412
rect 540 414 574 463
rect 614 580 664 649
rect 614 546 630 580
rect 614 482 664 546
rect 614 448 630 482
rect 614 432 664 448
rect 704 581 1130 615
rect 704 580 754 581
rect 704 546 720 580
rect 894 580 940 581
rect 704 497 754 546
rect 704 463 720 497
rect 704 414 754 463
rect 704 398 720 414
rect 574 380 720 398
rect 540 364 754 380
rect 794 513 810 547
rect 844 513 860 547
rect 794 479 860 513
rect 794 445 810 479
rect 844 445 860 479
rect 794 411 860 445
rect 894 546 900 580
rect 934 546 940 580
rect 1080 580 1130 581
rect 894 482 940 546
rect 894 448 900 482
rect 934 448 940 482
rect 894 432 940 448
rect 974 513 990 547
rect 1024 513 1041 547
rect 974 479 1041 513
rect 974 445 990 479
rect 1024 445 1041 479
rect 794 377 810 411
rect 844 398 860 411
rect 974 411 1041 445
rect 974 398 990 411
rect 844 377 990 398
rect 1024 377 1041 411
rect 794 364 1041 377
rect 1114 546 1130 580
rect 1080 497 1130 546
rect 1114 463 1130 497
rect 1080 414 1130 463
rect 1114 380 1130 414
rect 1080 364 1130 380
rect 472 314 966 330
rect 472 296 780 314
rect 764 280 780 296
rect 814 280 848 314
rect 882 280 916 314
rect 950 280 966 314
rect 764 264 966 280
rect 17 210 81 226
rect 17 176 47 210
rect 291 212 306 246
rect 340 212 355 246
rect 291 202 355 212
rect 17 120 81 176
rect 17 86 47 120
rect 17 70 81 86
rect 117 196 183 202
rect 117 162 133 196
rect 167 162 183 196
rect 117 116 183 162
rect 117 82 133 116
rect 167 82 183 116
rect 117 17 183 82
rect 219 186 355 202
rect 253 178 355 186
rect 253 152 306 178
rect 219 144 306 152
rect 340 144 355 178
rect 219 118 355 144
rect 253 110 355 118
rect 253 84 306 110
rect 219 76 306 84
rect 340 76 355 110
rect 219 60 355 76
rect 389 230 595 262
rect 1007 230 1041 364
rect 389 228 767 230
rect 389 210 423 228
rect 561 210 767 228
rect 389 120 423 176
rect 389 70 423 86
rect 459 188 525 194
rect 459 154 475 188
rect 509 154 525 188
rect 459 120 525 154
rect 459 86 475 120
rect 509 86 525 120
rect 459 17 525 86
rect 595 196 733 210
rect 561 120 595 176
rect 717 176 733 196
rect 561 70 595 86
rect 631 146 681 162
rect 631 112 647 146
rect 631 17 681 112
rect 717 120 767 176
rect 717 86 733 120
rect 803 196 1041 230
rect 803 181 869 196
rect 803 147 819 181
rect 853 147 869 181
rect 975 189 1041 196
rect 803 119 869 147
rect 905 133 939 162
rect 717 85 767 86
rect 975 155 991 189
rect 1025 155 1041 189
rect 975 119 1041 155
rect 1081 210 1131 226
rect 1115 176 1131 210
rect 1081 120 1131 176
rect 905 85 939 99
rect 1115 86 1131 120
rect 1081 85 1131 86
rect 717 51 1131 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
rlabel comment s 0 0 0 0 4 ebufn_4
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 991 390 1025 424 0 FreeSans 340 0 0 0 Z
port 7 nsew
flabel corelocali s 991 464 1025 498 0 FreeSans 340 0 0 0 Z
port 7 nsew
flabel corelocali s 223 242 257 276 0 FreeSans 340 0 0 0 TE_B
port 2 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 1152 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2060340
string GDS_START 2050860
<< end >>
