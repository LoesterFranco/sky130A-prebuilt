magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 79 47 109 177
rect 173 47 203 177
rect 280 47 310 131
rect 376 47 406 131
rect 472 47 502 131
rect 650 47 680 131
rect 754 47 784 131
<< pmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 282 369 318 497
rect 474 369 510 497
rect 570 369 606 497
rect 652 369 688 497
rect 746 369 782 497
<< ndiff >>
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 101 173 177
rect 109 67 126 101
rect 160 67 173 101
rect 109 47 173 67
rect 203 131 263 177
rect 203 93 280 131
rect 203 59 223 93
rect 257 59 280 93
rect 203 47 280 59
rect 310 47 376 131
rect 406 103 472 131
rect 406 69 416 103
rect 450 69 472 103
rect 406 47 472 69
rect 502 47 650 131
rect 680 101 754 131
rect 680 67 700 101
rect 734 67 754 101
rect 680 47 754 67
rect 784 101 839 131
rect 784 67 797 101
rect 831 67 839 101
rect 784 47 839 67
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 477 175 497
rect 117 443 129 477
rect 163 443 175 477
rect 117 409 175 443
rect 117 375 129 409
rect 163 375 175 409
rect 117 297 175 375
rect 211 485 282 497
rect 211 451 223 485
rect 257 451 282 485
rect 211 369 282 451
rect 318 369 474 497
rect 510 485 570 497
rect 510 451 522 485
rect 556 451 570 485
rect 510 369 570 451
rect 606 369 652 497
rect 688 485 746 497
rect 688 451 700 485
rect 734 451 746 485
rect 688 369 746 451
rect 782 485 838 497
rect 782 451 796 485
rect 830 451 838 485
rect 782 417 838 451
rect 782 383 796 417
rect 830 383 838 417
rect 782 369 838 383
rect 211 297 263 369
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 126 67 160 101
rect 223 59 257 93
rect 416 69 450 103
rect 700 67 734 101
rect 797 67 831 101
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 443 163 477
rect 129 375 163 409
rect 223 451 257 485
rect 522 451 556 485
rect 700 451 734 485
rect 796 451 830 485
rect 796 383 830 417
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 282 497 318 523
rect 474 497 510 523
rect 570 497 606 523
rect 652 497 688 523
rect 746 497 782 523
rect 282 354 318 369
rect 474 354 510 369
rect 570 354 606 369
rect 652 354 688 369
rect 746 354 782 369
rect 81 282 117 297
rect 175 282 211 297
rect 79 265 119 282
rect 173 265 213 282
rect 280 265 320 354
rect 79 249 238 265
rect 79 215 194 249
rect 228 215 238 249
rect 79 199 238 215
rect 280 249 334 265
rect 280 215 290 249
rect 324 215 334 249
rect 280 199 334 215
rect 376 203 430 219
rect 79 177 109 199
rect 173 177 203 199
rect 280 131 310 199
rect 376 169 386 203
rect 420 169 430 203
rect 376 153 430 169
rect 472 215 512 354
rect 568 323 608 354
rect 554 307 608 323
rect 554 273 564 307
rect 598 273 608 307
rect 554 257 608 273
rect 650 265 690 354
rect 744 265 784 354
rect 650 249 784 265
rect 650 215 673 249
rect 707 215 784 249
rect 472 205 556 215
rect 472 171 506 205
rect 540 171 556 205
rect 472 161 556 171
rect 650 199 784 215
rect 376 131 406 153
rect 472 131 502 161
rect 650 131 680 199
rect 754 131 784 199
rect 79 21 109 47
rect 173 21 203 47
rect 280 21 310 47
rect 376 21 406 47
rect 472 21 502 47
rect 650 21 680 47
rect 754 21 784 47
<< polycont >>
rect 194 215 228 249
rect 290 215 324 249
rect 386 169 420 203
rect 564 273 598 307
rect 673 215 707 249
rect 506 171 540 205
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 18 485 69 527
rect 18 451 35 485
rect 18 417 69 451
rect 18 383 35 417
rect 18 349 69 383
rect 18 315 35 349
rect 18 299 69 315
rect 103 477 175 493
rect 103 443 129 477
rect 163 443 175 477
rect 103 409 175 443
rect 223 485 257 527
rect 692 485 736 527
rect 223 435 257 451
rect 291 451 522 485
rect 556 451 572 485
rect 692 451 700 485
rect 734 451 736 485
rect 103 375 129 409
rect 163 375 175 409
rect 291 401 325 451
rect 692 435 736 451
rect 770 485 847 493
rect 770 451 796 485
rect 830 451 847 485
rect 770 417 847 451
rect 770 401 796 417
rect 103 319 175 375
rect 219 367 325 401
rect 359 383 796 401
rect 830 383 847 417
rect 359 367 847 383
rect 18 161 69 177
rect 18 127 35 161
rect 18 93 69 127
rect 18 59 35 93
rect 18 17 69 59
rect 103 101 160 319
rect 219 265 253 367
rect 359 333 393 367
rect 194 249 253 265
rect 228 215 253 249
rect 194 199 253 215
rect 287 299 393 333
rect 427 307 615 325
rect 287 249 331 299
rect 427 282 564 307
rect 425 273 564 282
rect 598 273 615 307
rect 425 265 615 273
rect 287 215 290 249
rect 324 215 331 249
rect 287 199 331 215
rect 384 256 615 265
rect 384 203 459 256
rect 671 249 709 325
rect 219 161 253 199
rect 384 169 386 203
rect 420 169 459 203
rect 219 127 341 161
rect 384 153 459 169
rect 506 205 615 221
rect 540 171 615 205
rect 506 155 615 171
rect 103 67 126 101
rect 307 119 341 127
rect 307 103 450 119
rect 103 51 160 67
rect 197 59 223 93
rect 257 59 273 93
rect 197 17 273 59
rect 307 69 416 103
rect 574 84 615 155
rect 671 215 673 249
rect 707 215 709 249
rect 671 151 709 215
rect 697 101 737 117
rect 307 53 450 69
rect 697 67 700 101
rect 734 67 737 101
rect 697 17 737 67
rect 797 101 847 367
rect 831 67 847 101
rect 797 51 847 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
flabel corelocali s 581 153 615 187 0 FreeSans 200 0 0 0 A1
port 2 nsew
flabel corelocali s 489 289 523 323 0 FreeSans 200 0 0 0 A0
port 1 nsew
flabel corelocali s 397 221 431 255 0 FreeSans 200 0 0 0 A0
port 1 nsew
flabel corelocali s 397 153 431 187 0 FreeSans 200 0 0 0 A0
port 1 nsew
flabel corelocali s 673 153 707 187 0 FreeSans 200 0 0 0 S
port 3 nsew
flabel corelocali s 581 85 615 119 0 FreeSans 200 0 0 0 A1
port 2 nsew
flabel corelocali s 121 425 155 459 0 FreeSans 200 0 0 0 X
port 8 nsew
flabel corelocali s 121 357 155 391 0 FreeSans 200 0 0 0 X
port 8 nsew
flabel corelocali s 581 289 615 323 0 FreeSans 200 0 0 0 A0
port 1 nsew
flabel corelocali s 673 289 707 323 0 FreeSans 200 0 0 0 S
port 3 nsew
flabel corelocali s 673 221 707 255 0 FreeSans 200 0 0 0 S
port 3 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
rlabel comment s 0 0 0 0 4 mux2_2
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2136170
string GDS_START 2128756
<< end >>
