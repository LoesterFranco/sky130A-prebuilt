magic
tech sky130A
magscale 1 2
timestamp 1599588232
<< locali >>
rect 121 332 359 376
rect 121 298 545 332
rect 313 162 420 262
rect 479 252 545 298
rect 587 288 653 430
rect 757 236 929 326
rect 757 184 812 236
rect 2403 70 2469 596
rect 2711 364 2767 596
rect 2733 226 2767 364
rect 2694 70 2767 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 23 444 211 595
rect 245 478 311 649
rect 419 520 511 596
rect 619 546 685 649
rect 733 524 799 596
rect 941 550 1007 649
rect 733 520 916 524
rect 419 512 589 520
rect 733 518 922 520
rect 733 517 926 518
rect 733 516 929 517
rect 1165 516 1215 545
rect 733 512 1215 516
rect 419 484 1215 512
rect 419 480 850 484
rect 911 483 1215 484
rect 914 482 1215 483
rect 918 480 1215 482
rect 419 478 846 480
rect 689 477 846 478
rect 923 477 1215 480
rect 1250 477 1371 545
rect 689 466 757 477
rect 23 410 539 444
rect 23 262 57 410
rect 473 366 539 410
rect 23 196 279 262
rect 23 70 73 196
rect 689 218 723 466
rect 867 439 901 450
rect 1165 443 1215 477
rect 784 432 833 438
rect 757 424 833 432
rect 757 390 799 424
rect 757 366 833 390
rect 867 360 997 439
rect 1031 391 1126 443
rect 1165 409 1303 443
rect 963 355 997 360
rect 1090 375 1126 391
rect 454 184 723 218
rect 963 291 1056 355
rect 1090 309 1235 375
rect 963 202 1009 291
rect 1090 257 1126 309
rect 1269 274 1303 409
rect 109 17 175 162
rect 221 85 271 162
rect 454 119 520 184
rect 846 168 1009 202
rect 1043 214 1126 257
rect 1160 240 1303 274
rect 1337 433 1371 477
rect 1405 469 1453 649
rect 1487 464 1553 549
rect 1487 433 1521 464
rect 1337 397 1521 433
rect 846 150 907 168
rect 612 85 682 150
rect 221 51 682 85
rect 718 17 776 150
rect 827 100 907 150
rect 941 17 1007 134
rect 1043 85 1124 214
rect 1160 199 1195 240
rect 1337 206 1371 397
rect 1159 119 1195 199
rect 1229 172 1371 206
rect 1405 218 1453 361
rect 1487 309 1521 397
rect 1555 424 1607 430
rect 1555 390 1567 424
rect 1601 390 1607 424
rect 1555 359 1607 390
rect 1647 343 1697 649
rect 1487 252 1663 309
rect 1737 283 1787 551
rect 1821 485 2019 551
rect 2061 532 2130 649
rect 2171 498 2237 577
rect 2274 539 2363 649
rect 1821 351 1865 485
rect 1901 315 1951 446
rect 1697 249 1787 283
rect 1821 269 1951 315
rect 1985 287 2019 485
rect 2053 464 2281 498
rect 2053 330 2105 464
rect 2139 424 2213 430
rect 2139 390 2143 424
rect 2177 390 2213 424
rect 2139 337 2213 390
rect 2247 360 2281 464
rect 2317 394 2363 539
rect 2247 326 2369 360
rect 1697 218 1731 249
rect 1405 184 1731 218
rect 1821 215 1887 269
rect 1985 235 2285 287
rect 1229 119 1294 172
rect 1410 116 1620 150
rect 1654 119 1731 184
rect 1765 181 1887 215
rect 1921 201 2285 235
rect 1410 85 1444 116
rect 1043 51 1444 85
rect 1586 85 1620 116
rect 1765 85 1799 181
rect 1921 147 1955 201
rect 1486 17 1552 82
rect 1586 51 1799 85
rect 1833 81 1955 147
rect 2033 17 2099 152
rect 2335 150 2369 326
rect 2191 116 2369 150
rect 2191 70 2257 116
rect 2302 17 2368 82
rect 2514 326 2571 596
rect 2609 364 2665 649
rect 2514 260 2697 326
rect 2514 91 2571 260
rect 2624 17 2658 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 799 390 833 424
rect 1567 390 1601 424
rect 2143 390 2177 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
<< metal1 >>
rect 0 683 2784 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 0 617 2784 649
rect 0 616 50 617
rect 787 424 845 430
rect 787 390 799 424
rect 833 421 845 424
rect 1555 424 1613 430
rect 1555 421 1567 424
rect 833 393 1567 421
rect 833 390 845 393
rect 787 384 845 390
rect 1555 390 1567 393
rect 1601 421 1613 424
rect 2131 424 2189 430
rect 2131 421 2143 424
rect 1601 393 2143 421
rect 1601 390 1613 393
rect 1555 384 1613 390
rect 2131 390 2143 393
rect 2177 390 2189 424
rect 2131 384 2189 390
rect 0 49 50 50
rect 0 17 2784 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
rect 0 -49 2784 -17
<< labels >>
rlabel locali s 313 162 420 262 6 D
port 1 nsew signal input
rlabel locali s 2733 226 2767 364 6 Q
port 2 nsew signal output
rlabel locali s 2711 364 2767 596 6 Q
port 2 nsew signal output
rlabel locali s 2694 70 2767 226 6 Q
port 2 nsew signal output
rlabel locali s 2403 70 2469 596 6 Q_N
port 3 nsew signal output
rlabel metal1 s 2131 421 2189 430 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 2131 384 2189 393 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 1555 421 1613 430 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 1555 384 1613 393 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 787 421 845 430 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 787 393 2189 421 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 787 384 845 393 6 RESET_B
port 4 nsew signal input
rlabel locali s 587 288 653 430 6 SCD
port 5 nsew signal input
rlabel locali s 479 252 545 298 6 SCE
port 6 nsew signal input
rlabel locali s 121 332 359 376 6 SCE
port 6 nsew signal input
rlabel locali s 121 298 545 332 6 SCE
port 6 nsew signal input
rlabel locali s 757 236 929 326 6 CLK
port 7 nsew clock input
rlabel locali s 757 184 812 236 6 CLK
port 7 nsew clock input
rlabel metal1 s 0 -49 2784 49 8 VGND
port 8 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 9 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 10 nsew power bidirectional
rlabel metal1 s 0 617 2784 715 6 VPWR
port 11 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2784 666
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1036430
string GDS_START 1014664
<< end >>
