magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1564 561
rect 123 413 157 527
rect 291 413 325 527
rect 1154 339 1188 493
rect 1222 378 1288 527
rect 1322 339 1356 493
rect 1390 378 1456 527
rect 1490 339 1547 493
rect 755 289 1547 339
rect 18 211 356 285
rect 390 211 721 285
rect 755 211 1188 255
rect 1222 177 1259 289
rect 1293 211 1547 255
rect 123 17 157 109
rect 291 17 325 109
rect 459 17 493 109
rect 627 17 661 109
rect 799 17 928 109
rect 1030 17 1120 109
rect 1222 129 1456 177
rect 0 -17 1564 17
<< obsli1 >>
rect 18 379 89 493
rect 191 379 257 493
rect 359 441 777 493
rect 359 379 425 441
rect 18 319 425 379
rect 459 353 493 407
rect 527 387 593 441
rect 816 407 1120 493
rect 627 373 1120 407
rect 627 353 721 373
rect 459 319 721 353
rect 18 143 1188 177
rect 18 51 89 143
rect 191 51 257 143
rect 359 51 425 143
rect 527 51 593 143
rect 695 51 761 143
rect 962 79 996 143
rect 1154 95 1188 143
rect 1490 95 1547 177
rect 1154 51 1547 95
<< metal1 >>
rect 0 496 1564 592
rect 0 -48 1564 48
<< labels >>
rlabel locali s 18 211 356 285 6 A1
port 1 nsew signal input
rlabel locali s 390 211 721 285 6 A2
port 2 nsew signal input
rlabel locali s 755 211 1188 255 6 A3
port 3 nsew signal input
rlabel locali s 1293 211 1547 255 6 B1
port 4 nsew signal input
rlabel locali s 1490 339 1547 493 6 Y
port 5 nsew signal output
rlabel locali s 1322 339 1356 493 6 Y
port 5 nsew signal output
rlabel locali s 1222 177 1259 289 6 Y
port 5 nsew signal output
rlabel locali s 1222 129 1456 177 6 Y
port 5 nsew signal output
rlabel locali s 1154 339 1188 493 6 Y
port 5 nsew signal output
rlabel locali s 755 289 1547 339 6 Y
port 5 nsew signal output
rlabel locali s 1030 17 1120 109 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 799 17 928 109 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 627 17 661 109 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 459 17 493 109 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 291 17 325 109 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 123 17 157 109 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 1564 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1564 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1390 378 1456 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1222 378 1288 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 291 413 325 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 123 413 157 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 1564 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 1564 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1564 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 954334
string GDS_START 939850
<< end >>
