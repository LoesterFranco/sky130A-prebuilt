magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 119 326 173 493
rect 307 326 361 493
rect 495 326 549 493
rect 683 326 737 493
rect 871 326 925 493
rect 1059 326 1113 493
rect 1247 326 1301 493
rect 1435 326 1489 493
rect 1623 326 1677 493
rect 23 292 1731 326
rect 23 173 57 292
rect 91 207 1585 258
rect 1620 173 1731 292
rect 23 139 1731 173
rect 401 51 455 139
rect 589 51 643 139
rect 777 51 831 139
rect 965 51 1019 139
rect 1153 51 1207 139
rect 1341 51 1395 139
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 19 360 85 527
rect 207 360 273 527
rect 395 360 461 527
rect 583 360 649 527
rect 771 360 837 527
rect 959 360 1025 527
rect 1147 360 1213 527
rect 1335 360 1401 527
rect 1523 360 1589 527
rect 1711 360 1777 527
rect 233 17 367 105
rect 489 17 555 105
rect 677 17 743 105
rect 865 17 931 105
rect 1053 17 1119 105
rect 1241 17 1307 105
rect 1429 17 1563 105
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
<< metal1 >>
rect 0 561 1840 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 0 496 1840 527
rect 0 17 1840 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
rect 0 -48 1840 -17
<< labels >>
rlabel locali s 91 207 1585 258 6 A
port 1 nsew signal input
rlabel locali s 1623 326 1677 493 6 Y
port 2 nsew signal output
rlabel locali s 1620 173 1731 292 6 Y
port 2 nsew signal output
rlabel locali s 1435 326 1489 493 6 Y
port 2 nsew signal output
rlabel locali s 1341 51 1395 139 6 Y
port 2 nsew signal output
rlabel locali s 1247 326 1301 493 6 Y
port 2 nsew signal output
rlabel locali s 1153 51 1207 139 6 Y
port 2 nsew signal output
rlabel locali s 1059 326 1113 493 6 Y
port 2 nsew signal output
rlabel locali s 965 51 1019 139 6 Y
port 2 nsew signal output
rlabel locali s 871 326 925 493 6 Y
port 2 nsew signal output
rlabel locali s 777 51 831 139 6 Y
port 2 nsew signal output
rlabel locali s 683 326 737 493 6 Y
port 2 nsew signal output
rlabel locali s 589 51 643 139 6 Y
port 2 nsew signal output
rlabel locali s 495 326 549 493 6 Y
port 2 nsew signal output
rlabel locali s 401 51 455 139 6 Y
port 2 nsew signal output
rlabel locali s 307 326 361 493 6 Y
port 2 nsew signal output
rlabel locali s 119 326 173 493 6 Y
port 2 nsew signal output
rlabel locali s 23 292 1731 326 6 Y
port 2 nsew signal output
rlabel locali s 23 173 57 292 6 Y
port 2 nsew signal output
rlabel locali s 23 139 1731 173 6 Y
port 2 nsew signal output
rlabel metal1 s 0 -48 1840 48 8 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 496 1840 592 6 VPWR
port 4 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1840 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3378224
string GDS_START 3365844
<< end >>
