magic
tech sky130A
magscale 1 2
timestamp 1599588209
<< nwell >>
rect -38 332 1670 704
<< pwell >>
rect 0 0 1632 49
<< scpmos >>
rect 86 398 116 566
rect 210 398 240 566
rect 426 392 456 560
rect 534 392 564 592
rect 612 392 642 592
rect 723 508 753 592
rect 854 508 884 592
rect 1018 368 1048 592
rect 1113 368 1143 592
rect 1213 368 1243 592
rect 1415 424 1445 592
rect 1516 368 1546 592
<< nmoslvt >>
rect 84 142 114 252
rect 196 104 226 252
rect 423 98 453 246
rect 541 80 571 208
rect 613 80 643 208
rect 745 124 775 208
rect 823 124 853 208
rect 1021 74 1051 222
rect 1099 74 1129 222
rect 1201 74 1231 222
rect 1399 74 1429 184
rect 1501 74 1531 222
<< ndiff >>
rect 27 214 84 252
rect 27 180 39 214
rect 73 180 84 214
rect 27 142 84 180
rect 114 240 196 252
rect 114 206 141 240
rect 175 206 196 240
rect 114 150 196 206
rect 114 142 141 150
rect 129 116 141 142
rect 175 116 196 150
rect 129 104 196 116
rect 226 240 299 252
rect 226 206 253 240
rect 287 206 299 240
rect 226 150 299 206
rect 226 116 253 150
rect 287 116 299 150
rect 226 104 299 116
rect 353 234 423 246
rect 353 200 371 234
rect 405 200 423 234
rect 353 98 423 200
rect 453 208 503 246
rect 964 210 1021 222
rect 453 98 541 208
rect 468 82 541 98
rect 468 48 480 82
rect 514 80 541 82
rect 571 80 613 208
rect 643 192 745 208
rect 643 158 677 192
rect 711 158 745 192
rect 643 124 745 158
rect 775 124 823 208
rect 853 183 910 208
rect 853 149 864 183
rect 898 149 910 183
rect 853 124 910 149
rect 964 176 976 210
rect 1010 176 1021 210
rect 643 80 693 124
rect 964 120 1021 176
rect 514 48 526 80
rect 468 36 526 48
rect 964 86 976 120
rect 1010 86 1021 120
rect 964 74 1021 86
rect 1051 74 1099 222
rect 1129 199 1201 222
rect 1129 165 1140 199
rect 1174 165 1201 199
rect 1129 116 1201 165
rect 1129 82 1140 116
rect 1174 82 1201 116
rect 1129 74 1201 82
rect 1231 210 1288 222
rect 1231 176 1242 210
rect 1276 176 1288 210
rect 1448 188 1501 222
rect 1448 184 1456 188
rect 1231 120 1288 176
rect 1231 86 1242 120
rect 1276 86 1288 120
rect 1231 74 1288 86
rect 1342 142 1399 184
rect 1342 108 1354 142
rect 1388 108 1399 142
rect 1342 74 1399 108
rect 1429 154 1456 184
rect 1490 154 1501 188
rect 1429 116 1501 154
rect 1429 82 1456 116
rect 1490 82 1501 116
rect 1429 74 1501 82
rect 1531 208 1605 222
rect 1531 174 1558 208
rect 1592 174 1605 208
rect 1531 120 1605 174
rect 1531 86 1558 120
rect 1592 86 1605 120
rect 1531 74 1605 86
<< pdiff >>
rect 134 596 192 608
rect 134 566 146 596
rect 27 554 86 566
rect 27 520 39 554
rect 73 520 86 554
rect 27 444 86 520
rect 27 410 39 444
rect 73 410 86 444
rect 27 398 86 410
rect 116 562 146 566
rect 180 566 192 596
rect 180 562 210 566
rect 116 398 210 562
rect 240 444 313 566
rect 474 580 534 592
rect 474 560 486 580
rect 240 410 260 444
rect 294 410 313 444
rect 240 398 313 410
rect 367 441 426 560
rect 367 407 379 441
rect 413 407 426 441
rect 367 392 426 407
rect 456 546 486 560
rect 520 546 534 580
rect 456 392 534 546
rect 564 392 612 592
rect 642 531 723 592
rect 642 497 657 531
rect 691 508 723 531
rect 753 508 854 592
rect 884 580 1018 592
rect 884 546 897 580
rect 931 546 966 580
rect 1000 546 1018 580
rect 884 508 1018 546
rect 691 497 705 508
rect 642 392 705 497
rect 965 368 1018 508
rect 1048 580 1113 592
rect 1048 546 1066 580
rect 1100 546 1113 580
rect 1048 497 1113 546
rect 1048 463 1066 497
rect 1100 463 1113 497
rect 1048 414 1113 463
rect 1048 380 1066 414
rect 1100 380 1113 414
rect 1048 368 1113 380
rect 1143 580 1213 592
rect 1143 546 1156 580
rect 1190 546 1213 580
rect 1143 462 1213 546
rect 1143 428 1156 462
rect 1190 428 1213 462
rect 1143 368 1213 428
rect 1243 580 1302 592
rect 1243 546 1256 580
rect 1290 546 1302 580
rect 1243 462 1302 546
rect 1243 428 1256 462
rect 1290 428 1302 462
rect 1243 368 1302 428
rect 1356 580 1415 592
rect 1356 546 1368 580
rect 1402 546 1415 580
rect 1356 470 1415 546
rect 1356 436 1368 470
rect 1402 436 1415 470
rect 1356 424 1415 436
rect 1445 580 1516 592
rect 1445 546 1458 580
rect 1492 546 1516 580
rect 1445 470 1516 546
rect 1445 436 1458 470
rect 1492 436 1516 470
rect 1445 424 1516 436
rect 1463 368 1516 424
rect 1546 580 1605 592
rect 1546 546 1559 580
rect 1593 546 1605 580
rect 1546 497 1605 546
rect 1546 463 1559 497
rect 1593 463 1605 497
rect 1546 414 1605 463
rect 1546 380 1559 414
rect 1593 380 1605 414
rect 1546 368 1605 380
<< ndiffc >>
rect 39 180 73 214
rect 141 206 175 240
rect 141 116 175 150
rect 253 206 287 240
rect 253 116 287 150
rect 371 200 405 234
rect 480 48 514 82
rect 677 158 711 192
rect 864 149 898 183
rect 976 176 1010 210
rect 976 86 1010 120
rect 1140 165 1174 199
rect 1140 82 1174 116
rect 1242 176 1276 210
rect 1242 86 1276 120
rect 1354 108 1388 142
rect 1456 154 1490 188
rect 1456 82 1490 116
rect 1558 174 1592 208
rect 1558 86 1592 120
<< pdiffc >>
rect 39 520 73 554
rect 39 410 73 444
rect 146 562 180 596
rect 260 410 294 444
rect 379 407 413 441
rect 486 546 520 580
rect 657 497 691 531
rect 897 546 931 580
rect 966 546 1000 580
rect 1066 546 1100 580
rect 1066 463 1100 497
rect 1066 380 1100 414
rect 1156 546 1190 580
rect 1156 428 1190 462
rect 1256 546 1290 580
rect 1256 428 1290 462
rect 1368 546 1402 580
rect 1368 436 1402 470
rect 1458 546 1492 580
rect 1458 436 1492 470
rect 1559 546 1593 580
rect 1559 463 1593 497
rect 1559 380 1593 414
<< poly >>
rect 86 566 116 592
rect 534 592 564 618
rect 612 592 642 618
rect 723 592 753 618
rect 854 592 884 618
rect 1018 592 1048 618
rect 1113 592 1143 618
rect 1213 592 1243 618
rect 1415 592 1445 618
rect 1516 592 1546 618
rect 210 566 240 592
rect 426 560 456 586
rect 86 383 116 398
rect 210 383 240 398
rect 723 493 753 508
rect 854 493 884 508
rect 720 476 756 493
rect 720 460 803 476
rect 851 464 887 493
rect 720 426 753 460
rect 787 426 803 460
rect 720 410 803 426
rect 845 448 911 464
rect 845 414 861 448
rect 895 414 911 448
rect 845 398 911 414
rect 83 356 119 383
rect 207 356 243 383
rect 426 377 456 392
rect 534 377 564 392
rect 612 377 642 392
rect 83 340 153 356
rect 83 306 103 340
rect 137 306 153 340
rect 83 290 153 306
rect 195 340 261 356
rect 195 306 211 340
rect 245 306 261 340
rect 195 290 261 306
rect 309 334 375 350
rect 309 300 325 334
rect 359 314 375 334
rect 423 314 459 377
rect 531 360 567 377
rect 501 344 567 360
rect 359 300 453 314
rect 84 252 114 290
rect 196 252 226 290
rect 309 284 453 300
rect 501 310 517 344
rect 551 310 567 344
rect 609 368 645 377
rect 609 338 775 368
rect 501 294 567 310
rect 84 116 114 142
rect 423 246 453 284
rect 537 253 567 294
rect 613 280 679 296
rect 196 78 226 104
rect 537 223 571 253
rect 541 208 571 223
rect 613 246 629 280
rect 663 246 679 280
rect 613 230 679 246
rect 613 208 643 230
rect 745 208 775 338
rect 845 253 875 398
rect 1415 409 1445 424
rect 1412 408 1448 409
rect 1399 378 1448 408
rect 1018 353 1048 368
rect 1113 353 1143 368
rect 1213 353 1243 368
rect 1015 336 1051 353
rect 917 320 1051 336
rect 917 286 933 320
rect 967 286 1051 320
rect 1110 310 1146 353
rect 1210 336 1246 353
rect 1201 320 1267 336
rect 917 270 1051 286
rect 823 223 875 253
rect 823 208 853 223
rect 1021 222 1051 270
rect 1093 294 1159 310
rect 1093 260 1109 294
rect 1143 260 1159 294
rect 1093 244 1159 260
rect 1201 286 1217 320
rect 1251 300 1267 320
rect 1399 300 1429 378
rect 1516 353 1546 368
rect 1513 330 1549 353
rect 1251 286 1429 300
rect 1201 270 1429 286
rect 1099 222 1129 244
rect 1201 222 1231 270
rect 423 72 453 98
rect 745 102 775 124
rect 715 86 781 102
rect 823 98 853 124
rect 541 54 571 80
rect 613 54 643 80
rect 715 52 731 86
rect 765 52 781 86
rect 1399 184 1429 270
rect 1477 314 1549 330
rect 1477 280 1493 314
rect 1527 280 1549 314
rect 1477 264 1549 280
rect 1501 222 1531 264
rect 715 36 781 52
rect 1021 48 1051 74
rect 1099 48 1129 74
rect 1201 48 1231 74
rect 1399 48 1429 74
rect 1501 48 1531 74
<< polycont >>
rect 753 426 787 460
rect 861 414 895 448
rect 103 306 137 340
rect 211 306 245 340
rect 325 300 359 334
rect 517 310 551 344
rect 629 246 663 280
rect 933 286 967 320
rect 1109 260 1143 294
rect 1217 286 1251 320
rect 731 52 765 86
rect 1493 280 1527 314
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 130 596 196 649
rect 19 554 89 570
rect 19 520 39 554
rect 73 520 89 554
rect 130 562 146 596
rect 180 562 196 596
rect 130 546 196 562
rect 470 580 537 649
rect 470 546 486 580
rect 520 546 537 580
rect 571 581 803 615
rect 19 512 89 520
rect 19 478 535 512
rect 19 444 89 478
rect 19 410 39 444
rect 73 410 89 444
rect 19 394 89 410
rect 237 410 260 444
rect 294 410 329 444
rect 237 394 329 410
rect 19 256 53 394
rect 87 340 161 356
rect 87 306 103 340
rect 137 306 161 340
rect 87 290 161 306
rect 195 340 261 356
rect 195 306 211 340
rect 245 306 261 340
rect 195 290 261 306
rect 295 350 329 394
rect 363 441 443 444
rect 363 407 379 441
rect 413 407 443 441
rect 363 388 443 407
rect 295 334 375 350
rect 295 300 325 334
rect 359 300 375 334
rect 295 284 375 300
rect 295 256 329 284
rect 19 214 89 256
rect 19 180 39 214
rect 73 180 89 214
rect 19 138 89 180
rect 125 240 191 256
rect 125 206 141 240
rect 175 206 191 240
rect 125 150 191 206
rect 125 116 141 150
rect 175 116 191 150
rect 125 17 191 116
rect 237 240 329 256
rect 409 260 443 388
rect 501 360 535 478
rect 571 428 605 581
rect 639 531 703 547
rect 639 497 657 531
rect 691 497 703 531
rect 639 481 703 497
rect 571 394 635 428
rect 501 344 567 360
rect 501 310 517 344
rect 551 310 567 344
rect 501 294 567 310
rect 601 296 635 394
rect 669 364 703 481
rect 737 460 803 581
rect 881 580 1016 649
rect 881 546 897 580
rect 931 546 966 580
rect 1000 546 1016 580
rect 881 530 1016 546
rect 1050 580 1116 596
rect 1050 546 1066 580
rect 1100 546 1116 580
rect 1050 497 1116 546
rect 1050 464 1066 497
rect 737 426 753 460
rect 787 426 803 460
rect 737 410 803 426
rect 845 463 1066 464
rect 1100 463 1116 497
rect 845 448 1116 463
rect 845 414 861 448
rect 895 414 1116 448
rect 845 398 1066 414
rect 1017 380 1066 398
rect 1100 380 1116 414
rect 1156 580 1206 649
rect 1190 546 1206 580
rect 1156 462 1206 546
rect 1190 428 1206 462
rect 1156 412 1206 428
rect 1240 580 1334 596
rect 1240 546 1256 580
rect 1290 546 1334 580
rect 1240 462 1334 546
rect 1240 428 1256 462
rect 1290 428 1334 462
rect 1240 412 1334 428
rect 1017 378 1116 380
rect 669 330 983 364
rect 601 280 679 296
rect 601 260 629 280
rect 409 250 629 260
rect 237 206 253 240
rect 287 206 329 240
rect 237 150 329 206
rect 365 246 629 250
rect 663 246 679 280
rect 365 234 679 246
rect 365 200 371 234
rect 405 226 679 234
rect 405 200 443 226
rect 365 184 443 200
rect 716 192 750 330
rect 917 320 983 330
rect 917 286 933 320
rect 967 286 983 320
rect 917 270 983 286
rect 1017 344 1266 378
rect 1017 226 1051 344
rect 1201 320 1266 344
rect 1085 294 1159 310
rect 1085 260 1109 294
rect 1143 260 1159 294
rect 1201 286 1217 320
rect 1251 286 1266 320
rect 1201 270 1266 286
rect 1085 236 1159 260
rect 1300 236 1334 412
rect 638 158 677 192
rect 711 158 750 192
rect 237 116 253 150
rect 287 116 598 150
rect 638 142 750 158
rect 848 183 914 212
rect 848 149 864 183
rect 898 149 914 183
rect 237 100 329 116
rect 564 102 598 116
rect 564 86 781 102
rect 464 48 480 82
rect 514 48 530 82
rect 564 52 731 86
rect 765 52 781 86
rect 564 51 781 52
rect 464 17 530 48
rect 848 17 914 149
rect 960 210 1051 226
rect 960 176 976 210
rect 1010 176 1051 210
rect 1226 210 1334 236
rect 960 120 1051 176
rect 960 86 976 120
rect 1010 86 1051 120
rect 960 70 1051 86
rect 1124 199 1190 202
rect 1124 165 1140 199
rect 1174 165 1190 199
rect 1124 116 1190 165
rect 1124 82 1140 116
rect 1174 82 1190 116
rect 1124 17 1190 82
rect 1226 176 1242 210
rect 1276 202 1334 210
rect 1368 580 1402 596
rect 1368 470 1402 546
rect 1368 330 1402 436
rect 1442 580 1508 649
rect 1442 546 1458 580
rect 1492 546 1508 580
rect 1442 470 1508 546
rect 1442 436 1458 470
rect 1492 436 1508 470
rect 1442 420 1508 436
rect 1543 580 1611 596
rect 1543 546 1559 580
rect 1593 546 1611 580
rect 1543 497 1611 546
rect 1543 463 1559 497
rect 1593 463 1611 497
rect 1543 414 1611 463
rect 1543 380 1559 414
rect 1593 380 1611 414
rect 1543 364 1611 380
rect 1368 314 1543 330
rect 1368 280 1493 314
rect 1527 280 1543 314
rect 1368 264 1543 280
rect 1276 176 1292 202
rect 1226 120 1292 176
rect 1368 168 1404 264
rect 1577 208 1611 364
rect 1226 86 1242 120
rect 1276 86 1292 120
rect 1226 70 1292 86
rect 1338 142 1404 168
rect 1338 108 1354 142
rect 1388 108 1404 142
rect 1338 70 1404 108
rect 1440 154 1456 188
rect 1490 154 1506 188
rect 1440 116 1506 154
rect 1440 82 1456 116
rect 1490 82 1506 116
rect 1440 17 1506 82
rect 1542 174 1558 208
rect 1592 174 1611 208
rect 1542 120 1611 174
rect 1542 86 1558 120
rect 1592 86 1611 120
rect 1542 70 1611 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dlrbp_1
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 1 nsew
flabel corelocali s 1567 94 1601 128 0 FreeSans 340 0 0 0 Q_N
port 9 nsew
flabel corelocali s 1567 168 1601 202 0 FreeSans 340 0 0 0 Q_N
port 9 nsew
flabel corelocali s 1279 464 1313 498 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 1279 538 1313 572 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 GATE
port 2 nsew
flabel corelocali s 1087 242 1121 276 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 1632 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3069844
string GDS_START 3057080
<< end >>
