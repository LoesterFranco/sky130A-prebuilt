magic
tech sky130A
magscale 1 2
timestamp 1601050058
<< locali >>
rect 17 195 87 325
rect 349 201 431 325
rect 717 193 783 213
rect 717 187 799 193
rect 717 153 765 187
rect 717 147 799 153
rect 1456 187 1565 213
rect 1456 153 1515 187
rect 1549 153 1565 187
rect 2040 326 2097 493
rect 1847 219 1938 265
rect 1456 147 1565 153
rect 2061 143 2097 326
rect 2040 51 2097 143
rect 2323 291 2375 493
rect 2333 165 2375 291
rect 2323 51 2375 165
<< viali >>
rect 765 153 799 187
rect 1515 153 1549 187
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2392 561
rect 35 393 69 493
rect 103 427 169 527
rect 35 359 168 393
rect 122 161 168 359
rect 35 127 168 161
rect 35 69 69 127
rect 103 17 169 93
rect 203 69 247 493
rect 286 427 357 527
rect 391 393 425 493
rect 467 450 633 484
rect 281 359 425 393
rect 281 165 315 359
rect 465 315 565 391
rect 281 127 425 165
rect 465 141 509 315
rect 599 281 633 450
rect 681 441 757 527
rect 817 407 851 475
rect 667 357 937 407
rect 975 383 1041 527
rect 1250 450 1416 484
rect 1464 451 1540 527
rect 667 315 717 357
rect 819 281 869 297
rect 599 247 869 281
rect 599 239 683 247
rect 545 129 615 203
rect 286 17 357 93
rect 391 61 425 127
rect 649 93 683 239
rect 825 231 869 247
rect 903 213 937 357
rect 971 283 1172 331
rect 1212 315 1259 397
rect 971 247 1037 283
rect 1307 261 1348 381
rect 1099 213 1165 247
rect 903 179 1165 213
rect 1213 225 1348 261
rect 1382 281 1416 450
rect 1588 417 1622 475
rect 1728 451 2006 527
rect 1450 383 2006 417
rect 1450 315 1500 383
rect 1382 247 1652 281
rect 1213 212 1281 225
rect 903 153 947 179
rect 881 119 947 153
rect 480 53 683 93
rect 717 17 751 105
rect 785 85 851 101
rect 981 85 1015 143
rect 1237 141 1281 212
rect 1382 93 1416 247
rect 1608 215 1652 247
rect 1686 168 1720 383
rect 1754 315 1911 349
rect 1754 222 1811 315
rect 1972 265 2006 383
rect 1767 185 1811 222
rect 1972 199 2025 265
rect 1686 167 1723 168
rect 1643 133 1723 167
rect 1767 151 1895 185
rect 785 51 1015 85
rect 1065 17 1135 93
rect 1260 53 1416 93
rect 1450 17 1515 105
rect 1549 85 1615 109
rect 1757 85 1791 117
rect 1549 51 1791 85
rect 1853 53 1895 151
rect 1945 17 2006 161
rect 2132 265 2195 483
rect 2231 353 2289 527
rect 2132 199 2299 265
rect 2132 51 2195 199
rect 2230 17 2289 109
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2392 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
<< metal1 >>
rect 0 561 2392 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2392 561
rect 0 496 2392 527
rect 753 187 811 193
rect 753 153 765 187
rect 799 184 811 187
rect 1503 187 1561 193
rect 1503 184 1515 187
rect 799 156 1515 184
rect 799 153 811 156
rect 753 147 811 153
rect 1503 153 1515 156
rect 1549 153 1561 187
rect 1503 147 1561 153
rect 0 17 2392 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2392 17
rect 0 -48 2392 -17
<< obsm1 >>
rect 201 388 259 397
rect 477 388 535 397
rect 1213 388 1271 397
rect 201 360 1271 388
rect 201 351 259 360
rect 477 351 535 360
rect 1213 351 1271 360
rect 1121 320 1179 329
rect 1759 320 1817 329
rect 1121 292 1817 320
rect 1121 283 1179 292
rect 1759 283 1817 292
rect 1213 252 1271 261
rect 584 224 1271 252
rect 584 193 627 224
rect 1213 215 1271 224
rect 110 184 168 193
rect 569 184 627 193
rect 110 156 627 184
rect 110 147 168 156
rect 569 147 627 156
<< labels >>
rlabel locali s 349 201 431 325 6 D
port 1 nsew signal input
rlabel locali s 2333 165 2375 291 6 Q
port 2 nsew signal output
rlabel locali s 2323 291 2375 493 6 Q
port 2 nsew signal output
rlabel locali s 2323 51 2375 165 6 Q
port 2 nsew signal output
rlabel locali s 2061 143 2097 326 6 Q_N
port 3 nsew signal output
rlabel locali s 2040 326 2097 493 6 Q_N
port 3 nsew signal output
rlabel locali s 2040 51 2097 143 6 Q_N
port 3 nsew signal output
rlabel locali s 1847 219 1938 265 6 RESET_B
port 4 nsew signal input
rlabel viali s 765 153 799 187 6 SET_B
port 5 nsew signal input
rlabel locali s 717 193 783 213 6 SET_B
port 5 nsew signal input
rlabel locali s 717 147 799 193 6 SET_B
port 5 nsew signal input
rlabel viali s 1515 153 1549 187 6 SET_B
port 5 nsew signal input
rlabel locali s 1456 147 1565 213 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1503 184 1561 193 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1503 147 1561 156 6 SET_B
port 5 nsew signal input
rlabel metal1 s 753 184 811 193 6 SET_B
port 5 nsew signal input
rlabel metal1 s 753 156 1561 184 6 SET_B
port 5 nsew signal input
rlabel metal1 s 753 147 811 156 6 SET_B
port 5 nsew signal input
rlabel locali s 17 195 87 325 6 CLK_N
port 6 nsew clock input
rlabel metal1 s 0 -48 2392 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 496 2392 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2392 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3319692
string GDS_START 3300142
<< end >>
