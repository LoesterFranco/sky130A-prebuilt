magic
tech sky130A
magscale 1 2
timestamp 1599588209
<< nwell >>
rect -38 332 1478 704
<< pwell >>
rect 0 0 1440 49
<< scpmos >>
rect 87 394 117 562
rect 211 394 241 562
rect 416 392 446 560
rect 540 392 570 592
rect 624 392 654 592
rect 763 508 793 592
rect 900 508 930 592
rect 1083 368 1113 568
rect 1207 368 1237 568
rect 1324 368 1354 592
<< nmoslvt >>
rect 84 136 114 246
rect 202 98 232 246
rect 430 82 460 230
rect 651 74 681 202
rect 729 74 759 202
rect 824 74 854 158
rect 909 74 939 158
rect 1109 74 1139 222
rect 1187 74 1217 222
rect 1305 74 1335 222
<< ndiff >>
rect 27 208 84 246
rect 27 174 39 208
rect 73 174 84 208
rect 27 136 84 174
rect 114 136 202 246
rect 129 98 202 136
rect 232 224 285 246
rect 232 190 243 224
rect 277 190 285 224
rect 232 98 285 190
rect 373 218 430 230
rect 373 184 385 218
rect 419 184 430 218
rect 129 82 187 98
rect 129 48 141 82
rect 175 48 187 82
rect 373 82 430 184
rect 460 202 510 230
rect 460 82 651 202
rect 129 36 187 48
rect 475 48 487 82
rect 521 48 590 82
rect 624 74 651 82
rect 681 74 729 202
rect 759 158 809 202
rect 1052 210 1109 222
rect 1052 176 1064 210
rect 1098 176 1109 210
rect 759 133 824 158
rect 759 99 779 133
rect 813 99 824 133
rect 759 74 824 99
rect 854 74 909 158
rect 939 120 998 158
rect 939 86 951 120
rect 985 86 998 120
rect 939 74 998 86
rect 1052 120 1109 176
rect 1052 86 1064 120
rect 1098 86 1109 120
rect 1052 74 1109 86
rect 1139 74 1187 222
rect 1217 197 1305 222
rect 1217 163 1244 197
rect 1278 163 1305 197
rect 1217 115 1305 163
rect 1217 81 1244 115
rect 1278 81 1305 115
rect 1217 74 1305 81
rect 1335 210 1408 222
rect 1335 176 1362 210
rect 1396 176 1408 210
rect 1335 120 1408 176
rect 1335 86 1362 120
rect 1396 86 1408 120
rect 1335 74 1408 86
rect 624 48 636 74
rect 1232 73 1290 74
rect 475 36 636 48
<< pdiff >>
rect 464 606 522 618
rect 135 562 193 563
rect 28 550 87 562
rect 28 516 40 550
rect 74 516 87 550
rect 28 440 87 516
rect 28 406 40 440
rect 74 406 87 440
rect 28 394 87 406
rect 117 551 211 562
rect 117 517 147 551
rect 181 517 211 551
rect 117 440 211 517
rect 117 406 147 440
rect 181 406 211 440
rect 117 394 211 406
rect 241 550 300 562
rect 464 572 476 606
rect 510 592 522 606
rect 510 572 540 592
rect 464 560 540 572
rect 241 516 254 550
rect 288 516 300 550
rect 241 440 300 516
rect 241 406 254 440
rect 288 406 300 440
rect 241 394 300 406
rect 357 446 416 560
rect 357 412 369 446
rect 403 412 416 446
rect 357 392 416 412
rect 446 392 540 560
rect 570 392 624 592
rect 654 508 763 592
rect 793 508 900 592
rect 930 568 983 592
rect 1255 582 1324 592
rect 1255 568 1267 582
rect 930 556 1083 568
rect 930 522 943 556
rect 977 522 1036 556
rect 1070 522 1083 556
rect 930 508 1083 522
rect 654 470 714 508
rect 654 436 668 470
rect 702 436 714 470
rect 654 392 714 436
rect 1030 368 1083 508
rect 1113 556 1207 568
rect 1113 522 1143 556
rect 1177 522 1207 556
rect 1113 485 1207 522
rect 1113 451 1143 485
rect 1177 451 1207 485
rect 1113 414 1207 451
rect 1113 380 1143 414
rect 1177 380 1207 414
rect 1113 368 1207 380
rect 1237 548 1267 568
rect 1301 548 1324 582
rect 1237 514 1324 548
rect 1237 480 1267 514
rect 1301 480 1324 514
rect 1237 446 1324 480
rect 1237 412 1267 446
rect 1301 412 1324 446
rect 1237 368 1324 412
rect 1354 580 1413 592
rect 1354 546 1367 580
rect 1401 546 1413 580
rect 1354 497 1413 546
rect 1354 463 1367 497
rect 1401 463 1413 497
rect 1354 414 1413 463
rect 1354 380 1367 414
rect 1401 380 1413 414
rect 1354 368 1413 380
<< ndiffc >>
rect 39 174 73 208
rect 243 190 277 224
rect 385 184 419 218
rect 141 48 175 82
rect 487 48 521 82
rect 590 48 624 82
rect 1064 176 1098 210
rect 779 99 813 133
rect 951 86 985 120
rect 1064 86 1098 120
rect 1244 163 1278 197
rect 1244 81 1278 115
rect 1362 176 1396 210
rect 1362 86 1396 120
<< pdiffc >>
rect 40 516 74 550
rect 40 406 74 440
rect 147 517 181 551
rect 147 406 181 440
rect 476 572 510 606
rect 254 516 288 550
rect 254 406 288 440
rect 369 412 403 446
rect 943 522 977 556
rect 1036 522 1070 556
rect 668 436 702 470
rect 1143 522 1177 556
rect 1143 451 1177 485
rect 1143 380 1177 414
rect 1267 548 1301 582
rect 1267 480 1301 514
rect 1267 412 1301 446
rect 1367 546 1401 580
rect 1367 463 1401 497
rect 1367 380 1401 414
<< poly >>
rect 87 562 117 588
rect 211 562 241 588
rect 416 560 446 586
rect 540 592 570 618
rect 624 592 654 618
rect 763 592 793 618
rect 900 592 930 618
rect 87 379 117 394
rect 211 379 241 394
rect 1083 568 1113 594
rect 1207 568 1237 594
rect 1324 592 1354 618
rect 763 493 793 508
rect 900 493 930 508
rect 760 472 796 493
rect 897 472 933 493
rect 760 456 849 472
rect 760 422 799 456
rect 833 422 849 456
rect 760 406 849 422
rect 897 456 963 472
rect 897 422 913 456
rect 947 422 963 456
rect 897 406 963 422
rect 84 356 120 379
rect 208 356 244 379
rect 416 377 446 392
rect 540 377 570 392
rect 624 377 654 392
rect 84 340 153 356
rect 84 306 103 340
rect 137 306 153 340
rect 84 290 153 306
rect 201 340 267 356
rect 201 306 217 340
rect 251 306 267 340
rect 413 334 449 377
rect 201 290 267 306
rect 315 318 449 334
rect 537 318 573 377
rect 621 355 657 377
rect 760 376 790 406
rect 84 246 114 290
rect 202 246 232 290
rect 315 284 331 318
rect 365 298 449 318
rect 507 302 573 318
rect 365 284 460 298
rect 315 268 460 284
rect 84 110 114 136
rect 430 230 460 268
rect 507 268 523 302
rect 557 268 573 302
rect 615 339 681 355
rect 615 305 631 339
rect 665 305 681 339
rect 615 289 681 305
rect 729 346 790 376
rect 507 252 573 268
rect 543 247 573 252
rect 202 72 232 98
rect 543 217 681 247
rect 651 202 681 217
rect 729 202 759 346
rect 801 288 867 304
rect 915 298 945 406
rect 1083 353 1113 368
rect 1207 353 1237 368
rect 1324 353 1354 368
rect 1080 345 1116 353
rect 801 254 817 288
rect 851 254 867 288
rect 801 238 867 254
rect 909 268 945 298
rect 993 315 1116 345
rect 993 310 1059 315
rect 1204 310 1240 353
rect 1321 330 1357 353
rect 1289 314 1357 330
rect 993 276 1009 310
rect 1043 276 1059 310
rect 430 56 460 82
rect 824 158 854 238
rect 909 158 939 268
rect 993 267 1059 276
rect 1181 294 1247 310
rect 993 237 1139 267
rect 1181 260 1197 294
rect 1231 260 1247 294
rect 1289 280 1305 314
rect 1339 280 1357 314
rect 1289 264 1357 280
rect 1181 244 1247 260
rect 1109 222 1139 237
rect 1187 222 1217 244
rect 1305 222 1335 264
rect 651 48 681 74
rect 729 48 759 74
rect 824 48 854 74
rect 909 48 939 74
rect 1109 48 1139 74
rect 1187 48 1217 74
rect 1305 48 1335 74
<< polycont >>
rect 799 422 833 456
rect 913 422 947 456
rect 103 306 137 340
rect 217 306 251 340
rect 331 284 365 318
rect 523 268 557 302
rect 631 305 665 339
rect 817 254 851 288
rect 1009 276 1043 310
rect 1197 260 1231 294
rect 1305 280 1339 314
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 19 550 90 566
rect 19 516 40 550
rect 74 516 90 550
rect 19 440 90 516
rect 19 406 40 440
rect 74 406 90 440
rect 19 390 90 406
rect 131 551 197 649
rect 460 606 526 649
rect 460 572 476 606
rect 510 572 526 606
rect 131 517 147 551
rect 181 517 197 551
rect 131 440 197 517
rect 131 406 147 440
rect 181 406 197 440
rect 131 390 197 406
rect 238 550 335 566
rect 238 516 254 550
rect 288 538 335 550
rect 927 556 1086 649
rect 1251 582 1317 649
rect 288 516 849 538
rect 238 504 849 516
rect 927 522 943 556
rect 977 522 1036 556
rect 1070 522 1086 556
rect 927 506 1086 522
rect 1127 556 1193 572
rect 1127 522 1143 556
rect 1177 522 1193 556
rect 238 440 335 504
rect 238 406 254 440
rect 288 406 335 440
rect 238 390 335 406
rect 19 250 53 390
rect 87 340 167 356
rect 87 306 103 340
rect 137 306 167 340
rect 87 290 167 306
rect 201 340 267 356
rect 201 306 217 340
rect 251 306 267 340
rect 201 290 267 306
rect 301 334 335 390
rect 369 446 449 470
rect 403 412 449 446
rect 651 436 668 470
rect 702 436 749 470
rect 369 402 449 412
rect 369 368 681 402
rect 301 318 381 334
rect 301 284 331 318
rect 365 284 381 318
rect 301 268 381 284
rect 301 250 335 268
rect 19 208 89 250
rect 19 174 39 208
rect 73 174 89 208
rect 213 224 335 250
rect 415 234 449 368
rect 615 339 681 368
rect 213 190 243 224
rect 277 190 335 224
rect 213 184 335 190
rect 369 218 449 234
rect 369 184 385 218
rect 419 184 449 218
rect 507 302 573 318
rect 507 268 523 302
rect 557 268 573 302
rect 19 150 89 174
rect 507 150 573 268
rect 615 305 631 339
rect 665 305 681 339
rect 715 372 749 436
rect 783 456 849 504
rect 1127 485 1193 522
rect 1127 472 1143 485
rect 783 422 799 456
rect 833 422 849 456
rect 783 406 849 422
rect 897 456 1143 472
rect 897 422 913 456
rect 947 451 1143 456
rect 1177 451 1193 485
rect 947 422 1193 451
rect 897 414 1193 422
rect 897 406 1143 414
rect 1093 380 1143 406
rect 1177 380 1193 414
rect 1251 548 1267 582
rect 1301 548 1317 582
rect 1251 514 1317 548
rect 1251 480 1267 514
rect 1301 480 1317 514
rect 1251 446 1317 480
rect 1251 412 1267 446
rect 1301 412 1317 446
rect 1351 580 1423 596
rect 1351 546 1367 580
rect 1401 546 1423 580
rect 1351 497 1423 546
rect 1351 463 1367 497
rect 1401 463 1423 497
rect 1351 414 1423 463
rect 1093 378 1193 380
rect 1351 380 1367 414
rect 1401 380 1423 414
rect 715 338 1014 372
rect 615 304 681 305
rect 980 326 1014 338
rect 1093 344 1317 378
rect 1351 364 1423 380
rect 980 310 1059 326
rect 615 288 867 304
rect 615 254 817 288
rect 851 254 867 288
rect 615 238 867 254
rect 980 276 1009 310
rect 1043 276 1059 310
rect 980 260 1059 276
rect 980 204 1014 260
rect 1093 226 1127 344
rect 1283 330 1317 344
rect 1283 314 1355 330
rect 1177 294 1247 310
rect 1177 260 1197 294
rect 1231 260 1247 294
rect 1283 280 1305 314
rect 1339 280 1355 314
rect 1283 264 1355 280
rect 1177 236 1247 260
rect 1389 226 1423 364
rect 19 116 573 150
rect 763 170 1014 204
rect 1048 210 1127 226
rect 1048 176 1064 210
rect 1098 176 1127 210
rect 1346 210 1423 226
rect 763 133 829 170
rect 763 99 779 133
rect 813 99 829 133
rect 125 48 141 82
rect 175 48 191 82
rect 125 17 191 48
rect 471 48 487 82
rect 521 48 590 82
rect 624 48 640 82
rect 763 70 829 99
rect 934 120 1002 136
rect 934 86 951 120
rect 985 86 1002 120
rect 471 17 640 48
rect 934 17 1002 86
rect 1048 120 1127 176
rect 1048 86 1064 120
rect 1098 86 1127 120
rect 1048 70 1127 86
rect 1228 197 1294 202
rect 1228 163 1244 197
rect 1278 163 1294 197
rect 1228 115 1294 163
rect 1228 81 1244 115
rect 1278 81 1294 115
rect 1228 17 1294 81
rect 1346 176 1362 210
rect 1396 176 1423 210
rect 1346 120 1423 176
rect 1346 86 1362 120
rect 1396 86 1423 120
rect 1346 70 1423 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 683 1440 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 0 617 1440 649
rect 0 17 1440 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -49 1440 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dlrtn_1
flabel pwell s 0 0 1440 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 0 617 1440 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 1440 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 1440 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 1 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew
flabel corelocali s 1183 242 1217 276 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew
flabel corelocali s 1375 390 1409 424 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 1375 464 1409 498 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 1375 538 1409 572 0 FreeSans 340 0 0 0 Q
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 1440 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3140018
string GDS_START 3129046
<< end >>
