magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 89 47 119 177
rect 165 47 195 177
rect 381 47 411 177
rect 487 47 517 177
rect 590 47 620 177
rect 684 47 714 177
<< pmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 373 297 409 497
rect 479 297 515 497
rect 582 297 618 497
rect 676 297 712 497
<< ndiff >>
rect 27 165 89 177
rect 27 131 35 165
rect 69 131 89 165
rect 27 97 89 131
rect 27 63 35 97
rect 69 63 89 97
rect 27 47 89 63
rect 119 47 165 177
rect 195 101 257 177
rect 195 67 215 101
rect 249 67 257 101
rect 195 47 257 67
rect 319 101 381 177
rect 319 67 327 101
rect 361 67 381 101
rect 319 47 381 67
rect 411 47 487 177
rect 517 97 590 177
rect 517 63 527 97
rect 561 63 590 97
rect 517 47 590 63
rect 620 101 684 177
rect 620 67 630 101
rect 664 67 684 101
rect 620 47 684 67
rect 714 165 793 177
rect 714 131 751 165
rect 785 131 793 165
rect 714 97 793 131
rect 714 63 751 97
rect 785 63 793 97
rect 714 47 793 63
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 409 175 497
rect 117 375 129 409
rect 163 375 175 409
rect 117 297 175 375
rect 211 485 265 497
rect 211 451 223 485
rect 257 451 265 485
rect 211 297 265 451
rect 319 477 373 497
rect 319 443 327 477
rect 361 443 373 477
rect 319 297 373 443
rect 409 477 479 497
rect 409 443 426 477
rect 460 443 479 477
rect 409 407 479 443
rect 409 373 426 407
rect 460 373 479 407
rect 409 297 479 373
rect 515 477 582 497
rect 515 443 536 477
rect 570 443 582 477
rect 515 409 582 443
rect 515 375 536 409
rect 570 375 582 409
rect 515 297 582 375
rect 618 477 676 497
rect 618 443 630 477
rect 664 443 676 477
rect 618 409 676 443
rect 618 375 630 409
rect 664 375 676 409
rect 618 297 676 375
rect 712 479 793 497
rect 712 445 751 479
rect 785 445 793 479
rect 712 411 793 445
rect 712 377 751 411
rect 785 377 793 411
rect 712 343 793 377
rect 712 309 751 343
rect 785 309 793 343
rect 712 297 793 309
<< ndiffc >>
rect 35 131 69 165
rect 35 63 69 97
rect 215 67 249 101
rect 327 67 361 101
rect 527 63 561 97
rect 630 67 664 101
rect 751 131 785 165
rect 751 63 785 97
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 375 163 409
rect 223 451 257 485
rect 327 443 361 477
rect 426 443 460 477
rect 426 373 460 407
rect 536 443 570 477
rect 536 375 570 409
rect 630 443 664 477
rect 630 375 664 409
rect 751 445 785 479
rect 751 377 785 411
rect 751 309 785 343
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 373 497 409 523
rect 479 497 515 523
rect 582 497 618 523
rect 676 497 712 523
rect 81 282 117 297
rect 175 282 211 297
rect 373 282 409 297
rect 479 282 515 297
rect 582 282 618 297
rect 676 282 712 297
rect 79 265 119 282
rect 173 265 213 282
rect 371 265 411 282
rect 477 265 517 282
rect 580 265 620 282
rect 674 265 714 282
rect 55 249 119 265
rect 55 215 65 249
rect 99 215 119 249
rect 55 199 119 215
rect 89 177 119 199
rect 165 249 233 265
rect 165 215 179 249
rect 213 215 233 249
rect 165 199 233 215
rect 328 249 411 265
rect 328 215 338 249
rect 372 215 411 249
rect 328 199 411 215
rect 453 249 517 265
rect 453 215 463 249
rect 497 215 517 249
rect 453 199 517 215
rect 559 249 714 265
rect 559 215 569 249
rect 603 215 714 249
rect 559 199 714 215
rect 165 177 195 199
rect 381 177 411 199
rect 487 177 517 199
rect 590 177 620 199
rect 684 177 714 199
rect 89 21 119 47
rect 165 21 195 47
rect 381 21 411 47
rect 487 21 517 47
rect 590 21 620 47
rect 684 21 714 47
<< polycont >>
rect 65 215 99 249
rect 179 215 213 249
rect 338 215 372 249
rect 463 215 497 249
rect 569 215 603 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 19 485 273 493
rect 19 451 35 485
rect 69 459 223 485
rect 69 451 85 459
rect 207 451 223 459
rect 257 451 273 485
rect 311 477 382 527
rect 19 417 85 451
rect 311 443 327 477
rect 361 443 382 477
rect 426 477 476 493
rect 460 443 476 477
rect 19 383 35 417
rect 69 383 85 417
rect 19 349 85 383
rect 129 409 175 425
rect 163 407 175 409
rect 426 407 476 443
rect 163 375 426 407
rect 129 373 426 375
rect 460 373 476 407
rect 520 477 586 527
rect 520 443 536 477
rect 570 443 586 477
rect 520 409 586 443
rect 520 375 536 409
rect 570 375 586 409
rect 630 477 712 493
rect 664 443 712 477
rect 630 409 712 443
rect 664 375 712 409
rect 129 359 476 373
rect 630 357 712 375
rect 19 315 35 349
rect 69 325 85 349
rect 69 315 603 325
rect 19 291 603 315
rect 18 249 125 255
rect 18 215 65 249
rect 99 215 125 249
rect 163 249 268 257
rect 163 215 179 249
rect 19 165 119 170
rect 19 131 35 165
rect 69 131 119 165
rect 213 135 268 249
rect 305 249 388 257
rect 305 215 338 249
rect 372 215 388 249
rect 432 249 523 255
rect 432 215 463 249
rect 497 215 523 249
rect 569 249 603 291
rect 305 135 364 215
rect 569 181 603 215
rect 425 147 603 181
rect 19 97 119 131
rect 425 101 459 147
rect 648 117 712 357
rect 751 479 785 527
rect 751 411 785 445
rect 751 343 785 377
rect 751 289 785 309
rect 19 63 35 97
rect 69 63 119 97
rect 19 17 119 63
rect 174 67 215 101
rect 249 67 327 101
rect 361 67 459 101
rect 174 51 459 67
rect 501 97 577 113
rect 501 63 527 97
rect 561 63 577 97
rect 501 17 577 63
rect 630 101 712 117
rect 664 67 712 101
rect 630 51 712 67
rect 751 165 785 197
rect 751 97 785 131
rect 751 17 785 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel corelocali s 315 221 349 255 0 FreeSans 200 0 0 0 A1
port 1 nsew
flabel corelocali s 484 221 518 255 0 FreeSans 200 0 0 0 A2
port 2 nsew
flabel corelocali s 671 425 705 459 0 FreeSans 200 0 0 0 X
port 9 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 200 0 0 0 B2
port 4 nsew
flabel corelocali s 213 221 247 255 0 FreeSans 200 0 0 0 B1
port 3 nsew
flabel corelocali s 313 153 347 187 0 FreeSans 200 0 0 0 A1
port 1 nsew
flabel corelocali s 217 153 251 187 0 FreeSans 200 0 0 0 B1
port 3 nsew
flabel corelocali s 670 357 704 391 0 FreeSans 200 0 0 0 X
port 9 nsew
flabel corelocali s 670 221 704 255 0 FreeSans 200 0 0 0 X
port 9 nsew
flabel corelocali s 671 289 705 323 0 FreeSans 200 0 0 0 X
port 9 nsew
flabel corelocali s 670 85 704 119 0 FreeSans 200 0 0 0 X
port 9 nsew
flabel corelocali s 671 153 705 187 0 FreeSans 200 0 0 0 X
port 9 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
rlabel comment s 0 0 0 0 4 a22o_2
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1266726
string GDS_START 1259122
<< end >>
