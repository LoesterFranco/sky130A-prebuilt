magic
tech sky130A
magscale 1 2
timestamp 1604502741
<< locali >>
rect 365 405 431 471
rect 25 236 117 310
rect 397 356 431 405
rect 397 225 475 356
rect 1629 310 1703 414
rect 1629 74 1690 310
rect 2028 364 2101 596
rect 2067 226 2101 364
rect 2033 70 2101 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 23 378 89 596
rect 129 412 179 649
rect 219 559 269 596
rect 315 593 407 649
rect 800 593 866 649
rect 1007 559 1241 593
rect 219 525 1041 559
rect 23 344 185 378
rect 219 363 288 525
rect 465 441 543 491
rect 151 310 185 344
rect 151 202 220 310
rect 254 297 363 363
rect 254 214 320 297
rect 509 248 543 441
rect 577 457 865 491
rect 577 316 611 457
rect 645 350 728 413
rect 577 282 660 316
rect 509 214 574 248
rect 23 180 220 202
rect 23 146 506 180
rect 23 70 89 146
rect 125 17 202 112
rect 372 17 438 112
rect 472 85 506 146
rect 540 119 574 214
rect 610 119 660 282
rect 694 190 728 350
rect 831 392 865 457
rect 907 436 973 491
rect 831 326 895 392
rect 929 290 963 436
rect 1007 290 1041 525
rect 1075 358 1141 525
rect 1175 392 1241 559
rect 1320 475 1386 649
rect 1432 482 1498 596
rect 1539 516 1605 649
rect 1719 516 1785 649
rect 1432 448 1803 482
rect 1432 426 1585 448
rect 1275 358 1517 392
rect 1075 334 1517 358
rect 1075 324 1309 334
rect 762 224 963 290
rect 997 224 1055 290
rect 1089 234 1169 290
rect 694 156 963 190
rect 694 85 728 156
rect 472 51 728 85
rect 806 17 874 122
rect 929 106 963 156
rect 1089 106 1123 234
rect 1203 190 1237 324
rect 1551 300 1585 426
rect 1343 266 1585 300
rect 1343 234 1493 266
rect 1157 140 1237 190
rect 929 51 1248 106
rect 1331 17 1397 200
rect 1443 74 1493 234
rect 1529 17 1595 230
rect 1737 264 1803 448
rect 1847 326 1897 572
rect 1938 364 1988 649
rect 2135 364 2185 649
rect 1847 260 2033 326
rect 1724 17 1790 230
rect 1847 108 1902 260
rect 1947 17 1997 226
rect 2135 17 2185 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
<< metal1 >>
rect 0 683 2208 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 0 617 2208 649
rect 0 17 2208 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
rect 0 -49 2208 -17
<< labels >>
rlabel locali s 397 356 431 405 6 D
port 1 nsew signal input
rlabel locali s 397 225 475 356 6 D
port 1 nsew signal input
rlabel locali s 365 405 431 471 6 D
port 1 nsew signal input
rlabel locali s 1629 310 1703 414 6 Q
port 2 nsew signal output
rlabel locali s 1629 74 1690 310 6 Q
port 2 nsew signal output
rlabel locali s 2067 226 2101 364 6 Q_N
port 3 nsew signal output
rlabel locali s 2033 70 2101 226 6 Q_N
port 3 nsew signal output
rlabel locali s 2028 364 2101 596 6 Q_N
port 3 nsew signal output
rlabel locali s 25 236 117 310 6 CLK
port 4 nsew clock input
rlabel metal1 s 0 -49 2208 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 617 2208 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2208 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3007460
string GDS_START 2991724
<< end >>
