magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1104 561
rect 23 387 89 527
rect 125 351 159 437
rect 195 387 261 527
rect 297 351 347 437
rect 29 317 347 351
rect 29 157 126 317
rect 383 303 433 527
rect 479 199 541 305
rect 727 455 793 527
rect 895 455 961 527
rect 729 302 987 336
rect 729 255 764 302
rect 937 258 987 302
rect 685 202 764 255
rect 798 202 903 255
rect 937 211 1020 258
rect 29 123 347 157
rect 21 17 89 89
rect 195 17 261 89
rect 382 17 537 89
rect 651 17 717 89
rect 989 17 1045 177
rect 0 -17 1104 17
<< obsli1 >>
rect 491 459 693 493
rect 491 339 525 459
rect 160 199 441 265
rect 407 157 441 199
rect 575 168 609 425
rect 657 404 693 459
rect 827 404 861 493
rect 1006 404 1072 479
rect 657 370 1072 404
rect 657 289 693 370
rect 1021 292 1072 370
rect 575 157 873 168
rect 407 134 873 157
rect 407 123 609 134
rect 575 51 609 123
rect 817 81 873 134
<< metal1 >>
rect 0 496 1104 592
rect 0 -48 1104 48
<< labels >>
rlabel locali s 798 202 903 255 6 A1
port 1 nsew signal input
rlabel locali s 937 258 987 302 6 A2
port 2 nsew signal input
rlabel locali s 937 211 1020 258 6 A2
port 2 nsew signal input
rlabel locali s 729 302 987 336 6 A2
port 2 nsew signal input
rlabel locali s 729 255 764 302 6 A2
port 2 nsew signal input
rlabel locali s 685 202 764 255 6 A2
port 2 nsew signal input
rlabel locali s 479 199 541 305 6 B1
port 3 nsew signal input
rlabel locali s 297 351 347 437 6 X
port 4 nsew signal output
rlabel locali s 125 351 159 437 6 X
port 4 nsew signal output
rlabel locali s 29 317 347 351 6 X
port 4 nsew signal output
rlabel locali s 29 157 126 317 6 X
port 4 nsew signal output
rlabel locali s 29 123 347 157 6 X
port 4 nsew signal output
rlabel locali s 989 17 1045 177 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 651 17 717 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 382 17 537 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 195 17 261 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 21 17 89 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 1104 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1104 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 895 455 961 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 727 455 793 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 383 303 433 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 195 387 261 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 23 387 89 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 1104 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 1104 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1104 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 4028982
string GDS_START 4020818
<< end >>
