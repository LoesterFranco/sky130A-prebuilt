magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 614 704
<< pwell >>
rect 0 0 576 49
<< scnmos >>
rect 79 47 497 202
<< scpmos >>
rect 79 368 497 619
<< ndiff >>
rect 27 190 79 202
rect 27 156 35 190
rect 69 156 79 190
rect 27 93 79 156
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 497 190 549 202
rect 497 156 507 190
rect 541 156 549 190
rect 497 93 549 156
rect 497 59 507 93
rect 541 59 549 93
rect 497 47 549 59
<< pdiff >>
rect 27 607 79 619
rect 27 573 35 607
rect 69 573 79 607
rect 27 510 79 573
rect 27 476 35 510
rect 69 476 79 510
rect 27 414 79 476
rect 27 380 35 414
rect 69 380 79 414
rect 27 368 79 380
rect 497 607 549 619
rect 497 573 507 607
rect 541 573 549 607
rect 497 510 549 573
rect 497 476 507 510
rect 541 476 549 510
rect 497 414 549 476
rect 497 380 507 414
rect 541 380 549 414
rect 497 368 549 380
<< ndiffc >>
rect 35 156 69 190
rect 35 59 69 93
rect 507 156 541 190
rect 507 59 541 93
<< pdiffc >>
rect 35 573 69 607
rect 35 476 69 510
rect 35 380 69 414
rect 507 573 541 607
rect 507 476 541 510
rect 507 380 541 414
<< poly >>
rect 79 619 497 645
rect 79 342 497 368
rect 79 320 216 342
rect 79 286 98 320
rect 132 286 166 320
rect 200 286 216 320
rect 79 270 216 286
rect 292 284 497 300
rect 292 250 308 284
rect 342 250 376 284
rect 410 250 444 284
rect 478 250 497 284
rect 292 228 497 250
rect 79 202 497 228
rect 79 21 497 47
<< polycont >>
rect 98 286 132 320
rect 166 286 200 320
rect 308 250 342 284
rect 376 250 410 284
rect 444 250 478 284
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 24 607 552 649
rect 24 573 35 607
rect 69 573 507 607
rect 541 573 552 607
rect 24 510 552 573
rect 24 476 35 510
rect 69 476 507 510
rect 541 476 552 510
rect 24 414 552 476
rect 24 380 35 414
rect 69 380 507 414
rect 541 380 552 414
rect 24 354 552 380
rect 24 286 98 320
rect 132 286 166 320
rect 200 286 239 320
rect 24 216 239 286
rect 273 284 552 354
rect 273 250 308 284
rect 342 250 376 284
rect 410 250 444 284
rect 478 250 552 284
rect 24 190 552 216
rect 24 156 35 190
rect 69 156 507 190
rect 541 156 552 190
rect 24 93 552 156
rect 24 59 35 93
rect 69 59 507 93
rect 541 59 552 93
rect 24 17 552 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
flabel pwell s 0 0 576 49 0 FreeSans 200 0 0 0 VNB
port 2 nsew
flabel nbase s 0 617 576 666 0 FreeSans 200 0 0 0 VPB
port 3 nsew
rlabel comment s 0 0 0 0 4 decaphe_6
flabel metal1 s 0 617 576 666 0 FreeSans 200 0 0 0 VPWR
port 4 nsew
flabel metal1 s 0 0 576 49 0 FreeSans 200 0 0 0 VGND
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 576 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2461774
string GDS_START 2458398
<< end >>
