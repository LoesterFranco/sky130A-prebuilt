magic
tech sky130A
magscale 1 2
timestamp 1604502741
<< locali >>
rect 87 244 167 378
rect 201 236 267 310
rect 1153 364 1225 596
rect 1191 230 1225 364
rect 1159 74 1225 230
rect 1543 70 1610 596
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 19 543 88 585
rect 128 577 194 649
rect 19 509 352 543
rect 19 412 88 509
rect 19 210 53 412
rect 234 378 284 475
rect 318 446 352 509
rect 386 522 436 564
rect 476 556 542 649
rect 386 488 820 522
rect 898 509 1007 649
rect 386 480 436 488
rect 318 412 575 446
rect 234 344 466 378
rect 301 294 466 344
rect 509 294 575 412
rect 609 296 643 488
rect 677 364 711 454
rect 754 410 820 488
rect 1041 464 1107 596
rect 863 398 1107 464
rect 677 330 1007 364
rect 19 108 90 210
rect 301 202 335 294
rect 609 238 703 296
rect 126 17 192 202
rect 226 150 335 202
rect 369 204 703 238
rect 369 184 435 204
rect 756 170 790 330
rect 941 248 1007 330
rect 1041 330 1107 398
rect 1259 420 1309 649
rect 1041 264 1155 330
rect 1041 214 1075 264
rect 1344 330 1410 596
rect 1454 364 1504 649
rect 1344 264 1464 330
rect 226 116 616 150
rect 662 136 790 170
rect 226 70 335 116
rect 582 102 616 116
rect 471 17 548 82
rect 582 51 815 102
rect 904 17 970 212
rect 1004 70 1075 214
rect 1259 17 1309 230
rect 1344 112 1411 264
rect 1457 17 1507 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
rlabel locali s 87 244 167 378 6 D
port 1 nsew signal input
rlabel locali s 1191 230 1225 364 6 Q
port 2 nsew signal output
rlabel locali s 1159 74 1225 230 6 Q
port 2 nsew signal output
rlabel locali s 1153 364 1225 596 6 Q
port 2 nsew signal output
rlabel locali s 1543 70 1610 596 6 Q_N
port 3 nsew signal output
rlabel locali s 201 236 267 310 6 GATE
port 4 nsew clock input
rlabel metal1 s 0 -49 1632 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 617 1632 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 2169540
string GDS_START 2156844
<< end >>
