magic
tech sky130A
magscale 1 2
timestamp 1599588232
<< locali >>
rect 169 236 263 356
rect 297 290 363 356
rect 496 370 553 596
rect 519 236 553 370
rect 217 114 263 134
rect 21 51 263 114
rect 439 202 553 236
rect 439 96 505 202
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 23 424 89 570
rect 123 458 189 649
rect 223 424 280 570
rect 314 458 462 649
rect 23 390 448 424
rect 23 148 96 390
rect 414 336 448 390
rect 414 270 480 336
rect 339 17 405 236
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
rlabel locali s 217 114 263 134 6 A
port 1 nsew signal input
rlabel locali s 21 51 263 114 6 A
port 1 nsew signal input
rlabel locali s 169 236 263 356 6 B
port 2 nsew signal input
rlabel locali s 297 290 363 356 6 C
port 3 nsew signal input
rlabel locali s 519 236 553 370 6 X
port 4 nsew signal output
rlabel locali s 496 370 553 596 6 X
port 4 nsew signal output
rlabel locali s 439 202 553 236 6 X
port 4 nsew signal output
rlabel locali s 439 96 505 202 6 X
port 4 nsew signal output
rlabel metal1 s 0 -49 576 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 6 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 617 576 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 576 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3242864
string GDS_START 3236850
<< end >>
