magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1840 561
rect 103 427 169 527
rect 18 195 88 325
rect 271 333 336 490
rect 370 435 420 527
rect 103 17 169 93
rect 283 123 375 333
rect 798 441 864 527
rect 991 435 1065 527
rect 1388 435 1438 527
rect 761 153 919 203
rect 309 17 375 89
rect 895 17 961 109
rect 1542 451 1608 527
rect 1421 207 1529 281
rect 1676 299 1737 527
rect 1771 289 1822 465
rect 1341 17 1379 105
rect 1481 127 1529 207
rect 1780 159 1822 289
rect 1676 17 1737 109
rect 1771 53 1822 159
rect 0 -17 1840 17
<< obsli1 >>
rect 18 393 69 493
rect 18 391 168 393
rect 18 359 131 391
rect 122 357 131 359
rect 165 357 168 391
rect 122 161 168 357
rect 18 127 168 161
rect 203 255 237 493
rect 454 427 504 493
rect 547 427 683 493
rect 454 401 488 427
rect 409 367 488 401
rect 522 391 615 393
rect 18 69 69 127
rect 203 69 237 221
rect 409 95 443 367
rect 522 357 581 391
rect 522 315 615 357
rect 477 255 547 277
rect 477 221 489 255
rect 523 221 547 255
rect 477 153 547 221
rect 581 197 615 315
rect 649 271 683 427
rect 717 407 751 475
rect 898 407 932 475
rect 717 373 932 407
rect 1099 401 1133 493
rect 1180 425 1354 493
rect 1021 367 1133 401
rect 1021 339 1055 367
rect 755 305 1055 339
rect 1194 357 1205 391
rect 1239 357 1286 391
rect 1194 333 1286 357
rect 649 237 987 271
rect 581 153 652 197
rect 686 95 720 237
rect 953 201 987 237
rect 1021 167 1055 305
rect 409 61 508 95
rect 549 61 720 95
rect 1003 89 1055 167
rect 1093 331 1286 333
rect 1320 349 1354 425
rect 1472 417 1506 475
rect 1472 383 1632 417
rect 1093 299 1228 331
rect 1320 315 1564 349
rect 1093 141 1135 299
rect 1320 297 1354 315
rect 1169 255 1239 265
rect 1169 221 1205 255
rect 1169 141 1239 221
rect 1273 263 1354 297
rect 1273 107 1307 263
rect 1341 173 1385 229
rect 1598 265 1632 383
rect 1598 259 1746 265
rect 1341 139 1447 173
rect 1003 55 1073 89
rect 1117 51 1307 107
rect 1413 93 1447 139
rect 1563 199 1746 259
rect 1563 164 1628 199
rect 1563 93 1627 164
rect 1413 59 1627 93
<< obsli1c >>
rect 131 357 165 391
rect 203 221 237 255
rect 581 357 615 391
rect 489 221 523 255
rect 1205 357 1239 391
rect 1205 221 1239 255
<< metal1 >>
rect 0 496 1840 592
rect 1409 193 1467 256
rect 749 184 879 193
rect 1409 184 1527 193
rect 749 156 1527 184
rect 749 147 879 156
rect 1469 147 1527 156
rect 0 -48 1840 48
<< obsm1 >>
rect 119 391 177 397
rect 119 357 131 391
rect 165 388 177 391
rect 569 391 627 397
rect 569 388 581 391
rect 165 360 581 388
rect 165 357 177 360
rect 119 351 177 357
rect 569 357 581 360
rect 615 388 627 391
rect 1193 391 1251 397
rect 1193 388 1205 391
rect 615 360 1205 388
rect 615 357 627 360
rect 569 351 627 357
rect 1193 357 1205 360
rect 1239 357 1251 391
rect 1193 351 1251 357
rect 191 255 249 261
rect 191 221 203 255
rect 237 252 249 255
rect 477 255 535 261
rect 477 252 489 255
rect 237 224 489 252
rect 237 221 249 224
rect 191 215 249 221
rect 477 221 489 224
rect 523 252 535 255
rect 1193 255 1251 261
rect 1193 252 1205 255
rect 523 224 1205 252
rect 523 221 535 224
rect 477 215 535 221
rect 1193 221 1205 224
rect 1239 221 1251 255
rect 1193 215 1251 221
<< labels >>
rlabel locali s 283 123 375 333 6 D
port 1 nsew signal input
rlabel locali s 271 333 336 490 6 D
port 1 nsew signal input
rlabel locali s 1780 159 1822 289 6 Q
port 2 nsew signal output
rlabel locali s 1771 289 1822 465 6 Q
port 2 nsew signal output
rlabel locali s 1771 53 1822 159 6 Q
port 2 nsew signal output
rlabel locali s 761 153 919 203 6 RESET_B
port 3 nsew signal input
rlabel locali s 1481 127 1529 207 6 RESET_B
port 3 nsew signal input
rlabel locali s 1421 207 1529 281 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 1469 147 1527 156 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 1409 193 1467 256 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 1409 184 1527 193 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 749 184 879 193 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 749 156 1527 184 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 749 147 879 156 6 RESET_B
port 3 nsew signal input
rlabel locali s 18 195 88 325 6 CLK_N
port 4 nsew clock input
rlabel locali s 1676 17 1737 109 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 1341 17 1379 105 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 895 17 961 109 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 309 17 375 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 103 17 169 93 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 1840 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1840 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 1676 299 1737 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 1542 451 1608 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 1388 435 1438 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 991 435 1065 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 798 441 864 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 370 435 420 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 103 427 169 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 1840 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 1840 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1840 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3369420
string GDS_START 3354318
<< end >>
