magic
tech sky130A
magscale 1 2
timestamp 1599588209
<< nwell >>
rect -38 332 902 704
<< pwell >>
rect 0 0 864 49
<< scpmos >>
rect 86 368 116 536
rect 193 368 223 568
rect 386 368 416 568
rect 494 368 524 568
rect 608 368 638 568
rect 732 368 762 592
<< nmoslvt >>
rect 84 112 114 222
rect 196 74 226 222
rect 274 74 304 222
rect 413 74 443 222
rect 605 74 635 222
rect 748 74 778 222
<< ndiff >>
rect 27 184 84 222
rect 27 150 39 184
rect 73 150 84 184
rect 27 112 84 150
rect 114 210 196 222
rect 114 176 128 210
rect 162 176 196 210
rect 114 120 196 176
rect 114 112 146 120
rect 129 86 146 112
rect 180 86 196 120
rect 129 74 196 86
rect 226 74 274 222
rect 304 128 413 222
rect 304 94 341 128
rect 375 94 413 128
rect 304 74 413 94
rect 443 74 605 222
rect 635 146 748 222
rect 635 112 675 146
rect 709 112 748 146
rect 635 74 748 112
rect 778 210 835 222
rect 778 176 789 210
rect 823 176 835 210
rect 778 120 835 176
rect 778 86 789 120
rect 823 86 835 120
rect 778 74 835 86
<< pdiff >>
rect 663 580 732 592
rect 663 568 675 580
rect 134 536 193 568
rect 27 524 86 536
rect 27 490 39 524
rect 73 490 86 524
rect 27 429 86 490
rect 27 395 39 429
rect 73 395 86 429
rect 27 368 86 395
rect 116 519 193 536
rect 116 485 146 519
rect 180 485 193 519
rect 116 368 193 485
rect 223 368 386 568
rect 416 531 494 568
rect 416 497 429 531
rect 463 497 494 531
rect 416 414 494 497
rect 416 380 429 414
rect 463 380 494 414
rect 416 368 494 380
rect 524 368 608 568
rect 638 546 675 568
rect 709 546 732 580
rect 638 497 732 546
rect 638 463 675 497
rect 709 463 732 497
rect 638 414 732 463
rect 638 380 675 414
rect 709 380 732 414
rect 638 368 732 380
rect 762 580 821 592
rect 762 546 775 580
rect 809 546 821 580
rect 762 497 821 546
rect 762 463 775 497
rect 809 463 821 497
rect 762 414 821 463
rect 762 380 775 414
rect 809 380 821 414
rect 762 368 821 380
<< ndiffc >>
rect 39 150 73 184
rect 128 176 162 210
rect 146 86 180 120
rect 341 94 375 128
rect 675 112 709 146
rect 789 176 823 210
rect 789 86 823 120
<< pdiffc >>
rect 39 490 73 524
rect 39 395 73 429
rect 146 485 180 519
rect 429 497 463 531
rect 429 380 463 414
rect 675 546 709 580
rect 675 463 709 497
rect 675 380 709 414
rect 775 546 809 580
rect 775 463 809 497
rect 775 380 809 414
<< poly >>
rect 193 568 223 594
rect 386 568 416 594
rect 494 568 524 594
rect 608 568 638 594
rect 732 592 762 618
rect 86 536 116 562
rect 86 353 116 368
rect 193 353 223 368
rect 386 353 416 368
rect 494 353 524 368
rect 608 353 638 368
rect 732 353 762 368
rect 83 336 119 353
rect 190 336 226 353
rect 83 320 226 336
rect 83 286 117 320
rect 151 286 226 320
rect 383 310 419 353
rect 491 310 527 353
rect 605 330 641 353
rect 605 314 671 330
rect 729 326 765 353
rect 83 270 226 286
rect 84 222 114 270
rect 196 222 226 270
rect 269 294 335 310
rect 269 260 285 294
rect 319 260 335 294
rect 269 244 335 260
rect 377 294 443 310
rect 377 260 393 294
rect 427 260 443 294
rect 377 244 443 260
rect 491 294 557 310
rect 491 260 507 294
rect 541 260 557 294
rect 491 244 557 260
rect 605 280 621 314
rect 655 280 671 314
rect 605 264 671 280
rect 713 310 779 326
rect 713 276 729 310
rect 763 276 779 310
rect 274 222 304 244
rect 413 222 443 244
rect 605 222 635 264
rect 713 260 779 276
rect 748 222 778 260
rect 84 86 114 112
rect 196 48 226 74
rect 274 48 304 74
rect 413 48 443 74
rect 605 48 635 74
rect 748 48 778 74
<< polycont >>
rect 117 286 151 320
rect 285 260 319 294
rect 393 260 427 294
rect 507 260 541 294
rect 621 280 655 314
rect 729 276 763 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 23 524 89 540
rect 23 490 39 524
rect 73 490 89 524
rect 23 446 89 490
rect 130 519 196 649
rect 130 485 146 519
rect 180 485 196 519
rect 130 480 196 485
rect 230 581 625 615
rect 230 446 264 581
rect 23 429 264 446
rect 23 395 39 429
rect 73 412 264 429
rect 413 531 479 547
rect 413 497 429 531
rect 463 497 479 531
rect 413 414 479 497
rect 73 395 89 412
rect 23 390 89 395
rect 23 226 57 390
rect 413 380 429 414
rect 463 380 479 414
rect 413 378 479 380
rect 101 320 167 356
rect 101 286 117 320
rect 151 286 167 320
rect 101 270 167 286
rect 201 344 479 378
rect 23 184 89 226
rect 23 150 39 184
rect 73 150 89 184
rect 23 108 89 150
rect 125 210 167 226
rect 125 176 128 210
rect 162 176 167 210
rect 125 136 167 176
rect 201 204 235 344
rect 591 330 625 581
rect 659 580 725 649
rect 659 546 675 580
rect 709 546 725 580
rect 659 497 725 546
rect 659 463 675 497
rect 709 463 725 497
rect 659 414 725 463
rect 659 380 675 414
rect 709 380 725 414
rect 659 364 725 380
rect 759 580 847 596
rect 759 546 775 580
rect 809 546 847 580
rect 759 497 847 546
rect 759 463 775 497
rect 809 463 847 497
rect 759 414 847 463
rect 759 380 775 414
rect 809 380 847 414
rect 759 364 847 380
rect 591 314 671 330
rect 269 294 337 310
rect 269 260 285 294
rect 319 260 337 294
rect 269 244 337 260
rect 201 170 269 204
rect 125 120 201 136
rect 125 86 146 120
rect 180 86 201 120
rect 125 17 201 86
rect 235 128 269 170
rect 303 196 337 244
rect 377 294 455 310
rect 377 260 393 294
rect 427 260 455 294
rect 377 236 455 260
rect 491 294 557 310
rect 491 260 507 294
rect 541 260 557 294
rect 591 280 621 314
rect 655 280 671 314
rect 591 264 671 280
rect 705 310 779 326
rect 705 276 729 310
rect 763 276 779 310
rect 491 196 557 260
rect 705 260 779 276
rect 705 230 739 260
rect 303 162 557 196
rect 591 196 739 230
rect 813 226 847 364
rect 773 210 847 226
rect 591 128 625 196
rect 773 176 789 210
rect 823 176 847 210
rect 235 94 341 128
rect 375 94 625 128
rect 235 78 625 94
rect 659 146 725 162
rect 659 112 675 146
rect 709 112 725 146
rect 659 17 725 112
rect 773 120 847 176
rect 773 86 789 120
rect 823 86 847 120
rect 773 70 847 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel comment s 0 0 0 0 4 mux2_1
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 799 390 833 424 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 799 464 833 498 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 799 538 833 572 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 S
port 3 nsew
flabel corelocali s 415 242 449 276 0 FreeSans 340 0 0 0 A0
port 1 nsew
flabel corelocali s 511 168 545 202 0 FreeSans 340 0 0 0 A1
port 2 nsew
flabel corelocali s 511 242 545 276 0 FreeSans 340 0 0 0 A1
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 864 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1903020
string GDS_START 1896158
<< end >>
