magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 25 238 119 372
rect 313 310 455 392
rect 597 310 663 376
rect 775 370 846 596
rect 812 236 846 370
rect 409 51 562 134
rect 775 96 846 236
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 23 440 89 596
rect 123 474 189 649
rect 329 507 519 649
rect 223 470 292 492
rect 553 470 619 596
rect 23 406 189 440
rect 223 426 619 470
rect 155 376 189 406
rect 519 420 619 426
rect 667 420 733 649
rect 155 310 251 376
rect 155 204 189 310
rect 519 276 553 420
rect 707 276 778 336
rect 23 170 189 204
rect 262 270 778 276
rect 262 242 741 270
rect 23 70 81 170
rect 115 17 175 136
rect 262 120 328 242
rect 675 17 741 208
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel locali s 25 238 119 372 6 A_N
port 1 nsew signal input
rlabel locali s 313 310 455 392 6 B
port 2 nsew signal input
rlabel locali s 409 51 562 134 6 C
port 3 nsew signal input
rlabel locali s 597 310 663 376 6 D
port 4 nsew signal input
rlabel locali s 812 236 846 370 6 X
port 5 nsew signal output
rlabel locali s 775 370 846 596 6 X
port 5 nsew signal output
rlabel locali s 775 96 846 236 6 X
port 5 nsew signal output
rlabel metal1 s 0 -49 864 49 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 617 864 715 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3202740
string GDS_START 3194918
<< end >>
