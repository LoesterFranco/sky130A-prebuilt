magic
tech sky130A
magscale 1 2
timestamp 1604502741
<< locali >>
rect 21 236 87 310
rect 121 260 236 578
rect 270 390 446 596
rect 270 226 304 390
rect 338 270 455 356
rect 489 260 555 356
rect 270 192 553 226
rect 487 70 553 192
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 26 364 76 649
rect 482 390 548 649
rect 23 17 89 202
rect 125 158 175 226
rect 125 124 453 158
rect 125 70 175 124
rect 211 17 351 90
rect 387 70 453 124
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
rlabel locali s 21 236 87 310 6 A1
port 1 nsew signal input
rlabel locali s 121 260 236 578 6 A2
port 2 nsew signal input
rlabel locali s 338 270 455 356 6 A3
port 3 nsew signal input
rlabel locali s 489 260 555 356 6 B1
port 4 nsew signal input
rlabel locali s 487 70 553 192 6 Y
port 5 nsew signal output
rlabel locali s 270 390 446 596 6 Y
port 5 nsew signal output
rlabel locali s 270 226 304 390 6 Y
port 5 nsew signal output
rlabel locali s 270 192 553 226 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -49 576 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 576 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 576 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 700518
string GDS_START 694474
<< end >>
