magic
tech sky130A
magscale 1 2
timestamp 1604502710
<< nwell >>
rect -38 332 134 704
<< psubdiff >>
rect 31 205 65 229
rect 31 122 65 171
rect 31 64 65 88
<< nsubdiff >>
rect 31 578 65 602
rect 31 492 65 544
rect 31 434 65 458
<< psubdiffcont >>
rect 31 171 65 205
rect 31 88 65 122
<< nsubdiffcont >>
rect 31 544 65 578
rect 31 458 65 492
<< locali >>
rect 0 649 31 683
rect 65 649 96 683
rect 18 578 78 613
rect 18 544 31 578
rect 65 544 78 578
rect 18 498 78 544
rect 18 458 31 498
rect 65 458 78 498
rect 18 378 78 458
rect 18 205 78 288
rect 18 171 31 205
rect 65 171 78 205
rect 18 122 78 171
rect 18 88 31 122
rect 65 88 78 122
rect 18 17 78 88
rect 0 -17 31 17
rect 65 -17 96 17
<< viali >>
rect 31 649 65 683
rect 31 492 65 498
rect 31 464 65 492
rect 31 -17 65 17
<< metal1 >>
rect 0 683 96 715
rect 0 649 31 683
rect 65 649 96 683
rect 0 617 96 649
rect 16 498 80 507
rect 16 464 31 498
rect 65 464 80 498
rect 16 455 80 464
rect 0 17 96 49
rect 0 -17 31 17
rect 65 -17 96 17
rect 0 -49 96 -17
<< labels >>
rlabel comment s 0 0 0 0 4 tapvgnd2_1
flabel metal1 s 31 464 65 498 0 FreeSans 340 0 0 0 VPB
port 2 nsew
flabel metal1 s 0 617 96 666 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel metal1 s 0 0 96 49 0 FreeSans 200 0 0 0 VGND
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 96 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 458216
string GDS_START 456312
<< end >>
