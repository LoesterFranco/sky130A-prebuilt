magic
tech sky130A
magscale 1 2
timestamp 1601050056
<< nwell >>
rect -38 332 1766 704
<< pwell >>
rect 0 0 1728 49
<< scpmos >>
rect 83 368 119 592
rect 173 368 209 592
rect 398 508 434 592
rect 505 429 541 513
rect 611 504 647 588
rect 695 504 731 588
rect 831 424 867 592
rect 986 424 1022 592
rect 1092 508 1128 592
rect 1217 508 1253 592
rect 1418 368 1454 568
rect 1519 368 1555 592
rect 1609 368 1645 592
<< nmoslvt >>
rect 84 74 114 222
rect 202 74 232 222
rect 497 119 527 203
rect 583 119 613 203
rect 678 101 708 185
rect 756 101 786 185
rect 924 75 954 185
rect 1010 75 1040 185
rect 1142 124 1172 208
rect 1220 124 1250 208
rect 1418 74 1448 184
rect 1528 74 1558 222
rect 1614 74 1644 222
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 131 202 222
rect 114 97 125 131
rect 159 97 202 131
rect 114 74 202 97
rect 232 189 307 222
rect 232 155 261 189
rect 295 155 307 189
rect 232 74 307 155
rect 385 119 497 203
rect 527 180 583 203
rect 527 146 538 180
rect 572 146 583 180
rect 527 119 583 146
rect 613 185 663 203
rect 1092 185 1142 208
rect 613 173 678 185
rect 613 139 628 173
rect 662 139 678 173
rect 613 119 678 139
rect 385 112 448 119
rect 385 78 399 112
rect 433 78 448 112
rect 628 101 678 119
rect 708 101 756 185
rect 786 101 924 185
rect 385 66 448 78
rect 801 88 924 101
rect 801 54 813 88
rect 847 75 924 88
rect 954 171 1010 185
rect 954 137 965 171
rect 999 137 1010 171
rect 954 75 1010 137
rect 1040 173 1142 185
rect 1040 139 1081 173
rect 1115 139 1142 173
rect 1040 124 1142 139
rect 1172 124 1220 208
rect 1250 183 1307 208
rect 1478 184 1528 222
rect 1250 149 1261 183
rect 1295 149 1307 183
rect 1250 124 1307 149
rect 1361 146 1418 184
rect 1040 75 1090 124
rect 1361 112 1373 146
rect 1407 112 1418 146
rect 847 54 859 75
rect 801 42 859 54
rect 1361 74 1418 112
rect 1448 120 1528 184
rect 1448 86 1464 120
rect 1498 86 1528 120
rect 1448 74 1528 86
rect 1558 210 1614 222
rect 1558 176 1569 210
rect 1603 176 1614 210
rect 1558 120 1614 176
rect 1558 86 1569 120
rect 1603 86 1614 120
rect 1558 74 1614 86
rect 1644 210 1701 222
rect 1644 176 1655 210
rect 1689 176 1701 210
rect 1644 120 1701 176
rect 1644 86 1655 120
rect 1689 86 1701 120
rect 1644 74 1701 86
<< pdiff >>
rect 319 627 383 639
rect 319 593 334 627
rect 368 593 383 627
rect 746 627 816 639
rect 319 592 383 593
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 510 83 546
rect 27 476 39 510
rect 73 476 83 510
rect 27 440 83 476
rect 27 406 39 440
rect 73 406 83 440
rect 27 368 83 406
rect 119 580 173 592
rect 119 546 129 580
rect 163 546 173 580
rect 119 508 173 546
rect 119 474 129 508
rect 163 474 173 508
rect 119 368 173 474
rect 209 580 265 592
rect 209 546 219 580
rect 253 546 265 580
rect 209 497 265 546
rect 319 508 398 592
rect 434 513 484 592
rect 746 593 764 627
rect 798 593 816 627
rect 746 592 816 593
rect 746 588 831 592
rect 561 513 611 588
rect 434 508 505 513
rect 209 463 219 497
rect 253 463 265 497
rect 209 414 265 463
rect 209 380 219 414
rect 253 380 265 414
rect 449 475 505 508
rect 449 441 461 475
rect 495 441 505 475
rect 449 429 505 441
rect 541 504 611 513
rect 647 504 695 588
rect 731 504 831 588
rect 541 488 596 504
rect 541 454 551 488
rect 585 454 596 488
rect 541 429 596 454
rect 209 368 265 380
rect 781 424 831 504
rect 867 475 986 592
rect 867 441 878 475
rect 912 441 986 475
rect 867 424 986 441
rect 1022 516 1092 592
rect 1022 482 1032 516
rect 1066 508 1092 516
rect 1128 508 1217 592
rect 1253 567 1308 592
rect 1469 568 1519 592
rect 1253 533 1263 567
rect 1297 533 1308 567
rect 1253 508 1308 533
rect 1362 556 1418 568
rect 1362 522 1374 556
rect 1408 522 1418 556
rect 1066 482 1077 508
rect 1022 424 1077 482
rect 1362 485 1418 522
rect 1362 451 1374 485
rect 1408 451 1418 485
rect 1362 414 1418 451
rect 1362 380 1374 414
rect 1408 380 1418 414
rect 1362 368 1418 380
rect 1454 556 1519 568
rect 1454 522 1464 556
rect 1498 522 1519 556
rect 1454 456 1519 522
rect 1454 422 1464 456
rect 1498 422 1519 456
rect 1454 368 1519 422
rect 1555 580 1609 592
rect 1555 546 1565 580
rect 1599 546 1609 580
rect 1555 512 1609 546
rect 1555 478 1565 512
rect 1599 478 1609 512
rect 1555 444 1609 478
rect 1555 410 1565 444
rect 1599 410 1609 444
rect 1555 368 1609 410
rect 1645 580 1701 592
rect 1645 546 1655 580
rect 1689 546 1701 580
rect 1645 497 1701 546
rect 1645 463 1655 497
rect 1689 463 1701 497
rect 1645 414 1701 463
rect 1645 380 1655 414
rect 1689 380 1701 414
rect 1645 368 1701 380
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 125 97 159 131
rect 261 155 295 189
rect 538 146 572 180
rect 628 139 662 173
rect 399 78 433 112
rect 813 54 847 88
rect 965 137 999 171
rect 1081 139 1115 173
rect 1261 149 1295 183
rect 1373 112 1407 146
rect 1464 86 1498 120
rect 1569 176 1603 210
rect 1569 86 1603 120
rect 1655 176 1689 210
rect 1655 86 1689 120
<< pdiffc >>
rect 334 593 368 627
rect 39 546 73 580
rect 39 476 73 510
rect 39 406 73 440
rect 129 546 163 580
rect 129 474 163 508
rect 219 546 253 580
rect 764 593 798 627
rect 219 463 253 497
rect 219 380 253 414
rect 461 441 495 475
rect 551 454 585 488
rect 878 441 912 475
rect 1032 482 1066 516
rect 1263 533 1297 567
rect 1374 522 1408 556
rect 1374 451 1408 485
rect 1374 380 1408 414
rect 1464 522 1498 556
rect 1464 422 1498 456
rect 1565 546 1599 580
rect 1565 478 1599 512
rect 1565 410 1599 444
rect 1655 546 1689 580
rect 1655 463 1689 497
rect 1655 380 1689 414
<< poly >>
rect 83 592 119 618
rect 173 592 209 618
rect 398 592 434 618
rect 611 588 647 614
rect 695 588 731 614
rect 831 592 867 618
rect 986 592 1022 618
rect 1092 592 1128 618
rect 1217 592 1253 618
rect 505 513 541 539
rect 398 476 434 508
rect 345 460 434 476
rect 345 426 361 460
rect 395 426 434 460
rect 345 410 434 426
rect 505 368 541 429
rect 611 417 647 504
rect 695 489 731 504
rect 695 459 766 489
rect 611 401 694 417
rect 611 381 644 401
rect 83 326 119 368
rect 35 310 119 326
rect 173 310 209 368
rect 280 338 541 368
rect 583 367 644 381
rect 678 367 694 401
rect 583 351 694 367
rect 280 320 352 338
rect 35 276 51 310
rect 85 276 119 310
rect 35 260 119 276
rect 161 294 232 310
rect 161 260 177 294
rect 211 260 232 294
rect 280 286 296 320
rect 330 286 352 320
rect 280 270 352 286
rect 84 222 114 260
rect 161 244 232 260
rect 202 222 232 244
rect 84 48 114 74
rect 202 48 232 74
rect 322 51 352 270
rect 400 280 466 296
rect 400 246 416 280
rect 450 260 466 280
rect 450 246 527 260
rect 400 230 527 246
rect 497 203 527 230
rect 583 203 613 351
rect 736 283 766 459
rect 1418 568 1454 594
rect 1519 592 1555 618
rect 1609 592 1645 618
rect 1092 476 1128 508
rect 1092 460 1175 476
rect 1092 426 1125 460
rect 1159 426 1175 460
rect 831 391 867 424
rect 808 375 929 391
rect 808 341 824 375
rect 858 341 929 375
rect 986 368 1022 424
rect 1092 410 1175 426
rect 1217 448 1253 508
rect 1217 432 1283 448
rect 1217 398 1233 432
rect 1267 398 1283 432
rect 986 344 1172 368
rect 808 325 929 341
rect 992 338 1172 344
rect 736 267 851 283
rect 736 253 801 267
rect 756 233 801 253
rect 835 233 851 267
rect 756 217 851 233
rect 899 230 929 325
rect 1010 280 1083 296
rect 1010 246 1033 280
rect 1067 246 1083 280
rect 1010 230 1083 246
rect 678 185 708 211
rect 756 185 786 217
rect 899 200 954 230
rect 924 185 954 200
rect 1010 185 1040 230
rect 1142 208 1172 338
rect 1217 364 1283 398
rect 1217 330 1233 364
rect 1267 330 1283 364
rect 1217 314 1283 330
rect 1220 208 1250 314
rect 1418 304 1454 368
rect 1519 336 1555 368
rect 1609 336 1645 368
rect 1382 288 1454 304
rect 1382 254 1398 288
rect 1432 254 1454 288
rect 1496 320 1644 336
rect 1496 286 1512 320
rect 1546 286 1644 320
rect 1496 270 1644 286
rect 1382 238 1454 254
rect 497 93 527 119
rect 583 93 613 119
rect 678 51 708 101
rect 756 75 786 101
rect 322 21 708 51
rect 1418 184 1448 238
rect 1528 222 1558 270
rect 1614 222 1644 270
rect 1142 102 1172 124
rect 1112 86 1178 102
rect 1220 98 1250 124
rect 924 49 954 75
rect 1010 49 1040 75
rect 1112 52 1128 86
rect 1162 52 1178 86
rect 1112 36 1178 52
rect 1418 48 1448 74
rect 1528 48 1558 74
rect 1614 48 1644 74
<< polycont >>
rect 361 426 395 460
rect 644 367 678 401
rect 51 276 85 310
rect 177 260 211 294
rect 296 286 330 320
rect 416 246 450 280
rect 1125 426 1159 460
rect 824 341 858 375
rect 1233 398 1267 432
rect 801 233 835 267
rect 1033 246 1067 280
rect 1233 330 1267 364
rect 1398 254 1432 288
rect 1512 286 1546 320
rect 1128 52 1162 86
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 23 580 89 596
rect 23 546 39 580
rect 73 546 89 580
rect 23 510 89 546
rect 23 476 39 510
rect 73 476 89 510
rect 23 440 89 476
rect 129 580 163 649
rect 315 627 387 649
rect 129 508 163 546
rect 129 458 163 474
rect 203 580 269 596
rect 315 593 334 627
rect 368 593 387 627
rect 742 627 820 649
rect 742 593 764 627
rect 798 593 820 627
rect 203 546 219 580
rect 253 559 269 580
rect 421 559 708 585
rect 964 581 1175 615
rect 964 559 998 581
rect 253 551 998 559
rect 253 546 455 551
rect 203 525 455 546
rect 674 525 998 551
rect 203 497 295 525
rect 203 463 219 497
rect 253 463 295 497
rect 23 406 39 440
rect 73 424 89 440
rect 73 406 169 424
rect 23 390 169 406
rect 25 310 101 356
rect 25 276 51 310
rect 85 276 101 310
rect 25 260 101 276
rect 135 310 169 390
rect 203 414 295 463
rect 203 380 219 414
rect 253 380 295 414
rect 345 460 411 476
rect 345 426 361 460
rect 395 426 411 460
rect 345 410 411 426
rect 203 344 295 380
rect 261 320 343 344
rect 135 294 227 310
rect 135 260 177 294
rect 211 260 227 294
rect 135 226 227 260
rect 23 210 227 226
rect 23 176 39 210
rect 73 192 227 210
rect 23 120 73 176
rect 23 86 39 120
rect 23 70 73 86
rect 109 131 159 158
rect 109 97 125 131
rect 109 17 159 97
rect 193 85 227 192
rect 261 286 296 320
rect 330 286 343 320
rect 261 270 343 286
rect 377 296 411 410
rect 445 475 511 491
rect 445 441 461 475
rect 495 441 511 475
rect 445 364 511 441
rect 551 488 591 517
rect 585 485 591 488
rect 585 454 827 485
rect 551 451 827 454
rect 551 425 591 451
rect 445 330 523 364
rect 377 280 455 296
rect 261 189 295 270
rect 377 246 416 280
rect 450 246 455 280
rect 377 230 455 246
rect 489 264 523 330
rect 557 332 591 425
rect 628 401 708 417
rect 628 367 644 401
rect 678 367 708 401
rect 628 366 708 367
rect 557 298 640 332
rect 489 230 572 264
rect 261 119 295 155
rect 329 162 504 196
rect 329 85 363 162
rect 193 51 363 85
rect 397 112 436 128
rect 397 78 399 112
rect 433 78 436 112
rect 397 17 436 78
rect 470 85 504 162
rect 538 180 572 230
rect 538 119 572 146
rect 606 189 640 298
rect 674 291 708 366
rect 793 391 827 451
rect 861 475 930 491
rect 861 441 878 475
rect 912 441 930 475
rect 861 425 930 441
rect 793 375 862 391
rect 793 341 824 375
rect 858 341 862 375
rect 793 325 862 341
rect 674 257 751 291
rect 896 283 930 425
rect 606 173 683 189
rect 606 139 628 173
rect 662 139 683 173
rect 606 123 683 139
rect 717 172 751 257
rect 785 267 930 283
rect 964 308 998 525
rect 1032 516 1066 547
rect 1032 376 1066 482
rect 1109 460 1175 581
rect 1247 567 1313 649
rect 1247 533 1263 567
rect 1297 533 1313 567
rect 1247 504 1313 533
rect 1358 556 1408 572
rect 1358 522 1374 556
rect 1109 426 1125 460
rect 1159 426 1175 460
rect 1358 485 1408 522
rect 1358 451 1374 485
rect 1109 410 1175 426
rect 1217 432 1283 448
rect 1217 398 1233 432
rect 1267 398 1283 432
rect 1032 342 1151 376
rect 964 280 1083 308
rect 964 274 1033 280
rect 785 233 801 267
rect 835 240 930 267
rect 1017 246 1033 274
rect 1067 246 1083 280
rect 835 233 983 240
rect 785 206 983 233
rect 1017 230 1083 246
rect 1117 280 1151 342
rect 1217 372 1283 398
rect 1358 414 1408 451
rect 1358 380 1374 414
rect 1448 556 1514 649
rect 1448 522 1464 556
rect 1498 522 1514 556
rect 1448 456 1514 522
rect 1448 422 1464 456
rect 1498 422 1514 456
rect 1448 406 1514 422
rect 1549 580 1621 596
rect 1549 546 1565 580
rect 1599 546 1621 580
rect 1549 512 1621 546
rect 1549 478 1565 512
rect 1599 478 1621 512
rect 1549 444 1621 478
rect 1549 410 1565 444
rect 1599 410 1621 444
rect 1549 406 1621 410
rect 1358 372 1408 380
rect 1217 364 1553 372
rect 1217 330 1233 364
rect 1267 338 1553 364
rect 1267 330 1283 338
rect 1217 314 1283 330
rect 1485 320 1553 338
rect 1382 288 1448 304
rect 1382 280 1398 288
rect 1117 254 1398 280
rect 1432 254 1448 288
rect 1117 246 1448 254
rect 949 189 983 206
rect 1117 189 1151 246
rect 1382 238 1448 246
rect 1485 286 1512 320
rect 1546 286 1553 320
rect 1485 270 1553 286
rect 717 138 915 172
rect 717 85 751 138
rect 470 51 751 85
rect 797 88 847 104
rect 797 54 813 88
rect 797 17 847 54
rect 881 85 915 138
rect 949 171 1015 189
rect 949 137 965 171
rect 999 137 1015 171
rect 1049 173 1151 189
rect 1049 139 1081 173
rect 1115 139 1151 173
rect 1245 183 1311 212
rect 1485 204 1519 270
rect 1587 226 1621 406
rect 1655 580 1705 649
rect 1689 546 1705 580
rect 1655 497 1705 546
rect 1689 463 1705 497
rect 1655 414 1705 463
rect 1689 380 1705 414
rect 1655 364 1705 380
rect 1245 149 1261 183
rect 1295 149 1311 183
rect 949 119 1015 137
rect 1112 86 1178 102
rect 1112 85 1128 86
rect 881 52 1128 85
rect 1162 52 1178 86
rect 881 51 1178 52
rect 1245 17 1311 149
rect 1357 170 1519 204
rect 1553 210 1621 226
rect 1553 176 1569 210
rect 1603 176 1621 210
rect 1357 146 1423 170
rect 1357 112 1373 146
rect 1407 112 1423 146
rect 1357 70 1423 112
rect 1460 120 1519 136
rect 1460 86 1464 120
rect 1498 86 1519 120
rect 1460 17 1519 86
rect 1553 120 1621 176
rect 1553 86 1569 120
rect 1603 86 1621 120
rect 1553 70 1621 86
rect 1655 210 1705 226
rect 1689 176 1705 210
rect 1655 120 1705 176
rect 1689 86 1705 120
rect 1655 17 1705 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
<< metal1 >>
rect 0 683 1728 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 0 617 1728 649
rect 0 17 1728 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
rect 0 -49 1728 -17
<< labels >>
flabel pwell s 0 0 1728 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 0 617 1728 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
rlabel comment s 0 0 0 0 4 dfxtp_2
flabel metal1 s 0 617 1728 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 1728 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 1567 464 1601 498 0 FreeSans 340 0 0 0 Q
port 7 nsew
flabel corelocali s 1567 538 1601 572 0 FreeSans 340 0 0 0 Q
port 7 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 415 242 449 276 0 FreeSans 340 0 0 0 D
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 1728 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 2926764
string GDS_START 2913780
<< end >>
