magic
tech sky130A
magscale 1 2
timestamp 1601050056
<< nwell >>
rect -38 332 710 704
<< pwell >>
rect 0 0 672 49
<< scpmos >>
rect 83 368 119 592
rect 183 368 219 592
rect 273 368 309 592
rect 369 368 405 592
rect 463 368 499 592
rect 553 368 589 592
<< nmoslvt >>
rect 84 74 114 222
rect 291 74 321 222
rect 391 74 421 222
<< ndiff >>
rect 27 202 84 222
rect 27 168 39 202
rect 73 168 84 202
rect 27 120 84 168
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 120 291 222
rect 114 86 139 120
rect 173 86 246 120
rect 280 86 291 120
rect 114 74 291 86
rect 321 194 391 222
rect 321 160 346 194
rect 380 160 391 194
rect 321 120 391 160
rect 321 86 346 120
rect 380 86 391 120
rect 321 74 391 86
rect 421 210 492 222
rect 421 176 446 210
rect 480 176 492 210
rect 421 120 492 176
rect 421 86 446 120
rect 480 86 492 120
rect 421 74 492 86
<< pdiff >>
rect 27 582 83 592
rect 27 548 39 582
rect 73 548 83 582
rect 27 514 83 548
rect 27 480 39 514
rect 73 480 83 514
rect 27 446 83 480
rect 27 412 39 446
rect 73 412 83 446
rect 27 368 83 412
rect 119 547 183 592
rect 119 513 139 547
rect 173 513 183 547
rect 119 479 183 513
rect 119 445 139 479
rect 173 445 183 479
rect 119 411 183 445
rect 119 377 139 411
rect 173 377 183 411
rect 119 368 183 377
rect 219 580 273 592
rect 219 546 229 580
rect 263 546 273 580
rect 219 497 273 546
rect 219 463 229 497
rect 263 463 273 497
rect 219 414 273 463
rect 219 380 229 414
rect 263 380 273 414
rect 219 368 273 380
rect 309 582 369 592
rect 309 548 319 582
rect 353 548 369 582
rect 309 514 369 548
rect 309 480 319 514
rect 353 480 369 514
rect 309 446 369 480
rect 309 412 319 446
rect 353 412 369 446
rect 309 368 369 412
rect 405 582 463 592
rect 405 548 419 582
rect 453 548 463 582
rect 405 514 463 548
rect 405 480 419 514
rect 453 480 463 514
rect 405 368 463 480
rect 499 582 553 592
rect 499 548 509 582
rect 543 548 553 582
rect 499 514 553 548
rect 499 480 509 514
rect 543 480 553 514
rect 499 446 553 480
rect 499 412 509 446
rect 543 412 553 446
rect 499 368 553 412
rect 589 580 645 592
rect 589 546 599 580
rect 633 546 645 580
rect 589 497 645 546
rect 589 463 599 497
rect 633 463 645 497
rect 589 414 645 463
rect 589 380 599 414
rect 633 380 645 414
rect 589 368 645 380
<< ndiffc >>
rect 39 168 73 202
rect 39 86 73 120
rect 139 86 173 120
rect 246 86 280 120
rect 346 160 380 194
rect 346 86 380 120
rect 446 176 480 210
rect 446 86 480 120
<< pdiffc >>
rect 39 548 73 582
rect 39 480 73 514
rect 39 412 73 446
rect 139 513 173 547
rect 139 445 173 479
rect 139 377 173 411
rect 229 546 263 580
rect 229 463 263 497
rect 229 380 263 414
rect 319 548 353 582
rect 319 480 353 514
rect 319 412 353 446
rect 419 548 453 582
rect 419 480 453 514
rect 509 548 543 582
rect 509 480 543 514
rect 509 412 543 446
rect 599 546 633 580
rect 599 463 633 497
rect 599 380 633 414
<< poly >>
rect 83 592 119 618
rect 183 592 219 618
rect 273 592 309 618
rect 369 592 405 618
rect 463 592 499 618
rect 553 592 589 618
rect 83 352 119 368
rect 183 352 219 368
rect 83 322 219 352
rect 129 294 219 322
rect 273 310 309 368
rect 129 274 145 294
rect 84 260 145 274
rect 179 260 219 294
rect 84 244 219 260
rect 261 294 327 310
rect 261 260 277 294
rect 311 260 327 294
rect 261 244 327 260
rect 369 267 405 368
rect 463 267 499 368
rect 553 345 589 368
rect 553 315 615 345
rect 585 310 615 315
rect 585 294 651 310
rect 84 222 114 244
rect 291 222 321 244
rect 369 237 537 267
rect 585 260 601 294
rect 635 260 651 294
rect 585 244 651 260
rect 391 222 421 237
rect 507 196 537 237
rect 507 180 596 196
rect 507 146 546 180
rect 580 146 596 180
rect 507 112 596 146
rect 507 78 546 112
rect 580 78 596 112
rect 84 48 114 74
rect 291 48 321 74
rect 391 48 421 74
rect 507 62 596 78
<< polycont >>
rect 145 260 179 294
rect 277 260 311 294
rect 601 260 635 294
rect 546 146 580 180
rect 546 78 580 112
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 23 582 263 615
rect 23 548 39 582
rect 73 581 263 582
rect 73 548 89 581
rect 23 514 89 548
rect 229 580 263 581
rect 23 480 39 514
rect 73 480 89 514
rect 23 446 89 480
rect 23 412 39 446
rect 73 412 89 446
rect 123 513 139 547
rect 173 513 189 547
rect 123 479 189 513
rect 123 445 139 479
rect 173 445 189 479
rect 123 411 189 445
rect 123 378 139 411
rect 23 377 139 378
rect 173 377 189 411
rect 23 344 189 377
rect 229 497 263 546
rect 229 414 263 463
rect 303 582 369 598
rect 303 548 319 582
rect 353 548 369 582
rect 303 514 369 548
rect 303 480 319 514
rect 353 480 369 514
rect 403 582 469 649
rect 403 548 419 582
rect 453 548 469 582
rect 403 514 469 548
rect 403 480 419 514
rect 453 480 469 514
rect 503 582 559 598
rect 503 548 509 582
rect 543 548 559 582
rect 503 514 559 548
rect 503 480 509 514
rect 543 480 559 514
rect 303 446 369 480
rect 503 446 559 480
rect 303 412 319 446
rect 353 412 509 446
rect 543 412 559 446
rect 593 580 649 596
rect 593 546 599 580
rect 633 546 649 580
rect 593 497 649 546
rect 593 463 599 497
rect 633 463 649 497
rect 593 414 649 463
rect 229 378 263 380
rect 593 380 599 414
rect 633 380 649 414
rect 593 378 649 380
rect 229 344 649 378
rect 23 202 71 344
rect 121 294 195 310
rect 121 260 145 294
rect 179 260 195 294
rect 121 236 195 260
rect 261 294 651 310
rect 261 260 277 294
rect 311 276 601 294
rect 311 260 327 276
rect 261 244 327 260
rect 585 260 601 276
rect 635 260 651 294
rect 585 236 651 260
rect 430 210 496 226
rect 330 202 396 210
rect 23 168 39 202
rect 73 194 396 202
rect 73 168 346 194
rect 23 120 89 168
rect 330 160 346 168
rect 380 160 396 194
rect 23 86 39 120
rect 73 86 89 120
rect 23 70 89 86
rect 123 120 296 130
rect 123 86 139 120
rect 173 86 246 120
rect 280 86 296 120
rect 123 17 296 86
rect 330 120 396 160
rect 330 86 346 120
rect 380 86 396 120
rect 330 70 396 86
rect 430 176 446 210
rect 480 176 496 210
rect 430 120 496 176
rect 430 86 446 120
rect 480 86 496 120
rect 430 17 496 86
rect 530 180 647 196
rect 530 146 546 180
rect 580 146 647 180
rect 530 112 647 146
rect 530 78 546 112
rect 580 78 647 112
rect 530 62 647 78
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
rlabel comment s 0 0 0 0 4 nor3_2
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 31 94 65 128 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 31 168 65 202 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 607 94 641 128 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 607 242 641 276 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 127 242 161 276 0 FreeSans 340 0 0 0 C
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 672 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1533656
string GDS_START 1526970
<< end >>
