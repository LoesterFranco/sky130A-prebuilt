magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 1382 704
<< pwell >>
rect 0 0 1344 49
<< scnmos >>
rect 84 115 114 225
rect 202 114 232 262
rect 456 74 486 222
rect 625 79 655 207
rect 703 79 733 207
rect 841 139 871 223
rect 919 139 949 223
rect 1031 95 1061 223
rect 1229 74 1259 222
<< pmoshvt >>
rect 87 419 117 587
rect 187 419 217 587
rect 428 392 458 560
rect 555 392 585 592
rect 639 392 669 592
rect 782 508 812 592
rect 866 508 896 592
rect 1026 392 1056 592
rect 1228 368 1258 592
<< ndiff >>
rect 152 225 202 262
rect 27 173 84 225
rect 27 139 39 173
rect 73 139 84 173
rect 27 115 84 139
rect 114 115 202 225
rect 129 114 202 115
rect 232 250 289 262
rect 232 216 243 250
rect 277 216 289 250
rect 232 114 289 216
rect 399 189 456 222
rect 399 155 411 189
rect 445 155 456 189
rect 129 82 187 114
rect 129 48 141 82
rect 175 48 187 82
rect 399 74 456 155
rect 486 207 536 222
rect 791 207 841 223
rect 486 195 625 207
rect 486 161 579 195
rect 613 161 625 195
rect 486 125 625 161
rect 486 91 579 125
rect 613 91 625 125
rect 486 79 625 91
rect 655 79 703 207
rect 733 195 841 207
rect 733 161 771 195
rect 805 161 841 195
rect 733 139 841 161
rect 871 139 919 223
rect 949 211 1031 223
rect 949 177 986 211
rect 1020 177 1031 211
rect 949 141 1031 177
rect 949 139 986 141
rect 733 79 783 139
rect 486 74 536 79
rect 974 107 986 139
rect 1020 107 1031 141
rect 974 95 1031 107
rect 1061 211 1118 223
rect 1061 177 1072 211
rect 1106 177 1118 211
rect 1061 141 1118 177
rect 1061 107 1072 141
rect 1106 107 1118 141
rect 1061 95 1118 107
rect 1172 210 1229 222
rect 1172 176 1184 210
rect 1218 176 1229 210
rect 1172 120 1229 176
rect 1172 86 1184 120
rect 1218 86 1229 120
rect 1172 74 1229 86
rect 1259 120 1317 222
rect 1259 86 1270 120
rect 1304 86 1317 120
rect 1259 74 1317 86
rect 129 36 187 48
<< pdiff >>
rect 476 606 537 618
rect 28 575 87 587
rect 28 541 40 575
rect 74 541 87 575
rect 28 465 87 541
rect 28 431 40 465
rect 74 431 87 465
rect 28 419 87 431
rect 117 575 187 587
rect 117 541 140 575
rect 174 541 187 575
rect 117 465 187 541
rect 117 431 140 465
rect 174 431 187 465
rect 117 419 187 431
rect 217 575 293 587
rect 217 541 247 575
rect 281 541 293 575
rect 476 572 489 606
rect 523 592 537 606
rect 523 572 555 592
rect 476 560 555 572
rect 217 465 293 541
rect 217 431 247 465
rect 281 431 293 465
rect 217 419 293 431
rect 369 438 428 560
rect 369 404 381 438
rect 415 404 428 438
rect 369 392 428 404
rect 458 392 555 560
rect 585 392 639 592
rect 669 539 782 592
rect 669 505 700 539
rect 734 508 782 539
rect 812 508 866 592
rect 896 567 1026 592
rect 896 533 910 567
rect 944 533 979 567
rect 1013 533 1026 567
rect 896 508 1026 533
rect 734 505 764 508
rect 669 447 764 505
rect 669 413 700 447
rect 734 413 764 447
rect 669 392 764 413
rect 967 392 1026 508
rect 1056 580 1115 592
rect 1056 546 1069 580
rect 1103 546 1115 580
rect 1056 509 1115 546
rect 1056 475 1069 509
rect 1103 475 1115 509
rect 1056 438 1115 475
rect 1056 404 1069 438
rect 1103 404 1115 438
rect 1056 392 1115 404
rect 1169 580 1228 592
rect 1169 546 1181 580
rect 1215 546 1228 580
rect 1169 497 1228 546
rect 1169 463 1181 497
rect 1215 463 1228 497
rect 1169 414 1228 463
rect 1169 380 1181 414
rect 1215 380 1228 414
rect 1169 368 1228 380
rect 1258 580 1317 592
rect 1258 546 1271 580
rect 1305 546 1317 580
rect 1258 497 1317 546
rect 1258 463 1271 497
rect 1305 463 1317 497
rect 1258 414 1317 463
rect 1258 380 1271 414
rect 1305 380 1317 414
rect 1258 368 1317 380
<< ndiffc >>
rect 39 139 73 173
rect 243 216 277 250
rect 411 155 445 189
rect 141 48 175 82
rect 579 161 613 195
rect 579 91 613 125
rect 771 161 805 195
rect 986 177 1020 211
rect 986 107 1020 141
rect 1072 177 1106 211
rect 1072 107 1106 141
rect 1184 176 1218 210
rect 1184 86 1218 120
rect 1270 86 1304 120
<< pdiffc >>
rect 40 541 74 575
rect 40 431 74 465
rect 140 541 174 575
rect 140 431 174 465
rect 247 541 281 575
rect 489 572 523 606
rect 247 431 281 465
rect 381 404 415 438
rect 700 505 734 539
rect 910 533 944 567
rect 979 533 1013 567
rect 700 413 734 447
rect 1069 546 1103 580
rect 1069 475 1103 509
rect 1069 404 1103 438
rect 1181 546 1215 580
rect 1181 463 1215 497
rect 1181 380 1215 414
rect 1271 546 1305 580
rect 1271 463 1305 497
rect 1271 380 1305 414
<< poly >>
rect 87 587 117 613
rect 187 587 217 613
rect 428 560 458 586
rect 555 592 585 618
rect 639 592 669 618
rect 782 592 812 618
rect 866 592 896 618
rect 1026 592 1056 618
rect 1228 592 1258 618
rect 87 404 117 419
rect 187 404 217 419
rect 84 313 120 404
rect 21 297 120 313
rect 184 366 220 404
rect 782 493 812 508
rect 866 493 896 508
rect 428 377 458 392
rect 555 377 585 392
rect 639 377 669 392
rect 184 350 255 366
rect 184 316 205 350
rect 239 316 255 350
rect 184 300 255 316
rect 311 338 377 354
rect 311 304 327 338
rect 361 336 377 338
rect 425 336 461 377
rect 361 304 461 336
rect 552 311 588 377
rect 636 360 672 377
rect 636 344 702 360
rect 779 357 815 493
rect 863 471 899 493
rect 863 455 949 471
rect 863 441 885 455
rect 869 421 885 441
rect 919 421 949 455
rect 869 405 949 421
rect 21 263 37 297
rect 71 283 120 297
rect 71 263 114 283
rect 21 247 114 263
rect 202 262 232 300
rect 311 270 461 304
rect 84 225 114 247
rect 84 89 114 115
rect 311 236 327 270
rect 361 267 461 270
rect 528 295 594 311
rect 361 237 486 267
rect 528 261 544 295
rect 578 261 594 295
rect 636 310 652 344
rect 686 310 702 344
rect 636 294 702 310
rect 746 341 868 357
rect 746 307 818 341
rect 852 307 868 341
rect 528 252 594 261
rect 746 291 868 307
rect 746 252 776 291
rect 528 245 655 252
rect 361 236 377 237
rect 311 202 377 236
rect 456 222 486 237
rect 564 222 655 245
rect 311 168 327 202
rect 361 168 377 202
rect 311 152 377 168
rect 202 88 232 114
rect 625 207 655 222
rect 703 222 776 252
rect 841 223 871 249
rect 919 223 949 405
rect 1026 377 1056 392
rect 1023 327 1059 377
rect 1228 353 1258 368
rect 997 311 1063 327
rect 1225 326 1261 353
rect 997 277 1013 311
rect 1047 277 1063 311
rect 997 261 1063 277
rect 1111 310 1261 326
rect 1111 276 1127 310
rect 1161 296 1261 310
rect 1161 276 1259 296
rect 1031 223 1061 261
rect 1111 260 1259 276
rect 703 207 733 222
rect 841 117 871 139
rect 805 101 871 117
rect 919 113 949 139
rect 456 48 486 74
rect 625 53 655 79
rect 703 53 733 79
rect 805 67 821 101
rect 855 67 871 101
rect 1229 222 1259 260
rect 1031 69 1061 95
rect 805 51 871 67
rect 1229 48 1259 74
<< polycont >>
rect 205 316 239 350
rect 327 304 361 338
rect 885 421 919 455
rect 37 263 71 297
rect 327 236 361 270
rect 544 261 578 295
rect 652 310 686 344
rect 818 307 852 341
rect 327 168 361 202
rect 1013 277 1047 311
rect 1127 276 1161 310
rect 821 67 855 101
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 24 575 90 591
rect 24 541 40 575
rect 74 541 90 575
rect 24 465 90 541
rect 24 431 40 465
rect 74 431 90 465
rect 24 381 90 431
rect 124 575 190 649
rect 472 606 541 649
rect 124 541 140 575
rect 174 541 190 575
rect 124 465 190 541
rect 124 431 140 465
rect 174 431 190 465
rect 124 415 190 431
rect 231 575 331 591
rect 231 541 247 575
rect 281 541 331 575
rect 472 572 489 606
rect 523 572 541 606
rect 472 556 541 572
rect 575 581 836 615
rect 231 522 331 541
rect 575 522 609 581
rect 231 488 609 522
rect 666 539 768 547
rect 666 505 700 539
rect 734 505 768 539
rect 231 465 331 488
rect 231 431 247 465
rect 281 431 331 465
rect 231 415 331 431
rect 24 347 155 381
rect 21 297 87 313
rect 21 263 37 297
rect 71 263 87 297
rect 21 236 87 263
rect 121 202 155 347
rect 189 350 263 366
rect 189 316 205 350
rect 239 316 263 350
rect 189 300 263 316
rect 297 354 331 415
rect 365 438 445 454
rect 365 404 381 438
rect 415 404 445 438
rect 666 447 768 505
rect 666 413 700 447
rect 365 388 445 404
rect 411 379 445 388
rect 297 338 377 354
rect 297 304 327 338
rect 361 304 377 338
rect 297 270 377 304
rect 297 266 327 270
rect 23 173 155 202
rect 227 250 327 266
rect 227 216 243 250
rect 277 236 327 250
rect 361 236 377 270
rect 277 216 377 236
rect 227 202 377 216
rect 227 200 327 202
rect 23 139 39 173
rect 73 166 155 173
rect 297 168 327 200
rect 361 168 377 202
rect 73 139 263 166
rect 297 152 377 168
rect 411 345 700 379
rect 411 189 461 345
rect 636 344 700 345
rect 445 155 461 189
rect 23 132 263 139
rect 23 111 89 132
rect 125 82 191 98
rect 125 48 141 82
rect 175 48 191 82
rect 229 85 263 132
rect 411 119 461 155
rect 495 295 594 311
rect 495 261 544 295
rect 578 261 594 295
rect 636 310 652 344
rect 686 310 700 344
rect 636 294 700 310
rect 495 245 594 261
rect 495 85 529 245
rect 229 51 529 85
rect 563 195 629 211
rect 563 161 579 195
rect 613 161 629 195
rect 563 125 629 161
rect 563 91 579 125
rect 613 91 629 125
rect 125 17 191 48
rect 563 17 629 91
rect 663 117 697 294
rect 734 211 768 447
rect 802 357 836 581
rect 894 567 1013 649
rect 894 533 910 567
rect 944 533 979 567
rect 894 505 1013 533
rect 1053 580 1131 596
rect 1053 546 1069 580
rect 1103 546 1131 580
rect 1053 509 1131 546
rect 1053 475 1069 509
rect 1103 475 1131 509
rect 1053 471 1131 475
rect 870 455 1131 471
rect 870 421 885 455
rect 919 438 1131 455
rect 919 421 1069 438
rect 870 405 1069 421
rect 1053 404 1069 405
rect 1103 404 1131 438
rect 1053 388 1131 404
rect 802 341 868 357
rect 802 307 818 341
rect 852 307 868 341
rect 802 291 868 307
rect 902 311 1063 327
rect 902 277 1013 311
rect 1047 277 1063 311
rect 902 261 1063 277
rect 1097 326 1131 388
rect 1165 580 1215 649
rect 1165 546 1181 580
rect 1165 497 1215 546
rect 1165 463 1181 497
rect 1165 414 1215 463
rect 1165 380 1181 414
rect 1165 364 1215 380
rect 1254 580 1321 596
rect 1254 546 1271 580
rect 1305 546 1321 580
rect 1254 497 1321 546
rect 1254 463 1271 497
rect 1305 463 1321 497
rect 1254 414 1321 463
rect 1254 380 1271 414
rect 1305 380 1321 414
rect 1097 310 1177 326
rect 1097 276 1127 310
rect 1161 276 1177 310
rect 902 211 936 261
rect 1097 260 1177 276
rect 1097 227 1131 260
rect 731 195 936 211
rect 731 161 771 195
rect 805 161 936 195
rect 970 211 1020 227
rect 970 177 986 211
rect 970 141 1020 177
rect 663 101 871 117
rect 663 67 821 101
rect 855 67 871 101
rect 663 51 871 67
rect 970 107 986 141
rect 970 17 1020 107
rect 1056 211 1131 227
rect 1056 177 1072 211
rect 1106 177 1131 211
rect 1056 141 1131 177
rect 1056 107 1072 141
rect 1106 107 1131 141
rect 1056 91 1131 107
rect 1168 210 1218 226
rect 1168 176 1184 210
rect 1168 120 1218 176
rect 1168 86 1184 120
rect 1168 17 1218 86
rect 1254 120 1321 380
rect 1254 86 1270 120
rect 1304 86 1321 120
rect 1254 70 1321 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
<< metal1 >>
rect 0 683 1344 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 0 617 1344 649
rect 0 17 1344 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
rect 0 -49 1344 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dlxtn_1
flabel pwell s 0 0 1344 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 0 617 1344 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 0 617 1344 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 1344 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 1279 94 1313 128 0 FreeSans 340 0 0 0 Q
port 7 nsew
flabel corelocali s 1279 168 1313 202 0 FreeSans 340 0 0 0 Q
port 7 nsew
flabel corelocali s 1279 242 1313 276 0 FreeSans 340 0 0 0 Q
port 7 nsew
flabel corelocali s 1279 316 1313 350 0 FreeSans 340 0 0 0 Q
port 7 nsew
flabel corelocali s 1279 390 1313 424 0 FreeSans 340 0 0 0 Q
port 7 nsew
flabel corelocali s 1279 464 1313 498 0 FreeSans 340 0 0 0 Q
port 7 nsew
flabel corelocali s 1279 538 1313 572 0 FreeSans 340 0 0 0 Q
port 7 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 D
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 1344 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2982588
string GDS_START 2971468
<< end >>
