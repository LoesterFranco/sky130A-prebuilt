magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 17 199 133 265
rect 2187 325 2237 425
rect 2375 325 2425 425
rect 2563 325 2613 425
rect 2751 325 2801 425
rect 2939 325 2989 425
rect 3127 325 3177 425
rect 3315 325 3365 425
rect 3503 325 3553 425
rect 2187 291 3661 325
rect 2130 215 3520 257
rect 17 51 63 199
rect 3554 181 3661 291
rect 665 145 3661 181
rect 665 51 741 145
rect 853 51 929 145
rect 1041 51 1117 145
rect 1229 51 1305 145
rect 1417 51 1493 145
rect 1605 51 1681 145
rect 1793 51 1869 145
rect 1981 51 2057 145
rect 2169 51 2245 145
rect 2357 51 2433 145
rect 2545 51 2621 145
rect 2733 51 2809 145
rect 2921 51 2997 145
rect 3109 51 3185 145
rect 3297 51 3373 145
rect 3485 51 3561 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3157 561
rect 3191 527 3249 561
rect 3283 527 3341 561
rect 3375 527 3433 561
rect 3467 527 3525 561
rect 3559 527 3617 561
rect 3651 527 3680 561
rect 60 299 103 527
rect 137 299 223 493
rect 177 257 223 299
rect 267 291 311 527
rect 345 257 431 493
rect 475 291 534 527
rect 575 333 639 493
rect 683 367 733 527
rect 777 333 827 493
rect 871 367 921 527
rect 965 333 1015 493
rect 1059 367 1109 527
rect 1153 333 1203 493
rect 1247 367 1297 527
rect 1341 333 1391 493
rect 1435 367 1485 527
rect 1529 333 1579 493
rect 1623 367 1673 527
rect 1717 333 1767 493
rect 1811 367 1861 527
rect 1905 333 1955 493
rect 1999 367 2049 527
rect 2093 459 3647 493
rect 2093 333 2143 459
rect 575 291 2143 333
rect 2281 359 2331 459
rect 2469 359 2519 459
rect 2657 359 2707 459
rect 2845 359 2895 459
rect 3033 359 3083 459
rect 3221 359 3271 459
rect 3409 359 3459 459
rect 3597 359 3647 459
rect 177 215 2096 257
rect 177 213 477 215
rect 97 17 173 165
rect 217 51 269 213
rect 313 17 373 179
rect 417 51 477 213
rect 521 17 631 181
rect 785 17 819 111
rect 973 17 1007 111
rect 1161 17 1195 111
rect 1349 17 1383 111
rect 1537 17 1571 111
rect 1725 17 1759 111
rect 1913 17 1947 111
rect 2101 17 2135 111
rect 2289 17 2323 111
rect 2477 17 2511 111
rect 2665 17 2699 111
rect 2853 17 2887 111
rect 3041 17 3075 111
rect 3229 17 3263 111
rect 3417 17 3451 111
rect 3605 17 3659 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3341 17
rect 3375 -17 3433 17
rect 3467 -17 3525 17
rect 3559 -17 3617 17
rect 3651 -17 3680 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 2881 527 2915 561
rect 2973 527 3007 561
rect 3065 527 3099 561
rect 3157 527 3191 561
rect 3249 527 3283 561
rect 3341 527 3375 561
rect 3433 527 3467 561
rect 3525 527 3559 561
rect 3617 527 3651 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
rect 2881 -17 2915 17
rect 2973 -17 3007 17
rect 3065 -17 3099 17
rect 3157 -17 3191 17
rect 3249 -17 3283 17
rect 3341 -17 3375 17
rect 3433 -17 3467 17
rect 3525 -17 3559 17
rect 3617 -17 3651 17
<< metal1 >>
rect 0 561 3680 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3157 561
rect 3191 527 3249 561
rect 3283 527 3341 561
rect 3375 527 3433 561
rect 3467 527 3525 561
rect 3559 527 3617 561
rect 3651 527 3680 561
rect 0 496 3680 527
rect 0 17 3680 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3341 17
rect 3375 -17 3433 17
rect 3467 -17 3525 17
rect 3559 -17 3617 17
rect 3651 -17 3680 17
rect 0 -48 3680 -17
<< labels >>
rlabel locali s 17 199 133 265 6 A
port 1 nsew signal input
rlabel locali s 17 51 63 199 6 A
port 1 nsew signal input
rlabel locali s 2130 215 3520 257 6 SLEEP
port 2 nsew signal input
rlabel locali s 3554 181 3661 291 6 X
port 3 nsew signal output
rlabel locali s 3503 325 3553 425 6 X
port 3 nsew signal output
rlabel locali s 3485 51 3561 145 6 X
port 3 nsew signal output
rlabel locali s 3315 325 3365 425 6 X
port 3 nsew signal output
rlabel locali s 3297 51 3373 145 6 X
port 3 nsew signal output
rlabel locali s 3127 325 3177 425 6 X
port 3 nsew signal output
rlabel locali s 3109 51 3185 145 6 X
port 3 nsew signal output
rlabel locali s 2939 325 2989 425 6 X
port 3 nsew signal output
rlabel locali s 2921 51 2997 145 6 X
port 3 nsew signal output
rlabel locali s 2751 325 2801 425 6 X
port 3 nsew signal output
rlabel locali s 2733 51 2809 145 6 X
port 3 nsew signal output
rlabel locali s 2563 325 2613 425 6 X
port 3 nsew signal output
rlabel locali s 2545 51 2621 145 6 X
port 3 nsew signal output
rlabel locali s 2375 325 2425 425 6 X
port 3 nsew signal output
rlabel locali s 2357 51 2433 145 6 X
port 3 nsew signal output
rlabel locali s 2187 325 2237 425 6 X
port 3 nsew signal output
rlabel locali s 2187 291 3661 325 6 X
port 3 nsew signal output
rlabel locali s 2169 51 2245 145 6 X
port 3 nsew signal output
rlabel locali s 1981 51 2057 145 6 X
port 3 nsew signal output
rlabel locali s 1793 51 1869 145 6 X
port 3 nsew signal output
rlabel locali s 1605 51 1681 145 6 X
port 3 nsew signal output
rlabel locali s 1417 51 1493 145 6 X
port 3 nsew signal output
rlabel locali s 1229 51 1305 145 6 X
port 3 nsew signal output
rlabel locali s 1041 51 1117 145 6 X
port 3 nsew signal output
rlabel locali s 853 51 929 145 6 X
port 3 nsew signal output
rlabel locali s 665 145 3661 181 6 X
port 3 nsew signal output
rlabel locali s 665 51 741 145 6 X
port 3 nsew signal output
rlabel metal1 s 0 -48 3680 48 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 496 3680 592 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 3680 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2669582
string GDS_START 2644260
<< end >>
