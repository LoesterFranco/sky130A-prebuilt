magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 356 1862 704
rect -38 332 296 356
rect 574 332 1862 356
<< pwell >>
rect 0 0 1824 49
<< scnmos >>
rect 84 126 114 236
rect 223 88 253 236
rect 426 120 456 268
rect 529 74 559 202
rect 610 74 640 202
rect 725 74 755 158
rect 797 74 827 158
rect 995 74 1025 202
rect 1082 74 1112 202
rect 1168 74 1198 202
rect 1254 74 1284 202
rect 1452 74 1482 222
rect 1538 74 1568 222
rect 1624 74 1654 222
rect 1710 74 1740 222
<< pmoshvt >>
rect 86 394 116 562
rect 210 394 240 562
rect 423 392 453 560
rect 532 392 562 592
rect 610 392 640 592
rect 717 508 747 592
rect 842 508 872 592
rect 995 368 1025 536
rect 1085 368 1115 536
rect 1185 368 1215 536
rect 1285 368 1315 536
rect 1392 368 1422 592
rect 1482 368 1512 592
rect 1582 368 1612 592
rect 1686 368 1716 592
<< ndiff >>
rect 364 256 426 268
rect 27 198 84 236
rect 27 164 39 198
rect 73 164 84 198
rect 27 126 84 164
rect 114 172 223 236
rect 114 138 152 172
rect 186 138 223 172
rect 114 126 223 138
rect 129 88 223 126
rect 253 224 310 236
rect 253 190 264 224
rect 298 190 310 224
rect 253 134 310 190
rect 253 100 264 134
rect 298 100 310 134
rect 364 222 378 256
rect 412 222 426 256
rect 364 120 426 222
rect 456 202 506 268
rect 456 120 529 202
rect 253 88 310 100
rect 471 86 483 120
rect 517 86 529 120
rect 471 74 529 86
rect 559 74 610 202
rect 640 169 710 202
rect 640 135 657 169
rect 691 158 710 169
rect 1395 210 1452 222
rect 938 190 995 202
rect 691 135 725 158
rect 640 74 725 135
rect 755 74 797 158
rect 827 133 884 158
rect 827 99 838 133
rect 872 99 884 133
rect 827 74 884 99
rect 938 156 950 190
rect 984 156 995 190
rect 938 120 995 156
rect 938 86 950 120
rect 984 86 995 120
rect 938 74 995 86
rect 1025 174 1082 202
rect 1025 140 1036 174
rect 1070 140 1082 174
rect 1025 74 1082 140
rect 1112 188 1168 202
rect 1112 154 1123 188
rect 1157 154 1168 188
rect 1112 116 1168 154
rect 1112 82 1123 116
rect 1157 82 1168 116
rect 1112 74 1168 82
rect 1198 120 1254 202
rect 1198 86 1209 120
rect 1243 86 1254 120
rect 1198 74 1254 86
rect 1284 189 1341 202
rect 1284 155 1295 189
rect 1329 155 1341 189
rect 1284 119 1341 155
rect 1284 85 1295 119
rect 1329 85 1341 119
rect 1284 74 1341 85
rect 1395 176 1407 210
rect 1441 176 1452 210
rect 1395 123 1452 176
rect 1395 89 1407 123
rect 1441 89 1452 123
rect 1395 74 1452 89
rect 1482 210 1538 222
rect 1482 176 1493 210
rect 1527 176 1538 210
rect 1482 123 1538 176
rect 1482 89 1493 123
rect 1527 89 1538 123
rect 1482 74 1538 89
rect 1568 123 1624 222
rect 1568 89 1579 123
rect 1613 89 1624 123
rect 1568 74 1624 89
rect 1654 210 1710 222
rect 1654 176 1665 210
rect 1699 176 1710 210
rect 1654 123 1710 176
rect 1654 89 1665 123
rect 1699 89 1710 123
rect 1654 74 1710 89
rect 1740 123 1797 222
rect 1740 89 1751 123
rect 1785 89 1797 123
rect 1740 74 1797 89
<< pdiff >>
rect 134 592 192 604
rect 134 562 146 592
rect 27 550 86 562
rect 27 516 39 550
rect 73 516 86 550
rect 27 440 86 516
rect 27 406 39 440
rect 73 406 86 440
rect 27 394 86 406
rect 116 558 146 562
rect 180 562 192 592
rect 180 558 210 562
rect 116 394 210 558
rect 240 440 310 562
rect 471 578 532 592
rect 471 560 483 578
rect 240 406 258 440
rect 292 406 310 440
rect 240 394 310 406
rect 364 439 423 560
rect 364 405 376 439
rect 410 405 423 439
rect 364 392 423 405
rect 453 544 483 560
rect 517 544 532 578
rect 453 392 532 544
rect 562 392 610 592
rect 640 531 717 592
rect 640 497 653 531
rect 687 508 717 531
rect 747 508 842 592
rect 872 580 977 592
rect 872 546 908 580
rect 942 546 977 580
rect 1333 580 1392 592
rect 872 536 977 546
rect 1333 546 1345 580
rect 1379 546 1392 580
rect 1333 536 1392 546
rect 872 508 995 536
rect 687 497 699 508
rect 640 392 699 497
rect 942 368 995 508
rect 1025 524 1085 536
rect 1025 490 1038 524
rect 1072 490 1085 524
rect 1025 410 1085 490
rect 1025 376 1038 410
rect 1072 376 1085 410
rect 1025 368 1085 376
rect 1115 524 1185 536
rect 1115 490 1138 524
rect 1172 490 1185 524
rect 1115 431 1185 490
rect 1115 397 1138 431
rect 1172 397 1185 431
rect 1115 368 1185 397
rect 1215 524 1285 536
rect 1215 490 1238 524
rect 1272 490 1285 524
rect 1215 414 1285 490
rect 1215 380 1238 414
rect 1272 380 1285 414
rect 1215 368 1285 380
rect 1315 500 1392 536
rect 1315 466 1345 500
rect 1379 466 1392 500
rect 1315 426 1392 466
rect 1315 392 1345 426
rect 1379 392 1392 426
rect 1315 368 1392 392
rect 1422 580 1482 592
rect 1422 546 1435 580
rect 1469 546 1482 580
rect 1422 497 1482 546
rect 1422 463 1435 497
rect 1469 463 1482 497
rect 1422 414 1482 463
rect 1422 380 1435 414
rect 1469 380 1482 414
rect 1422 368 1482 380
rect 1512 580 1582 592
rect 1512 546 1535 580
rect 1569 546 1582 580
rect 1512 462 1582 546
rect 1512 428 1535 462
rect 1569 428 1582 462
rect 1512 368 1582 428
rect 1612 580 1686 592
rect 1612 546 1635 580
rect 1669 546 1686 580
rect 1612 497 1686 546
rect 1612 463 1635 497
rect 1669 463 1686 497
rect 1612 414 1686 463
rect 1612 380 1635 414
rect 1669 380 1686 414
rect 1612 368 1686 380
rect 1716 580 1781 592
rect 1716 546 1735 580
rect 1769 546 1781 580
rect 1716 462 1781 546
rect 1716 428 1735 462
rect 1769 428 1781 462
rect 1716 368 1781 428
<< ndiffc >>
rect 39 164 73 198
rect 152 138 186 172
rect 264 190 298 224
rect 264 100 298 134
rect 378 222 412 256
rect 483 86 517 120
rect 657 135 691 169
rect 838 99 872 133
rect 950 156 984 190
rect 950 86 984 120
rect 1036 140 1070 174
rect 1123 154 1157 188
rect 1123 82 1157 116
rect 1209 86 1243 120
rect 1295 155 1329 189
rect 1295 85 1329 119
rect 1407 176 1441 210
rect 1407 89 1441 123
rect 1493 176 1527 210
rect 1493 89 1527 123
rect 1579 89 1613 123
rect 1665 176 1699 210
rect 1665 89 1699 123
rect 1751 89 1785 123
<< pdiffc >>
rect 39 516 73 550
rect 39 406 73 440
rect 146 558 180 592
rect 258 406 292 440
rect 376 405 410 439
rect 483 544 517 578
rect 653 497 687 531
rect 908 546 942 580
rect 1345 546 1379 580
rect 1038 490 1072 524
rect 1038 376 1072 410
rect 1138 490 1172 524
rect 1138 397 1172 431
rect 1238 490 1272 524
rect 1238 380 1272 414
rect 1345 466 1379 500
rect 1345 392 1379 426
rect 1435 546 1469 580
rect 1435 463 1469 497
rect 1435 380 1469 414
rect 1535 546 1569 580
rect 1535 428 1569 462
rect 1635 546 1669 580
rect 1635 463 1669 497
rect 1635 380 1669 414
rect 1735 546 1769 580
rect 1735 428 1769 462
<< poly >>
rect 532 592 562 618
rect 610 592 640 618
rect 717 592 747 618
rect 842 592 872 618
rect 1392 592 1422 618
rect 1482 592 1512 618
rect 1582 592 1612 618
rect 1686 592 1716 618
rect 86 562 116 588
rect 210 562 240 588
rect 423 560 453 586
rect 86 379 116 394
rect 210 379 240 394
rect 995 536 1025 562
rect 1085 536 1115 562
rect 1185 536 1215 562
rect 1285 536 1315 562
rect 717 493 747 508
rect 842 493 872 508
rect 714 476 750 493
rect 839 476 875 493
rect 714 460 797 476
rect 714 426 747 460
rect 781 426 797 460
rect 714 410 797 426
rect 839 460 905 476
rect 839 426 855 460
rect 889 426 905 460
rect 839 410 905 426
rect 83 356 119 379
rect 207 356 243 379
rect 423 377 453 392
rect 532 377 562 392
rect 610 377 640 392
rect 420 356 456 377
rect 529 360 565 377
rect 44 340 119 356
rect 44 306 60 340
rect 94 306 119 340
rect 44 290 119 306
rect 200 340 266 356
rect 200 306 216 340
rect 250 306 266 340
rect 200 290 266 306
rect 314 340 456 356
rect 314 306 330 340
rect 364 306 456 340
rect 314 290 456 306
rect 499 344 565 360
rect 499 310 515 344
rect 549 310 565 344
rect 607 368 643 377
rect 607 338 755 368
rect 499 294 565 310
rect 725 311 755 338
rect 725 295 830 311
rect 84 236 114 290
rect 223 236 253 290
rect 426 268 456 290
rect 84 100 114 126
rect 529 202 559 294
rect 607 274 673 290
rect 607 240 623 274
rect 657 240 673 274
rect 607 224 673 240
rect 725 261 780 295
rect 814 261 830 295
rect 725 245 830 261
rect 610 202 640 224
rect 426 94 456 120
rect 223 62 253 88
rect 725 158 755 245
rect 872 203 902 410
rect 995 353 1025 368
rect 1085 353 1115 368
rect 1185 353 1215 368
rect 1285 353 1315 368
rect 1392 353 1422 368
rect 1482 353 1512 368
rect 1582 353 1612 368
rect 1686 353 1716 368
rect 992 336 1028 353
rect 944 320 1028 336
rect 944 286 960 320
rect 994 300 1028 320
rect 1082 300 1118 353
rect 994 286 1118 300
rect 1182 290 1218 353
rect 1282 290 1318 353
rect 944 270 1118 286
rect 797 173 902 203
rect 995 202 1025 270
rect 1082 240 1118 270
rect 1168 274 1318 290
rect 1168 240 1193 274
rect 1227 240 1261 274
rect 1295 240 1318 274
rect 1389 326 1425 353
rect 1479 326 1515 353
rect 1579 326 1615 353
rect 1683 326 1719 353
rect 1389 310 1719 326
rect 1389 276 1465 310
rect 1499 276 1533 310
rect 1567 276 1601 310
rect 1635 276 1669 310
rect 1703 290 1719 310
rect 1703 276 1740 290
rect 1389 260 1740 276
rect 1082 202 1112 240
rect 1168 224 1318 240
rect 1168 202 1198 224
rect 1254 202 1284 224
rect 1452 222 1482 260
rect 1538 222 1568 260
rect 1624 222 1654 260
rect 1710 222 1740 260
rect 797 158 827 173
rect 529 48 559 74
rect 610 48 640 74
rect 725 48 755 74
rect 797 48 827 74
rect 995 48 1025 74
rect 1082 48 1112 74
rect 1168 48 1198 74
rect 1254 48 1284 74
rect 1452 48 1482 74
rect 1538 48 1568 74
rect 1624 48 1654 74
rect 1710 48 1740 74
<< polycont >>
rect 747 426 781 460
rect 855 426 889 460
rect 60 306 94 340
rect 216 306 250 340
rect 330 306 364 340
rect 515 310 549 344
rect 623 240 657 274
rect 780 261 814 295
rect 960 286 994 320
rect 1193 240 1227 274
rect 1261 240 1295 274
rect 1465 276 1499 310
rect 1533 276 1567 310
rect 1601 276 1635 310
rect 1669 276 1703 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 130 592 196 649
rect 23 550 89 566
rect 23 516 39 550
rect 73 516 89 550
rect 130 558 146 592
rect 180 558 196 592
rect 130 542 196 558
rect 467 578 533 649
rect 467 544 483 578
rect 517 544 533 578
rect 467 542 533 544
rect 569 581 797 615
rect 23 508 89 516
rect 23 474 533 508
rect 23 440 171 474
rect 23 406 39 440
rect 73 406 171 440
rect 23 390 171 406
rect 237 406 258 440
rect 292 406 326 440
rect 237 390 326 406
rect 360 439 448 440
rect 360 405 376 439
rect 410 405 448 439
rect 360 404 448 405
rect 25 340 103 356
rect 25 306 60 340
rect 94 306 103 340
rect 25 290 103 306
rect 137 256 171 390
rect 292 356 326 390
rect 205 340 258 356
rect 205 306 216 340
rect 250 306 258 340
rect 205 290 258 306
rect 292 340 380 356
rect 292 306 330 340
rect 364 306 380 340
rect 292 290 380 306
rect 23 222 171 256
rect 292 240 326 290
rect 414 256 448 404
rect 499 360 533 474
rect 569 428 603 581
rect 637 531 693 547
rect 637 497 653 531
rect 687 497 693 531
rect 637 481 693 497
rect 569 394 625 428
rect 499 344 557 360
rect 499 310 515 344
rect 549 310 557 344
rect 499 294 557 310
rect 591 290 625 394
rect 659 379 693 481
rect 731 460 797 581
rect 869 580 981 649
rect 869 546 908 580
rect 942 546 981 580
rect 869 530 981 546
rect 1022 524 1088 540
rect 1022 496 1038 524
rect 731 426 747 460
rect 781 426 797 460
rect 731 413 797 426
rect 839 490 1038 496
rect 1072 490 1088 524
rect 839 460 1088 490
rect 839 426 855 460
rect 889 426 1088 460
rect 839 413 1088 426
rect 1038 410 1088 413
rect 659 345 1004 379
rect 591 274 668 290
rect 591 256 623 274
rect 248 224 326 240
rect 23 198 89 222
rect 23 164 39 198
rect 73 164 89 198
rect 248 190 264 224
rect 298 190 326 224
rect 360 222 378 256
rect 412 240 623 256
rect 657 240 668 274
rect 412 222 668 240
rect 248 188 326 190
rect 23 122 89 164
rect 136 172 202 188
rect 136 138 152 172
rect 186 138 202 172
rect 136 17 202 138
rect 248 154 601 188
rect 702 185 736 345
rect 944 320 1004 345
rect 248 134 326 154
rect 248 100 264 134
rect 298 100 326 134
rect 248 84 326 100
rect 467 86 483 120
rect 517 86 533 120
rect 467 17 533 86
rect 567 85 601 154
rect 635 169 736 185
rect 635 135 657 169
rect 691 135 736 169
rect 635 119 736 135
rect 770 295 830 311
rect 770 261 780 295
rect 814 261 830 295
rect 944 286 960 320
rect 994 286 1004 320
rect 944 270 1004 286
rect 1072 376 1088 410
rect 1122 524 1188 649
rect 1329 580 1395 649
rect 1329 546 1345 580
rect 1379 546 1395 580
rect 1122 490 1138 524
rect 1172 490 1188 524
rect 1122 431 1188 490
rect 1122 397 1138 431
rect 1172 397 1188 431
rect 1122 392 1188 397
rect 1222 524 1288 540
rect 1222 490 1238 524
rect 1272 490 1288 524
rect 1222 414 1288 490
rect 1038 358 1088 376
rect 1222 380 1238 414
rect 1272 380 1288 414
rect 1329 500 1395 546
rect 1329 466 1345 500
rect 1379 466 1395 500
rect 1329 426 1395 466
rect 1329 392 1345 426
rect 1379 392 1395 426
rect 1435 580 1485 596
rect 1469 546 1485 580
rect 1435 497 1485 546
rect 1469 463 1485 497
rect 1435 414 1485 463
rect 1519 580 1585 649
rect 1519 546 1535 580
rect 1569 546 1585 580
rect 1519 462 1585 546
rect 1519 428 1535 462
rect 1569 428 1585 462
rect 1619 580 1685 596
rect 1619 546 1635 580
rect 1669 546 1685 580
rect 1619 497 1685 546
rect 1619 463 1635 497
rect 1669 463 1685 497
rect 1222 358 1288 380
rect 1469 394 1485 414
rect 1619 414 1685 463
rect 1719 580 1785 649
rect 1719 546 1735 580
rect 1769 546 1785 580
rect 1719 462 1785 546
rect 1719 428 1735 462
rect 1769 428 1785 462
rect 1619 394 1635 414
rect 1469 380 1635 394
rect 1669 394 1685 414
rect 1669 380 1799 394
rect 1435 360 1799 380
rect 1038 326 1387 358
rect 1038 324 1719 326
rect 770 245 830 261
rect 770 85 804 245
rect 934 190 1000 206
rect 1038 190 1072 324
rect 1353 310 1719 324
rect 1177 274 1319 290
rect 1177 240 1193 274
rect 1227 240 1261 274
rect 1295 240 1319 274
rect 1353 276 1465 310
rect 1499 276 1533 310
rect 1567 276 1601 310
rect 1635 276 1669 310
rect 1703 276 1719 310
rect 1353 260 1719 276
rect 1177 224 1319 240
rect 1753 226 1799 360
rect 1391 210 1443 226
rect 567 51 804 85
rect 838 133 888 162
rect 872 99 888 133
rect 838 17 888 99
rect 934 156 950 190
rect 984 156 1000 190
rect 934 120 1000 156
rect 1036 174 1072 190
rect 1070 140 1072 174
rect 1036 124 1072 140
rect 1107 189 1345 190
rect 1107 188 1295 189
rect 1107 154 1123 188
rect 1157 155 1295 188
rect 1329 155 1345 189
rect 1157 154 1345 155
rect 934 86 950 120
rect 984 90 1000 120
rect 1107 116 1157 154
rect 1107 90 1123 116
rect 984 86 1123 90
rect 934 82 1123 86
rect 934 56 1157 82
rect 1193 86 1209 120
rect 1243 86 1259 120
rect 1193 17 1259 86
rect 1293 119 1345 154
rect 1293 85 1295 119
rect 1329 85 1345 119
rect 1293 69 1345 85
rect 1391 176 1407 210
rect 1441 176 1443 210
rect 1391 123 1443 176
rect 1391 89 1407 123
rect 1441 89 1443 123
rect 1391 17 1443 89
rect 1477 210 1799 226
rect 1477 176 1493 210
rect 1527 176 1665 210
rect 1699 176 1799 210
rect 1477 123 1529 176
rect 1477 89 1493 123
rect 1527 89 1529 123
rect 1477 73 1529 89
rect 1563 123 1629 142
rect 1563 89 1579 123
rect 1613 89 1629 123
rect 1563 17 1629 89
rect 1663 123 1701 176
rect 1663 89 1665 123
rect 1699 89 1701 123
rect 1663 73 1701 89
rect 1735 123 1801 142
rect 1735 89 1751 123
rect 1785 89 1801 123
rect 1735 17 1801 89
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
<< metal1 >>
rect 0 683 1824 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 0 617 1824 649
rect 0 17 1824 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
rect 0 -49 1824 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dlrtp_4
flabel pwell s 0 0 1824 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 1824 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 1824 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 1824 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 D
port 1 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 GATE
port 2 nsew
flabel corelocali s 1183 242 1217 276 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew
flabel corelocali s 1279 242 1313 276 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew
flabel corelocali s 1759 242 1793 276 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 1759 316 1793 350 0 FreeSans 340 0 0 0 Q
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 1824 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3034352
string GDS_START 3020624
<< end >>
