magic
tech sky130A
magscale 1 2
timestamp 1599588238
<< locali >>
rect 25 200 104 439
rect 409 339 455 356
rect 362 262 455 339
rect 1852 362 1990 597
rect 1912 70 1990 362
rect 2215 364 2287 596
rect 2253 226 2287 364
rect 2213 70 2287 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2304 683
rect 23 504 73 649
rect 113 526 169 596
rect 203 550 269 649
rect 405 550 471 649
rect 113 516 178 526
rect 281 516 393 518
rect 613 516 669 538
rect 113 504 669 516
rect 703 505 854 539
rect 888 533 957 649
rect 998 508 1065 536
rect 138 484 669 504
rect 138 482 306 484
rect 378 482 669 484
rect 138 462 285 482
rect 629 471 669 482
rect 802 499 854 505
rect 989 499 1065 508
rect 138 166 172 462
rect 319 428 365 450
rect 206 424 260 428
rect 206 390 223 424
rect 257 390 260 424
rect 206 226 260 390
rect 294 373 365 428
rect 495 416 595 448
rect 629 437 768 471
rect 495 413 600 416
rect 495 412 604 413
rect 495 408 605 412
rect 495 403 610 408
rect 495 373 700 403
rect 294 228 328 373
rect 583 365 700 373
rect 589 359 700 365
rect 495 310 561 339
rect 489 298 561 310
rect 595 315 700 359
rect 489 228 555 298
rect 595 278 632 315
rect 294 195 555 228
rect 589 241 632 278
rect 734 274 768 437
rect 294 194 512 195
rect 34 132 172 166
rect 34 74 100 132
rect 206 17 256 166
rect 294 119 384 194
rect 589 161 623 241
rect 666 240 768 274
rect 802 465 1065 499
rect 666 207 707 240
rect 418 17 484 160
rect 522 85 623 161
rect 657 119 707 207
rect 802 206 836 465
rect 978 456 1021 465
rect 741 119 836 206
rect 870 218 926 431
rect 978 323 1012 456
rect 1046 424 1122 431
rect 1046 390 1087 424
rect 1121 390 1122 424
rect 1046 365 1122 390
rect 1156 348 1206 649
rect 978 289 1112 323
rect 1246 314 1296 551
rect 1340 473 1533 539
rect 1046 257 1112 289
rect 1149 280 1296 314
rect 1330 373 1465 439
rect 1149 218 1183 280
rect 1330 246 1364 373
rect 1499 319 1533 473
rect 1567 467 1612 649
rect 1652 467 1728 546
rect 1567 424 1660 433
rect 1601 390 1660 424
rect 1567 367 1660 390
rect 1694 387 1728 467
rect 1762 421 1805 649
rect 1694 353 1794 387
rect 870 184 1183 218
rect 1217 180 1364 246
rect 1398 285 1726 319
rect 1217 150 1251 180
rect 870 116 1251 150
rect 1398 146 1432 285
rect 1666 253 1726 285
rect 1486 214 1552 246
rect 1760 214 1794 353
rect 1486 180 1794 214
rect 870 85 904 116
rect 522 51 904 85
rect 999 17 1065 82
rect 1285 80 1432 146
rect 1507 17 1599 136
rect 1697 70 1794 180
rect 1828 17 1878 226
rect 2038 326 2088 595
rect 2122 364 2181 649
rect 2038 260 2219 326
rect 2038 70 2088 260
rect 2129 17 2179 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2304 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 223 390 257 424
rect 1087 390 1121 424
rect 1567 390 1601 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
<< metal1 >>
rect 0 683 2304 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2304 683
rect 0 617 2304 649
rect 211 424 269 430
rect 211 390 223 424
rect 257 421 269 424
rect 1075 424 1133 430
rect 1075 421 1087 424
rect 257 393 1087 421
rect 257 390 269 393
rect 211 384 269 390
rect 1075 390 1087 393
rect 1121 421 1133 424
rect 1555 424 1613 430
rect 1555 421 1567 424
rect 1121 393 1567 421
rect 1121 390 1133 393
rect 1075 384 1133 390
rect 1555 390 1567 393
rect 1601 390 1613 424
rect 1555 384 1613 390
rect 0 17 2304 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2304 17
rect 0 -49 2304 -17
<< labels >>
rlabel locali s 25 200 104 439 6 D
port 1 nsew signal input
rlabel locali s 2253 226 2287 364 6 Q
port 2 nsew signal output
rlabel locali s 2215 364 2287 596 6 Q
port 2 nsew signal output
rlabel locali s 2213 70 2287 226 6 Q
port 2 nsew signal output
rlabel locali s 1912 70 1990 362 6 Q_N
port 3 nsew signal output
rlabel locali s 1852 362 1990 597 6 Q_N
port 3 nsew signal output
rlabel metal1 s 1555 421 1613 430 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 1555 384 1613 393 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 1075 421 1133 430 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 1075 384 1133 393 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 211 421 269 430 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 211 393 1613 421 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 211 384 269 393 6 RESET_B
port 4 nsew signal input
rlabel locali s 409 339 455 356 6 CLK
port 5 nsew clock input
rlabel locali s 362 262 455 339 6 CLK
port 5 nsew clock input
rlabel metal1 s 0 -49 2304 49 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 617 2304 715 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2304 666
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2549030
string GDS_START 2530424
<< end >>
