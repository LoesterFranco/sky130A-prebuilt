magic
tech sky130A
magscale 1 2
timestamp 1601050082
<< locali >>
rect 21 256 87 326
rect 121 290 509 356
rect 713 394 747 596
rect 877 394 943 596
rect 713 360 1031 394
rect 551 256 611 310
rect 21 222 611 256
rect 21 56 87 222
rect 985 226 1031 360
rect 210 54 276 188
rect 713 192 1031 226
rect 713 70 747 192
rect 881 70 931 192
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 23 384 73 649
rect 113 508 163 592
rect 203 542 466 592
rect 500 508 566 592
rect 113 474 566 508
rect 113 390 163 474
rect 500 458 566 474
rect 607 458 673 649
rect 299 424 365 440
rect 299 390 679 424
rect 645 326 679 390
rect 787 428 837 649
rect 983 428 1033 649
rect 645 260 937 326
rect 645 188 679 260
rect 310 154 679 188
rect 310 70 376 154
rect 410 17 476 120
rect 510 70 576 154
rect 610 17 676 120
rect 783 17 833 158
rect 967 17 1033 158
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 683 1056 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 0 617 1056 649
rect 0 17 1056 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -49 1056 -17
<< labels >>
rlabel locali s 551 256 611 310 6 A
port 1 nsew signal input
rlabel locali s 21 256 87 326 6 A
port 1 nsew signal input
rlabel locali s 21 222 611 256 6 A
port 1 nsew signal input
rlabel locali s 21 56 87 222 6 A
port 1 nsew signal input
rlabel locali s 121 290 509 356 6 B
port 2 nsew signal input
rlabel locali s 210 54 276 188 6 C
port 3 nsew signal input
rlabel locali s 985 226 1031 360 6 X
port 4 nsew signal output
rlabel locali s 881 70 931 192 6 X
port 4 nsew signal output
rlabel locali s 877 394 943 596 6 X
port 4 nsew signal output
rlabel locali s 713 394 747 596 6 X
port 4 nsew signal output
rlabel locali s 713 360 1031 394 6 X
port 4 nsew signal output
rlabel locali s 713 192 1031 226 6 X
port 4 nsew signal output
rlabel locali s 713 70 747 192 6 X
port 4 nsew signal output
rlabel metal1 s 0 -49 1056 49 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1056 715 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1056 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 975548
string GDS_START 966112
<< end >>
