magic
tech sky130A
magscale 1 2
timestamp 1599588218
<< nwell >>
rect -38 332 1478 704
<< pwell >>
rect 0 0 1440 49
<< scpmos >>
rect 83 392 119 592
rect 347 392 383 592
rect 549 368 585 592
rect 639 368 675 592
rect 739 368 775 592
rect 839 368 875 592
rect 1041 368 1077 592
rect 1131 368 1167 592
rect 1231 368 1267 592
rect 1321 368 1357 592
<< nmoslvt >>
rect 158 74 188 202
rect 281 124 311 252
rect 553 74 583 222
rect 639 74 669 222
rect 766 74 796 222
rect 852 74 882 222
rect 952 74 982 222
rect 1038 74 1068 222
rect 1231 74 1261 222
rect 1326 74 1356 222
<< ndiff >>
rect 225 202 281 252
rect 101 190 158 202
rect 101 156 113 190
rect 147 156 158 190
rect 101 122 158 156
rect 101 88 113 122
rect 147 88 158 122
rect 101 74 158 88
rect 188 124 281 202
rect 311 244 389 252
rect 311 210 341 244
rect 375 210 389 244
rect 311 124 389 210
rect 188 107 261 124
rect 188 74 215 107
rect 203 73 215 74
rect 249 73 261 107
rect 203 61 261 73
rect 443 92 553 222
rect 443 58 473 92
rect 507 74 553 92
rect 583 152 639 222
rect 583 118 594 152
rect 628 118 639 152
rect 583 74 639 118
rect 669 84 766 222
rect 669 74 700 84
rect 507 58 538 74
rect 443 46 538 58
rect 684 50 700 74
rect 734 74 766 84
rect 796 210 852 222
rect 796 176 807 210
rect 841 176 852 210
rect 796 120 852 176
rect 796 86 807 120
rect 841 86 852 120
rect 796 74 852 86
rect 882 152 952 222
rect 882 118 907 152
rect 941 118 952 152
rect 882 74 952 118
rect 982 210 1038 222
rect 982 176 993 210
rect 1027 176 1038 210
rect 982 120 1038 176
rect 982 86 993 120
rect 1027 86 1038 120
rect 982 74 1038 86
rect 1068 152 1231 222
rect 1068 118 1079 152
rect 1113 118 1186 152
rect 1220 118 1231 152
rect 1068 74 1231 118
rect 1261 210 1326 222
rect 1261 176 1281 210
rect 1315 176 1326 210
rect 1261 120 1326 176
rect 1261 86 1281 120
rect 1315 86 1326 120
rect 1261 74 1326 86
rect 1356 210 1413 222
rect 1356 176 1367 210
rect 1401 176 1413 210
rect 1356 120 1413 176
rect 1356 86 1367 120
rect 1401 86 1413 120
rect 1356 74 1413 86
rect 734 50 751 74
rect 684 38 751 50
<< pdiff >>
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 512 83 546
rect 27 478 39 512
rect 73 478 83 512
rect 27 444 83 478
rect 27 410 39 444
rect 73 410 83 444
rect 27 392 83 410
rect 119 580 347 592
rect 119 546 129 580
rect 163 546 216 580
rect 250 546 303 580
rect 337 546 347 580
rect 119 512 347 546
rect 119 478 129 512
rect 163 478 216 512
rect 250 478 303 512
rect 337 478 347 512
rect 119 444 347 478
rect 119 410 129 444
rect 163 410 216 444
rect 250 410 303 444
rect 337 410 347 444
rect 119 392 347 410
rect 383 580 439 592
rect 383 546 393 580
rect 427 546 439 580
rect 383 512 439 546
rect 383 478 393 512
rect 427 478 439 512
rect 383 444 439 478
rect 383 410 393 444
rect 427 410 439 444
rect 383 392 439 410
rect 493 580 549 592
rect 493 546 505 580
rect 539 546 549 580
rect 493 496 549 546
rect 493 462 505 496
rect 539 462 549 496
rect 493 420 549 462
rect 493 386 505 420
rect 539 386 549 420
rect 493 368 549 386
rect 585 531 639 592
rect 585 497 595 531
rect 629 497 639 531
rect 585 420 639 497
rect 585 386 595 420
rect 629 386 639 420
rect 585 368 639 386
rect 675 580 739 592
rect 675 546 695 580
rect 729 546 739 580
rect 675 488 739 546
rect 675 454 695 488
rect 729 454 739 488
rect 675 368 739 454
rect 775 556 839 592
rect 775 522 795 556
rect 829 522 839 556
rect 775 368 839 522
rect 875 540 931 592
rect 875 506 885 540
rect 919 506 931 540
rect 875 472 931 506
rect 875 438 885 472
rect 919 438 931 472
rect 875 368 931 438
rect 985 531 1041 592
rect 985 497 997 531
rect 1031 497 1041 531
rect 985 414 1041 497
rect 985 380 997 414
rect 1031 380 1041 414
rect 985 368 1041 380
rect 1077 580 1131 592
rect 1077 546 1087 580
rect 1121 546 1131 580
rect 1077 508 1131 546
rect 1077 474 1087 508
rect 1121 474 1131 508
rect 1077 368 1131 474
rect 1167 580 1231 592
rect 1167 546 1187 580
rect 1221 546 1231 580
rect 1167 503 1231 546
rect 1167 469 1187 503
rect 1221 469 1231 503
rect 1167 424 1231 469
rect 1167 390 1187 424
rect 1221 390 1231 424
rect 1167 368 1231 390
rect 1267 580 1321 592
rect 1267 546 1277 580
rect 1311 546 1321 580
rect 1267 508 1321 546
rect 1267 474 1277 508
rect 1311 474 1321 508
rect 1267 368 1321 474
rect 1357 580 1413 592
rect 1357 546 1367 580
rect 1401 546 1413 580
rect 1357 503 1413 546
rect 1357 469 1367 503
rect 1401 469 1413 503
rect 1357 424 1413 469
rect 1357 390 1367 424
rect 1401 390 1413 424
rect 1357 368 1413 390
<< ndiffc >>
rect 113 156 147 190
rect 113 88 147 122
rect 341 210 375 244
rect 215 73 249 107
rect 473 58 507 92
rect 594 118 628 152
rect 700 50 734 84
rect 807 176 841 210
rect 807 86 841 120
rect 907 118 941 152
rect 993 176 1027 210
rect 993 86 1027 120
rect 1079 118 1113 152
rect 1186 118 1220 152
rect 1281 176 1315 210
rect 1281 86 1315 120
rect 1367 176 1401 210
rect 1367 86 1401 120
<< pdiffc >>
rect 39 546 73 580
rect 39 478 73 512
rect 39 410 73 444
rect 129 546 163 580
rect 216 546 250 580
rect 303 546 337 580
rect 129 478 163 512
rect 216 478 250 512
rect 303 478 337 512
rect 129 410 163 444
rect 216 410 250 444
rect 303 410 337 444
rect 393 546 427 580
rect 393 478 427 512
rect 393 410 427 444
rect 505 546 539 580
rect 505 462 539 496
rect 505 386 539 420
rect 595 497 629 531
rect 595 386 629 420
rect 695 546 729 580
rect 695 454 729 488
rect 795 522 829 556
rect 885 506 919 540
rect 885 438 919 472
rect 997 497 1031 531
rect 997 380 1031 414
rect 1087 546 1121 580
rect 1087 474 1121 508
rect 1187 546 1221 580
rect 1187 469 1221 503
rect 1187 390 1221 424
rect 1277 546 1311 580
rect 1277 474 1311 508
rect 1367 546 1401 580
rect 1367 469 1401 503
rect 1367 390 1401 424
<< poly >>
rect 83 592 119 618
rect 347 592 383 618
rect 549 592 585 618
rect 639 592 675 618
rect 739 592 775 618
rect 839 592 875 618
rect 1041 592 1077 618
rect 1131 592 1167 618
rect 1231 592 1267 618
rect 1321 592 1357 618
rect 83 360 119 392
rect 347 360 383 392
rect 83 344 239 360
rect 83 310 121 344
rect 155 310 189 344
rect 223 310 239 344
rect 83 294 239 310
rect 281 344 383 360
rect 281 310 315 344
rect 349 310 383 344
rect 549 336 585 368
rect 639 336 675 368
rect 739 336 775 368
rect 839 336 875 368
rect 1041 336 1077 368
rect 1131 336 1167 368
rect 1231 336 1267 368
rect 1321 336 1357 368
rect 281 294 383 310
rect 431 320 675 336
rect 158 202 188 294
rect 281 252 311 294
rect 431 286 447 320
rect 481 286 515 320
rect 549 286 583 320
rect 617 300 675 320
rect 723 320 875 336
rect 617 286 669 300
rect 431 270 669 286
rect 723 286 739 320
rect 773 300 875 320
rect 952 320 1161 336
rect 773 286 882 300
rect 723 270 882 286
rect 553 222 583 270
rect 639 222 669 270
rect 766 222 796 270
rect 852 222 882 270
rect 952 286 988 320
rect 1022 286 1111 320
rect 1145 286 1161 320
rect 952 270 1161 286
rect 1231 320 1396 336
rect 1231 286 1278 320
rect 1312 286 1346 320
rect 1380 286 1396 320
rect 1231 270 1396 286
rect 952 222 982 270
rect 1038 222 1068 270
rect 1231 222 1261 270
rect 1326 222 1356 270
rect 158 48 188 74
rect 281 48 311 124
rect 553 48 583 74
rect 639 48 669 74
rect 766 48 796 74
rect 852 48 882 74
rect 952 48 982 74
rect 1038 48 1068 74
rect 1231 48 1261 74
rect 1326 48 1356 74
<< polycont >>
rect 121 310 155 344
rect 189 310 223 344
rect 315 310 349 344
rect 447 286 481 320
rect 515 286 549 320
rect 583 286 617 320
rect 739 286 773 320
rect 988 286 1022 320
rect 1111 286 1145 320
rect 1278 286 1312 320
rect 1346 286 1380 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 23 580 89 596
rect 23 546 39 580
rect 73 546 89 580
rect 23 512 89 546
rect 23 478 39 512
rect 73 478 89 512
rect 23 444 89 478
rect 23 410 39 444
rect 73 410 89 444
rect 23 394 89 410
rect 123 580 343 649
rect 123 546 129 580
rect 163 546 216 580
rect 250 546 303 580
rect 337 546 343 580
rect 123 512 343 546
rect 123 478 129 512
rect 163 478 216 512
rect 250 478 303 512
rect 337 478 343 512
rect 123 444 343 478
rect 123 410 129 444
rect 163 410 216 444
rect 250 410 303 444
rect 337 410 343 444
rect 123 394 343 410
rect 377 580 443 596
rect 377 546 393 580
rect 427 546 443 580
rect 377 512 443 546
rect 377 478 393 512
rect 427 478 443 512
rect 377 444 443 478
rect 377 410 393 444
rect 427 428 443 444
rect 499 581 745 615
rect 499 580 555 581
rect 499 546 505 580
rect 539 546 555 580
rect 679 580 745 581
rect 499 496 555 546
rect 499 462 505 496
rect 539 462 555 496
rect 427 410 465 428
rect 377 394 465 410
rect 23 260 57 394
rect 105 344 263 360
rect 105 310 121 344
rect 155 310 189 344
rect 223 310 263 344
rect 105 294 263 310
rect 299 344 365 360
rect 299 310 315 344
rect 349 310 365 344
rect 299 294 365 310
rect 431 336 465 394
rect 499 420 555 462
rect 499 386 505 420
rect 539 386 555 420
rect 499 370 555 386
rect 595 531 645 547
rect 629 497 645 531
rect 595 420 645 497
rect 679 546 695 580
rect 729 546 745 580
rect 679 488 745 546
rect 779 581 1137 615
rect 779 556 835 581
rect 779 522 795 556
rect 829 522 835 556
rect 1071 580 1137 581
rect 779 506 835 522
rect 869 540 935 547
rect 869 506 885 540
rect 919 506 935 540
rect 679 454 695 488
rect 729 472 745 488
rect 869 472 935 506
rect 729 454 885 472
rect 679 438 885 454
rect 919 438 935 472
rect 981 531 1031 547
rect 981 497 997 531
rect 629 404 645 420
rect 981 424 1031 497
rect 1071 546 1087 580
rect 1121 546 1137 580
rect 1071 508 1137 546
rect 1071 474 1087 508
rect 1121 474 1137 508
rect 1071 458 1137 474
rect 1171 580 1237 596
rect 1171 546 1187 580
rect 1221 546 1237 580
rect 1171 503 1237 546
rect 1171 469 1187 503
rect 1221 469 1237 503
rect 1171 424 1237 469
rect 1277 580 1311 649
rect 1277 508 1311 546
rect 1277 458 1311 474
rect 1351 580 1417 596
rect 1351 546 1367 580
rect 1401 546 1417 580
rect 1351 503 1417 546
rect 1351 469 1367 503
rect 1401 469 1417 503
rect 1351 424 1417 469
rect 981 414 1187 424
rect 629 386 857 404
rect 595 370 857 386
rect 823 356 857 370
rect 981 380 997 414
rect 1031 390 1187 414
rect 1221 390 1367 424
rect 1401 390 1417 424
rect 981 364 1031 380
rect 431 320 633 336
rect 431 286 447 320
rect 481 286 515 320
rect 549 286 583 320
rect 617 286 633 320
rect 431 270 633 286
rect 723 320 789 336
rect 723 286 739 320
rect 773 286 789 320
rect 723 270 789 286
rect 823 310 935 356
rect 1081 327 1223 356
rect 972 320 1223 327
rect 431 260 465 270
rect 23 226 163 260
rect 97 190 163 226
rect 324 244 465 260
rect 324 210 341 244
rect 375 210 465 244
rect 723 236 757 270
rect 823 236 857 310
rect 972 286 988 320
rect 1022 286 1111 320
rect 1145 286 1223 320
rect 972 270 1223 286
rect 1262 320 1415 356
rect 1262 286 1278 320
rect 1312 286 1346 320
rect 1380 286 1415 320
rect 1262 270 1415 286
rect 97 156 113 190
rect 147 176 163 190
rect 499 202 757 236
rect 791 210 1315 236
rect 499 176 533 202
rect 147 156 533 176
rect 791 176 807 210
rect 841 202 993 210
rect 841 176 857 202
rect 791 168 857 176
rect 1027 202 1281 210
rect 1027 176 1043 202
rect 97 142 533 156
rect 578 152 857 168
rect 97 122 163 142
rect 97 88 113 122
rect 147 88 163 122
rect 578 118 594 152
rect 628 134 857 152
rect 628 118 644 134
rect 97 72 163 88
rect 198 107 303 108
rect 198 73 215 107
rect 249 73 303 107
rect 198 17 303 73
rect 439 92 542 108
rect 439 58 473 92
rect 507 58 542 92
rect 578 70 644 118
rect 791 120 857 134
rect 680 84 755 100
rect 439 17 542 58
rect 680 50 700 84
rect 734 50 755 84
rect 791 86 807 120
rect 841 86 857 120
rect 791 70 857 86
rect 891 152 957 168
rect 891 118 907 152
rect 941 118 957 152
rect 680 17 755 50
rect 891 17 957 118
rect 993 120 1043 176
rect 1265 176 1281 202
rect 1027 86 1043 120
rect 993 70 1043 86
rect 1077 152 1231 168
rect 1077 118 1079 152
rect 1113 118 1186 152
rect 1220 118 1231 152
rect 1077 17 1231 118
rect 1265 120 1315 176
rect 1265 86 1281 120
rect 1265 70 1315 86
rect 1351 210 1417 226
rect 1351 176 1367 210
rect 1401 176 1417 210
rect 1351 120 1417 176
rect 1351 86 1367 120
rect 1401 86 1417 120
rect 1351 17 1417 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 683 1440 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 0 617 1440 649
rect 0 17 1440 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -49 1440 -17
<< labels >>
flabel pwell s 0 0 1440 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nwell s 0 617 1440 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
rlabel comment s 0 0 0 0 4 nor4bb_2
flabel metal1 s 0 617 1440 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 1440 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 C_N
port 3 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 C_N
port 3 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 D_N
port 4 nsew
flabel corelocali s 1279 316 1313 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 1375 316 1409 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 1087 316 1121 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 1183 316 1217 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 Y
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 1440 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1573848
string GDS_START 1562212
<< end >>
