magic
tech sky130A
magscale 1 2
timestamp 1601050058
<< locali >>
rect 575 357 627 493
rect 17 215 115 255
rect 153 215 248 257
rect 204 135 248 215
rect 297 215 363 257
rect 297 135 339 215
rect 397 208 479 269
rect 593 117 627 357
rect 575 51 627 117
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 18 449 85 493
rect 286 451 357 527
rect 18 325 69 449
rect 119 417 165 425
rect 391 417 441 493
rect 119 377 441 417
rect 119 359 156 377
rect 274 375 441 377
rect 491 371 541 527
rect 187 337 253 343
rect 187 325 547 337
rect 18 303 559 325
rect 18 291 253 303
rect 519 296 559 303
rect 18 17 109 170
rect 525 181 559 296
rect 505 157 559 181
rect 390 148 559 157
rect 390 123 541 148
rect 390 93 424 123
rect 164 51 424 93
rect 475 17 541 89
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 297 215 363 257 6 A1
port 1 nsew signal input
rlabel locali s 297 135 339 215 6 A1
port 1 nsew signal input
rlabel locali s 397 208 479 269 6 A2
port 2 nsew signal input
rlabel locali s 204 135 248 215 6 B1
port 3 nsew signal input
rlabel locali s 153 215 248 257 6 B1
port 3 nsew signal input
rlabel locali s 17 215 115 255 6 B2
port 4 nsew signal input
rlabel locali s 593 117 627 357 6 X
port 5 nsew signal output
rlabel locali s 575 357 627 493 6 X
port 5 nsew signal output
rlabel locali s 575 51 627 117 6 X
port 5 nsew signal output
rlabel metal1 s 0 -48 644 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 4134734
string GDS_START 4128146
<< end >>
