magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1288 561
rect 103 427 169 527
rect 17 197 66 325
rect 103 17 169 93
rect 391 367 454 527
rect 292 191 358 265
rect 764 427 822 527
rect 860 427 916 527
rect 1022 427 1185 527
rect 900 199 1087 265
rect 375 17 441 89
rect 748 17 814 106
rect 1019 17 1185 97
rect 1219 83 1271 491
rect 0 -17 1288 17
<< obsli1 >>
rect 35 393 69 493
rect 35 359 156 393
rect 122 323 156 359
rect 122 280 156 289
rect 203 391 248 493
rect 203 357 214 391
rect 203 337 248 357
rect 122 214 168 280
rect 122 161 156 214
rect 35 127 156 161
rect 35 69 69 127
rect 203 69 237 337
rect 291 333 357 483
rect 580 451 730 485
rect 494 391 551 401
rect 528 357 551 391
rect 291 299 428 333
rect 394 219 428 299
rect 494 271 551 357
rect 585 323 653 399
rect 585 289 586 323
rect 620 289 653 323
rect 585 283 653 289
rect 394 157 468 219
rect 585 207 619 283
rect 696 265 730 451
rect 950 373 988 493
rect 764 307 1185 373
rect 696 249 866 265
rect 307 153 468 157
rect 307 123 428 153
rect 543 141 619 207
rect 666 205 866 249
rect 307 69 341 123
rect 666 107 700 205
rect 1121 165 1185 307
rect 568 73 700 107
rect 848 131 1185 165
rect 848 51 918 131
<< obsli1c >>
rect 122 289 156 323
rect 214 357 248 391
rect 494 357 528 391
rect 586 289 620 323
<< metal1 >>
rect 0 496 1288 592
rect 0 -48 1288 48
<< obsm1 >>
rect 202 391 260 397
rect 202 357 214 391
rect 248 388 260 391
rect 482 391 540 397
rect 482 388 494 391
rect 248 360 494 388
rect 248 357 260 360
rect 202 351 260 357
rect 482 357 494 360
rect 528 357 540 391
rect 482 351 540 357
rect 110 323 168 329
rect 110 289 122 323
rect 156 320 168 323
rect 574 323 632 329
rect 574 320 586 323
rect 156 292 586 320
rect 156 289 168 292
rect 110 283 168 289
rect 574 289 586 292
rect 620 289 632 323
rect 574 283 632 289
<< labels >>
rlabel locali s 292 191 358 265 6 D
port 1 nsew signal input
rlabel locali s 1219 83 1271 491 6 Q
port 2 nsew signal output
rlabel locali s 900 199 1087 265 6 RESET_B
port 3 nsew signal input
rlabel locali s 17 197 66 325 6 GATE_N
port 4 nsew clock input
rlabel locali s 1019 17 1185 97 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 748 17 814 106 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 375 17 441 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 103 17 169 93 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 1288 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1288 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 1022 427 1185 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 860 427 916 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 764 427 822 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 391 367 454 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 103 427 169 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 1288 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 1288 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1288 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2637530
string GDS_START 2625950
<< end >>
