magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 191 275 263 356
rect 747 270 881 356
rect 1369 270 1435 356
rect 1550 368 1619 596
rect 1585 234 1619 368
rect 1553 88 1619 234
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 17 458 89 577
rect 129 461 185 649
rect 219 581 735 615
rect 17 213 65 458
rect 219 424 275 581
rect 99 390 275 424
rect 309 513 521 547
rect 669 542 735 581
rect 891 547 957 649
rect 1107 581 1442 615
rect 1107 547 1173 581
rect 99 247 149 390
rect 309 276 343 513
rect 377 344 421 479
rect 455 378 521 513
rect 567 508 613 524
rect 1214 513 1264 547
rect 917 508 1264 513
rect 567 479 1264 508
rect 567 474 951 479
rect 567 375 629 474
rect 679 390 851 440
rect 377 310 551 344
rect 679 341 713 390
rect 115 241 149 247
rect 17 77 81 213
rect 115 207 269 241
rect 309 233 477 276
rect 117 17 183 173
rect 219 85 269 207
rect 325 153 391 199
rect 427 187 477 233
rect 511 257 551 310
rect 631 275 713 341
rect 511 191 597 257
rect 679 225 713 275
rect 679 191 818 225
rect 917 193 951 474
rect 985 395 1067 445
rect 1214 395 1264 479
rect 985 261 1031 395
rect 1301 390 1374 500
rect 1408 424 1442 581
rect 1476 458 1510 649
rect 1408 390 1516 424
rect 1301 361 1335 390
rect 1065 295 1335 361
rect 985 227 1232 261
rect 917 157 1032 193
rect 511 153 1032 157
rect 325 123 1032 153
rect 325 119 545 123
rect 640 85 706 89
rect 219 51 706 85
rect 854 17 920 89
rect 966 70 1032 123
rect 1066 85 1132 193
rect 1166 119 1232 227
rect 1278 234 1335 295
rect 1482 334 1516 390
rect 1482 268 1551 334
rect 1482 236 1516 268
rect 1278 200 1344 234
rect 1378 202 1516 236
rect 1656 364 1706 649
rect 1378 166 1412 202
rect 1266 132 1412 166
rect 1266 85 1300 132
rect 1446 98 1517 168
rect 1066 51 1300 85
rect 1380 17 1517 98
rect 1655 17 1705 250
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
<< metal1 >>
rect 0 683 1728 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 0 617 1728 649
rect 0 17 1728 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
rect 0 -49 1728 -17
<< obsm1 >>
rect 19 273 77 282
rect 307 273 365 282
rect 19 245 365 273
rect 19 236 77 245
rect 307 236 365 245
rect 499 273 557 282
rect 979 273 1037 282
rect 499 245 1037 273
rect 499 236 557 245
rect 979 236 1037 245
<< labels >>
rlabel locali s 191 275 263 356 6 A
port 1 nsew signal input
rlabel locali s 747 270 881 356 6 B
port 2 nsew signal input
rlabel locali s 1369 270 1435 356 6 C
port 3 nsew signal input
rlabel locali s 1585 234 1619 368 6 X
port 4 nsew signal output
rlabel locali s 1553 88 1619 234 6 X
port 4 nsew signal output
rlabel locali s 1550 368 1619 596 6 X
port 4 nsew signal output
rlabel metal1 s 0 -49 1728 49 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1728 715 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1728 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 615708
string GDS_START 602552
<< end >>
