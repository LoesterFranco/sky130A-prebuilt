magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 27 391 69 493
rect 223 391 257 493
rect 27 357 257 391
rect 27 165 69 357
rect 27 131 179 165
rect 213 149 326 255
rect 489 249 534 323
rect 447 215 534 249
rect 575 83 629 265
rect 663 85 730 325
rect 833 199 901 326
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 103 425 179 527
rect 327 459 549 493
rect 327 357 361 459
rect 405 389 471 423
rect 515 393 549 459
rect 583 428 659 527
rect 735 393 769 493
rect 405 323 455 389
rect 515 359 769 393
rect 803 383 880 527
rect 107 289 455 323
rect 107 199 151 289
rect 360 169 408 289
rect 360 135 541 169
rect 18 17 85 93
rect 197 17 348 89
rect 481 59 541 135
rect 803 17 880 161
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
rlabel locali s 575 83 629 265 6 A1
port 1 nsew signal input
rlabel locali s 663 85 730 325 6 A2
port 2 nsew signal input
rlabel locali s 833 199 901 326 6 A3
port 3 nsew signal input
rlabel locali s 489 249 534 323 6 B1
port 4 nsew signal input
rlabel locali s 447 215 534 249 6 B1
port 4 nsew signal input
rlabel locali s 213 149 326 255 6 B2
port 5 nsew signal input
rlabel locali s 223 391 257 493 6 X
port 6 nsew signal output
rlabel locali s 27 391 69 493 6 X
port 6 nsew signal output
rlabel locali s 27 357 257 391 6 X
port 6 nsew signal output
rlabel locali s 27 165 69 357 6 X
port 6 nsew signal output
rlabel locali s 27 131 179 165 6 X
port 6 nsew signal output
rlabel metal1 s 0 -48 920 48 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 496 920 592 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 920 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1432050
string GDS_START 1423652
<< end >>
