magic
tech sky130A
magscale 1 2
timestamp 1599588238
<< locali >>
rect 25 226 110 360
rect 167 226 263 360
rect 679 364 751 596
rect 503 236 569 310
rect 717 226 751 364
rect 678 70 751 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 23 394 89 649
rect 211 498 277 596
rect 311 532 377 649
rect 579 532 645 649
rect 211 464 645 498
rect 211 394 357 464
rect 323 206 357 394
rect 395 364 538 430
rect 395 244 461 364
rect 611 330 645 464
rect 23 158 289 192
rect 23 70 89 158
rect 123 17 189 124
rect 223 70 289 158
rect 323 70 389 206
rect 427 202 461 244
rect 611 264 683 330
rect 427 136 544 202
rect 578 17 644 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel locali s 25 226 110 360 6 A1
port 1 nsew signal input
rlabel locali s 167 226 263 360 6 A2
port 2 nsew signal input
rlabel locali s 503 236 569 310 6 B1_N
port 3 nsew signal input
rlabel locali s 717 226 751 364 6 X
port 4 nsew signal output
rlabel locali s 679 364 751 596 6 X
port 4 nsew signal output
rlabel locali s 678 70 751 226 6 X
port 4 nsew signal output
rlabel metal1 s 0 -49 768 49 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 617 768 715 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1406212
string GDS_START 1398884
<< end >>
