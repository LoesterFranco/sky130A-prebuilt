magic
tech sky130A
magscale 1 2
timestamp 1604502729
<< locali >>
rect 113 364 190 430
rect 155 226 189 364
rect 283 270 359 430
rect 397 294 463 430
rect 505 236 577 310
rect 679 260 745 356
rect 123 70 189 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 23 532 89 649
rect 214 532 319 649
rect 553 498 645 596
rect 45 464 645 498
rect 45 330 79 464
rect 45 264 121 330
rect 553 388 645 464
rect 679 390 745 649
rect 611 226 645 388
rect 23 17 89 226
rect 223 17 289 226
rect 323 188 389 226
rect 611 192 745 226
rect 323 158 570 188
rect 323 154 645 158
rect 323 70 389 154
rect 423 17 502 120
rect 536 92 645 154
rect 679 70 745 192
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel locali s 283 270 359 430 6 A1
port 1 nsew signal input
rlabel locali s 397 294 463 430 6 A2
port 2 nsew signal input
rlabel locali s 505 236 577 310 6 A3
port 3 nsew signal input
rlabel locali s 679 260 745 356 6 B1
port 4 nsew signal input
rlabel locali s 155 226 189 364 6 X
port 5 nsew signal output
rlabel locali s 123 70 189 226 6 X
port 5 nsew signal output
rlabel locali s 113 364 190 430 6 X
port 5 nsew signal output
rlabel metal1 s 0 -49 768 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 768 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1376772
string GDS_START 1369958
<< end >>
