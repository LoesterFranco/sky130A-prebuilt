magic
tech sky130A
magscale 1 2
timestamp 1601050047
<< nwell >>
rect -38 332 3398 704
rect 2684 310 3060 332
<< pwell >>
rect 0 0 3360 49
<< scpmos >>
rect 86 464 116 592
rect 182 464 212 592
rect 266 464 296 592
rect 356 464 386 592
rect 557 464 587 592
rect 759 368 789 592
rect 849 368 879 592
rect 1051 497 1081 581
rect 1129 497 1159 581
rect 1236 453 1266 581
rect 1498 424 1528 592
rect 1582 424 1612 592
rect 1672 424 1702 592
rect 1873 424 1903 592
rect 1951 424 1981 592
rect 2058 508 2088 592
rect 2136 508 2166 592
rect 2355 392 2385 592
rect 2479 392 2509 592
rect 2563 392 2593 592
rect 2773 464 2803 592
rect 2935 368 2965 592
rect 3137 384 3167 552
rect 3244 368 3274 592
<< nmoslvt >>
rect 89 119 119 203
rect 167 119 197 203
rect 275 119 305 203
rect 353 119 383 203
rect 521 119 551 203
rect 719 82 749 230
rect 837 82 867 230
rect 1121 119 1151 203
rect 1193 119 1223 203
rect 1279 119 1309 203
rect 1507 119 1537 229
rect 1613 119 1643 229
rect 1734 119 1764 229
rect 1846 119 1876 229
rect 1924 119 1954 229
rect 2134 119 2164 203
rect 2242 119 2272 203
rect 2362 74 2392 222
rect 2448 74 2478 222
rect 2554 74 2584 222
rect 2792 138 2822 222
rect 2942 74 2972 222
rect 3140 74 3170 184
rect 3242 74 3272 222
<< ndiff >>
rect 662 218 719 230
rect 32 178 89 203
rect 32 144 44 178
rect 78 144 89 178
rect 32 119 89 144
rect 119 119 167 203
rect 197 178 275 203
rect 197 144 208 178
rect 242 144 275 178
rect 197 119 275 144
rect 305 119 353 203
rect 383 171 521 203
rect 383 137 394 171
rect 428 137 521 171
rect 383 119 521 137
rect 551 180 608 203
rect 551 146 562 180
rect 596 146 608 180
rect 551 119 608 146
rect 662 184 674 218
rect 708 184 719 218
rect 662 82 719 184
rect 749 82 837 230
rect 867 218 954 230
rect 867 184 893 218
rect 927 184 954 218
rect 867 82 954 184
rect 1064 178 1121 203
rect 1064 144 1076 178
rect 1110 144 1121 178
rect 1064 119 1121 144
rect 1151 119 1193 203
rect 1223 180 1279 203
rect 1223 146 1234 180
rect 1268 146 1279 180
rect 1223 119 1279 146
rect 1309 170 1380 203
rect 1309 136 1335 170
rect 1369 136 1380 170
rect 1309 119 1380 136
rect 1434 124 1507 229
rect 764 48 776 82
rect 810 48 822 82
rect 764 36 822 48
rect 1434 90 1446 124
rect 1480 119 1507 124
rect 1537 188 1613 229
rect 1537 154 1568 188
rect 1602 154 1613 188
rect 1537 119 1613 154
rect 1643 188 1734 229
rect 1643 154 1668 188
rect 1702 154 1734 188
rect 1643 119 1734 154
rect 1764 186 1846 229
rect 1764 152 1775 186
rect 1809 152 1846 186
rect 1764 119 1846 152
rect 1876 119 1924 229
rect 1954 203 2112 229
rect 2312 203 2362 222
rect 1954 191 2134 203
rect 1954 157 1965 191
rect 1999 157 2066 191
rect 2100 157 2134 191
rect 1954 119 2134 157
rect 2164 119 2242 203
rect 2272 119 2362 203
rect 1480 90 1492 119
rect 1434 78 1492 90
rect 2287 82 2362 119
rect 2287 48 2300 82
rect 2334 74 2362 82
rect 2392 192 2448 222
rect 2392 158 2403 192
rect 2437 158 2448 192
rect 2392 116 2448 158
rect 2392 82 2403 116
rect 2437 82 2448 116
rect 2392 74 2448 82
rect 2478 172 2554 222
rect 2478 138 2509 172
rect 2543 138 2554 172
rect 2478 74 2554 138
rect 2584 108 2657 222
rect 2735 197 2792 222
rect 2735 163 2747 197
rect 2781 163 2792 197
rect 2735 138 2792 163
rect 2822 138 2942 222
rect 2871 120 2942 138
rect 2584 74 2611 108
rect 2645 74 2657 108
rect 2871 86 2890 120
rect 2924 86 2942 120
rect 2871 74 2942 86
rect 2972 210 3029 222
rect 2972 176 2983 210
rect 3017 176 3029 210
rect 3185 194 3242 222
rect 3185 184 3197 194
rect 2972 120 3029 176
rect 2972 86 2983 120
rect 3017 86 3029 120
rect 2972 74 3029 86
rect 3083 146 3140 184
rect 3083 112 3095 146
rect 3129 112 3140 146
rect 3083 74 3140 112
rect 3170 160 3197 184
rect 3231 160 3242 194
rect 3170 120 3242 160
rect 3170 86 3197 120
rect 3231 86 3242 120
rect 3170 74 3242 86
rect 3272 194 3329 222
rect 3272 160 3283 194
rect 3317 160 3329 194
rect 3272 120 3329 160
rect 3272 86 3283 120
rect 3317 86 3329 120
rect 3272 74 3329 86
rect 2334 48 2347 74
rect 2599 62 2657 74
rect 2287 36 2347 48
<< pdiff >>
rect 2184 628 2242 639
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 510 86 546
rect 27 476 39 510
rect 73 476 86 510
rect 27 464 86 476
rect 116 579 182 592
rect 116 545 129 579
rect 163 545 182 579
rect 116 511 182 545
rect 116 477 129 511
rect 163 477 182 511
rect 116 464 182 477
rect 212 464 266 592
rect 296 520 356 592
rect 296 486 309 520
rect 343 486 356 520
rect 296 464 356 486
rect 386 580 444 592
rect 386 546 399 580
rect 433 546 444 580
rect 386 510 444 546
rect 386 476 399 510
rect 433 476 444 510
rect 386 464 444 476
rect 498 580 557 592
rect 498 546 510 580
rect 544 546 557 580
rect 498 510 557 546
rect 498 476 510 510
rect 544 476 557 510
rect 498 464 557 476
rect 587 580 646 592
rect 587 546 600 580
rect 634 546 646 580
rect 587 510 646 546
rect 587 476 600 510
rect 634 476 646 510
rect 587 464 646 476
rect 700 580 759 592
rect 700 546 712 580
rect 746 546 759 580
rect 700 510 759 546
rect 700 476 712 510
rect 746 476 759 510
rect 700 440 759 476
rect 700 406 712 440
rect 746 406 759 440
rect 700 368 759 406
rect 789 580 849 592
rect 789 546 802 580
rect 836 546 849 580
rect 789 508 849 546
rect 789 474 802 508
rect 836 474 849 508
rect 789 368 849 474
rect 879 580 938 592
rect 2184 594 2196 628
rect 2230 594 2242 628
rect 2403 628 2461 639
rect 2184 592 2242 594
rect 2403 594 2415 628
rect 2449 594 2461 628
rect 2403 592 2461 594
rect 879 546 892 580
rect 926 546 938 580
rect 879 499 938 546
rect 879 465 892 499
rect 926 465 938 499
rect 992 556 1051 581
rect 992 522 1004 556
rect 1038 522 1051 556
rect 992 497 1051 522
rect 1081 497 1129 581
rect 1159 515 1236 581
rect 1159 497 1189 515
rect 879 418 938 465
rect 879 384 892 418
rect 926 384 938 418
rect 879 368 938 384
rect 1177 481 1189 497
rect 1223 481 1236 515
rect 1177 453 1236 481
rect 1266 521 1335 581
rect 1266 487 1289 521
rect 1323 487 1335 521
rect 1266 453 1335 487
rect 1405 573 1498 592
rect 1405 539 1450 573
rect 1484 539 1498 573
rect 1405 424 1498 539
rect 1528 424 1582 592
rect 1612 580 1672 592
rect 1612 546 1625 580
rect 1659 546 1672 580
rect 1612 424 1672 546
rect 1702 580 1760 592
rect 1702 546 1715 580
rect 1749 546 1760 580
rect 1702 512 1760 546
rect 1702 478 1715 512
rect 1749 478 1760 512
rect 1702 424 1760 478
rect 1814 544 1873 592
rect 1814 510 1826 544
rect 1860 510 1873 544
rect 1814 424 1873 510
rect 1903 424 1951 592
rect 1981 580 2058 592
rect 1981 546 1994 580
rect 2028 546 2058 580
rect 1981 508 2058 546
rect 2088 508 2136 592
rect 2166 508 2242 592
rect 2296 578 2355 592
rect 2296 544 2308 578
rect 2342 544 2355 578
rect 1981 472 2040 508
rect 1981 438 1994 472
rect 2028 438 2040 472
rect 1981 424 2040 438
rect 2296 392 2355 544
rect 2385 392 2479 592
rect 2509 392 2563 592
rect 2593 580 2652 592
rect 2593 546 2606 580
rect 2640 546 2652 580
rect 2593 462 2652 546
rect 2593 428 2606 462
rect 2640 428 2652 462
rect 2593 392 2652 428
rect 2720 464 2773 592
rect 2803 554 2935 592
rect 2803 520 2816 554
rect 2850 520 2888 554
rect 2922 520 2935 554
rect 2803 464 2935 520
rect 2720 404 2750 464
rect 2720 392 2822 404
rect 2720 358 2757 392
rect 2791 358 2822 392
rect 2720 346 2822 358
rect 2882 368 2935 464
rect 2965 580 3024 592
rect 2965 546 2978 580
rect 3012 546 3024 580
rect 3185 580 3244 592
rect 3185 552 3197 580
rect 2965 497 3024 546
rect 2965 463 2978 497
rect 3012 463 3024 497
rect 2965 414 3024 463
rect 2965 380 2978 414
rect 3012 380 3024 414
rect 3078 540 3137 552
rect 3078 506 3090 540
rect 3124 506 3137 540
rect 3078 430 3137 506
rect 3078 396 3090 430
rect 3124 396 3137 430
rect 3078 384 3137 396
rect 3167 546 3197 552
rect 3231 546 3244 580
rect 3167 505 3244 546
rect 3167 471 3197 505
rect 3231 471 3244 505
rect 3167 430 3244 471
rect 3167 396 3197 430
rect 3231 396 3244 430
rect 3167 384 3244 396
rect 2965 368 3024 380
rect 3185 368 3244 384
rect 3274 580 3333 592
rect 3274 546 3287 580
rect 3321 546 3333 580
rect 3274 497 3333 546
rect 3274 463 3287 497
rect 3321 463 3333 497
rect 3274 414 3333 463
rect 3274 380 3287 414
rect 3321 380 3333 414
rect 3274 368 3333 380
<< ndiffc >>
rect 44 144 78 178
rect 208 144 242 178
rect 394 137 428 171
rect 562 146 596 180
rect 674 184 708 218
rect 893 184 927 218
rect 1076 144 1110 178
rect 1234 146 1268 180
rect 1335 136 1369 170
rect 776 48 810 82
rect 1446 90 1480 124
rect 1568 154 1602 188
rect 1668 154 1702 188
rect 1775 152 1809 186
rect 1965 157 1999 191
rect 2066 157 2100 191
rect 2300 48 2334 82
rect 2403 158 2437 192
rect 2403 82 2437 116
rect 2509 138 2543 172
rect 2747 163 2781 197
rect 2611 74 2645 108
rect 2890 86 2924 120
rect 2983 176 3017 210
rect 2983 86 3017 120
rect 3095 112 3129 146
rect 3197 160 3231 194
rect 3197 86 3231 120
rect 3283 160 3317 194
rect 3283 86 3317 120
<< pdiffc >>
rect 39 546 73 580
rect 39 476 73 510
rect 129 545 163 579
rect 129 477 163 511
rect 309 486 343 520
rect 399 546 433 580
rect 399 476 433 510
rect 510 546 544 580
rect 510 476 544 510
rect 600 546 634 580
rect 600 476 634 510
rect 712 546 746 580
rect 712 476 746 510
rect 712 406 746 440
rect 802 546 836 580
rect 802 474 836 508
rect 2196 594 2230 628
rect 2415 594 2449 628
rect 892 546 926 580
rect 892 465 926 499
rect 1004 522 1038 556
rect 892 384 926 418
rect 1189 481 1223 515
rect 1289 487 1323 521
rect 1450 539 1484 573
rect 1625 546 1659 580
rect 1715 546 1749 580
rect 1715 478 1749 512
rect 1826 510 1860 544
rect 1994 546 2028 580
rect 2308 544 2342 578
rect 1994 438 2028 472
rect 2606 546 2640 580
rect 2606 428 2640 462
rect 2816 520 2850 554
rect 2888 520 2922 554
rect 2757 358 2791 392
rect 2978 546 3012 580
rect 2978 463 3012 497
rect 2978 380 3012 414
rect 3090 506 3124 540
rect 3090 396 3124 430
rect 3197 546 3231 580
rect 3197 471 3231 505
rect 3197 396 3231 430
rect 3287 546 3321 580
rect 3287 463 3321 497
rect 3287 380 3321 414
<< poly >>
rect 86 592 116 618
rect 182 592 212 618
rect 266 592 296 618
rect 356 592 386 618
rect 557 592 587 618
rect 759 592 789 618
rect 849 592 879 618
rect 86 449 116 464
rect 182 449 212 464
rect 266 449 296 464
rect 356 449 386 464
rect 557 449 587 464
rect 83 375 119 449
rect 179 375 215 449
rect 266 423 299 449
rect 44 359 119 375
rect 44 325 60 359
rect 94 325 119 359
rect 44 291 119 325
rect 44 257 60 291
rect 94 257 119 291
rect 44 241 119 257
rect 161 359 227 375
rect 161 325 177 359
rect 211 325 227 359
rect 161 291 227 325
rect 269 362 299 423
rect 353 440 389 449
rect 554 440 590 449
rect 353 410 441 440
rect 554 410 646 440
rect 411 362 441 410
rect 269 346 363 362
rect 269 312 313 346
rect 347 312 363 346
rect 269 296 363 312
rect 411 346 568 362
rect 411 312 518 346
rect 552 312 568 346
rect 411 296 568 312
rect 161 257 177 291
rect 211 257 227 291
rect 161 241 227 257
rect 89 203 119 241
rect 167 203 197 241
rect 275 203 305 296
rect 411 248 441 296
rect 616 248 646 410
rect 1051 581 1081 607
rect 1129 581 1159 607
rect 1236 581 1266 607
rect 1498 592 1528 618
rect 1582 592 1612 618
rect 1672 592 1702 618
rect 1873 592 1903 618
rect 1951 592 1981 618
rect 2058 592 2088 618
rect 2136 592 2166 618
rect 2355 592 2385 618
rect 2479 592 2509 618
rect 2563 592 2593 618
rect 2773 592 2803 618
rect 2935 592 2965 618
rect 3244 592 3274 618
rect 1051 482 1081 497
rect 1129 482 1159 497
rect 1048 459 1084 482
rect 977 443 1084 459
rect 977 409 993 443
rect 1027 429 1084 443
rect 1027 409 1043 429
rect 759 353 789 368
rect 849 353 879 368
rect 756 336 792 353
rect 694 320 792 336
rect 846 334 882 353
rect 977 351 1043 409
rect 1126 381 1162 482
rect 1236 438 1266 453
rect 1085 365 1162 381
rect 694 286 710 320
rect 744 286 792 320
rect 694 270 792 286
rect 834 318 900 334
rect 834 284 850 318
rect 884 284 900 318
rect 353 218 441 248
rect 521 218 646 248
rect 719 230 749 270
rect 834 268 900 284
rect 977 273 1007 351
rect 1085 331 1101 365
rect 1135 351 1162 365
rect 1204 408 1269 438
rect 2058 493 2088 508
rect 2136 493 2166 508
rect 2055 436 2091 493
rect 2133 476 2169 493
rect 2133 460 2199 476
rect 1498 409 1528 424
rect 1582 409 1612 424
rect 1672 409 1702 424
rect 1873 409 1903 424
rect 1951 409 1981 424
rect 1135 331 1151 351
rect 1085 315 1151 331
rect 837 230 867 268
rect 977 243 1151 273
rect 1204 248 1234 408
rect 1384 369 1450 385
rect 1276 344 1342 360
rect 1276 310 1292 344
rect 1326 310 1342 344
rect 1276 294 1342 310
rect 1384 335 1400 369
rect 1434 335 1450 369
rect 1384 301 1450 335
rect 353 203 383 218
rect 521 203 551 218
rect 89 93 119 119
rect 167 51 197 119
rect 275 93 305 119
rect 353 93 383 119
rect 521 51 551 119
rect 1121 203 1151 243
rect 1193 218 1234 248
rect 1193 203 1223 218
rect 1279 203 1309 294
rect 1384 267 1400 301
rect 1434 281 1450 301
rect 1495 281 1531 409
rect 1579 324 1615 409
rect 1669 402 1705 409
rect 1669 376 1798 402
rect 1870 392 1906 409
rect 1669 372 1748 376
rect 1732 342 1748 372
rect 1782 342 1798 376
rect 1732 326 1798 342
rect 1840 376 1906 392
rect 1840 342 1856 376
rect 1890 342 1906 376
rect 1840 326 1906 342
rect 1948 388 1984 409
rect 1948 372 2014 388
rect 1948 338 1964 372
rect 1998 338 2014 372
rect 1579 308 1686 324
rect 1434 267 1537 281
rect 1384 251 1537 267
rect 1579 274 1636 308
rect 1670 274 1686 308
rect 1579 258 1686 274
rect 1507 229 1537 251
rect 1613 229 1643 258
rect 1734 229 1764 326
rect 1846 229 1876 326
rect 1948 322 2014 338
rect 2056 274 2086 436
rect 2133 426 2149 460
rect 2183 440 2199 460
rect 2183 426 2272 440
rect 2133 410 2272 426
rect 1924 244 2086 274
rect 2134 299 2200 315
rect 2134 265 2150 299
rect 2184 265 2200 299
rect 2134 249 2200 265
rect 1924 229 1954 244
rect 1121 93 1151 119
rect 719 56 749 82
rect 167 21 551 51
rect 837 51 867 82
rect 1193 51 1223 119
rect 1279 93 1309 119
rect 2134 203 2164 249
rect 2242 203 2272 410
rect 2773 449 2803 464
rect 2770 419 2867 449
rect 2355 377 2385 392
rect 2479 377 2509 392
rect 2563 377 2593 392
rect 2352 360 2388 377
rect 2326 344 2392 360
rect 2326 310 2342 344
rect 2376 310 2392 344
rect 2476 310 2512 377
rect 2560 360 2596 377
rect 2326 294 2392 310
rect 2362 222 2392 294
rect 2440 294 2512 310
rect 2440 260 2456 294
rect 2490 280 2512 294
rect 2554 344 2688 360
rect 2554 310 2570 344
rect 2604 310 2638 344
rect 2672 310 2688 344
rect 2837 310 2867 419
rect 3137 552 3167 578
rect 3137 369 3167 384
rect 2935 353 2965 368
rect 2932 326 2968 353
rect 2921 314 2987 326
rect 3134 314 3170 369
rect 3244 353 3274 368
rect 2921 310 3170 314
rect 3241 310 3277 353
rect 2554 294 2688 310
rect 2792 294 2879 310
rect 2490 260 2506 280
rect 2440 244 2506 260
rect 2448 222 2478 244
rect 2554 222 2584 294
rect 2792 260 2829 294
rect 2863 260 2879 294
rect 2921 276 2937 310
rect 2971 276 3170 310
rect 2921 260 3170 276
rect 2792 244 2879 260
rect 2792 222 2822 244
rect 2942 222 2972 260
rect 1507 93 1537 119
rect 1613 93 1643 119
rect 1734 93 1764 119
rect 1846 93 1876 119
rect 1924 51 1954 119
rect 2134 93 2164 119
rect 2242 93 2272 119
rect 837 21 1954 51
rect 2792 112 2822 138
rect 3140 184 3170 260
rect 3212 294 3278 310
rect 3212 260 3228 294
rect 3262 260 3278 294
rect 3212 244 3278 260
rect 3242 222 3272 244
rect 2362 48 2392 74
rect 2448 48 2478 74
rect 2554 48 2584 74
rect 2942 48 2972 74
rect 3140 48 3170 74
rect 3242 48 3272 74
<< polycont >>
rect 60 325 94 359
rect 60 257 94 291
rect 177 325 211 359
rect 313 312 347 346
rect 518 312 552 346
rect 177 257 211 291
rect 993 409 1027 443
rect 710 286 744 320
rect 850 284 884 318
rect 1101 331 1135 365
rect 1292 310 1326 344
rect 1400 335 1434 369
rect 1400 267 1434 301
rect 1748 342 1782 376
rect 1856 342 1890 376
rect 1964 338 1998 372
rect 1636 274 1670 308
rect 2149 426 2183 460
rect 2150 265 2184 299
rect 2342 310 2376 344
rect 2456 260 2490 294
rect 2570 310 2604 344
rect 2638 310 2672 344
rect 2829 260 2863 294
rect 2937 276 2971 310
rect 3228 260 3262 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3360 683
rect 23 580 79 596
rect 23 546 39 580
rect 73 546 79 580
rect 23 510 79 546
rect 23 476 39 510
rect 73 476 79 510
rect 113 579 179 649
rect 113 545 129 579
rect 163 545 179 579
rect 113 511 179 545
rect 113 477 129 511
rect 163 477 179 511
rect 213 581 449 615
rect 23 443 79 476
rect 213 443 247 581
rect 383 580 449 581
rect 293 520 343 547
rect 293 486 309 520
rect 293 460 343 486
rect 383 546 399 580
rect 433 546 449 580
rect 383 510 449 546
rect 383 476 399 510
rect 433 476 449 510
rect 383 464 449 476
rect 494 580 544 649
rect 494 546 510 580
rect 494 510 544 546
rect 494 476 510 510
rect 494 460 544 476
rect 578 580 650 596
rect 578 546 600 580
rect 634 546 650 580
rect 578 510 650 546
rect 578 476 600 510
rect 634 476 650 510
rect 578 460 650 476
rect 696 580 746 596
rect 696 546 712 580
rect 696 510 746 546
rect 696 476 712 510
rect 23 409 247 443
rect 309 430 343 460
rect 309 396 431 430
rect 25 359 110 375
rect 25 325 60 359
rect 94 325 110 359
rect 25 291 110 325
rect 25 257 60 291
rect 94 257 110 291
rect 25 241 110 257
rect 161 359 263 375
rect 161 325 177 359
rect 211 325 263 359
rect 161 291 263 325
rect 297 346 363 362
rect 297 312 313 346
rect 347 312 363 346
rect 297 296 363 312
rect 161 257 177 291
rect 211 257 263 291
rect 397 262 431 396
rect 578 362 612 460
rect 696 440 746 476
rect 786 580 836 649
rect 786 546 802 580
rect 786 508 836 546
rect 786 474 802 508
rect 786 458 836 474
rect 876 580 956 596
rect 876 546 892 580
rect 926 546 956 580
rect 876 499 956 546
rect 876 465 892 499
rect 926 465 956 499
rect 1004 556 1054 649
rect 1038 522 1054 556
rect 1004 493 1054 522
rect 1088 581 1501 615
rect 696 406 712 440
rect 746 406 828 424
rect 696 390 828 406
rect 502 346 612 362
rect 502 312 518 346
rect 552 312 612 346
rect 502 296 612 312
rect 161 241 263 257
rect 297 228 512 262
rect 297 207 331 228
rect 28 178 94 207
rect 28 144 44 178
rect 78 144 94 178
rect 28 17 94 144
rect 192 178 331 207
rect 192 144 208 178
rect 242 173 331 178
rect 242 144 258 173
rect 192 115 258 144
rect 378 171 444 194
rect 378 137 394 171
rect 428 137 444 171
rect 378 17 444 137
rect 478 85 512 228
rect 546 180 612 296
rect 694 320 760 356
rect 694 286 710 320
rect 744 286 760 320
rect 694 270 760 286
rect 794 334 828 390
rect 876 418 956 465
rect 1088 459 1122 581
rect 1385 573 1501 581
rect 876 384 892 418
rect 926 384 956 418
rect 990 443 1122 459
rect 1173 515 1239 547
rect 1173 481 1189 515
rect 1223 481 1239 515
rect 1173 449 1239 481
rect 1273 521 1339 547
rect 1385 539 1450 573
rect 1484 564 1501 573
rect 1625 580 1659 649
rect 1484 539 1586 564
rect 1385 530 1586 539
rect 1625 530 1659 546
rect 1699 580 1766 596
rect 1699 546 1715 580
rect 1749 546 1766 580
rect 1273 487 1289 521
rect 1323 496 1339 521
rect 1552 496 1586 530
rect 1699 512 1766 546
rect 1699 496 1715 512
rect 1323 487 1518 496
rect 1273 462 1518 487
rect 990 409 993 443
rect 1027 425 1122 443
rect 1205 428 1239 449
rect 1027 409 1043 425
rect 990 393 1043 409
rect 1205 394 1450 428
rect 876 368 956 384
rect 922 344 956 368
rect 1081 365 1151 381
rect 1081 350 1101 365
rect 1135 360 1151 365
rect 1384 369 1450 394
rect 1081 344 1087 350
rect 794 318 888 334
rect 794 284 850 318
rect 884 284 888 318
rect 794 268 888 284
rect 922 316 1087 344
rect 1135 344 1342 360
rect 1135 331 1292 344
rect 1121 316 1292 331
rect 922 310 1292 316
rect 1326 310 1342 344
rect 794 234 828 268
rect 922 234 958 310
rect 1276 294 1342 310
rect 1384 335 1400 369
rect 1434 335 1450 369
rect 1384 301 1450 335
rect 658 218 828 234
rect 658 184 674 218
rect 708 184 828 218
rect 862 218 958 234
rect 862 184 893 218
rect 927 184 958 218
rect 992 241 1194 275
rect 1384 267 1400 301
rect 1434 267 1450 301
rect 1384 260 1450 267
rect 546 146 562 180
rect 596 146 612 180
rect 992 150 1026 241
rect 546 119 612 146
rect 646 116 1026 150
rect 1060 178 1126 207
rect 1060 144 1076 178
rect 1110 144 1126 178
rect 646 85 680 116
rect 478 51 680 85
rect 760 48 776 82
rect 810 48 826 82
rect 760 17 826 48
rect 1060 17 1126 144
rect 1160 85 1194 241
rect 1234 226 1450 260
rect 1234 180 1284 226
rect 1484 192 1518 462
rect 1268 146 1284 180
rect 1234 119 1284 146
rect 1319 170 1518 192
rect 1319 136 1335 170
rect 1369 158 1518 170
rect 1552 478 1715 496
rect 1749 478 1766 512
rect 1810 544 1876 649
rect 2180 628 2246 649
rect 1810 510 1826 544
rect 1860 510 1876 544
rect 1810 494 1876 510
rect 1978 580 2044 596
rect 2180 594 2196 628
rect 2230 594 2246 628
rect 2399 628 2465 649
rect 1978 546 1994 580
rect 2028 546 2044 580
rect 2292 578 2358 596
rect 2399 594 2415 628
rect 2449 594 2465 628
rect 2292 560 2308 578
rect 1552 462 1766 478
rect 1552 216 1586 462
rect 1732 460 1766 462
rect 1978 472 2044 546
rect 1657 424 1698 428
rect 1732 426 1906 460
rect 1657 390 1663 424
rect 1697 392 1698 424
rect 1697 390 1798 392
rect 1657 376 1798 390
rect 1657 358 1748 376
rect 1732 342 1748 358
rect 1782 342 1798 376
rect 1732 326 1798 342
rect 1840 376 1906 426
rect 1978 438 1994 472
rect 2028 456 2044 472
rect 2133 544 2308 560
rect 2342 560 2358 578
rect 2590 580 2656 596
rect 2590 560 2606 580
rect 2342 546 2606 560
rect 2640 546 2656 580
rect 2342 544 2656 546
rect 2133 526 2656 544
rect 2133 460 2199 526
rect 2028 438 2082 456
rect 1978 422 2082 438
rect 1840 342 1856 376
rect 1890 342 1906 376
rect 1840 326 1906 342
rect 1945 372 2014 388
rect 1945 350 1964 372
rect 1620 308 1686 324
rect 1620 274 1636 308
rect 1670 292 1686 308
rect 1945 316 1951 350
rect 1998 338 2014 372
rect 2048 379 2082 422
rect 2133 426 2149 460
rect 2183 426 2199 460
rect 2133 413 2199 426
rect 2234 458 2556 492
rect 2234 379 2268 458
rect 2048 345 2268 379
rect 1985 316 2014 338
rect 1945 311 2014 316
rect 1945 299 2200 311
rect 1670 274 1911 292
rect 1620 258 1911 274
rect 1552 188 1618 216
rect 1369 136 1385 158
rect 1319 85 1385 136
rect 1552 154 1568 188
rect 1602 154 1618 188
rect 1160 51 1385 85
rect 1430 90 1446 124
rect 1480 90 1496 124
rect 1552 119 1618 154
rect 1652 188 1718 216
rect 1652 154 1668 188
rect 1702 154 1718 188
rect 1430 85 1496 90
rect 1652 85 1718 154
rect 1430 51 1718 85
rect 1759 186 1825 216
rect 1759 152 1775 186
rect 1809 152 1825 186
rect 1759 17 1825 152
rect 1877 107 1911 258
rect 1945 265 2150 299
rect 2184 265 2200 299
rect 1945 252 2200 265
rect 2234 218 2268 345
rect 2326 390 2335 424
rect 2369 390 2392 424
rect 2326 344 2392 390
rect 2522 378 2556 458
rect 2590 476 2656 526
rect 2800 554 2938 649
rect 2800 520 2816 554
rect 2850 520 2888 554
rect 2922 520 2938 554
rect 2800 510 2938 520
rect 2978 580 3055 596
rect 3012 546 3055 580
rect 3181 580 3231 649
rect 2978 497 3055 546
rect 2590 462 2944 476
rect 2590 428 2606 462
rect 2640 442 2944 462
rect 2640 428 2656 442
rect 2590 412 2656 428
rect 2722 392 2826 408
rect 2522 344 2688 378
rect 2326 310 2342 344
rect 2376 310 2392 344
rect 2554 310 2570 344
rect 2604 310 2638 344
rect 2672 310 2688 344
rect 2326 294 2392 310
rect 2440 294 2506 310
rect 2554 294 2688 310
rect 2722 358 2757 392
rect 2791 358 2826 392
rect 2440 260 2456 294
rect 2490 260 2506 294
rect 2722 260 2756 358
rect 2910 326 2944 442
rect 3012 463 3055 497
rect 2978 414 3055 463
rect 3012 380 3055 414
rect 2978 364 3055 380
rect 2910 310 2987 326
rect 2815 294 2876 310
rect 2815 260 2829 294
rect 2863 260 2876 294
rect 1949 191 2268 218
rect 1949 157 1965 191
rect 1999 157 2066 191
rect 2100 184 2268 191
rect 2302 226 2781 260
rect 2815 238 2876 260
rect 2910 276 2937 310
rect 2971 276 2987 310
rect 2910 260 2987 276
rect 2100 157 2116 184
rect 1949 141 2116 157
rect 2302 150 2336 226
rect 2747 197 2781 226
rect 2910 204 2944 260
rect 3021 226 3055 364
rect 2150 116 2336 150
rect 2387 158 2403 192
rect 2437 158 2453 192
rect 2387 116 2453 158
rect 2493 172 2713 192
rect 2493 138 2509 172
rect 2543 158 2713 172
rect 2543 138 2559 158
rect 2493 119 2559 138
rect 2150 107 2184 116
rect 1877 73 2184 107
rect 2387 82 2403 116
rect 2437 85 2453 116
rect 2595 108 2645 124
rect 2595 85 2611 108
rect 2437 82 2611 85
rect 2283 48 2300 82
rect 2334 48 2351 82
rect 2387 74 2611 82
rect 2387 51 2645 74
rect 2679 100 2713 158
rect 2747 134 2781 163
rect 2815 170 2944 204
rect 2983 210 3055 226
rect 3017 176 3055 210
rect 2815 100 2849 170
rect 2679 66 2849 100
rect 2883 120 2947 136
rect 2883 86 2890 120
rect 2924 86 2947 120
rect 2283 17 2351 48
rect 2883 17 2947 86
rect 2983 120 3055 176
rect 3017 86 3055 120
rect 2983 70 3055 86
rect 3090 540 3140 556
rect 3124 506 3140 540
rect 3090 430 3140 506
rect 3124 396 3140 430
rect 3090 310 3140 396
rect 3181 546 3197 580
rect 3181 505 3231 546
rect 3181 471 3197 505
rect 3181 430 3231 471
rect 3181 396 3197 430
rect 3181 380 3231 396
rect 3271 580 3343 596
rect 3271 546 3287 580
rect 3321 546 3343 580
rect 3271 497 3343 546
rect 3271 463 3287 497
rect 3321 463 3343 497
rect 3271 414 3343 463
rect 3271 380 3287 414
rect 3321 380 3343 414
rect 3271 364 3343 380
rect 3090 294 3275 310
rect 3090 260 3228 294
rect 3262 260 3275 294
rect 3090 244 3275 260
rect 3090 146 3145 244
rect 3309 210 3343 364
rect 3090 112 3095 146
rect 3129 112 3145 146
rect 3090 70 3145 112
rect 3181 194 3231 210
rect 3181 160 3197 194
rect 3181 120 3231 160
rect 3181 86 3197 120
rect 3181 17 3231 86
rect 3267 194 3343 210
rect 3267 160 3283 194
rect 3317 160 3343 194
rect 3267 120 3343 160
rect 3267 86 3283 120
rect 3317 86 3343 120
rect 3267 70 3343 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3360 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 3199 649 3233 683
rect 3295 649 3329 683
rect 1087 331 1101 350
rect 1101 331 1121 350
rect 1087 316 1121 331
rect 1663 390 1697 424
rect 1951 338 1964 350
rect 1964 338 1985 350
rect 1951 316 1985 338
rect 2335 390 2369 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
<< metal1 >>
rect 0 683 3360 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3360 683
rect 0 617 3360 649
rect 1651 424 1709 430
rect 1651 390 1663 424
rect 1697 421 1709 424
rect 2323 424 2381 430
rect 2323 421 2335 424
rect 1697 393 2335 421
rect 1697 390 1709 393
rect 1651 384 1709 390
rect 2323 390 2335 393
rect 2369 390 2381 424
rect 2323 384 2381 390
rect 1075 350 1133 356
rect 1075 316 1087 350
rect 1121 347 1133 350
rect 1939 350 1997 356
rect 1939 347 1951 350
rect 1121 319 1951 347
rect 1121 316 1133 319
rect 1075 310 1133 316
rect 1939 316 1951 319
rect 1985 316 1997 350
rect 1939 310 1997 316
rect 0 17 3360 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3360 17
rect 0 -49 3360 -17
<< labels >>
rlabel comment s 0 0 0 0 4 sdfbbn_1
flabel pwell s 0 0 3360 49 0 FreeSans 200 0 0 0 VNB
port 8 nsew
flabel nbase s 0 617 3360 666 0 FreeSans 200 0 0 0 VPB
port 9 nsew
flabel metal1 s 2335 390 2369 424 0 FreeSans 340 0 0 0 SET_B
port 6 nsew
flabel metal1 s 0 617 3360 666 0 FreeSans 340 0 0 0 VPWR
port 10 nsew
flabel metal1 s 0 0 3360 49 0 FreeSans 340 0 0 0 VGND
port 7 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 SCD
port 4 nsew
flabel corelocali s 3007 390 3041 424 0 FreeSans 340 0 0 0 Q_N
port 12 nsew
flabel corelocali s 3007 464 3041 498 0 FreeSans 340 0 0 0 Q_N
port 12 nsew
flabel corelocali s 3007 538 3041 572 0 FreeSans 340 0 0 0 Q_N
port 12 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 CLK_N
port 1 nsew
flabel corelocali s 2815 242 2849 276 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew
flabel corelocali s 3295 390 3329 424 0 FreeSans 340 0 0 0 Q
port 11 nsew
flabel corelocali s 3295 464 3329 498 0 FreeSans 340 0 0 0 Q
port 11 nsew
flabel corelocali s 3295 538 3329 572 0 FreeSans 340 0 0 0 Q
port 11 nsew
<< properties >>
string FIXED_BBOX 0 0 3360 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 964808
string GDS_START 940362
<< end >>
