magic
tech sky130A
magscale 1 2
timestamp 1604502705
<< nwell >>
rect -38 332 614 704
<< pwell >>
rect 0 0 576 49
<< scnmos >>
rect 125 112 155 222
rect 233 74 263 222
rect 327 74 357 222
rect 441 74 471 222
<< pmoshvt >>
rect 116 368 146 536
rect 230 368 260 592
rect 314 368 344 592
rect 428 368 458 592
<< ndiff >>
rect 27 186 125 222
rect 27 152 80 186
rect 114 152 125 186
rect 27 112 125 152
rect 155 199 233 222
rect 155 165 182 199
rect 216 165 233 199
rect 155 120 233 165
rect 155 112 182 120
rect 170 86 182 112
rect 216 86 233 120
rect 170 74 233 86
rect 263 210 327 222
rect 263 176 282 210
rect 316 176 327 210
rect 263 120 327 176
rect 263 86 282 120
rect 316 86 327 120
rect 263 74 327 86
rect 357 152 441 222
rect 357 118 382 152
rect 416 118 441 152
rect 357 74 441 118
rect 471 210 528 222
rect 471 176 482 210
rect 516 176 528 210
rect 471 120 528 176
rect 471 86 482 120
rect 516 86 528 120
rect 471 74 528 86
<< pdiff >>
rect 171 580 230 592
rect 171 546 183 580
rect 217 546 230 580
rect 171 536 230 546
rect 57 524 116 536
rect 57 490 69 524
rect 103 490 116 524
rect 57 414 116 490
rect 57 380 69 414
rect 103 380 116 414
rect 57 368 116 380
rect 146 508 230 536
rect 146 474 183 508
rect 217 474 230 508
rect 146 368 230 474
rect 260 368 314 592
rect 344 368 428 592
rect 458 580 517 592
rect 458 546 471 580
rect 505 546 517 580
rect 458 508 517 546
rect 458 474 471 508
rect 505 474 517 508
rect 458 368 517 474
<< ndiffc >>
rect 80 152 114 186
rect 182 165 216 199
rect 182 86 216 120
rect 282 176 316 210
rect 282 86 316 120
rect 382 118 416 152
rect 482 176 516 210
rect 482 86 516 120
<< pdiffc >>
rect 183 546 217 580
rect 69 490 103 524
rect 69 380 103 414
rect 183 474 217 508
rect 471 546 505 580
rect 471 474 505 508
<< poly >>
rect 230 592 260 618
rect 314 592 344 618
rect 428 592 458 618
rect 116 536 146 562
rect 116 353 146 368
rect 230 353 260 368
rect 314 353 344 368
rect 428 353 458 368
rect 113 310 149 353
rect 227 336 263 353
rect 197 320 263 336
rect 89 294 155 310
rect 89 260 105 294
rect 139 260 155 294
rect 197 286 213 320
rect 247 286 263 320
rect 197 270 263 286
rect 311 336 347 353
rect 425 336 461 353
rect 311 320 377 336
rect 311 286 327 320
rect 361 286 377 320
rect 311 270 377 286
rect 425 320 491 336
rect 425 286 441 320
rect 475 286 491 320
rect 425 270 491 286
rect 89 244 155 260
rect 125 222 155 244
rect 233 222 263 270
rect 327 222 357 270
rect 441 222 471 270
rect 125 86 155 112
rect 233 48 263 74
rect 327 48 357 74
rect 441 48 471 74
<< polycont >>
rect 105 260 139 294
rect 213 286 247 320
rect 327 286 361 320
rect 441 286 475 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 167 580 233 649
rect 167 546 183 580
rect 217 546 233 580
rect 21 524 119 540
rect 21 490 69 524
rect 103 490 119 524
rect 21 424 119 490
rect 167 508 233 546
rect 167 474 183 508
rect 217 474 233 508
rect 167 458 233 474
rect 455 580 559 596
rect 455 546 471 580
rect 505 546 559 580
rect 455 508 559 546
rect 455 474 471 508
rect 505 474 559 508
rect 455 458 559 474
rect 21 414 459 424
rect 21 380 69 414
rect 103 390 459 414
rect 103 380 119 390
rect 21 364 119 380
rect 21 202 55 364
rect 197 320 263 356
rect 89 294 163 310
rect 89 260 105 294
rect 139 260 163 294
rect 197 286 213 320
rect 247 286 263 320
rect 197 270 263 286
rect 311 320 377 356
rect 311 286 327 320
rect 361 286 377 320
rect 311 270 377 286
rect 425 336 459 390
rect 425 320 491 336
rect 425 286 441 320
rect 475 286 491 320
rect 425 270 491 286
rect 89 236 163 260
rect 525 236 559 458
rect 266 210 559 236
rect 21 186 130 202
rect 21 152 80 186
rect 114 152 130 186
rect 21 136 130 152
rect 166 199 232 202
rect 166 165 182 199
rect 216 165 232 199
rect 166 120 232 165
rect 166 86 182 120
rect 216 86 232 120
rect 166 17 232 86
rect 266 176 282 210
rect 316 202 482 210
rect 316 176 332 202
rect 266 120 332 176
rect 466 176 482 202
rect 516 176 559 210
rect 266 86 282 120
rect 316 86 332 120
rect 266 70 332 86
rect 366 152 432 168
rect 366 118 382 152
rect 416 118 432 152
rect 366 17 432 118
rect 466 120 559 176
rect 466 86 482 120
rect 516 86 559 120
rect 466 70 559 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
rlabel comment s 0 0 0 0 4 nor3b_1
flabel pwell s 0 0 576 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 576 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 576 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 576 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 511 94 545 128 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 511 168 545 202 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 127 242 161 276 0 FreeSans 340 0 0 0 C_N
port 3 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 B
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 576 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1962180
string GDS_START 1956974
<< end >>
