magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 1050 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 89 47 119 131
rect 184 47 214 177
rect 278 47 308 177
rect 473 47 503 131
rect 572 47 602 131
rect 669 47 699 131
rect 753 47 783 131
rect 891 47 921 131
<< pmoshvt >>
rect 81 413 117 497
rect 186 297 222 497
rect 280 297 316 497
rect 465 413 501 497
rect 565 413 601 497
rect 661 413 697 497
rect 755 413 791 497
rect 883 413 919 497
<< ndiff >>
rect 134 131 184 177
rect 27 101 89 131
rect 27 67 35 101
rect 69 67 89 101
rect 27 47 89 67
rect 119 93 184 131
rect 119 59 129 93
rect 163 59 184 93
rect 119 47 184 59
rect 214 101 278 177
rect 214 67 234 101
rect 268 67 278 101
rect 214 47 278 67
rect 308 93 367 177
rect 308 59 325 93
rect 359 59 367 93
rect 308 47 367 59
rect 421 101 473 131
rect 421 67 429 101
rect 463 67 473 101
rect 421 47 473 67
rect 503 47 572 131
rect 602 47 669 131
rect 699 47 753 131
rect 783 101 891 131
rect 783 67 837 101
rect 871 67 891 101
rect 783 47 891 67
rect 921 101 973 131
rect 921 67 931 101
rect 965 67 973 101
rect 921 47 973 67
<< pdiff >>
rect 27 477 81 497
rect 27 443 35 477
rect 69 443 81 477
rect 27 413 81 443
rect 117 485 186 497
rect 117 451 129 485
rect 163 451 186 485
rect 117 413 186 451
rect 134 297 186 413
rect 222 343 280 497
rect 222 309 234 343
rect 268 309 280 343
rect 222 297 280 309
rect 316 485 465 497
rect 316 451 344 485
rect 378 451 412 485
rect 446 451 465 485
rect 316 413 465 451
rect 501 477 565 497
rect 501 443 519 477
rect 553 443 565 477
rect 501 413 565 443
rect 601 485 661 497
rect 601 451 613 485
rect 647 451 661 485
rect 601 413 661 451
rect 697 477 755 497
rect 697 443 709 477
rect 743 443 755 477
rect 697 413 755 443
rect 791 485 883 497
rect 791 451 837 485
rect 871 451 883 485
rect 791 413 883 451
rect 919 477 973 497
rect 919 443 931 477
rect 965 443 973 477
rect 919 413 973 443
rect 316 297 444 413
<< ndiffc >>
rect 35 67 69 101
rect 129 59 163 93
rect 234 67 268 101
rect 325 59 359 93
rect 429 67 463 101
rect 837 67 871 101
rect 931 67 965 101
<< pdiffc >>
rect 35 443 69 477
rect 129 451 163 485
rect 234 309 268 343
rect 344 451 378 485
rect 412 451 446 485
rect 519 443 553 477
rect 613 451 647 485
rect 709 443 743 477
rect 837 451 871 485
rect 931 443 965 477
<< poly >>
rect 81 497 117 523
rect 186 497 222 523
rect 280 497 316 523
rect 465 497 501 523
rect 565 497 601 523
rect 661 497 697 523
rect 755 497 791 523
rect 883 497 919 523
rect 81 398 117 413
rect 79 265 119 398
rect 465 398 501 413
rect 565 398 601 413
rect 661 398 697 413
rect 755 398 791 413
rect 883 398 919 413
rect 186 282 222 297
rect 280 282 316 297
rect 21 249 119 265
rect 21 215 32 249
rect 66 215 119 249
rect 21 199 119 215
rect 89 131 119 199
rect 184 265 224 282
rect 278 265 318 282
rect 463 265 503 398
rect 563 346 603 398
rect 545 330 603 346
rect 545 296 559 330
rect 593 296 603 330
rect 545 280 603 296
rect 184 249 347 265
rect 184 215 303 249
rect 337 215 347 249
rect 184 199 347 215
rect 399 249 503 265
rect 399 215 409 249
rect 443 215 503 249
rect 399 199 503 215
rect 184 177 214 199
rect 278 177 308 199
rect 473 131 503 199
rect 572 131 602 280
rect 659 221 699 398
rect 645 205 699 221
rect 645 171 655 205
rect 689 171 699 205
rect 645 155 699 171
rect 669 131 699 155
rect 753 281 793 398
rect 753 265 807 281
rect 753 231 763 265
rect 797 231 807 265
rect 753 215 807 231
rect 881 219 921 398
rect 753 131 783 215
rect 861 203 921 219
rect 861 169 871 203
rect 905 169 921 203
rect 861 153 921 169
rect 891 131 921 153
rect 89 21 119 47
rect 184 21 214 47
rect 278 21 308 47
rect 473 21 503 47
rect 572 21 602 47
rect 669 21 699 47
rect 753 21 783 47
rect 891 21 921 47
<< polycont >>
rect 32 215 66 249
rect 559 296 593 330
rect 303 215 337 249
rect 409 215 443 249
rect 655 171 689 205
rect 763 231 797 265
rect 871 169 905 203
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 35 477 69 493
rect 103 485 179 527
rect 103 451 129 485
rect 163 451 179 485
rect 328 485 462 527
rect 328 451 344 485
rect 378 451 412 485
rect 446 451 462 485
rect 519 477 553 493
rect 35 411 69 443
rect 587 485 665 527
rect 587 451 613 485
rect 647 451 665 485
rect 709 477 743 493
rect 519 417 553 443
rect 821 485 887 527
rect 821 451 837 485
rect 871 451 887 485
rect 931 477 983 493
rect 709 417 743 443
rect 965 443 983 477
rect 931 417 983 443
rect 35 377 415 411
rect 30 249 66 327
rect 30 215 32 249
rect 30 199 66 215
rect 100 161 144 377
rect 35 127 144 161
rect 213 309 234 343
rect 268 309 284 343
rect 35 101 69 127
rect 213 101 268 309
rect 381 265 415 377
rect 477 383 743 417
rect 777 383 983 417
rect 303 249 347 265
rect 337 215 347 249
rect 303 161 347 215
rect 381 249 443 265
rect 381 215 409 249
rect 381 199 443 215
rect 477 161 521 383
rect 777 349 821 383
rect 559 330 821 349
rect 593 315 821 330
rect 593 296 603 315
rect 559 280 603 296
rect 741 265 801 281
rect 303 127 521 161
rect 654 205 707 255
rect 654 171 655 205
rect 689 171 707 205
rect 35 51 69 67
rect 103 59 129 93
rect 163 59 179 93
rect 103 17 179 59
rect 213 67 234 101
rect 429 101 463 127
rect 213 51 268 67
rect 302 59 325 93
rect 359 59 378 93
rect 302 17 378 59
rect 654 84 707 171
rect 741 231 763 265
rect 797 231 801 265
rect 741 85 801 231
rect 835 203 905 261
rect 835 169 871 203
rect 835 153 905 169
rect 949 117 983 383
rect 837 101 887 117
rect 429 51 463 67
rect 871 67 887 101
rect 837 17 887 67
rect 931 101 983 117
rect 965 67 983 101
rect 931 51 983 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
flabel corelocali s 30 289 64 323 0 FreeSans 200 0 0 0 A_N
port 1 nsew
flabel corelocali s 654 85 688 119 0 FreeSans 200 0 0 0 C
port 3 nsew
flabel corelocali s 835 153 869 187 0 FreeSans 200 0 0 0 B_N
port 2 nsew
flabel corelocali s 654 153 688 187 0 FreeSans 200 0 0 0 C
port 3 nsew
flabel corelocali s 231 238 231 238 0 FreeSans 200 0 0 0 X
port 9 nsew
flabel corelocali s 231 306 231 306 0 FreeSans 200 0 0 0 X
port 9 nsew
flabel corelocali s 654 221 688 255 0 FreeSans 200 0 0 0 C
port 3 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 200 0 0 0 A_N
port 1 nsew
flabel corelocali s 231 170 231 170 0 FreeSans 200 0 0 0 X
port 9 nsew
flabel corelocali s 757 85 791 119 0 FreeSans 200 0 0 0 D
port 4 nsew
rlabel comment s 0 0 0 0 4 and4bb_2
<< properties >>
string FIXED_BBOX 0 0 1012 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1614398
string GDS_START 1606206
<< end >>
