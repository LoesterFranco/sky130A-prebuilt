magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 86 153 166 327
rect 202 309 472 343
rect 202 164 268 309
rect 202 130 456 164
rect 234 51 268 130
rect 422 51 456 130
rect 581 199 639 265
rect 673 128 768 265
rect 1187 199 1269 324
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 17 417 69 493
rect 103 451 179 527
rect 302 451 378 527
rect 490 451 566 527
rect 736 451 802 527
rect 962 451 1164 527
rect 1219 417 1253 493
rect 17 383 988 417
rect 17 117 52 383
rect 506 309 910 343
rect 506 249 540 309
rect 954 275 988 383
rect 302 215 540 249
rect 17 51 69 117
rect 124 17 190 94
rect 302 17 378 94
rect 506 157 540 215
rect 506 123 639 157
rect 816 241 988 275
rect 1072 383 1253 417
rect 816 199 860 241
rect 1072 165 1106 383
rect 595 94 639 123
rect 942 94 1012 162
rect 1072 131 1253 165
rect 494 17 560 89
rect 595 60 1012 94
rect 1077 17 1143 93
rect 1219 51 1253 131
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
rlabel locali s 1187 199 1269 324 6 A_N
port 1 nsew signal input
rlabel locali s 86 153 166 327 6 B_N
port 2 nsew signal input
rlabel locali s 673 128 768 265 6 C
port 3 nsew signal input
rlabel locali s 581 199 639 265 6 D
port 4 nsew signal input
rlabel locali s 422 51 456 130 6 X
port 5 nsew signal output
rlabel locali s 234 51 268 130 6 X
port 5 nsew signal output
rlabel locali s 202 309 472 343 6 X
port 5 nsew signal output
rlabel locali s 202 164 268 309 6 X
port 5 nsew signal output
rlabel locali s 202 130 456 164 6 X
port 5 nsew signal output
rlabel metal1 s 0 -48 1288 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 1288 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1288 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1623500
string GDS_START 1614458
<< end >>
