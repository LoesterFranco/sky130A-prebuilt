magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 552 561
rect 19 459 253 493
rect 19 325 85 459
rect 187 451 253 459
rect 287 451 362 527
rect 472 371 525 527
rect 323 325 535 333
rect 19 299 535 325
rect 19 289 368 299
rect 25 153 115 255
rect 153 215 248 255
rect 198 135 248 215
rect 298 215 368 255
rect 298 135 340 215
rect 402 199 467 265
rect 501 165 535 299
rect 389 131 535 165
rect 19 17 109 119
rect 389 101 425 131
rect 164 51 425 101
rect 461 17 527 97
rect 0 -17 552 17
<< obsli1 >>
rect 119 417 165 425
rect 119 407 242 417
rect 391 407 425 433
rect 119 367 425 407
rect 119 359 295 367
<< metal1 >>
rect 0 496 552 592
rect 0 -48 552 48
<< labels >>
rlabel locali s 298 215 368 255 6 A1
port 1 nsew signal input
rlabel locali s 298 135 340 215 6 A1
port 1 nsew signal input
rlabel locali s 402 199 467 265 6 A2
port 2 nsew signal input
rlabel locali s 198 135 248 215 6 B1
port 3 nsew signal input
rlabel locali s 153 215 248 255 6 B1
port 3 nsew signal input
rlabel locali s 25 153 115 255 6 B2
port 4 nsew signal input
rlabel locali s 501 165 535 299 6 Y
port 5 nsew signal output
rlabel locali s 389 131 535 165 6 Y
port 5 nsew signal output
rlabel locali s 389 101 425 131 6 Y
port 5 nsew signal output
rlabel locali s 323 325 535 333 6 Y
port 5 nsew signal output
rlabel locali s 187 451 253 459 6 Y
port 5 nsew signal output
rlabel locali s 164 51 425 101 6 Y
port 5 nsew signal output
rlabel locali s 19 459 253 493 6 Y
port 5 nsew signal output
rlabel locali s 19 325 85 459 6 Y
port 5 nsew signal output
rlabel locali s 19 299 535 325 6 Y
port 5 nsew signal output
rlabel locali s 19 289 368 299 6 Y
port 5 nsew signal output
rlabel locali s 461 17 527 97 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 19 17 109 119 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 552 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 552 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 472 371 525 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 287 451 362 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 552 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 552 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 552 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 4156938
string GDS_START 4151324
<< end >>
