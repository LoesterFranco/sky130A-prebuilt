magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 17 294 75 491
rect 17 53 75 162
<< obsli1 >>
rect 0 527 29 561
rect 63 527 92 561
rect 0 -17 29 17
rect 63 -17 92 17
<< obsli1c >>
rect 29 527 63 561
rect 29 -17 63 17
<< metal1 >>
rect 0 561 92 592
rect 0 527 29 561
rect 63 527 92 561
rect 0 496 92 527
rect 0 17 92 48
rect 0 -17 29 17
rect 63 -17 92 17
rect 0 -48 92 -17
<< labels >>
rlabel locali s 17 53 75 162 6 VNB
port 1 nsew
rlabel locali s 17 294 75 491 6 VPB
port 2 nsew
rlabel metal1 s 0 -48 92 48 8 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 496 92 592 6 VPWR
port 4 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE WELLTAP
string FIXED_BBOX 0 0 92 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 952044
string GDS_START 950176
<< end >>
