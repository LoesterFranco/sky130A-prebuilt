magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 2706 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 89 47 119 131
rect 183 47 213 131
rect 381 47 411 131
rect 499 47 529 131
rect 581 47 611 131
rect 687 47 717 131
rect 763 47 793 131
rect 971 47 1001 119
rect 1087 47 1117 119
rect 1185 47 1215 131
rect 1351 47 1381 175
rect 1452 47 1482 119
rect 1585 47 1615 119
rect 1686 47 1716 131
rect 1884 47 1914 177
rect 2002 47 2032 177
rect 2096 47 2126 177
rect 2296 47 2326 131
rect 2463 47 2493 177
rect 2557 47 2587 177
<< pmoshvt >>
rect 81 363 117 491
rect 175 363 211 491
rect 373 369 409 497
rect 467 369 503 497
rect 568 369 604 497
rect 662 369 698 497
rect 765 369 801 497
rect 972 413 1008 497
rect 1075 413 1111 497
rect 1181 413 1217 497
rect 1323 347 1359 497
rect 1428 413 1464 497
rect 1522 413 1558 497
rect 1655 413 1691 497
rect 1876 297 1912 497
rect 1994 297 2030 497
rect 2088 297 2124 497
rect 2288 369 2324 497
rect 2455 297 2491 497
rect 2549 297 2585 497
<< ndiff >>
rect 27 119 89 131
rect 27 85 35 119
rect 69 85 89 119
rect 27 47 89 85
rect 119 93 183 131
rect 119 59 129 93
rect 163 59 183 93
rect 119 47 183 59
rect 213 119 265 131
rect 213 85 223 119
rect 257 85 265 119
rect 213 47 265 85
rect 319 89 381 131
rect 319 55 331 89
rect 365 55 381 89
rect 319 47 381 55
rect 411 89 499 131
rect 411 55 445 89
rect 479 55 499 89
rect 411 47 499 55
rect 529 47 581 131
rect 611 89 687 131
rect 611 55 632 89
rect 666 55 687 89
rect 611 47 687 55
rect 717 47 763 131
rect 793 93 861 131
rect 1291 131 1351 175
rect 1135 119 1185 131
rect 793 59 819 93
rect 853 59 861 93
rect 793 47 861 59
rect 915 107 971 119
rect 915 73 923 107
rect 957 73 971 107
rect 915 47 971 73
rect 1001 107 1087 119
rect 1001 73 1033 107
rect 1067 73 1087 107
rect 1001 47 1087 73
rect 1117 47 1185 119
rect 1215 101 1351 131
rect 1215 67 1269 101
rect 1303 67 1351 101
rect 1215 47 1351 67
rect 1381 119 1431 175
rect 1822 162 1884 177
rect 1630 119 1686 131
rect 1381 107 1452 119
rect 1381 73 1397 107
rect 1431 73 1452 107
rect 1381 47 1452 73
rect 1482 107 1585 119
rect 1482 73 1519 107
rect 1553 73 1585 107
rect 1482 47 1585 73
rect 1615 47 1686 119
rect 1716 107 1768 131
rect 1716 73 1726 107
rect 1760 73 1768 107
rect 1716 47 1768 73
rect 1822 128 1830 162
rect 1864 128 1884 162
rect 1822 94 1884 128
rect 1822 60 1830 94
rect 1864 60 1884 94
rect 1822 47 1884 60
rect 1914 123 2002 177
rect 1914 89 1936 123
rect 1970 89 2002 123
rect 1914 47 2002 89
rect 2032 169 2096 177
rect 2032 135 2042 169
rect 2076 135 2096 169
rect 2032 101 2096 135
rect 2032 67 2042 101
rect 2076 67 2096 101
rect 2032 47 2096 67
rect 2126 122 2180 177
rect 2341 161 2463 177
rect 2341 131 2380 161
rect 2126 88 2138 122
rect 2172 88 2180 122
rect 2126 47 2180 88
rect 2234 119 2296 131
rect 2234 85 2242 119
rect 2276 85 2296 119
rect 2234 47 2296 85
rect 2326 127 2380 131
rect 2414 127 2463 161
rect 2326 93 2463 127
rect 2326 59 2380 93
rect 2414 59 2463 93
rect 2326 47 2463 59
rect 2493 143 2557 177
rect 2493 109 2503 143
rect 2537 109 2557 143
rect 2493 47 2557 109
rect 2587 161 2639 177
rect 2587 127 2597 161
rect 2631 127 2639 161
rect 2587 93 2639 127
rect 2587 59 2597 93
rect 2631 59 2639 93
rect 2587 47 2639 59
<< pdiff >>
rect 27 477 81 491
rect 27 443 35 477
rect 69 443 81 477
rect 27 409 81 443
rect 27 375 35 409
rect 69 375 81 409
rect 27 363 81 375
rect 117 461 175 491
rect 117 427 129 461
rect 163 427 175 461
rect 117 363 175 427
rect 211 477 265 491
rect 211 443 223 477
rect 257 443 265 477
rect 211 409 265 443
rect 211 375 223 409
rect 257 375 265 409
rect 211 363 265 375
rect 319 452 373 497
rect 319 418 327 452
rect 361 418 373 452
rect 319 369 373 418
rect 409 483 467 497
rect 409 449 421 483
rect 455 449 467 483
rect 409 369 467 449
rect 503 369 568 497
rect 604 483 662 497
rect 604 449 616 483
rect 650 449 662 483
rect 604 369 662 449
rect 698 369 765 497
rect 801 483 860 497
rect 801 449 818 483
rect 852 449 860 483
rect 801 369 860 449
rect 918 472 972 497
rect 918 438 926 472
rect 960 438 972 472
rect 918 413 972 438
rect 1008 472 1075 497
rect 1008 438 1025 472
rect 1059 438 1075 472
rect 1008 413 1075 438
rect 1111 413 1181 497
rect 1217 485 1323 497
rect 1217 451 1277 485
rect 1311 451 1323 485
rect 1217 417 1323 451
rect 1217 413 1277 417
rect 1234 383 1277 413
rect 1311 383 1323 417
rect 1234 347 1323 383
rect 1359 477 1428 497
rect 1359 443 1371 477
rect 1405 443 1428 477
rect 1359 413 1428 443
rect 1464 467 1522 497
rect 1464 433 1476 467
rect 1510 433 1522 467
rect 1464 413 1522 433
rect 1558 413 1655 497
rect 1691 477 1768 497
rect 1691 443 1725 477
rect 1759 443 1768 477
rect 1691 413 1768 443
rect 1822 485 1876 497
rect 1822 451 1830 485
rect 1864 451 1876 485
rect 1822 417 1876 451
rect 1359 347 1411 413
rect 1822 383 1830 417
rect 1864 383 1876 417
rect 1822 349 1876 383
rect 1822 315 1830 349
rect 1864 315 1876 349
rect 1822 297 1876 315
rect 1912 455 1994 497
rect 1912 421 1936 455
rect 1970 421 1994 455
rect 1912 375 1994 421
rect 1912 341 1936 375
rect 1970 341 1994 375
rect 1912 297 1994 341
rect 2030 475 2088 497
rect 2030 441 2042 475
rect 2076 441 2088 475
rect 2030 407 2088 441
rect 2030 373 2042 407
rect 2076 373 2088 407
rect 2030 339 2088 373
rect 2030 305 2042 339
rect 2076 305 2088 339
rect 2030 297 2088 305
rect 2124 485 2180 497
rect 2124 451 2138 485
rect 2172 451 2180 485
rect 2124 373 2180 451
rect 2124 339 2138 373
rect 2172 339 2180 373
rect 2234 485 2288 497
rect 2234 451 2242 485
rect 2276 451 2288 485
rect 2234 417 2288 451
rect 2234 383 2242 417
rect 2276 383 2288 417
rect 2234 369 2288 383
rect 2324 485 2455 497
rect 2324 451 2380 485
rect 2414 451 2455 485
rect 2324 417 2455 451
rect 2324 383 2380 417
rect 2414 383 2455 417
rect 2324 369 2455 383
rect 2124 297 2180 339
rect 2341 349 2455 369
rect 2341 315 2380 349
rect 2414 315 2455 349
rect 2341 297 2455 315
rect 2491 449 2549 497
rect 2491 415 2503 449
rect 2537 415 2549 449
rect 2491 381 2549 415
rect 2491 347 2503 381
rect 2537 347 2549 381
rect 2491 297 2549 347
rect 2585 485 2639 497
rect 2585 451 2597 485
rect 2631 451 2639 485
rect 2585 417 2639 451
rect 2585 383 2597 417
rect 2631 383 2639 417
rect 2585 349 2639 383
rect 2585 315 2597 349
rect 2631 315 2639 349
rect 2585 297 2639 315
<< ndiffc >>
rect 35 85 69 119
rect 129 59 163 93
rect 223 85 257 119
rect 331 55 365 89
rect 445 55 479 89
rect 632 55 666 89
rect 819 59 853 93
rect 923 73 957 107
rect 1033 73 1067 107
rect 1269 67 1303 101
rect 1397 73 1431 107
rect 1519 73 1553 107
rect 1726 73 1760 107
rect 1830 128 1864 162
rect 1830 60 1864 94
rect 1936 89 1970 123
rect 2042 135 2076 169
rect 2042 67 2076 101
rect 2138 88 2172 122
rect 2242 85 2276 119
rect 2380 127 2414 161
rect 2380 59 2414 93
rect 2503 109 2537 143
rect 2597 127 2631 161
rect 2597 59 2631 93
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 129 427 163 461
rect 223 443 257 477
rect 223 375 257 409
rect 327 418 361 452
rect 421 449 455 483
rect 616 449 650 483
rect 818 449 852 483
rect 926 438 960 472
rect 1025 438 1059 472
rect 1277 451 1311 485
rect 1277 383 1311 417
rect 1371 443 1405 477
rect 1476 433 1510 467
rect 1725 443 1759 477
rect 1830 451 1864 485
rect 1830 383 1864 417
rect 1830 315 1864 349
rect 1936 421 1970 455
rect 1936 341 1970 375
rect 2042 441 2076 475
rect 2042 373 2076 407
rect 2042 305 2076 339
rect 2138 451 2172 485
rect 2138 339 2172 373
rect 2242 451 2276 485
rect 2242 383 2276 417
rect 2380 451 2414 485
rect 2380 383 2414 417
rect 2380 315 2414 349
rect 2503 415 2537 449
rect 2503 347 2537 381
rect 2597 451 2631 485
rect 2597 383 2631 417
rect 2597 315 2631 349
<< poly >>
rect 81 491 117 517
rect 175 491 211 517
rect 373 497 409 523
rect 467 497 503 523
rect 568 497 604 523
rect 662 497 698 523
rect 765 497 801 523
rect 972 497 1008 523
rect 1075 497 1111 523
rect 1181 497 1217 523
rect 1323 497 1359 523
rect 1428 497 1464 523
rect 1522 497 1558 523
rect 1655 497 1691 523
rect 1876 497 1912 523
rect 1994 497 2030 523
rect 2088 497 2124 523
rect 2288 497 2324 523
rect 2455 497 2491 523
rect 2549 497 2585 523
rect 972 398 1008 413
rect 1075 398 1111 413
rect 1181 398 1217 413
rect 970 375 1010 398
rect 1073 381 1113 398
rect 81 348 117 363
rect 175 348 211 363
rect 373 354 409 369
rect 467 354 503 369
rect 568 354 604 369
rect 662 354 698 369
rect 765 354 801 369
rect 955 365 1031 375
rect 47 318 119 348
rect 47 265 77 318
rect 173 274 213 348
rect 371 331 411 354
rect 465 331 505 354
rect 566 337 606 354
rect 660 337 700 354
rect 356 321 505 331
rect 356 287 372 321
rect 406 301 505 321
rect 551 321 615 337
rect 406 287 432 301
rect 356 277 432 287
rect 551 287 561 321
rect 595 287 615 321
rect 23 249 77 265
rect 23 215 33 249
rect 67 215 77 249
rect 129 264 213 274
rect 129 230 145 264
rect 179 230 213 264
rect 129 220 213 230
rect 23 199 77 215
rect 47 176 77 199
rect 47 146 119 176
rect 89 131 119 146
rect 183 131 213 220
rect 381 131 411 277
rect 551 271 615 287
rect 657 321 721 337
rect 657 287 667 321
rect 701 287 721 321
rect 657 271 721 287
rect 763 304 803 354
rect 955 331 971 365
rect 1005 331 1031 365
rect 955 321 1031 331
rect 1073 365 1137 381
rect 1073 331 1083 365
rect 1117 331 1137 365
rect 1073 315 1137 331
rect 763 288 827 304
rect 463 225 529 235
rect 463 191 479 225
rect 513 191 529 225
rect 463 181 529 191
rect 499 131 529 181
rect 581 131 611 271
rect 763 254 773 288
rect 807 254 827 288
rect 1073 279 1113 315
rect 763 238 827 254
rect 971 249 1113 279
rect 653 207 717 223
rect 653 173 663 207
rect 697 173 717 207
rect 653 157 717 173
rect 687 131 717 157
rect 763 131 793 238
rect 971 119 1001 249
rect 1179 213 1219 398
rect 1428 398 1464 413
rect 1522 398 1558 413
rect 1655 398 1691 413
rect 1323 332 1359 347
rect 1321 309 1361 332
rect 1426 315 1466 398
rect 1520 375 1560 398
rect 1653 381 1693 398
rect 1519 365 1595 375
rect 1519 331 1535 365
rect 1569 331 1595 365
rect 1519 321 1595 331
rect 1653 365 1741 381
rect 1653 331 1697 365
rect 1731 331 1741 365
rect 1653 315 1741 331
rect 1261 299 1361 309
rect 1261 265 1277 299
rect 1311 265 1361 299
rect 1261 255 1361 265
rect 1321 220 1361 255
rect 1413 299 1477 315
rect 1413 265 1423 299
rect 1457 279 1477 299
rect 1457 265 1615 279
rect 1413 249 1615 265
rect 1053 191 1117 207
rect 1053 157 1063 191
rect 1097 157 1117 191
rect 1179 203 1269 213
rect 1179 183 1219 203
rect 1053 141 1117 157
rect 1087 119 1117 141
rect 1185 169 1219 183
rect 1253 169 1269 203
rect 1321 190 1381 220
rect 1351 175 1381 190
rect 1452 191 1523 207
rect 1185 159 1269 169
rect 1185 131 1215 159
rect 1452 157 1479 191
rect 1513 157 1523 191
rect 1452 141 1523 157
rect 1452 119 1482 141
rect 1585 119 1615 249
rect 1686 131 1716 315
rect 2288 354 2324 369
rect 1876 282 1912 297
rect 1994 282 2030 297
rect 2088 282 2124 297
rect 1874 265 1914 282
rect 1992 265 2032 282
rect 2086 265 2126 282
rect 2286 265 2326 354
rect 2455 282 2491 297
rect 2549 282 2585 297
rect 2453 265 2493 282
rect 2547 265 2587 282
rect 1765 249 1914 265
rect 1765 215 1775 249
rect 1809 215 1914 249
rect 1765 199 1914 215
rect 1956 249 2326 265
rect 1956 215 1966 249
rect 2000 215 2326 249
rect 1956 199 2326 215
rect 2424 249 2587 265
rect 2424 215 2434 249
rect 2468 215 2587 249
rect 2424 199 2587 215
rect 1884 177 1914 199
rect 2002 177 2032 199
rect 2096 177 2126 199
rect 2296 131 2326 199
rect 2463 177 2493 199
rect 2557 177 2587 199
rect 89 21 119 47
rect 183 21 213 47
rect 381 21 411 47
rect 499 21 529 47
rect 581 21 611 47
rect 687 21 717 47
rect 763 21 793 47
rect 971 21 1001 47
rect 1087 21 1117 47
rect 1185 21 1215 47
rect 1351 21 1381 47
rect 1452 21 1482 47
rect 1585 21 1615 47
rect 1686 21 1716 47
rect 1884 21 1914 47
rect 2002 21 2032 47
rect 2096 21 2126 47
rect 2296 21 2326 47
rect 2463 21 2493 47
rect 2557 21 2587 47
<< polycont >>
rect 372 287 406 321
rect 561 287 595 321
rect 33 215 67 249
rect 145 230 179 264
rect 667 287 701 321
rect 971 331 1005 365
rect 1083 331 1117 365
rect 479 191 513 225
rect 773 254 807 288
rect 663 173 697 207
rect 1535 331 1569 365
rect 1697 331 1731 365
rect 1277 265 1311 299
rect 1423 265 1457 299
rect 1063 157 1097 191
rect 1219 169 1253 203
rect 1479 157 1513 191
rect 1775 215 1809 249
rect 1966 215 2000 249
rect 2434 215 2468 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2668 561
rect 35 477 69 493
rect 35 409 69 443
rect 103 461 179 527
rect 103 427 129 461
rect 163 427 179 461
rect 223 477 257 493
rect 223 409 257 443
rect 69 391 179 393
rect 69 375 139 391
rect 35 359 139 375
rect 133 357 139 359
rect 173 357 179 391
rect 19 249 89 325
rect 19 215 33 249
rect 67 215 89 249
rect 19 195 89 215
rect 133 264 179 357
rect 133 230 145 264
rect 133 194 179 230
rect 133 161 172 194
rect 35 127 172 161
rect 35 119 69 127
rect 223 119 257 375
rect 35 69 69 85
rect 103 59 129 93
rect 163 59 179 93
rect 223 69 257 85
rect 304 452 361 489
rect 304 418 327 452
rect 395 483 471 527
rect 818 483 852 527
rect 395 449 421 483
rect 455 449 471 483
rect 575 449 616 483
rect 650 449 774 483
rect 304 415 361 418
rect 304 372 706 415
rect 304 89 338 372
rect 372 321 406 337
rect 372 157 406 287
rect 450 225 484 372
rect 667 337 706 372
rect 740 399 774 449
rect 818 433 852 449
rect 903 472 960 488
rect 1277 485 1311 527
rect 903 438 926 472
rect 999 438 1025 472
rect 1059 438 1243 472
rect 903 414 960 438
rect 903 399 937 414
rect 740 365 937 399
rect 1067 391 1165 402
rect 551 321 625 337
rect 551 287 561 321
rect 595 287 625 321
rect 551 271 625 287
rect 667 321 711 337
rect 701 287 711 321
rect 667 271 711 287
rect 763 288 869 331
rect 763 254 773 288
rect 807 254 869 288
rect 450 191 479 225
rect 513 191 539 225
rect 663 207 707 223
rect 763 211 869 254
rect 697 173 707 207
rect 903 177 937 365
rect 663 157 707 173
rect 372 123 707 157
rect 741 143 937 177
rect 741 89 775 143
rect 103 17 179 59
rect 304 55 331 89
rect 365 55 381 89
rect 304 51 381 55
rect 429 55 445 89
rect 479 55 495 89
rect 610 55 632 89
rect 666 55 775 89
rect 819 93 859 109
rect 853 59 859 93
rect 903 107 937 143
rect 971 365 1029 381
rect 1005 331 1029 365
rect 1067 365 1123 391
rect 1067 331 1083 365
rect 1117 357 1123 365
rect 1157 357 1165 391
rect 1117 331 1165 357
rect 971 207 1029 331
rect 1199 315 1243 438
rect 1277 417 1311 451
rect 1277 367 1311 383
rect 1345 477 1405 493
rect 1345 443 1371 477
rect 1703 477 1764 527
rect 1345 427 1405 443
rect 1450 433 1476 467
rect 1510 433 1657 467
rect 1199 299 1311 315
rect 1199 297 1277 299
rect 1141 265 1277 297
rect 1141 263 1311 265
rect 971 191 1097 207
rect 971 187 1063 191
rect 971 153 1029 187
rect 1063 153 1097 157
rect 971 141 1097 153
rect 1141 107 1175 263
rect 1277 249 1311 263
rect 1219 213 1253 219
rect 1345 213 1389 427
rect 1423 391 1471 393
rect 1423 357 1435 391
rect 1469 357 1471 391
rect 1423 299 1471 357
rect 1457 265 1471 299
rect 1423 249 1471 265
rect 1505 365 1579 381
rect 1505 331 1535 365
rect 1569 331 1579 365
rect 1505 315 1579 331
rect 1219 203 1389 213
rect 1505 207 1543 315
rect 1623 281 1657 433
rect 1703 443 1725 477
rect 1759 443 1764 477
rect 1703 427 1764 443
rect 1814 485 1880 491
rect 1814 451 1830 485
rect 1864 451 1880 485
rect 1814 417 1880 451
rect 1814 383 1830 417
rect 1864 383 1880 417
rect 1814 381 1880 383
rect 1697 365 1880 381
rect 1731 349 1880 365
rect 1731 331 1830 349
rect 1697 315 1830 331
rect 1864 315 1880 349
rect 1914 455 1998 527
rect 1914 421 1936 455
rect 1970 421 1998 455
rect 1914 375 1998 421
rect 1914 341 1936 375
rect 1970 341 1998 375
rect 1914 325 1998 341
rect 2042 475 2098 491
rect 2076 441 2098 475
rect 2042 407 2098 441
rect 2076 373 2098 407
rect 2042 339 2098 373
rect 1253 169 1389 203
rect 1219 153 1389 169
rect 903 73 923 107
rect 957 73 973 107
rect 1017 73 1033 107
rect 1067 73 1175 107
rect 1235 101 1309 117
rect 429 17 495 55
rect 819 17 859 59
rect 1235 67 1269 101
rect 1303 67 1309 101
rect 1345 107 1389 153
rect 1423 191 1543 207
rect 1423 187 1479 191
rect 1423 153 1437 187
rect 1471 157 1479 187
rect 1513 157 1543 191
rect 1471 153 1543 157
rect 1423 141 1543 153
rect 1587 265 1657 281
rect 1843 265 1880 315
rect 2076 305 2098 339
rect 2138 485 2172 527
rect 2338 485 2459 527
rect 2138 373 2172 451
rect 2138 323 2172 339
rect 2226 451 2242 485
rect 2276 451 2292 485
rect 2226 417 2292 451
rect 2226 383 2242 417
rect 2276 383 2292 417
rect 1587 249 1809 265
rect 1587 215 1775 249
rect 1587 199 1809 215
rect 1843 249 2000 265
rect 1843 215 1966 249
rect 1843 199 2000 215
rect 1587 107 1631 199
rect 1843 165 1880 199
rect 1807 162 1880 165
rect 1807 128 1830 162
rect 1864 128 1880 162
rect 2042 169 2098 305
rect 1345 73 1397 107
rect 1431 73 1447 107
rect 1503 73 1519 107
rect 1553 73 1631 107
rect 1676 107 1760 123
rect 1676 73 1726 107
rect 1235 17 1309 67
rect 1676 17 1760 73
rect 1807 94 1880 128
rect 1807 60 1830 94
rect 1864 60 1880 94
rect 1914 123 1998 139
rect 1914 89 1936 123
rect 1970 89 1998 123
rect 1914 17 1998 89
rect 2076 135 2098 169
rect 2226 265 2292 383
rect 2338 451 2380 485
rect 2414 451 2459 485
rect 2597 485 2631 527
rect 2338 417 2459 451
rect 2338 383 2380 417
rect 2414 383 2459 417
rect 2338 349 2459 383
rect 2338 315 2380 349
rect 2414 315 2459 349
rect 2338 299 2459 315
rect 2503 449 2557 465
rect 2537 415 2557 449
rect 2503 381 2557 415
rect 2537 347 2557 381
rect 2226 249 2468 265
rect 2226 215 2434 249
rect 2226 199 2468 215
rect 2042 101 2098 135
rect 2076 67 2098 101
rect 2042 51 2098 67
rect 2136 122 2182 138
rect 2136 88 2138 122
rect 2172 88 2182 122
rect 2136 17 2182 88
rect 2226 119 2276 199
rect 2226 85 2242 119
rect 2226 69 2276 85
rect 2333 127 2380 161
rect 2414 127 2459 161
rect 2333 93 2459 127
rect 2333 59 2380 93
rect 2414 59 2459 93
rect 2333 17 2459 59
rect 2503 143 2557 347
rect 2597 417 2631 451
rect 2597 349 2631 383
rect 2597 279 2631 315
rect 2537 109 2557 143
rect 2503 53 2557 109
rect 2597 161 2631 191
rect 2597 93 2631 127
rect 2597 17 2631 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2668 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 139 357 173 391
rect 223 85 257 119
rect 1123 357 1157 391
rect 1029 153 1063 187
rect 1435 357 1469 391
rect 1437 153 1471 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
<< metal1 >>
rect 0 561 2668 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2668 561
rect 0 496 2668 527
rect 127 391 185 397
rect 127 357 139 391
rect 173 388 185 391
rect 1111 391 1169 397
rect 1111 388 1123 391
rect 173 360 1123 388
rect 173 357 185 360
rect 127 351 185 357
rect 1111 357 1123 360
rect 1157 388 1169 391
rect 1423 391 1481 397
rect 1423 388 1435 391
rect 1157 360 1435 388
rect 1157 357 1169 360
rect 1111 351 1169 357
rect 1423 357 1435 360
rect 1469 357 1481 391
rect 1423 351 1481 357
rect 1017 187 1075 193
rect 1017 153 1029 187
rect 1063 184 1075 187
rect 1425 187 1483 193
rect 1425 184 1437 187
rect 1063 156 1437 184
rect 1063 153 1075 156
rect 1017 147 1075 153
rect 1425 153 1437 156
rect 1471 153 1483 187
rect 1425 147 1483 153
rect 201 119 269 125
rect 201 85 223 119
rect 257 116 269 119
rect 1017 116 1045 147
rect 257 88 1045 116
rect 257 85 269 88
rect 201 79 269 85
rect 0 17 2668 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2668 17
rect 0 -48 2668 -17
<< labels >>
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel corelocali s 2513 289 2547 323 0 FreeSans 400 0 0 0 Q_N
port 10 nsew
flabel corelocali s 2053 85 2087 119 0 FreeSans 200 0 0 0 Q
port 9 nsew
flabel corelocali s 29 221 63 255 0 FreeSans 400 0 0 0 CLK
port 1 nsew
flabel corelocali s 673 153 707 187 0 FreeSans 300 0 0 0 SCE
port 4 nsew
flabel corelocali s 581 289 615 323 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel corelocali s 765 221 799 255 0 FreeSans 300 0 0 0 SCD
port 3 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel nbase s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
port 7 nsew
rlabel comment s 0 0 0 0 4 sdfxbp_2
<< properties >>
string FIXED_BBOX 0 0 2668 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 321516
string GDS_START 302866
<< end >>
