magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 2481 325 2531 425
rect 2669 325 2719 425
rect 2857 325 2907 425
rect 3045 325 3095 425
rect 2481 291 3095 325
rect 81 215 759 257
rect 849 215 1527 257
rect 1689 215 2367 257
rect 2481 181 2563 291
rect 2597 215 3071 257
rect 113 145 3103 181
rect 113 51 179 145
rect 301 51 367 145
rect 489 51 555 145
rect 677 51 743 145
rect 865 51 931 145
rect 1053 51 1119 145
rect 1241 51 1307 145
rect 1429 51 1495 145
rect 1721 51 1787 145
rect 1909 51 1975 145
rect 2097 51 2163 145
rect 2285 51 2351 145
rect 2473 51 2539 145
rect 2661 51 2727 145
rect 2849 51 2915 145
rect 3037 51 3103 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3157 561
rect 3191 527 3220 561
rect 19 325 85 493
rect 121 359 171 527
rect 215 325 265 493
rect 309 359 359 527
rect 403 325 453 493
rect 497 359 547 527
rect 591 325 641 493
rect 685 359 735 527
rect 779 459 1589 493
rect 779 325 829 459
rect 19 291 829 325
rect 873 325 923 425
rect 967 359 1017 459
rect 1061 325 1111 425
rect 1155 359 1205 459
rect 1249 325 1299 425
rect 1343 359 1393 459
rect 1437 325 1487 425
rect 1531 359 1589 459
rect 1627 459 3199 493
rect 1627 359 1685 459
rect 1729 325 1779 425
rect 1815 359 1873 459
rect 1917 325 1967 425
rect 2011 359 2061 459
rect 2105 325 2155 425
rect 2199 359 2249 459
rect 2293 325 2343 425
rect 873 291 2343 325
rect 2387 291 2437 459
rect 2575 359 2625 459
rect 2763 359 2813 459
rect 2951 359 3001 459
rect 3139 293 3199 459
rect 27 17 79 181
rect 213 17 267 111
rect 401 17 455 111
rect 589 17 643 111
rect 777 17 831 111
rect 965 17 1019 111
rect 1153 17 1207 111
rect 1341 17 1395 111
rect 1529 17 1687 111
rect 1821 17 1875 111
rect 2009 17 2063 111
rect 2197 17 2251 111
rect 2385 17 2439 111
rect 2573 17 2627 111
rect 2761 17 2815 111
rect 2949 17 3003 111
rect 3137 17 3193 181
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3220 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 2881 527 2915 561
rect 2973 527 3007 561
rect 3065 527 3099 561
rect 3157 527 3191 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
rect 2881 -17 2915 17
rect 2973 -17 3007 17
rect 3065 -17 3099 17
rect 3157 -17 3191 17
<< metal1 >>
rect 0 561 3220 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3157 561
rect 3191 527 3220 561
rect 0 496 3220 527
rect 0 17 3220 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3220 17
rect 0 -48 3220 -17
<< labels >>
rlabel locali s 81 215 759 257 6 A
port 1 nsew signal input
rlabel locali s 849 215 1527 257 6 B
port 2 nsew signal input
rlabel locali s 1689 215 2367 257 6 C
port 3 nsew signal input
rlabel locali s 2597 215 3071 257 6 D
port 4 nsew signal input
rlabel locali s 3045 325 3095 425 6 Y
port 5 nsew signal output
rlabel locali s 3037 51 3103 145 6 Y
port 5 nsew signal output
rlabel locali s 2857 325 2907 425 6 Y
port 5 nsew signal output
rlabel locali s 2849 51 2915 145 6 Y
port 5 nsew signal output
rlabel locali s 2669 325 2719 425 6 Y
port 5 nsew signal output
rlabel locali s 2661 51 2727 145 6 Y
port 5 nsew signal output
rlabel locali s 2481 325 2531 425 6 Y
port 5 nsew signal output
rlabel locali s 2481 291 3095 325 6 Y
port 5 nsew signal output
rlabel locali s 2481 181 2563 291 6 Y
port 5 nsew signal output
rlabel locali s 2473 51 2539 145 6 Y
port 5 nsew signal output
rlabel locali s 2285 51 2351 145 6 Y
port 5 nsew signal output
rlabel locali s 2097 51 2163 145 6 Y
port 5 nsew signal output
rlabel locali s 1909 51 1975 145 6 Y
port 5 nsew signal output
rlabel locali s 1721 51 1787 145 6 Y
port 5 nsew signal output
rlabel locali s 1429 51 1495 145 6 Y
port 5 nsew signal output
rlabel locali s 1241 51 1307 145 6 Y
port 5 nsew signal output
rlabel locali s 1053 51 1119 145 6 Y
port 5 nsew signal output
rlabel locali s 865 51 931 145 6 Y
port 5 nsew signal output
rlabel locali s 677 51 743 145 6 Y
port 5 nsew signal output
rlabel locali s 489 51 555 145 6 Y
port 5 nsew signal output
rlabel locali s 301 51 367 145 6 Y
port 5 nsew signal output
rlabel locali s 113 145 3103 181 6 Y
port 5 nsew signal output
rlabel locali s 113 51 179 145 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -48 3220 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 3220 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 3220 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3520610
string GDS_START 3497104
<< end >>
