magic
tech sky130A
magscale 1 2
timestamp 1599588232
<< locali >>
rect 123 394 189 547
rect 323 394 389 547
rect 123 378 389 394
rect 123 360 647 378
rect 25 326 71 356
rect 323 344 647 360
rect 25 260 218 326
rect 301 236 455 310
rect 489 236 555 310
rect 601 247 647 344
rect 697 270 875 356
rect 601 202 641 247
rect 1157 236 1223 310
rect 291 168 641 202
rect 291 119 357 168
rect 603 119 641 168
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 23 581 480 615
rect 23 390 89 581
rect 223 428 289 581
rect 423 446 480 581
rect 514 480 656 649
rect 690 446 747 596
rect 781 458 850 649
rect 423 424 747 446
rect 884 424 975 596
rect 423 412 975 424
rect 1009 412 1075 649
rect 681 390 975 412
rect 909 378 975 390
rect 1109 378 1175 596
rect 909 344 1175 378
rect 23 192 255 226
rect 23 70 73 192
rect 109 17 175 158
rect 221 85 255 192
rect 391 85 457 134
rect 221 51 457 85
rect 503 85 569 134
rect 675 85 741 226
rect 775 202 1123 236
rect 775 119 841 202
rect 875 85 941 168
rect 503 51 941 85
rect 987 17 1037 168
rect 1073 70 1123 202
rect 1159 17 1225 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
<< metal1 >>
rect 0 683 1248 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 0 617 1248 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 1248 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
rect 0 -49 1248 -17
<< labels >>
rlabel locali s 489 236 555 310 6 A1
port 1 nsew signal input
rlabel locali s 697 270 875 356 6 A2
port 2 nsew signal input
rlabel locali s 1157 236 1223 310 6 A3
port 3 nsew signal input
rlabel locali s 301 236 455 310 6 B1
port 4 nsew signal input
rlabel locali s 25 326 71 356 6 B2
port 5 nsew signal input
rlabel locali s 25 260 218 326 6 B2
port 5 nsew signal input
rlabel locali s 603 119 641 168 6 Y
port 6 nsew signal output
rlabel locali s 601 247 647 344 6 Y
port 6 nsew signal output
rlabel locali s 601 202 641 247 6 Y
port 6 nsew signal output
rlabel locali s 323 394 389 547 6 Y
port 6 nsew signal output
rlabel locali s 323 344 647 360 6 Y
port 6 nsew signal output
rlabel locali s 291 168 641 202 6 Y
port 6 nsew signal output
rlabel locali s 291 119 357 168 6 Y
port 6 nsew signal output
rlabel locali s 123 394 189 547 6 Y
port 6 nsew signal output
rlabel locali s 123 378 389 394 6 Y
port 6 nsew signal output
rlabel locali s 123 360 647 378 6 Y
port 6 nsew signal output
rlabel metal1 s 0 -49 1248 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 8 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 9 nsew power bidirectional
rlabel metal1 s 0 617 1248 715 6 VPWR
port 10 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1248 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3875768
string GDS_START 3865274
<< end >>
