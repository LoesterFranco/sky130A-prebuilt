magic
tech sky130A
magscale 1 2
timestamp 1599588209
<< nwell >>
rect -38 332 2054 704
<< pwell >>
rect 0 0 2016 49
<< scpmos >>
rect 86 424 116 592
rect 176 424 206 592
rect 266 424 296 592
rect 356 424 386 592
rect 500 368 530 592
rect 600 368 630 592
rect 690 368 720 592
rect 780 368 810 592
rect 870 368 900 592
rect 960 368 990 592
rect 1060 368 1090 592
rect 1150 368 1180 592
rect 1240 368 1270 592
rect 1330 368 1360 592
rect 1440 368 1470 592
rect 1530 368 1560 592
rect 1630 368 1660 592
rect 1720 368 1750 592
rect 1810 368 1840 592
rect 1900 368 1930 592
<< nmoslvt >>
rect 84 114 114 262
rect 202 114 232 262
rect 431 74 461 222
rect 538 74 568 222
rect 626 74 656 222
rect 712 74 742 222
rect 798 74 828 222
rect 884 74 914 222
rect 970 74 1000 222
rect 1088 74 1118 222
rect 1286 74 1316 222
rect 1372 74 1402 222
rect 1458 74 1488 222
rect 1544 74 1574 222
rect 1630 74 1660 222
rect 1716 74 1746 222
rect 1802 74 1832 222
rect 1902 74 1932 222
<< ndiff >>
rect 27 240 84 262
rect 27 206 39 240
rect 73 206 84 240
rect 27 160 84 206
rect 27 126 39 160
rect 73 126 84 160
rect 27 114 84 126
rect 114 114 202 262
rect 232 250 296 262
rect 232 216 246 250
rect 280 216 296 250
rect 232 114 296 216
rect 374 192 431 222
rect 374 158 386 192
rect 420 158 431 192
rect 374 120 431 158
rect 129 82 187 114
rect 129 48 141 82
rect 175 48 187 82
rect 374 86 386 120
rect 420 86 431 120
rect 374 74 431 86
rect 461 180 538 222
rect 461 146 480 180
rect 514 146 538 180
rect 461 74 538 146
rect 568 122 626 222
rect 568 88 580 122
rect 614 88 626 122
rect 568 74 626 88
rect 656 189 712 222
rect 656 155 667 189
rect 701 155 712 189
rect 656 74 712 155
rect 742 144 798 222
rect 742 110 753 144
rect 787 110 798 144
rect 742 74 798 110
rect 828 116 884 222
rect 828 82 839 116
rect 873 82 884 116
rect 828 74 884 82
rect 914 184 970 222
rect 914 150 925 184
rect 959 150 970 184
rect 914 74 970 150
rect 1000 116 1088 222
rect 1000 82 1027 116
rect 1061 82 1088 116
rect 1000 74 1088 82
rect 1118 160 1175 222
rect 1118 126 1129 160
rect 1163 126 1175 160
rect 1118 74 1175 126
rect 1229 189 1286 222
rect 1229 155 1241 189
rect 1275 155 1286 189
rect 1229 74 1286 155
rect 1316 133 1372 222
rect 1316 99 1327 133
rect 1361 99 1372 133
rect 1316 74 1372 99
rect 1402 189 1458 222
rect 1402 155 1413 189
rect 1447 155 1458 189
rect 1402 74 1458 155
rect 1488 133 1544 222
rect 1488 99 1499 133
rect 1533 99 1544 133
rect 1488 74 1544 99
rect 1574 210 1630 222
rect 1574 176 1585 210
rect 1619 176 1630 210
rect 1574 120 1630 176
rect 1574 86 1585 120
rect 1619 86 1630 120
rect 1574 74 1630 86
rect 1660 131 1716 222
rect 1660 97 1671 131
rect 1705 97 1716 131
rect 1660 74 1716 97
rect 1746 210 1802 222
rect 1746 176 1757 210
rect 1791 176 1802 210
rect 1746 120 1802 176
rect 1746 86 1757 120
rect 1791 86 1802 120
rect 1746 74 1802 86
rect 1832 131 1902 222
rect 1832 97 1843 131
rect 1877 97 1902 131
rect 1832 74 1902 97
rect 1932 210 1989 222
rect 1932 176 1943 210
rect 1977 176 1989 210
rect 1932 120 1989 176
rect 1932 86 1943 120
rect 1977 86 1989 120
rect 1932 74 1989 86
rect 1015 70 1073 74
rect 129 36 187 48
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 508 86 546
rect 27 474 39 508
rect 73 474 86 508
rect 27 424 86 474
rect 116 580 176 592
rect 116 546 129 580
rect 163 546 176 580
rect 116 470 176 546
rect 116 436 129 470
rect 163 436 176 470
rect 116 424 176 436
rect 206 584 266 592
rect 206 550 219 584
rect 253 550 266 584
rect 206 516 266 550
rect 206 482 219 516
rect 253 482 266 516
rect 206 424 266 482
rect 296 580 356 592
rect 296 546 309 580
rect 343 546 356 580
rect 296 470 356 546
rect 296 436 309 470
rect 343 436 356 470
rect 296 424 356 436
rect 386 584 500 592
rect 386 550 417 584
rect 451 550 500 584
rect 386 516 500 550
rect 386 482 417 516
rect 451 482 500 516
rect 386 424 500 482
rect 447 368 500 424
rect 530 582 600 592
rect 530 548 543 582
rect 577 548 600 582
rect 530 514 600 548
rect 530 480 543 514
rect 577 480 600 514
rect 530 446 600 480
rect 530 412 543 446
rect 577 412 600 446
rect 530 368 600 412
rect 630 584 690 592
rect 630 550 643 584
rect 677 550 690 584
rect 630 516 690 550
rect 630 482 643 516
rect 677 482 690 516
rect 630 368 690 482
rect 720 582 780 592
rect 720 548 733 582
rect 767 548 780 582
rect 720 514 780 548
rect 720 480 733 514
rect 767 480 780 514
rect 720 446 780 480
rect 720 412 733 446
rect 767 412 780 446
rect 720 368 780 412
rect 810 584 870 592
rect 810 550 823 584
rect 857 550 870 584
rect 810 516 870 550
rect 810 482 823 516
rect 857 482 870 516
rect 810 368 870 482
rect 900 580 960 592
rect 900 546 913 580
rect 947 546 960 580
rect 900 500 960 546
rect 900 466 913 500
rect 947 466 960 500
rect 900 420 960 466
rect 900 386 913 420
rect 947 386 960 420
rect 900 368 960 386
rect 990 580 1060 592
rect 990 546 1013 580
rect 1047 546 1060 580
rect 990 488 1060 546
rect 990 454 1013 488
rect 1047 454 1060 488
rect 990 368 1060 454
rect 1090 580 1150 592
rect 1090 546 1103 580
rect 1137 546 1150 580
rect 1090 497 1150 546
rect 1090 463 1103 497
rect 1137 463 1150 497
rect 1090 414 1150 463
rect 1090 380 1103 414
rect 1137 380 1150 414
rect 1090 368 1150 380
rect 1180 580 1240 592
rect 1180 546 1193 580
rect 1227 546 1240 580
rect 1180 482 1240 546
rect 1180 448 1193 482
rect 1227 448 1240 482
rect 1180 368 1240 448
rect 1270 580 1330 592
rect 1270 546 1283 580
rect 1317 546 1330 580
rect 1270 497 1330 546
rect 1270 463 1283 497
rect 1317 463 1330 497
rect 1270 414 1330 463
rect 1270 380 1283 414
rect 1317 380 1330 414
rect 1270 368 1330 380
rect 1360 580 1440 592
rect 1360 546 1383 580
rect 1417 546 1440 580
rect 1360 508 1440 546
rect 1360 474 1383 508
rect 1417 474 1440 508
rect 1360 368 1440 474
rect 1470 580 1530 592
rect 1470 546 1483 580
rect 1517 546 1530 580
rect 1470 497 1530 546
rect 1470 463 1483 497
rect 1517 463 1530 497
rect 1470 414 1530 463
rect 1470 380 1483 414
rect 1517 380 1530 414
rect 1470 368 1530 380
rect 1560 580 1630 592
rect 1560 546 1573 580
rect 1607 546 1630 580
rect 1560 508 1630 546
rect 1560 474 1573 508
rect 1607 474 1630 508
rect 1560 368 1630 474
rect 1660 580 1720 592
rect 1660 546 1673 580
rect 1707 546 1720 580
rect 1660 510 1720 546
rect 1660 476 1673 510
rect 1707 476 1720 510
rect 1660 440 1720 476
rect 1660 406 1673 440
rect 1707 406 1720 440
rect 1660 368 1720 406
rect 1750 580 1810 592
rect 1750 546 1763 580
rect 1797 546 1810 580
rect 1750 508 1810 546
rect 1750 474 1763 508
rect 1797 474 1810 508
rect 1750 368 1810 474
rect 1840 580 1900 592
rect 1840 546 1853 580
rect 1887 546 1900 580
rect 1840 510 1900 546
rect 1840 476 1853 510
rect 1887 476 1900 510
rect 1840 440 1900 476
rect 1840 406 1853 440
rect 1887 406 1900 440
rect 1840 368 1900 406
rect 1930 580 1989 592
rect 1930 546 1943 580
rect 1977 546 1989 580
rect 1930 510 1989 546
rect 1930 476 1943 510
rect 1977 476 1989 510
rect 1930 440 1989 476
rect 1930 406 1943 440
rect 1977 406 1989 440
rect 1930 368 1989 406
<< ndiffc >>
rect 39 206 73 240
rect 39 126 73 160
rect 246 216 280 250
rect 386 158 420 192
rect 141 48 175 82
rect 386 86 420 120
rect 480 146 514 180
rect 580 88 614 122
rect 667 155 701 189
rect 753 110 787 144
rect 839 82 873 116
rect 925 150 959 184
rect 1027 82 1061 116
rect 1129 126 1163 160
rect 1241 155 1275 189
rect 1327 99 1361 133
rect 1413 155 1447 189
rect 1499 99 1533 133
rect 1585 176 1619 210
rect 1585 86 1619 120
rect 1671 97 1705 131
rect 1757 176 1791 210
rect 1757 86 1791 120
rect 1843 97 1877 131
rect 1943 176 1977 210
rect 1943 86 1977 120
<< pdiffc >>
rect 39 546 73 580
rect 39 474 73 508
rect 129 546 163 580
rect 129 436 163 470
rect 219 550 253 584
rect 219 482 253 516
rect 309 546 343 580
rect 309 436 343 470
rect 417 550 451 584
rect 417 482 451 516
rect 543 548 577 582
rect 543 480 577 514
rect 543 412 577 446
rect 643 550 677 584
rect 643 482 677 516
rect 733 548 767 582
rect 733 480 767 514
rect 733 412 767 446
rect 823 550 857 584
rect 823 482 857 516
rect 913 546 947 580
rect 913 466 947 500
rect 913 386 947 420
rect 1013 546 1047 580
rect 1013 454 1047 488
rect 1103 546 1137 580
rect 1103 463 1137 497
rect 1103 380 1137 414
rect 1193 546 1227 580
rect 1193 448 1227 482
rect 1283 546 1317 580
rect 1283 463 1317 497
rect 1283 380 1317 414
rect 1383 546 1417 580
rect 1383 474 1417 508
rect 1483 546 1517 580
rect 1483 463 1517 497
rect 1483 380 1517 414
rect 1573 546 1607 580
rect 1573 474 1607 508
rect 1673 546 1707 580
rect 1673 476 1707 510
rect 1673 406 1707 440
rect 1763 546 1797 580
rect 1763 474 1797 508
rect 1853 546 1887 580
rect 1853 476 1887 510
rect 1853 406 1887 440
rect 1943 546 1977 580
rect 1943 476 1977 510
rect 1943 406 1977 440
<< poly >>
rect 86 592 116 618
rect 176 592 206 618
rect 266 592 296 618
rect 356 592 386 618
rect 500 592 530 618
rect 600 592 630 618
rect 690 592 720 618
rect 780 592 810 618
rect 870 592 900 618
rect 960 592 990 618
rect 1060 592 1090 618
rect 1150 592 1180 618
rect 1240 592 1270 618
rect 1330 592 1360 618
rect 1440 592 1470 618
rect 1530 592 1560 618
rect 1630 592 1660 618
rect 1720 592 1750 618
rect 1810 592 1840 618
rect 1900 592 1930 618
rect 86 409 116 424
rect 176 409 206 424
rect 266 409 296 424
rect 356 409 386 424
rect 83 379 209 409
rect 263 393 299 409
rect 353 393 386 409
rect 84 340 154 379
rect 84 306 104 340
rect 138 306 154 340
rect 263 363 383 393
rect 263 360 359 363
rect 263 331 309 360
rect 84 290 154 306
rect 202 326 309 331
rect 343 326 359 360
rect 500 353 530 368
rect 600 353 630 368
rect 690 353 720 368
rect 780 353 810 368
rect 870 353 900 368
rect 960 353 990 368
rect 1060 353 1090 368
rect 1150 353 1180 368
rect 1240 353 1270 368
rect 1330 353 1360 368
rect 1440 353 1470 368
rect 1530 353 1560 368
rect 1630 353 1660 368
rect 1720 353 1750 368
rect 1810 353 1840 368
rect 1900 353 1930 368
rect 497 345 533 353
rect 597 345 633 353
rect 687 345 723 353
rect 777 345 813 353
rect 202 301 359 326
rect 431 315 813 345
rect 867 336 903 353
rect 957 336 993 353
rect 1057 336 1093 353
rect 1147 336 1183 353
rect 867 320 1183 336
rect 84 262 114 290
rect 202 262 232 301
rect 431 294 742 315
rect 431 260 447 294
rect 481 260 515 294
rect 549 260 583 294
rect 617 265 742 294
rect 867 286 883 320
rect 917 286 951 320
rect 985 286 1019 320
rect 1053 306 1183 320
rect 1237 330 1273 353
rect 1327 330 1363 353
rect 1437 330 1473 353
rect 1527 330 1563 353
rect 1237 314 1563 330
rect 1053 286 1118 306
rect 867 267 1118 286
rect 617 260 656 265
rect 431 244 656 260
rect 431 222 461 244
rect 538 222 568 244
rect 626 222 656 244
rect 712 222 742 265
rect 798 237 1118 267
rect 1237 280 1268 314
rect 1302 280 1336 314
rect 1370 280 1404 314
rect 1438 280 1472 314
rect 1506 294 1563 314
rect 1627 326 1663 353
rect 1717 326 1753 353
rect 1807 326 1843 353
rect 1897 326 1933 353
rect 1627 310 1986 326
rect 1627 296 1664 310
rect 1506 280 1574 294
rect 1237 264 1574 280
rect 798 222 828 237
rect 884 222 914 237
rect 970 222 1000 237
rect 1088 222 1118 237
rect 1286 222 1316 264
rect 1372 222 1402 264
rect 1458 222 1488 264
rect 1544 222 1574 264
rect 1630 276 1664 296
rect 1698 276 1732 310
rect 1766 276 1800 310
rect 1834 276 1868 310
rect 1902 276 1936 310
rect 1970 276 1986 310
rect 1630 260 1986 276
rect 1630 222 1660 260
rect 1716 222 1746 260
rect 1802 222 1832 260
rect 1902 222 1932 260
rect 84 88 114 114
rect 202 88 232 114
rect 431 48 461 74
rect 538 48 568 74
rect 626 48 656 74
rect 712 48 742 74
rect 798 48 828 74
rect 884 48 914 74
rect 970 48 1000 74
rect 1088 48 1118 74
rect 1286 48 1316 74
rect 1372 48 1402 74
rect 1458 48 1488 74
rect 1544 48 1574 74
rect 1630 48 1660 74
rect 1716 48 1746 74
rect 1802 48 1832 74
rect 1902 48 1932 74
<< polycont >>
rect 104 306 138 340
rect 309 326 343 360
rect 447 260 481 294
rect 515 260 549 294
rect 583 260 617 294
rect 883 286 917 320
rect 951 286 985 320
rect 1019 286 1053 320
rect 1268 280 1302 314
rect 1336 280 1370 314
rect 1404 280 1438 314
rect 1472 280 1506 314
rect 1664 276 1698 310
rect 1732 276 1766 310
rect 1800 276 1834 310
rect 1868 276 1902 310
rect 1936 276 1970 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 23 580 89 649
rect 23 546 39 580
rect 73 546 89 580
rect 23 508 89 546
rect 23 474 39 508
rect 73 474 89 508
rect 23 458 89 474
rect 129 580 163 596
rect 129 470 163 546
rect 203 584 269 649
rect 203 550 219 584
rect 253 550 269 584
rect 203 516 269 550
rect 203 482 219 516
rect 253 482 269 516
rect 203 478 269 482
rect 303 580 359 596
rect 303 546 309 580
rect 343 546 359 580
rect 303 470 359 546
rect 401 584 467 649
rect 401 550 417 584
rect 451 550 467 584
rect 401 516 467 550
rect 401 482 417 516
rect 451 482 467 516
rect 401 478 467 482
rect 505 582 593 598
rect 505 548 543 582
rect 577 548 593 582
rect 505 514 593 548
rect 505 480 543 514
rect 577 480 593 514
rect 627 584 693 649
rect 627 550 643 584
rect 677 550 693 584
rect 627 516 693 550
rect 627 482 643 516
rect 677 482 693 516
rect 627 480 693 482
rect 727 582 773 598
rect 727 548 733 582
rect 767 548 773 582
rect 727 514 773 548
rect 727 480 733 514
rect 767 480 773 514
rect 807 584 873 649
rect 807 550 823 584
rect 857 550 873 584
rect 807 516 873 550
rect 807 482 823 516
rect 857 482 873 516
rect 807 480 873 482
rect 907 580 963 596
rect 907 546 913 580
rect 947 546 963 580
rect 907 500 963 546
rect 303 444 309 470
rect 129 424 163 436
rect 20 390 163 424
rect 225 436 309 444
rect 343 444 359 470
rect 505 446 593 480
rect 727 446 773 480
rect 907 466 913 500
rect 947 466 963 500
rect 907 446 963 466
rect 343 436 427 444
rect 225 410 427 436
rect 505 412 543 446
rect 577 412 733 446
rect 767 420 963 446
rect 997 580 1063 649
rect 997 546 1013 580
rect 1047 546 1063 580
rect 997 488 1063 546
rect 997 454 1013 488
rect 1047 454 1063 488
rect 997 438 1063 454
rect 1103 580 1137 596
rect 1103 497 1137 546
rect 767 412 913 420
rect 20 256 54 390
rect 88 340 167 356
rect 88 306 104 340
rect 138 306 167 340
rect 88 290 167 306
rect 225 266 259 410
rect 393 378 427 410
rect 897 386 913 412
rect 947 404 963 420
rect 1103 414 1137 463
rect 1177 580 1227 649
rect 1177 546 1193 580
rect 1177 482 1227 546
rect 1177 448 1193 482
rect 1177 432 1227 448
rect 1267 580 1333 596
rect 1267 546 1283 580
rect 1317 546 1333 580
rect 1267 497 1333 546
rect 1267 463 1283 497
rect 1317 463 1333 497
rect 947 386 1103 404
rect 897 380 1103 386
rect 1267 424 1333 463
rect 1367 580 1433 649
rect 1367 546 1383 580
rect 1417 546 1433 580
rect 1367 508 1433 546
rect 1367 474 1383 508
rect 1417 474 1433 508
rect 1367 458 1433 474
rect 1467 580 1533 596
rect 1467 546 1483 580
rect 1517 546 1533 580
rect 1467 497 1533 546
rect 1467 463 1483 497
rect 1517 463 1533 497
rect 1467 424 1533 463
rect 1573 580 1623 649
rect 1607 546 1623 580
rect 1573 508 1623 546
rect 1607 474 1623 508
rect 1573 458 1623 474
rect 1657 580 1723 596
rect 1657 546 1673 580
rect 1707 546 1723 580
rect 1657 510 1723 546
rect 1657 476 1673 510
rect 1707 476 1723 510
rect 1657 440 1723 476
rect 1763 580 1797 649
rect 1763 508 1797 546
rect 1763 458 1797 474
rect 1837 580 1903 596
rect 1837 546 1853 580
rect 1887 546 1903 580
rect 1837 510 1903 546
rect 1837 476 1853 510
rect 1887 476 1903 510
rect 1657 424 1673 440
rect 1267 414 1673 424
rect 1267 398 1283 414
rect 1137 380 1283 398
rect 1317 390 1483 414
rect 1317 380 1333 390
rect 293 360 359 376
rect 293 326 309 360
rect 343 326 359 360
rect 393 344 863 378
rect 897 370 1333 380
rect 293 310 359 326
rect 829 336 863 344
rect 1103 364 1333 370
rect 1467 380 1483 390
rect 1517 406 1673 414
rect 1707 424 1723 440
rect 1837 440 1903 476
rect 1837 424 1853 440
rect 1707 406 1853 424
rect 1887 406 1903 440
rect 1517 390 1903 406
rect 1943 580 1993 649
rect 1977 546 1993 580
rect 1943 510 1993 546
rect 1977 476 1993 510
rect 1943 440 1993 476
rect 1977 406 1993 440
rect 1943 390 1993 406
rect 1517 380 1533 390
rect 1467 364 1533 380
rect 829 320 1069 336
rect 431 294 633 310
rect 431 276 447 294
rect 20 240 89 256
rect 20 206 39 240
rect 73 206 89 240
rect 20 166 89 206
rect 225 250 284 266
rect 225 216 246 250
rect 280 216 284 250
rect 225 200 284 216
rect 318 260 447 276
rect 481 260 515 294
rect 549 260 583 294
rect 617 260 633 294
rect 829 286 883 320
rect 917 286 951 320
rect 985 286 1019 320
rect 1053 286 1069 320
rect 318 242 633 260
rect 1103 252 1137 364
rect 1369 330 1415 356
rect 1237 314 1522 330
rect 1237 280 1268 314
rect 1302 280 1336 314
rect 1370 280 1404 314
rect 1438 280 1472 314
rect 1506 280 1522 314
rect 1237 264 1522 280
rect 1653 310 1991 356
rect 1653 276 1664 310
rect 1698 276 1732 310
rect 1766 276 1800 310
rect 1834 276 1868 310
rect 1902 276 1936 310
rect 1970 276 1991 310
rect 1653 260 1991 276
rect 318 166 352 242
rect 667 218 1137 252
rect 1225 226 1619 230
rect 667 208 701 218
rect 20 160 352 166
rect 20 126 39 160
rect 73 132 352 160
rect 386 192 420 208
rect 73 126 89 132
rect 20 110 89 126
rect 386 120 420 158
rect 125 82 191 98
rect 125 48 141 82
rect 175 48 191 82
rect 464 189 701 208
rect 464 180 667 189
rect 464 146 480 180
rect 514 174 667 180
rect 514 146 530 174
rect 464 119 530 146
rect 1225 210 1993 226
rect 1225 196 1585 210
rect 1225 189 1275 196
rect 564 122 630 140
rect 386 85 420 86
rect 564 88 580 122
rect 614 88 630 122
rect 667 119 701 155
rect 737 150 925 184
rect 959 160 1179 184
rect 959 150 1129 160
rect 737 144 787 150
rect 564 85 630 88
rect 737 110 753 144
rect 1113 126 1129 150
rect 1163 126 1179 160
rect 1113 119 1179 126
rect 1225 155 1241 189
rect 1413 189 1447 196
rect 1225 119 1275 155
rect 1311 133 1377 162
rect 737 85 787 110
rect 386 51 787 85
rect 823 82 839 116
rect 873 82 1027 116
rect 1061 85 1077 116
rect 1311 99 1327 133
rect 1361 99 1377 133
rect 1619 192 1757 210
rect 1413 119 1447 155
rect 1483 133 1549 162
rect 1311 85 1377 99
rect 1483 99 1499 133
rect 1533 99 1549 133
rect 1483 85 1549 99
rect 1061 82 1549 85
rect 823 51 1549 82
rect 1585 120 1619 176
rect 1791 192 1943 210
rect 1585 70 1619 86
rect 1655 131 1721 158
rect 1655 97 1671 131
rect 1705 97 1721 131
rect 125 17 191 48
rect 1655 17 1721 97
rect 1757 120 1791 176
rect 1927 176 1943 192
rect 1977 176 1993 210
rect 1757 70 1791 86
rect 1827 131 1893 158
rect 1827 97 1843 131
rect 1877 97 1893 131
rect 1827 17 1893 97
rect 1927 120 1993 176
rect 1927 86 1943 120
rect 1977 86 1993 120
rect 1927 70 1993 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
rlabel comment s 0 0 0 0 4 nand4bb_4
flabel pwell s 0 0 2016 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nwell s 0 617 2016 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 2016 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 2016 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 1375 316 1409 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 1663 316 1697 350 0 FreeSans 340 0 0 0 D
port 4 nsew
flabel corelocali s 1759 316 1793 350 0 FreeSans 340 0 0 0 D
port 4 nsew
flabel corelocali s 1855 316 1889 350 0 FreeSans 340 0 0 0 D
port 4 nsew
flabel corelocali s 1951 316 1985 350 0 FreeSans 340 0 0 0 D
port 4 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 B_N
port 2 nsew
flabel corelocali s 511 464 545 498 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 511 538 545 572 0 FreeSans 340 0 0 0 Y
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 2016 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1511178
string GDS_START 1495272
<< end >>
