magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 1670 704
<< pwell >>
rect 0 0 1632 49
<< scnmos >>
rect 83 98 113 246
rect 169 98 199 246
rect 285 98 315 246
rect 371 98 401 246
rect 486 98 516 246
rect 572 98 602 246
rect 808 74 838 222
rect 894 74 924 222
rect 980 74 1010 222
rect 1066 74 1096 222
rect 1261 74 1291 222
rect 1347 74 1377 222
rect 1433 74 1463 222
rect 1519 74 1549 222
<< pmoshvt >>
rect 86 392 116 592
rect 186 392 216 592
rect 388 368 418 592
rect 478 368 508 592
rect 568 368 598 592
rect 658 368 688 592
rect 762 392 792 592
rect 891 392 921 592
rect 1026 392 1056 592
rect 1116 392 1146 592
rect 1226 392 1256 592
rect 1326 392 1356 592
rect 1426 392 1456 592
rect 1516 392 1546 592
<< ndiff >>
rect 27 234 83 246
rect 27 200 38 234
rect 72 200 83 234
rect 27 144 83 200
rect 27 110 38 144
rect 72 110 83 144
rect 27 98 83 110
rect 113 234 169 246
rect 113 200 124 234
rect 158 200 169 234
rect 113 144 169 200
rect 113 110 124 144
rect 158 110 169 144
rect 113 98 169 110
rect 199 98 285 246
rect 315 234 371 246
rect 315 200 326 234
rect 360 200 371 234
rect 315 98 371 200
rect 401 98 486 246
rect 516 234 572 246
rect 516 200 527 234
rect 561 200 572 234
rect 516 98 572 200
rect 602 98 673 246
rect 214 92 270 98
rect 214 58 225 92
rect 259 58 270 92
rect 416 92 471 98
rect 214 46 270 58
rect 416 58 427 92
rect 461 58 471 92
rect 617 82 673 98
rect 416 46 471 58
rect 617 48 627 82
rect 661 48 673 82
rect 751 190 808 222
rect 751 156 763 190
rect 797 156 808 190
rect 751 74 808 156
rect 838 120 894 222
rect 838 86 849 120
rect 883 86 894 120
rect 838 74 894 86
rect 924 214 980 222
rect 924 180 935 214
rect 969 180 980 214
rect 924 116 980 180
rect 924 82 935 116
rect 969 82 980 116
rect 924 74 980 82
rect 1010 204 1066 222
rect 1010 170 1021 204
rect 1055 170 1066 204
rect 1010 74 1066 170
rect 1096 188 1151 222
rect 1096 154 1107 188
rect 1141 154 1151 188
rect 1096 120 1151 154
rect 1096 86 1107 120
rect 1141 86 1151 120
rect 1096 74 1151 86
rect 1205 188 1261 222
rect 1205 154 1216 188
rect 1250 154 1261 188
rect 1205 120 1261 154
rect 1205 86 1216 120
rect 1250 86 1261 120
rect 1205 74 1261 86
rect 1291 174 1347 222
rect 1291 140 1302 174
rect 1336 140 1347 174
rect 1291 74 1347 140
rect 1377 210 1433 222
rect 1377 176 1388 210
rect 1422 176 1433 210
rect 1377 120 1433 176
rect 1377 86 1388 120
rect 1422 86 1433 120
rect 1377 74 1433 86
rect 1463 184 1519 222
rect 1463 150 1474 184
rect 1508 150 1519 184
rect 1463 116 1519 150
rect 1463 82 1474 116
rect 1508 82 1519 116
rect 1463 74 1519 82
rect 1549 210 1605 222
rect 1549 176 1560 210
rect 1594 176 1605 210
rect 1549 120 1605 176
rect 1549 86 1560 120
rect 1594 86 1605 120
rect 1549 74 1605 86
rect 617 36 673 48
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 510 86 546
rect 27 476 39 510
rect 73 476 86 510
rect 27 440 86 476
rect 27 406 39 440
rect 73 406 86 440
rect 27 392 86 406
rect 116 531 186 592
rect 116 497 139 531
rect 173 497 186 531
rect 116 440 186 497
rect 116 406 139 440
rect 173 406 186 440
rect 116 392 186 406
rect 216 580 275 592
rect 216 546 229 580
rect 263 546 275 580
rect 216 509 275 546
rect 216 475 229 509
rect 263 475 275 509
rect 216 438 275 475
rect 216 404 229 438
rect 263 404 275 438
rect 216 392 275 404
rect 329 568 388 592
rect 329 534 341 568
rect 375 534 388 568
rect 329 368 388 534
rect 418 421 478 592
rect 418 387 431 421
rect 465 387 478 421
rect 418 368 478 387
rect 508 568 568 592
rect 508 534 521 568
rect 555 534 568 568
rect 508 368 568 534
rect 598 419 658 592
rect 598 385 611 419
rect 645 385 658 419
rect 598 368 658 385
rect 688 570 762 592
rect 688 536 703 570
rect 737 536 762 570
rect 688 392 762 536
rect 792 580 891 592
rect 792 546 825 580
rect 859 546 891 580
rect 792 508 891 546
rect 792 474 825 508
rect 859 474 891 508
rect 792 440 891 474
rect 792 406 825 440
rect 859 406 891 440
rect 792 392 891 406
rect 921 580 1026 592
rect 921 546 956 580
rect 990 546 1026 580
rect 921 492 1026 546
rect 921 458 956 492
rect 990 458 1026 492
rect 921 392 1026 458
rect 1056 580 1116 592
rect 1056 546 1069 580
rect 1103 546 1116 580
rect 1056 510 1116 546
rect 1056 476 1069 510
rect 1103 476 1116 510
rect 1056 440 1116 476
rect 1056 406 1069 440
rect 1103 406 1116 440
rect 1056 392 1116 406
rect 1146 580 1226 592
rect 1146 546 1169 580
rect 1203 546 1226 580
rect 1146 500 1226 546
rect 1146 466 1169 500
rect 1203 466 1226 500
rect 1146 392 1226 466
rect 1256 580 1326 592
rect 1256 546 1269 580
rect 1303 546 1326 580
rect 1256 510 1326 546
rect 1256 476 1269 510
rect 1303 476 1326 510
rect 1256 440 1326 476
rect 1256 406 1269 440
rect 1303 406 1326 440
rect 1256 392 1326 406
rect 1356 580 1426 592
rect 1356 546 1369 580
rect 1403 546 1426 580
rect 1356 500 1426 546
rect 1356 466 1369 500
rect 1403 466 1426 500
rect 1356 392 1426 466
rect 1456 580 1516 592
rect 1456 546 1469 580
rect 1503 546 1516 580
rect 1456 510 1516 546
rect 1456 476 1469 510
rect 1503 476 1516 510
rect 1456 440 1516 476
rect 1456 406 1469 440
rect 1503 406 1516 440
rect 1456 392 1516 406
rect 1546 580 1605 592
rect 1546 546 1559 580
rect 1593 546 1605 580
rect 1546 510 1605 546
rect 1546 476 1559 510
rect 1593 476 1605 510
rect 1546 440 1605 476
rect 1546 406 1559 440
rect 1593 406 1605 440
rect 1546 392 1605 406
rect 688 368 741 392
<< ndiffc >>
rect 38 200 72 234
rect 38 110 72 144
rect 124 200 158 234
rect 124 110 158 144
rect 326 200 360 234
rect 527 200 561 234
rect 225 58 259 92
rect 427 58 461 92
rect 627 48 661 82
rect 763 156 797 190
rect 849 86 883 120
rect 935 180 969 214
rect 935 82 969 116
rect 1021 170 1055 204
rect 1107 154 1141 188
rect 1107 86 1141 120
rect 1216 154 1250 188
rect 1216 86 1250 120
rect 1302 140 1336 174
rect 1388 176 1422 210
rect 1388 86 1422 120
rect 1474 150 1508 184
rect 1474 82 1508 116
rect 1560 176 1594 210
rect 1560 86 1594 120
<< pdiffc >>
rect 39 546 73 580
rect 39 476 73 510
rect 39 406 73 440
rect 139 497 173 531
rect 139 406 173 440
rect 229 546 263 580
rect 229 475 263 509
rect 229 404 263 438
rect 341 534 375 568
rect 431 387 465 421
rect 521 534 555 568
rect 611 385 645 419
rect 703 536 737 570
rect 825 546 859 580
rect 825 474 859 508
rect 825 406 859 440
rect 956 546 990 580
rect 956 458 990 492
rect 1069 546 1103 580
rect 1069 476 1103 510
rect 1069 406 1103 440
rect 1169 546 1203 580
rect 1169 466 1203 500
rect 1269 546 1303 580
rect 1269 476 1303 510
rect 1269 406 1303 440
rect 1369 546 1403 580
rect 1369 466 1403 500
rect 1469 546 1503 580
rect 1469 476 1503 510
rect 1469 406 1503 440
rect 1559 546 1593 580
rect 1559 476 1593 510
rect 1559 406 1593 440
<< poly >>
rect 86 592 116 618
rect 186 592 216 618
rect 388 592 418 618
rect 478 592 508 618
rect 568 592 598 618
rect 658 592 688 618
rect 762 592 792 618
rect 891 592 921 618
rect 1026 592 1056 618
rect 1116 592 1146 618
rect 1226 592 1256 618
rect 1326 592 1356 618
rect 1426 592 1456 618
rect 1516 592 1546 618
rect 86 377 116 392
rect 186 377 216 392
rect 83 356 119 377
rect 44 351 119 356
rect 183 351 219 377
rect 762 377 792 392
rect 891 377 921 392
rect 1026 377 1056 392
rect 1116 377 1146 392
rect 1226 377 1256 392
rect 1326 377 1356 392
rect 1426 377 1456 392
rect 1516 377 1546 392
rect 388 353 418 368
rect 478 353 508 368
rect 568 353 598 368
rect 658 353 688 368
rect 759 356 795 377
rect 888 356 924 377
rect 1023 356 1059 377
rect 1113 356 1149 377
rect 44 340 219 351
rect 44 306 60 340
rect 94 306 219 340
rect 385 334 421 353
rect 475 334 511 353
rect 565 334 601 353
rect 655 334 691 353
rect 44 290 219 306
rect 275 318 691 334
rect 83 246 113 290
rect 169 246 199 290
rect 275 284 291 318
rect 325 284 359 318
rect 393 284 427 318
rect 461 284 691 318
rect 759 340 924 356
rect 759 306 789 340
rect 823 306 924 340
rect 759 290 924 306
rect 275 268 691 284
rect 285 246 315 268
rect 371 246 401 268
rect 486 246 516 268
rect 572 246 602 268
rect 808 222 838 290
rect 894 222 924 290
rect 980 340 1149 356
rect 980 306 996 340
rect 1030 326 1149 340
rect 1223 356 1259 377
rect 1323 356 1359 377
rect 1423 356 1459 377
rect 1513 356 1549 377
rect 1223 340 1377 356
rect 1030 306 1096 326
rect 980 290 1096 306
rect 1223 306 1239 340
rect 1273 306 1307 340
rect 1341 306 1377 340
rect 1223 290 1377 306
rect 1423 340 1549 356
rect 1423 306 1481 340
rect 1515 306 1549 340
rect 1423 290 1549 306
rect 980 222 1010 290
rect 1066 222 1096 290
rect 1261 222 1291 290
rect 1347 222 1377 290
rect 1433 222 1463 290
rect 1519 222 1549 290
rect 83 72 113 98
rect 169 72 199 98
rect 285 72 315 98
rect 371 72 401 98
rect 486 72 516 98
rect 572 72 602 98
rect 808 48 838 74
rect 894 48 924 74
rect 980 48 1010 74
rect 1066 48 1096 74
rect 1261 48 1291 74
rect 1347 48 1377 74
rect 1433 48 1463 74
rect 1519 48 1549 74
<< polycont >>
rect 60 306 94 340
rect 291 284 325 318
rect 359 284 393 318
rect 427 284 461 318
rect 789 306 823 340
rect 996 306 1030 340
rect 1239 306 1273 340
rect 1307 306 1341 340
rect 1481 306 1515 340
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 23 581 279 615
rect 23 580 89 581
rect 23 546 39 580
rect 73 546 89 580
rect 213 580 279 581
rect 23 510 89 546
rect 23 476 39 510
rect 73 476 89 510
rect 23 440 89 476
rect 23 406 39 440
rect 73 406 89 440
rect 23 390 89 406
rect 123 531 178 547
rect 123 497 139 531
rect 173 497 178 531
rect 123 440 178 497
rect 123 406 139 440
rect 173 406 178 440
rect 123 390 178 406
rect 25 340 110 356
rect 25 306 60 340
rect 94 306 110 340
rect 25 290 110 306
rect 144 334 178 390
rect 213 546 229 580
rect 263 546 279 580
rect 213 509 279 546
rect 325 568 391 649
rect 325 534 341 568
rect 375 534 391 568
rect 325 526 391 534
rect 505 568 571 649
rect 505 534 521 568
rect 555 534 571 568
rect 505 526 571 534
rect 685 570 755 649
rect 685 536 703 570
rect 737 536 755 570
rect 685 530 755 536
rect 809 580 875 596
rect 809 546 825 580
rect 859 546 875 580
rect 213 475 229 509
rect 263 492 279 509
rect 809 508 875 546
rect 809 492 825 508
rect 263 475 825 492
rect 213 474 825 475
rect 859 474 875 508
rect 213 458 875 474
rect 927 580 1019 649
rect 927 546 956 580
rect 990 546 1019 580
rect 927 492 1019 546
rect 927 458 956 492
rect 990 458 1019 492
rect 1053 580 1119 596
rect 1053 546 1069 580
rect 1103 546 1119 580
rect 1053 510 1119 546
rect 1053 476 1069 510
rect 1103 476 1119 510
rect 213 438 279 458
rect 213 404 229 438
rect 263 404 279 438
rect 809 440 875 458
rect 213 388 279 404
rect 415 421 661 424
rect 415 387 431 421
rect 465 419 661 421
rect 465 387 611 419
rect 415 385 611 387
rect 645 385 661 419
rect 809 406 825 440
rect 859 424 875 440
rect 1053 440 1119 476
rect 1153 580 1219 649
rect 1153 546 1169 580
rect 1203 546 1219 580
rect 1153 500 1219 546
rect 1153 466 1169 500
rect 1203 466 1219 500
rect 1153 458 1219 466
rect 1253 580 1319 596
rect 1253 546 1269 580
rect 1303 546 1319 580
rect 1253 510 1319 546
rect 1253 476 1269 510
rect 1303 476 1319 510
rect 1053 424 1069 440
rect 859 406 1069 424
rect 1103 424 1119 440
rect 1253 440 1319 476
rect 1353 580 1419 649
rect 1353 546 1369 580
rect 1403 546 1419 580
rect 1353 500 1419 546
rect 1353 466 1369 500
rect 1403 466 1419 500
rect 1353 458 1419 466
rect 1453 580 1519 596
rect 1453 546 1469 580
rect 1503 546 1519 580
rect 1453 510 1519 546
rect 1453 476 1469 510
rect 1503 476 1519 510
rect 1253 424 1269 440
rect 1103 406 1269 424
rect 1303 424 1319 440
rect 1453 440 1519 476
rect 1453 424 1469 440
rect 1303 406 1469 424
rect 1503 406 1519 440
rect 809 390 1519 406
rect 1559 580 1609 649
rect 1593 546 1609 580
rect 1559 510 1609 546
rect 1593 476 1609 510
rect 1559 440 1609 476
rect 1593 406 1609 440
rect 1559 390 1609 406
rect 415 368 661 385
rect 144 318 477 334
rect 144 284 291 318
rect 325 284 359 318
rect 393 284 427 318
rect 461 284 477 318
rect 144 268 477 284
rect 144 250 245 268
rect 22 234 72 250
rect 22 200 38 234
rect 22 144 72 200
rect 22 110 38 144
rect 22 17 72 110
rect 108 234 245 250
rect 511 234 661 368
rect 697 340 839 356
rect 697 306 789 340
rect 823 306 839 340
rect 697 290 839 306
rect 980 340 1127 356
rect 980 306 996 340
rect 1030 306 1127 340
rect 980 290 1127 306
rect 1177 340 1415 356
rect 1177 306 1239 340
rect 1273 306 1307 340
rect 1341 306 1415 340
rect 1177 290 1415 306
rect 1465 340 1607 356
rect 1465 306 1481 340
rect 1515 306 1607 340
rect 1465 290 1607 306
rect 108 200 124 234
rect 158 200 245 234
rect 310 200 326 234
rect 360 200 527 234
rect 561 200 661 234
rect 763 214 969 230
rect 108 166 245 200
rect 763 190 935 214
rect 108 144 729 166
rect 108 110 124 144
rect 158 132 729 144
rect 797 180 935 190
rect 797 156 969 180
rect 763 154 969 156
rect 1005 222 1336 256
rect 1005 204 1057 222
rect 1005 170 1021 204
rect 1055 170 1057 204
rect 1005 154 1057 170
rect 1091 154 1107 188
rect 1141 154 1157 188
rect 763 140 797 154
rect 158 110 174 132
rect 108 94 174 110
rect 209 92 275 98
rect 209 58 225 92
rect 259 58 275 92
rect 209 17 275 58
rect 411 92 477 98
rect 411 58 427 92
rect 461 58 477 92
rect 411 17 477 58
rect 611 82 661 98
rect 611 48 627 82
rect 695 85 729 132
rect 935 120 969 154
rect 1091 120 1157 154
rect 833 86 849 120
rect 883 86 899 120
rect 833 85 899 86
rect 695 51 899 85
rect 935 116 1107 120
rect 969 86 1107 116
rect 1141 86 1157 120
rect 969 82 1157 86
rect 935 66 1157 82
rect 1200 154 1216 188
rect 1250 154 1266 188
rect 1200 120 1266 154
rect 1200 86 1216 120
rect 1250 86 1266 120
rect 1302 174 1336 222
rect 1302 119 1336 140
rect 1372 222 1610 256
rect 1372 210 1422 222
rect 1372 176 1388 210
rect 1558 210 1610 222
rect 1372 120 1422 176
rect 1200 85 1266 86
rect 1372 86 1388 120
rect 1372 85 1422 86
rect 1200 51 1422 85
rect 1458 184 1524 188
rect 1458 150 1474 184
rect 1508 150 1524 184
rect 1458 116 1524 150
rect 1458 82 1474 116
rect 1508 82 1524 116
rect 611 17 661 48
rect 1458 17 1524 82
rect 1558 176 1560 210
rect 1594 176 1610 210
rect 1558 120 1610 176
rect 1558 86 1560 120
rect 1594 86 1610 120
rect 1558 70 1610 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a41o_4
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nwell s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 X
port 10 nsew
flabel corelocali s 1183 316 1217 350 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 1279 316 1313 350 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 1375 316 1409 350 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 1471 316 1505 350 0 FreeSans 340 0 0 0 A4
port 4 nsew
flabel corelocali s 1567 316 1601 350 0 FreeSans 340 0 0 0 A4
port 4 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 B1
port 5 nsew
flabel corelocali s 607 390 641 424 0 FreeSans 340 0 0 0 X
port 10 nsew
flabel corelocali s 607 242 641 276 0 FreeSans 340 0 0 0 X
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 1632 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3781754
string GDS_START 3768376
<< end >>
