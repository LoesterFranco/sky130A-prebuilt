magic
tech sky130A
magscale 1 2
timestamp 1601050082
<< locali >>
rect 91 212 167 356
rect 313 290 417 356
rect 895 290 973 356
rect 1015 236 1127 302
rect 1315 236 1415 310
rect 2969 364 3048 596
rect 3172 364 3247 596
rect 2969 124 3003 364
rect 3213 230 3247 364
rect 3175 74 3247 230
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3264 683
rect 23 492 89 596
rect 191 526 241 649
rect 275 581 445 615
rect 275 492 309 581
rect 23 458 309 492
rect 23 162 57 458
rect 343 424 377 547
rect 411 496 445 581
rect 479 530 529 649
rect 637 496 709 596
rect 411 462 709 496
rect 205 390 533 424
rect 205 256 271 390
rect 467 305 533 390
rect 575 305 641 428
rect 675 269 709 462
rect 205 222 408 256
rect 23 96 132 162
rect 230 17 296 178
rect 342 109 408 222
rect 606 235 709 269
rect 743 581 957 615
rect 743 460 793 581
rect 442 17 508 201
rect 606 109 672 235
rect 743 201 777 460
rect 827 458 889 547
rect 923 492 957 581
rect 991 526 1041 649
rect 1143 496 1209 594
rect 1255 530 1321 649
rect 1533 530 1599 649
rect 1633 546 1804 596
rect 1633 496 1667 546
rect 1838 512 1904 596
rect 2016 546 2082 649
rect 2235 546 2301 649
rect 1143 492 1667 496
rect 923 462 1667 492
rect 1808 478 1904 512
rect 1938 478 2519 512
rect 2553 504 2639 596
rect 2728 530 2846 649
rect 923 458 1242 462
rect 827 424 861 458
rect 706 109 777 201
rect 811 390 1174 424
rect 811 213 861 390
rect 1113 358 1174 390
rect 811 121 948 213
rect 1208 202 1242 458
rect 1345 364 1505 428
rect 1411 362 1505 364
rect 1471 202 1505 362
rect 1555 330 1589 462
rect 1717 428 1774 476
rect 1623 364 1774 428
rect 1555 296 1706 330
rect 811 82 861 121
rect 982 17 1048 202
rect 1148 121 1242 202
rect 1276 17 1310 202
rect 1346 168 1505 202
rect 1346 70 1412 168
rect 1458 17 1524 134
rect 1560 85 1610 226
rect 1656 119 1706 296
rect 1740 85 1774 364
rect 1808 358 1842 478
rect 1938 444 1972 478
rect 1876 392 1972 444
rect 2123 410 2214 444
rect 2080 358 2146 366
rect 1808 324 2146 358
rect 1808 190 1842 324
rect 2080 306 2146 324
rect 2180 304 2214 410
rect 2485 360 2519 478
rect 2605 377 2639 504
rect 2886 476 2920 596
rect 2692 411 2920 476
rect 2809 384 2920 411
rect 1876 224 1938 290
rect 1972 272 2038 290
rect 2180 272 2348 304
rect 1972 238 2348 272
rect 2390 260 2451 360
rect 2485 294 2571 360
rect 2605 343 2775 377
rect 2613 260 2679 309
rect 1898 204 1938 224
rect 1808 124 1864 190
rect 1898 170 2146 204
rect 1898 85 1938 170
rect 1560 51 1938 85
rect 2013 17 2078 136
rect 2112 85 2146 170
rect 2180 119 2214 238
rect 2390 226 2679 260
rect 2741 306 2775 343
rect 2741 240 2852 306
rect 2390 204 2424 226
rect 2248 170 2424 204
rect 2741 188 2775 240
rect 2886 206 2920 384
rect 2248 85 2282 170
rect 2458 154 2775 188
rect 2112 51 2282 85
rect 2316 17 2366 136
rect 2458 70 2524 154
rect 2638 17 2807 120
rect 2841 85 2920 206
rect 3088 364 3138 649
rect 3037 264 3179 330
rect 3037 85 3071 264
rect 2841 51 3071 85
rect 3105 17 3139 230
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3264 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 3199 649 3233 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
<< metal1 >>
rect 0 683 3264 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3264 683
rect 0 617 3264 649
rect 0 17 3264 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3264 17
rect 0 -49 3264 -17
<< obsm1 >>
rect 595 421 653 430
rect 2803 421 2861 430
rect 595 393 2861 421
rect 595 384 653 393
rect 2803 384 2861 393
<< labels >>
rlabel locali s 91 212 167 356 6 D
port 1 nsew signal input
rlabel locali s 313 290 417 356 6 DE
port 2 nsew signal input
rlabel locali s 2969 364 3048 596 6 Q
port 3 nsew signal output
rlabel locali s 2969 124 3003 364 6 Q
port 3 nsew signal output
rlabel locali s 3213 230 3247 364 6 Q_N
port 4 nsew signal output
rlabel locali s 3175 74 3247 230 6 Q_N
port 4 nsew signal output
rlabel locali s 3172 364 3247 596 6 Q_N
port 4 nsew signal output
rlabel locali s 1015 236 1127 302 6 SCD
port 5 nsew signal input
rlabel locali s 895 290 973 356 6 SCE
port 6 nsew signal input
rlabel locali s 1315 236 1415 310 6 CLK
port 7 nsew clock input
rlabel metal1 s 0 -49 3264 49 8 VGND
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 617 3264 715 6 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 3264 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 476332
string GDS_START 453500
<< end >>
