magic
tech sky130A
magscale 1 2
timestamp 1599588209
<< nwell >>
rect -38 332 1862 704
<< pwell >>
rect 0 0 1824 49
<< scpmos >>
rect 174 368 204 536
rect 264 368 294 536
rect 371 368 401 592
rect 543 368 573 592
rect 835 368 865 592
rect 925 368 955 592
rect 1174 368 1204 592
rect 1340 368 1370 592
rect 1604 368 1634 592
rect 1698 368 1728 592
<< nmoslvt >>
rect 84 74 114 222
rect 282 74 312 222
rect 368 74 398 222
rect 454 74 484 222
rect 540 74 570 222
rect 626 74 656 222
rect 712 74 742 222
rect 798 74 828 222
rect 884 74 914 222
rect 1082 74 1112 222
rect 1168 74 1198 222
rect 1254 74 1284 222
rect 1343 74 1373 222
rect 1429 74 1459 222
rect 1515 74 1545 222
rect 1601 74 1631 222
rect 1710 74 1740 222
<< ndiff >>
rect 27 207 84 222
rect 27 173 39 207
rect 73 173 84 207
rect 27 158 84 173
rect 34 74 84 158
rect 114 132 164 222
rect 232 138 282 222
rect 114 120 171 132
rect 114 86 125 120
rect 159 86 171 120
rect 114 74 171 86
rect 225 123 282 138
rect 225 89 237 123
rect 271 89 282 123
rect 225 74 282 89
rect 312 210 368 222
rect 312 176 323 210
rect 357 176 368 210
rect 312 74 368 176
rect 398 123 454 222
rect 398 89 409 123
rect 443 89 454 123
rect 398 74 454 89
rect 484 189 540 222
rect 484 155 495 189
rect 529 155 540 189
rect 484 74 540 155
rect 570 144 626 222
rect 570 110 581 144
rect 615 110 626 144
rect 570 74 626 110
rect 656 116 712 222
rect 656 82 667 116
rect 701 82 712 116
rect 656 74 712 82
rect 742 184 798 222
rect 742 150 753 184
rect 787 150 798 184
rect 742 74 798 150
rect 828 116 884 222
rect 828 82 839 116
rect 873 82 884 116
rect 828 74 884 82
rect 914 196 964 222
rect 1025 207 1082 222
rect 914 184 971 196
rect 914 150 925 184
rect 959 150 971 184
rect 1025 173 1037 207
rect 1071 173 1082 207
rect 1025 158 1082 173
rect 914 138 971 150
rect 914 74 964 138
rect 1032 74 1082 158
rect 1112 120 1168 222
rect 1112 86 1123 120
rect 1157 86 1168 120
rect 1112 74 1168 86
rect 1198 207 1254 222
rect 1198 173 1209 207
rect 1243 173 1254 207
rect 1198 74 1254 173
rect 1284 136 1343 222
rect 1284 102 1295 136
rect 1329 102 1343 136
rect 1284 74 1343 102
rect 1373 207 1429 222
rect 1373 173 1384 207
rect 1418 173 1429 207
rect 1373 120 1429 173
rect 1373 86 1384 120
rect 1418 86 1429 120
rect 1373 74 1429 86
rect 1459 140 1515 222
rect 1459 106 1470 140
rect 1504 106 1515 140
rect 1459 74 1515 106
rect 1545 207 1601 222
rect 1545 173 1556 207
rect 1590 173 1601 207
rect 1545 120 1601 173
rect 1545 86 1556 120
rect 1590 86 1601 120
rect 1545 74 1601 86
rect 1631 140 1710 222
rect 1631 106 1646 140
rect 1680 106 1710 140
rect 1631 74 1710 106
rect 1740 210 1797 222
rect 1740 176 1751 210
rect 1785 176 1797 210
rect 1740 120 1797 176
rect 1740 86 1751 120
rect 1785 86 1797 120
rect 1740 74 1797 86
<< pdiff >>
rect 312 580 371 592
rect 312 546 324 580
rect 358 546 371 580
rect 312 536 371 546
rect 105 524 174 536
rect 105 490 117 524
rect 151 490 174 524
rect 105 440 174 490
rect 105 406 117 440
rect 151 406 174 440
rect 105 368 174 406
rect 204 524 264 536
rect 204 490 217 524
rect 251 490 264 524
rect 204 414 264 490
rect 204 380 217 414
rect 251 380 264 414
rect 204 368 264 380
rect 294 500 371 536
rect 294 466 324 500
rect 358 466 371 500
rect 294 420 371 466
rect 294 386 324 420
rect 358 386 371 420
rect 294 368 371 386
rect 401 580 543 592
rect 401 546 414 580
rect 448 546 496 580
rect 530 546 543 580
rect 401 500 543 546
rect 401 466 414 500
rect 448 466 496 500
rect 530 466 543 500
rect 401 420 543 466
rect 401 386 414 420
rect 448 386 496 420
rect 530 386 543 420
rect 401 368 543 386
rect 573 580 835 592
rect 573 546 586 580
rect 620 546 685 580
rect 719 546 788 580
rect 822 546 835 580
rect 573 492 835 546
rect 573 458 586 492
rect 620 458 685 492
rect 719 458 788 492
rect 822 458 835 492
rect 573 368 835 458
rect 865 580 925 592
rect 865 546 878 580
rect 912 546 925 580
rect 865 497 925 546
rect 865 463 878 497
rect 912 463 925 497
rect 865 414 925 463
rect 865 380 878 414
rect 912 380 925 414
rect 865 368 925 380
rect 955 580 1174 592
rect 955 546 968 580
rect 1002 546 1052 580
rect 1086 546 1127 580
rect 1161 546 1174 580
rect 955 492 1174 546
rect 955 458 968 492
rect 1002 458 1052 492
rect 1086 458 1127 492
rect 1161 458 1174 492
rect 955 368 1174 458
rect 1204 580 1340 592
rect 1204 546 1217 580
rect 1251 546 1293 580
rect 1327 546 1340 580
rect 1204 503 1340 546
rect 1204 469 1217 503
rect 1251 469 1293 503
rect 1327 469 1340 503
rect 1204 424 1340 469
rect 1204 390 1217 424
rect 1251 390 1293 424
rect 1327 390 1340 424
rect 1204 368 1340 390
rect 1370 580 1604 592
rect 1370 546 1383 580
rect 1417 546 1467 580
rect 1501 546 1557 580
rect 1591 546 1604 580
rect 1370 492 1604 546
rect 1370 458 1383 492
rect 1417 458 1467 492
rect 1501 458 1557 492
rect 1591 458 1604 492
rect 1370 368 1604 458
rect 1634 580 1698 592
rect 1634 546 1651 580
rect 1685 546 1698 580
rect 1634 503 1698 546
rect 1634 469 1651 503
rect 1685 469 1698 503
rect 1634 424 1698 469
rect 1634 390 1651 424
rect 1685 390 1698 424
rect 1634 368 1698 390
rect 1728 580 1797 592
rect 1728 546 1741 580
rect 1775 546 1797 580
rect 1728 510 1797 546
rect 1728 476 1741 510
rect 1775 476 1797 510
rect 1728 440 1797 476
rect 1728 406 1741 440
rect 1775 406 1797 440
rect 1728 368 1797 406
<< ndiffc >>
rect 39 173 73 207
rect 125 86 159 120
rect 237 89 271 123
rect 323 176 357 210
rect 409 89 443 123
rect 495 155 529 189
rect 581 110 615 144
rect 667 82 701 116
rect 753 150 787 184
rect 839 82 873 116
rect 925 150 959 184
rect 1037 173 1071 207
rect 1123 86 1157 120
rect 1209 173 1243 207
rect 1295 102 1329 136
rect 1384 173 1418 207
rect 1384 86 1418 120
rect 1470 106 1504 140
rect 1556 173 1590 207
rect 1556 86 1590 120
rect 1646 106 1680 140
rect 1751 176 1785 210
rect 1751 86 1785 120
<< pdiffc >>
rect 324 546 358 580
rect 117 490 151 524
rect 117 406 151 440
rect 217 490 251 524
rect 217 380 251 414
rect 324 466 358 500
rect 324 386 358 420
rect 414 546 448 580
rect 496 546 530 580
rect 414 466 448 500
rect 496 466 530 500
rect 414 386 448 420
rect 496 386 530 420
rect 586 546 620 580
rect 685 546 719 580
rect 788 546 822 580
rect 586 458 620 492
rect 685 458 719 492
rect 788 458 822 492
rect 878 546 912 580
rect 878 463 912 497
rect 878 380 912 414
rect 968 546 1002 580
rect 1052 546 1086 580
rect 1127 546 1161 580
rect 968 458 1002 492
rect 1052 458 1086 492
rect 1127 458 1161 492
rect 1217 546 1251 580
rect 1293 546 1327 580
rect 1217 469 1251 503
rect 1293 469 1327 503
rect 1217 390 1251 424
rect 1293 390 1327 424
rect 1383 546 1417 580
rect 1467 546 1501 580
rect 1557 546 1591 580
rect 1383 458 1417 492
rect 1467 458 1501 492
rect 1557 458 1591 492
rect 1651 546 1685 580
rect 1651 469 1685 503
rect 1651 390 1685 424
rect 1741 546 1775 580
rect 1741 476 1775 510
rect 1741 406 1775 440
<< poly >>
rect 371 592 401 618
rect 543 592 573 618
rect 835 592 865 618
rect 925 592 955 618
rect 1174 592 1204 618
rect 1340 592 1370 618
rect 1604 592 1634 618
rect 1698 592 1728 618
rect 174 536 204 562
rect 264 536 294 562
rect 174 353 204 368
rect 264 353 294 368
rect 371 353 401 368
rect 543 353 573 368
rect 835 353 865 368
rect 925 353 955 368
rect 1174 353 1204 368
rect 1340 353 1370 368
rect 1604 353 1634 368
rect 1698 353 1728 368
rect 171 345 207 353
rect 261 345 297 353
rect 33 315 297 345
rect 368 336 404 353
rect 540 336 573 353
rect 832 336 868 353
rect 368 320 570 336
rect 33 310 207 315
rect 33 276 49 310
rect 83 276 117 310
rect 151 276 207 310
rect 33 260 207 276
rect 368 286 384 320
rect 418 286 452 320
rect 486 286 520 320
rect 554 286 570 320
rect 368 267 570 286
rect 84 222 114 260
rect 282 237 570 267
rect 282 222 312 237
rect 368 222 398 237
rect 454 222 484 237
rect 540 222 570 237
rect 626 331 868 336
rect 922 331 958 353
rect 1171 336 1207 353
rect 1337 336 1373 353
rect 626 320 958 331
rect 626 286 642 320
rect 676 286 710 320
rect 744 286 778 320
rect 812 286 958 320
rect 626 270 958 286
rect 1082 320 1373 336
rect 1082 286 1119 320
rect 1153 286 1187 320
rect 1221 286 1255 320
rect 1289 286 1323 320
rect 1357 286 1373 320
rect 1601 326 1637 353
rect 1695 326 1731 353
rect 1601 310 1803 326
rect 1601 290 1617 310
rect 1082 270 1373 286
rect 626 222 656 270
rect 712 222 742 270
rect 798 222 828 270
rect 884 222 914 270
rect 1082 222 1112 270
rect 1168 222 1198 270
rect 1254 222 1284 270
rect 1343 222 1373 270
rect 1429 276 1617 290
rect 1651 276 1685 310
rect 1719 276 1753 310
rect 1787 276 1803 310
rect 1429 260 1803 276
rect 1429 222 1459 260
rect 1515 222 1545 260
rect 1601 222 1631 260
rect 1710 222 1740 260
rect 84 48 114 74
rect 282 48 312 74
rect 368 48 398 74
rect 454 48 484 74
rect 540 48 570 74
rect 626 48 656 74
rect 712 48 742 74
rect 798 48 828 74
rect 884 48 914 74
rect 1082 48 1112 74
rect 1168 48 1198 74
rect 1254 48 1284 74
rect 1343 48 1373 74
rect 1429 48 1459 74
rect 1515 48 1545 74
rect 1601 48 1631 74
rect 1710 48 1740 74
<< polycont >>
rect 49 276 83 310
rect 117 276 151 310
rect 384 286 418 320
rect 452 286 486 320
rect 520 286 554 320
rect 642 286 676 320
rect 710 286 744 320
rect 778 286 812 320
rect 1119 286 1153 320
rect 1187 286 1221 320
rect 1255 286 1289 320
rect 1323 286 1357 320
rect 1617 276 1651 310
rect 1685 276 1719 310
rect 1753 276 1787 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 101 524 167 649
rect 308 580 374 649
rect 308 546 324 580
rect 358 546 374 580
rect 101 490 117 524
rect 151 490 167 524
rect 101 440 167 490
rect 101 406 117 440
rect 151 406 167 440
rect 101 390 167 406
rect 201 524 267 540
rect 201 490 217 524
rect 251 490 267 524
rect 201 414 267 490
rect 201 380 217 414
rect 251 380 267 414
rect 25 310 167 356
rect 25 276 49 310
rect 83 276 117 310
rect 151 276 167 310
rect 25 260 167 276
rect 201 336 267 380
rect 308 500 374 546
rect 308 466 324 500
rect 358 466 374 500
rect 308 420 374 466
rect 308 386 324 420
rect 358 386 374 420
rect 308 370 374 386
rect 410 580 534 596
rect 410 546 414 580
rect 448 546 496 580
rect 530 546 534 580
rect 410 500 534 546
rect 410 466 414 500
rect 448 466 496 500
rect 530 466 534 500
rect 410 424 534 466
rect 570 580 838 649
rect 570 546 586 580
rect 620 546 685 580
rect 719 546 788 580
rect 822 546 838 580
rect 570 492 838 546
rect 570 458 586 492
rect 620 458 685 492
rect 719 458 788 492
rect 822 458 838 492
rect 874 580 918 596
rect 874 546 878 580
rect 912 546 918 580
rect 874 497 918 546
rect 874 463 878 497
rect 912 463 918 497
rect 874 424 918 463
rect 952 580 1177 649
rect 952 546 968 580
rect 1002 546 1052 580
rect 1086 546 1127 580
rect 1161 546 1177 580
rect 952 492 1177 546
rect 952 458 968 492
rect 1002 458 1052 492
rect 1086 458 1127 492
rect 1161 458 1177 492
rect 1213 580 1332 596
rect 1213 546 1217 580
rect 1251 546 1293 580
rect 1327 546 1332 580
rect 1213 503 1332 546
rect 1213 469 1217 503
rect 1251 469 1293 503
rect 1327 469 1332 503
rect 1213 424 1332 469
rect 1367 580 1607 649
rect 1367 546 1383 580
rect 1417 546 1467 580
rect 1501 546 1557 580
rect 1591 546 1607 580
rect 1367 492 1607 546
rect 1367 458 1383 492
rect 1417 458 1467 492
rect 1501 458 1557 492
rect 1591 458 1607 492
rect 1643 580 1701 596
rect 1643 546 1651 580
rect 1685 546 1701 580
rect 1643 503 1701 546
rect 1643 469 1651 503
rect 1685 469 1701 503
rect 1643 424 1701 469
rect 410 420 1217 424
rect 410 386 414 420
rect 448 386 496 420
rect 530 414 1217 420
rect 530 390 878 414
rect 530 386 536 390
rect 410 370 536 386
rect 862 380 878 390
rect 912 390 1217 414
rect 1251 390 1293 424
rect 1327 390 1651 424
rect 1685 390 1701 424
rect 1735 580 1791 649
rect 1735 546 1741 580
rect 1775 546 1791 580
rect 1735 510 1791 546
rect 1735 476 1741 510
rect 1775 476 1791 510
rect 1735 440 1791 476
rect 1735 406 1741 440
rect 1775 406 1791 440
rect 1735 390 1791 406
rect 912 380 935 390
rect 862 364 935 380
rect 201 320 570 336
rect 201 286 384 320
rect 418 286 452 320
rect 486 286 520 320
rect 554 286 570 320
rect 626 320 828 356
rect 626 286 642 320
rect 676 286 710 320
rect 744 286 778 320
rect 812 286 828 320
rect 201 226 267 286
rect 889 252 935 364
rect 985 320 1511 356
rect 985 286 1119 320
rect 1153 286 1187 320
rect 1221 286 1255 320
rect 1289 286 1323 320
rect 1357 286 1511 320
rect 985 270 1511 286
rect 1561 310 1803 356
rect 1561 276 1617 310
rect 1651 276 1685 310
rect 1719 276 1753 310
rect 1787 276 1803 310
rect 1561 260 1803 276
rect 479 226 935 252
rect 1193 226 1434 236
rect 23 207 267 226
rect 23 173 39 207
rect 73 192 267 207
rect 307 218 935 226
rect 307 210 545 218
rect 73 173 89 192
rect 307 176 323 210
rect 357 189 545 210
rect 357 176 495 189
rect 23 154 89 173
rect 479 155 495 176
rect 529 155 545 189
rect 1021 210 1801 226
rect 1021 207 1751 210
rect 221 123 287 142
rect 109 86 125 120
rect 159 86 175 120
rect 109 17 175 86
rect 221 89 237 123
rect 271 89 287 123
rect 221 85 287 89
rect 393 123 443 142
rect 393 89 409 123
rect 479 119 545 155
rect 581 150 753 184
rect 787 150 925 184
rect 959 150 975 184
rect 1021 173 1037 207
rect 1071 192 1209 207
rect 1071 173 1087 192
rect 1021 154 1087 173
rect 1193 173 1209 192
rect 1243 202 1384 207
rect 1193 154 1243 173
rect 1418 192 1556 207
rect 1418 173 1420 192
rect 581 144 615 150
rect 393 85 443 89
rect 1121 120 1159 142
rect 1279 136 1345 168
rect 1279 120 1295 136
rect 1107 116 1123 120
rect 581 85 615 110
rect 221 51 615 85
rect 651 82 667 116
rect 701 82 839 116
rect 873 86 1123 116
rect 1157 102 1295 120
rect 1329 102 1345 136
rect 1157 86 1345 102
rect 873 82 1345 86
rect 651 66 1345 82
rect 1384 120 1420 173
rect 1554 173 1556 192
rect 1590 192 1751 207
rect 1590 173 1592 192
rect 1418 86 1420 120
rect 1384 70 1420 86
rect 1454 140 1520 156
rect 1454 106 1470 140
rect 1504 106 1520 140
rect 1454 17 1520 106
rect 1554 120 1592 173
rect 1735 176 1751 192
rect 1785 176 1801 210
rect 1554 86 1556 120
rect 1590 86 1592 120
rect 1554 70 1592 86
rect 1626 140 1701 156
rect 1626 106 1646 140
rect 1680 106 1701 140
rect 1626 17 1701 106
rect 1735 120 1801 176
rect 1735 86 1751 120
rect 1785 86 1801 120
rect 1735 70 1801 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
<< metal1 >>
rect 0 683 1824 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 0 617 1824 649
rect 0 17 1824 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
rect 0 -49 1824 -17
<< labels >>
rlabel comment s 0 0 0 0 4 nand4b_4
flabel pwell s 0 0 1824 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nwell s 0 617 1824 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 1824 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 1824 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 1087 316 1121 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 1183 316 1217 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 1279 316 1313 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 1375 316 1409 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 1471 316 1505 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 895 242 929 276 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 1567 316 1601 350 0 FreeSans 340 0 0 0 D
port 4 nsew
flabel corelocali s 1663 316 1697 350 0 FreeSans 340 0 0 0 D
port 4 nsew
flabel corelocali s 1759 316 1793 350 0 FreeSans 340 0 0 0 D
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 1824 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1476954
string GDS_START 1462946
<< end >>
