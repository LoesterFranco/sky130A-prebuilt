magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 20 199 81 323
rect 115 171 179 423
rect 213 257 257 323
rect 937 257 983 331
rect 213 207 387 257
rect 562 207 714 257
rect 778 207 983 257
rect 115 131 679 171
rect 115 51 177 131
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 29 457 483 491
rect 29 357 81 457
rect 235 451 483 457
rect 235 357 273 451
rect 307 331 383 415
rect 427 367 483 451
rect 527 367 573 527
rect 619 331 673 493
rect 719 367 765 527
rect 811 331 865 493
rect 911 367 957 527
rect 307 291 865 331
rect 29 17 79 163
rect 725 127 967 171
rect 725 95 759 127
rect 211 17 287 95
rect 403 17 479 95
rect 517 53 759 95
rect 795 17 871 91
rect 917 53 967 127
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
rlabel locali s 562 207 714 257 6 A1
port 1 nsew signal input
rlabel locali s 937 257 983 331 6 A2
port 2 nsew signal input
rlabel locali s 778 207 983 257 6 A2
port 2 nsew signal input
rlabel locali s 213 257 257 323 6 B1
port 3 nsew signal input
rlabel locali s 213 207 387 257 6 B1
port 3 nsew signal input
rlabel locali s 20 199 81 323 6 C1
port 4 nsew signal input
rlabel locali s 115 171 179 423 6 Y
port 5 nsew signal output
rlabel locali s 115 131 679 171 6 Y
port 5 nsew signal output
rlabel locali s 115 51 177 131 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -48 1012 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 1012 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1012 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1115742
string GDS_START 1106622
<< end >>
