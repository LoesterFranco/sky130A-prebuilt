magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 1574 704
<< pwell >>
rect 0 0 1536 49
<< scnmos >>
rect 140 82 170 210
rect 226 82 256 210
rect 312 82 342 210
rect 398 82 428 210
rect 493 82 523 230
rect 579 82 609 230
rect 674 85 704 233
rect 760 85 790 233
rect 858 105 888 233
rect 944 105 974 233
rect 1146 117 1176 245
rect 1232 117 1262 245
rect 1330 117 1360 245
rect 1416 117 1446 245
<< pmoshvt >>
rect 124 392 154 592
rect 214 392 244 592
rect 304 392 334 592
rect 394 392 424 592
rect 588 368 618 592
rect 678 368 708 592
rect 768 368 798 592
rect 858 368 888 592
rect 961 392 991 592
rect 1051 392 1081 592
rect 1141 392 1171 592
rect 1231 392 1261 592
rect 1327 392 1357 592
rect 1417 392 1447 592
<< ndiff >>
rect 624 230 674 233
rect 443 210 493 230
rect 87 128 140 210
rect 87 94 95 128
rect 129 94 140 128
rect 87 82 140 94
rect 170 198 226 210
rect 170 164 181 198
rect 215 164 226 198
rect 170 128 226 164
rect 170 94 181 128
rect 215 94 226 128
rect 170 82 226 94
rect 256 192 312 210
rect 256 158 267 192
rect 301 158 312 192
rect 256 124 312 158
rect 256 90 267 124
rect 301 90 312 124
rect 256 82 312 90
rect 342 198 398 210
rect 342 164 353 198
rect 387 164 398 198
rect 342 128 398 164
rect 342 94 353 128
rect 387 94 398 128
rect 342 82 398 94
rect 428 176 493 210
rect 428 142 439 176
rect 473 142 493 176
rect 428 82 493 142
rect 523 214 579 230
rect 523 180 534 214
rect 568 180 579 214
rect 523 128 579 180
rect 523 94 534 128
rect 568 94 579 128
rect 523 82 579 94
rect 609 138 674 230
rect 609 104 624 138
rect 658 104 674 138
rect 609 85 674 104
rect 704 214 760 233
rect 704 180 715 214
rect 749 180 760 214
rect 704 131 760 180
rect 704 97 715 131
rect 749 97 760 131
rect 704 85 760 97
rect 790 214 858 233
rect 790 180 801 214
rect 835 180 858 214
rect 790 131 858 180
rect 790 97 801 131
rect 835 105 858 131
rect 888 152 944 233
rect 888 118 899 152
rect 933 118 944 152
rect 888 105 944 118
rect 974 221 1027 233
rect 974 187 985 221
rect 1019 187 1027 221
rect 974 105 1027 187
rect 1081 117 1146 245
rect 1176 237 1232 245
rect 1176 203 1187 237
rect 1221 203 1232 237
rect 1176 117 1232 203
rect 1262 232 1330 245
rect 1262 198 1273 232
rect 1307 198 1330 232
rect 1262 117 1330 198
rect 1360 163 1416 245
rect 1360 129 1371 163
rect 1405 129 1416 163
rect 1360 117 1416 129
rect 1446 233 1499 245
rect 1446 199 1457 233
rect 1491 199 1499 233
rect 1446 163 1499 199
rect 1446 129 1457 163
rect 1491 129 1499 163
rect 1446 117 1499 129
rect 835 97 843 105
rect 790 85 843 97
rect 609 82 659 85
rect 1081 85 1131 117
rect 1081 51 1089 85
rect 1123 51 1131 85
rect 1081 39 1131 51
<< pdiff >>
rect 69 577 124 592
rect 69 543 77 577
rect 111 543 124 577
rect 69 392 124 543
rect 154 438 214 592
rect 154 404 167 438
rect 201 404 214 438
rect 154 392 214 404
rect 244 577 304 592
rect 244 543 257 577
rect 291 543 304 577
rect 244 392 304 543
rect 334 521 394 592
rect 334 487 347 521
rect 381 487 394 521
rect 334 392 394 487
rect 424 573 479 592
rect 424 539 437 573
rect 471 539 479 573
rect 424 392 479 539
rect 533 573 588 592
rect 533 539 541 573
rect 575 539 588 573
rect 533 368 588 539
rect 618 414 678 592
rect 618 380 631 414
rect 665 380 678 414
rect 618 368 678 380
rect 708 573 768 592
rect 708 539 721 573
rect 755 539 768 573
rect 708 368 768 539
rect 798 414 858 592
rect 798 380 811 414
rect 845 380 858 414
rect 798 368 858 380
rect 888 573 961 592
rect 888 539 901 573
rect 935 539 961 573
rect 888 392 961 539
rect 991 580 1051 592
rect 991 546 1004 580
rect 1038 546 1051 580
rect 991 508 1051 546
rect 991 474 1004 508
rect 1038 474 1051 508
rect 991 392 1051 474
rect 1081 578 1141 592
rect 1081 544 1094 578
rect 1128 544 1141 578
rect 1081 392 1141 544
rect 1171 580 1231 592
rect 1171 546 1184 580
rect 1218 546 1231 580
rect 1171 510 1231 546
rect 1171 476 1184 510
rect 1218 476 1231 510
rect 1171 440 1231 476
rect 1171 406 1184 440
rect 1218 406 1231 440
rect 1171 392 1231 406
rect 1261 580 1327 592
rect 1261 546 1277 580
rect 1311 546 1327 580
rect 1261 508 1327 546
rect 1261 474 1277 508
rect 1311 474 1327 508
rect 1261 392 1327 474
rect 1357 580 1417 592
rect 1357 546 1370 580
rect 1404 546 1417 580
rect 1357 510 1417 546
rect 1357 476 1370 510
rect 1404 476 1417 510
rect 1357 440 1417 476
rect 1357 406 1370 440
rect 1404 406 1417 440
rect 1357 392 1417 406
rect 1447 580 1502 592
rect 1447 546 1460 580
rect 1494 546 1502 580
rect 1447 510 1502 546
rect 1447 476 1460 510
rect 1494 476 1502 510
rect 1447 440 1502 476
rect 1447 406 1460 440
rect 1494 406 1502 440
rect 1447 392 1502 406
rect 888 368 943 392
<< ndiffc >>
rect 95 94 129 128
rect 181 164 215 198
rect 181 94 215 128
rect 267 158 301 192
rect 267 90 301 124
rect 353 164 387 198
rect 353 94 387 128
rect 439 142 473 176
rect 534 180 568 214
rect 534 94 568 128
rect 624 104 658 138
rect 715 180 749 214
rect 715 97 749 131
rect 801 180 835 214
rect 801 97 835 131
rect 899 118 933 152
rect 985 187 1019 221
rect 1187 203 1221 237
rect 1273 198 1307 232
rect 1371 129 1405 163
rect 1457 199 1491 233
rect 1457 129 1491 163
rect 1089 51 1123 85
<< pdiffc >>
rect 77 543 111 577
rect 167 404 201 438
rect 257 543 291 577
rect 347 487 381 521
rect 437 539 471 573
rect 541 539 575 573
rect 631 380 665 414
rect 721 539 755 573
rect 811 380 845 414
rect 901 539 935 573
rect 1004 546 1038 580
rect 1004 474 1038 508
rect 1094 544 1128 578
rect 1184 546 1218 580
rect 1184 476 1218 510
rect 1184 406 1218 440
rect 1277 546 1311 580
rect 1277 474 1311 508
rect 1370 546 1404 580
rect 1370 476 1404 510
rect 1370 406 1404 440
rect 1460 546 1494 580
rect 1460 476 1494 510
rect 1460 406 1494 440
<< poly >>
rect 124 592 154 618
rect 214 592 244 618
rect 304 592 334 618
rect 394 592 424 618
rect 588 592 618 618
rect 678 592 708 618
rect 768 592 798 618
rect 858 592 888 618
rect 961 592 991 618
rect 1051 592 1081 618
rect 1141 592 1171 618
rect 1231 592 1261 618
rect 1327 592 1357 618
rect 1417 592 1447 618
rect 124 377 154 392
rect 214 377 244 392
rect 304 377 334 392
rect 394 377 424 392
rect 121 360 157 377
rect 211 360 247 377
rect 99 344 247 360
rect 99 310 115 344
rect 149 318 247 344
rect 301 360 337 377
rect 391 360 427 377
rect 961 377 991 392
rect 1051 377 1081 392
rect 1141 377 1171 392
rect 1231 377 1261 392
rect 1327 377 1357 392
rect 1417 377 1447 392
rect 301 344 427 360
rect 588 353 618 368
rect 678 353 708 368
rect 768 353 798 368
rect 858 353 888 368
rect 585 350 621 353
rect 675 350 711 353
rect 765 350 801 353
rect 855 350 891 353
rect 149 310 256 318
rect 99 288 256 310
rect 301 310 323 344
rect 357 324 427 344
rect 357 310 428 324
rect 301 294 428 310
rect 140 210 170 288
rect 226 210 256 288
rect 312 210 342 294
rect 398 210 428 294
rect 493 320 891 350
rect 958 350 994 377
rect 1048 350 1084 377
rect 958 334 1084 350
rect 493 314 801 320
rect 958 314 1009 334
rect 493 280 527 314
rect 561 280 595 314
rect 629 280 663 314
rect 697 280 731 314
rect 765 280 801 314
rect 493 264 801 280
rect 944 300 1009 314
rect 1043 300 1084 334
rect 944 284 1084 300
rect 1138 356 1174 377
rect 1228 356 1264 377
rect 1324 356 1360 377
rect 1414 356 1450 377
rect 1138 340 1282 356
rect 1138 306 1232 340
rect 1266 306 1282 340
rect 1324 340 1515 356
rect 1324 320 1465 340
rect 1138 290 1282 306
rect 1330 306 1465 320
rect 1499 306 1515 340
rect 1330 290 1515 306
rect 944 278 974 284
rect 493 230 523 264
rect 579 230 609 264
rect 674 233 704 264
rect 760 233 790 264
rect 858 248 974 278
rect 858 233 888 248
rect 944 233 974 248
rect 1146 245 1176 290
rect 1232 245 1262 290
rect 1330 245 1360 290
rect 1416 245 1446 290
rect 140 56 170 82
rect 226 56 256 82
rect 312 56 342 82
rect 398 56 428 82
rect 493 56 523 82
rect 579 56 609 82
rect 674 59 704 85
rect 760 59 790 85
rect 858 79 888 105
rect 944 79 974 105
rect 1146 91 1176 117
rect 1232 91 1262 117
rect 1330 91 1360 117
rect 1416 91 1446 117
<< polycont >>
rect 115 310 149 344
rect 323 310 357 344
rect 527 280 561 314
rect 595 280 629 314
rect 663 280 697 314
rect 731 280 765 314
rect 1009 300 1043 334
rect 1232 306 1266 340
rect 1465 306 1499 340
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 241 596 487 615
rect 61 581 487 596
rect 61 577 307 581
rect 61 543 77 577
rect 111 543 257 577
rect 291 543 307 577
rect 421 573 487 581
rect 61 540 307 543
rect 347 521 381 547
rect 421 539 437 573
rect 471 539 487 573
rect 421 532 487 539
rect 525 573 591 649
rect 525 539 541 573
rect 575 539 591 573
rect 525 532 591 539
rect 705 573 771 649
rect 705 539 721 573
rect 755 539 771 573
rect 705 532 771 539
rect 885 573 951 649
rect 885 539 901 573
rect 935 539 951 573
rect 885 532 951 539
rect 988 580 1054 596
rect 988 546 1004 580
rect 1038 546 1054 580
rect 25 472 301 506
rect 25 208 59 472
rect 151 404 167 438
rect 201 404 233 438
rect 99 344 165 360
rect 99 310 115 344
rect 149 310 165 344
rect 99 294 165 310
rect 199 260 233 404
rect 267 428 301 472
rect 988 508 1054 546
rect 1094 578 1144 649
rect 1128 544 1144 578
rect 1094 526 1144 544
rect 1184 580 1218 596
rect 988 498 1004 508
rect 381 487 1004 498
rect 347 474 1004 487
rect 1038 492 1054 508
rect 1184 510 1218 546
rect 1038 476 1184 492
rect 1038 474 1218 476
rect 347 464 1218 474
rect 347 462 381 464
rect 988 458 1218 464
rect 1258 580 1330 649
rect 1258 546 1277 580
rect 1311 546 1330 580
rect 1258 508 1330 546
rect 1258 474 1277 508
rect 1311 474 1330 508
rect 1258 458 1330 474
rect 1370 580 1404 596
rect 1370 510 1404 546
rect 1184 440 1218 458
rect 505 428 861 430
rect 267 414 861 428
rect 267 394 631 414
rect 505 380 631 394
rect 665 380 811 414
rect 845 380 861 414
rect 505 364 861 380
rect 895 390 1143 424
rect 1370 440 1404 476
rect 1218 406 1370 424
rect 1184 390 1404 406
rect 1444 580 1510 649
rect 1444 546 1460 580
rect 1494 546 1510 580
rect 1444 510 1510 546
rect 1444 476 1460 510
rect 1494 476 1510 510
rect 1444 440 1510 476
rect 1444 406 1460 440
rect 1494 406 1510 440
rect 1444 390 1510 406
rect 307 344 373 360
rect 307 310 323 344
rect 357 310 373 344
rect 895 330 929 390
rect 307 294 373 310
rect 411 314 929 330
rect 411 280 527 314
rect 561 280 595 314
rect 629 280 663 314
rect 697 280 731 314
rect 765 296 929 314
rect 985 334 1059 356
rect 985 300 1009 334
rect 1043 300 1059 334
rect 765 280 781 296
rect 985 284 1059 300
rect 411 264 781 280
rect 411 260 465 264
rect 181 226 465 260
rect 1109 253 1143 390
rect 1177 340 1415 356
rect 1177 306 1232 340
rect 1266 306 1415 340
rect 1177 290 1415 306
rect 1449 340 1515 356
rect 1449 306 1465 340
rect 1499 306 1515 340
rect 1449 290 1515 306
rect 1109 237 1221 253
rect 835 230 1035 237
rect 25 202 71 208
rect 25 168 31 202
rect 65 168 71 202
rect 25 162 71 168
rect 181 198 217 226
rect 215 164 217 198
rect 351 198 387 226
rect 181 128 217 164
rect 79 94 95 128
rect 129 94 145 128
rect 79 17 145 94
rect 215 94 217 128
rect 181 78 217 94
rect 251 158 267 192
rect 301 158 317 192
rect 251 124 317 158
rect 251 90 267 124
rect 301 90 317 124
rect 251 17 317 90
rect 351 164 353 198
rect 507 214 749 230
rect 507 202 534 214
rect 351 128 387 164
rect 351 94 353 128
rect 351 78 387 94
rect 423 176 473 192
rect 423 142 439 176
rect 423 17 473 142
rect 507 168 511 202
rect 568 196 715 214
rect 568 180 584 196
rect 545 168 584 180
rect 507 128 584 168
rect 699 180 715 196
rect 507 94 534 128
rect 568 94 584 128
rect 507 78 584 94
rect 620 138 663 162
rect 620 104 624 138
rect 658 104 663 138
rect 620 17 663 104
rect 699 131 749 180
rect 699 97 715 131
rect 699 81 749 97
rect 785 221 1035 230
rect 785 214 985 221
rect 785 180 801 214
rect 835 187 985 214
rect 1019 187 1035 221
rect 1109 203 1187 237
rect 1109 187 1221 203
rect 1257 233 1507 249
rect 1257 232 1457 233
rect 1257 198 1273 232
rect 1307 199 1457 232
rect 1491 199 1507 233
rect 1307 198 1507 199
rect 1257 197 1507 198
rect 785 131 835 180
rect 1457 163 1507 197
rect 1355 153 1371 163
rect 785 97 801 131
rect 883 152 1371 153
rect 883 118 899 152
rect 933 129 1371 152
rect 1405 129 1421 163
rect 933 119 1421 129
rect 1491 129 1507 163
rect 933 118 949 119
rect 883 101 949 118
rect 785 17 835 97
rect 1457 85 1507 129
rect 1073 51 1089 85
rect 1123 51 1507 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 31 168 65 202
rect 511 180 534 202
rect 534 180 545 202
rect 511 168 545 180
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 19 202 77 208
rect 19 168 31 202
rect 65 199 77 202
rect 499 202 557 208
rect 499 199 511 202
rect 65 171 511 199
rect 65 168 77 171
rect 19 162 77 168
rect 499 168 511 171
rect 545 168 557 202
rect 499 162 557 168
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a311o_4
flabel pwell s 0 0 1536 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nwell s 0 617 1536 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 10 nsew
flabel metal1 s 0 617 1536 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 1536 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 C1
port 5 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 B1
port 4 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 1471 316 1505 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 1183 316 1217 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 1279 316 1313 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 1375 316 1409 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 1536 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3594508
string GDS_START 3582222
<< end >>
