magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 301 333 367 492
rect 489 333 555 492
rect 677 333 743 492
rect 301 299 815 333
rect 17 143 79 265
rect 749 181 815 299
rect 301 147 815 181
rect 301 51 367 147
rect 489 51 555 147
rect 677 51 743 147
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 19 299 79 527
rect 113 265 179 493
rect 213 299 267 527
rect 401 367 455 527
rect 589 367 643 527
rect 777 367 831 527
rect 113 215 678 265
rect 29 17 79 109
rect 113 53 179 215
rect 213 17 267 122
rect 401 17 455 113
rect 589 17 643 113
rect 777 17 831 113
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
rlabel locali s 17 143 79 265 6 A
port 1 nsew signal input
rlabel locali s 749 181 815 299 6 X
port 2 nsew signal output
rlabel locali s 677 333 743 492 6 X
port 2 nsew signal output
rlabel locali s 677 51 743 147 6 X
port 2 nsew signal output
rlabel locali s 489 333 555 492 6 X
port 2 nsew signal output
rlabel locali s 489 51 555 147 6 X
port 2 nsew signal output
rlabel locali s 301 333 367 492 6 X
port 2 nsew signal output
rlabel locali s 301 299 815 333 6 X
port 2 nsew signal output
rlabel locali s 301 147 815 181 6 X
port 2 nsew signal output
rlabel locali s 301 51 367 147 6 X
port 2 nsew signal output
rlabel metal1 s 0 -48 920 48 8 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 496 920 592 6 VPWR
port 4 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 920 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3353952
string GDS_START 3346728
<< end >>
