magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 235 333 311 493
rect 435 333 501 493
rect 235 299 627 333
rect 85 199 164 265
rect 202 199 266 265
rect 300 192 352 265
rect 308 153 352 192
rect 386 153 445 265
rect 575 167 627 299
rect 555 51 627 167
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 17 319 101 385
rect 17 165 51 319
rect 151 299 201 527
rect 345 367 400 527
rect 575 367 618 527
rect 17 131 274 165
rect 479 199 541 265
rect 17 89 94 131
rect 240 119 274 131
rect 479 119 520 199
rect 133 17 206 97
rect 240 85 520 119
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 85 199 164 265 6 A_N
port 1 nsew signal input
rlabel locali s 386 153 445 265 6 B
port 2 nsew signal input
rlabel locali s 308 153 352 192 6 C
port 3 nsew signal input
rlabel locali s 300 192 352 265 6 C
port 3 nsew signal input
rlabel locali s 202 199 266 265 6 D
port 4 nsew signal input
rlabel locali s 575 167 627 299 6 Y
port 5 nsew signal output
rlabel locali s 555 51 627 167 6 Y
port 5 nsew signal output
rlabel locali s 435 333 501 493 6 Y
port 5 nsew signal output
rlabel locali s 235 333 311 493 6 Y
port 5 nsew signal output
rlabel locali s 235 299 627 333 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -48 644 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2321804
string GDS_START 2315926
<< end >>
