magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1196 561
rect 19 360 85 493
rect 119 326 153 487
rect 188 360 254 493
rect 288 326 322 487
rect 356 360 422 493
rect 456 326 490 487
rect 524 360 590 493
rect 624 326 658 487
rect 692 360 758 493
rect 792 326 826 487
rect 860 360 926 493
rect 960 326 994 487
rect 1028 360 1094 493
rect 23 292 1088 326
rect 23 173 57 292
rect 91 207 973 258
rect 1034 173 1088 292
rect 23 139 1088 173
rect 207 17 273 105
rect 307 56 345 139
rect 379 17 445 105
rect 479 56 517 139
rect 551 17 617 105
rect 651 56 689 139
rect 723 17 789 105
rect 823 56 861 139
rect 895 17 961 105
rect 0 -17 1196 17
<< metal1 >>
rect 0 496 1196 592
rect 14 428 1182 468
rect 14 416 72 428
rect 186 416 244 428
rect 366 416 424 428
rect 542 416 600 428
rect 687 416 745 428
rect 859 416 917 428
rect 1039 416 1097 428
rect 0 -48 1196 48
<< labels >>
rlabel locali s 91 207 973 258 6 A
port 1 nsew signal input
rlabel locali s 1034 173 1088 292 6 Y
port 2 nsew signal output
rlabel locali s 960 326 994 487 6 Y
port 2 nsew signal output
rlabel locali s 823 56 861 139 6 Y
port 2 nsew signal output
rlabel locali s 792 326 826 487 6 Y
port 2 nsew signal output
rlabel locali s 651 56 689 139 6 Y
port 2 nsew signal output
rlabel locali s 624 326 658 487 6 Y
port 2 nsew signal output
rlabel locali s 479 56 517 139 6 Y
port 2 nsew signal output
rlabel locali s 456 326 490 487 6 Y
port 2 nsew signal output
rlabel locali s 307 56 345 139 6 Y
port 2 nsew signal output
rlabel locali s 288 326 322 487 6 Y
port 2 nsew signal output
rlabel locali s 119 326 153 487 6 Y
port 2 nsew signal output
rlabel locali s 23 292 1088 326 6 Y
port 2 nsew signal output
rlabel locali s 23 173 57 292 6 Y
port 2 nsew signal output
rlabel locali s 23 139 1088 173 6 Y
port 2 nsew signal output
rlabel locali s 19 360 85 493 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 188 360 254 493 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 356 360 422 493 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 524 360 590 493 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 692 360 758 493 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 860 360 926 493 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 1028 360 1094 493 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 1039 416 1097 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 859 416 917 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 687 416 745 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 542 416 600 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 366 416 424 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 186 416 244 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 14 428 1182 468 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 14 416 72 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 895 17 961 105 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 723 17 789 105 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 551 17 617 105 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 379 17 445 105 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 207 17 273 105 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 1196 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1196 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 527 1196 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 1196 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2272554
string GDS_START 2262086
<< end >>
