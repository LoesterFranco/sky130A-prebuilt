magic
tech sky130A
magscale 1 2
timestamp 1604502741
<< locali >>
rect 85 236 161 310
rect 392 365 458 431
rect 872 581 1066 615
rect 872 331 906 581
rect 1032 467 1066 581
rect 1208 581 1490 615
rect 1208 467 1242 581
rect 1032 433 1242 467
rect 846 282 912 331
rect 1456 382 1490 581
rect 1456 360 1703 382
rect 1456 348 1714 360
rect 1648 294 1714 348
rect 2224 364 2292 596
rect 2047 196 2116 330
rect 2258 226 2292 364
rect 2213 70 2292 226
rect 2505 70 2572 596
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2592 683
rect 17 378 107 596
rect 141 412 207 649
rect 17 344 229 378
rect 17 202 51 344
rect 195 260 229 344
rect 263 317 313 596
rect 361 485 482 649
rect 516 459 591 551
rect 263 251 523 317
rect 263 226 297 251
rect 17 70 89 202
rect 123 17 189 202
rect 225 70 297 226
rect 557 217 591 459
rect 331 17 381 213
rect 417 183 591 217
rect 625 359 686 467
rect 788 393 838 649
rect 625 325 812 359
rect 940 399 990 547
rect 1100 501 1174 649
rect 1308 456 1374 547
rect 1308 422 1422 456
rect 940 365 1204 399
rect 417 121 467 183
rect 625 149 659 325
rect 515 83 659 149
rect 693 180 744 291
rect 778 248 812 325
rect 1170 317 1204 365
rect 1288 322 1354 388
rect 949 251 1020 317
rect 949 248 983 251
rect 778 214 983 248
rect 1062 236 1128 317
rect 1170 251 1236 317
rect 1170 202 1204 251
rect 1017 180 1204 202
rect 693 168 1204 180
rect 693 146 1067 168
rect 1003 119 1067 146
rect 1238 134 1286 217
rect 712 17 831 112
rect 883 85 965 112
rect 1102 85 1168 134
rect 883 51 1168 85
rect 1212 17 1286 134
rect 1320 85 1354 322
rect 1388 314 1422 422
rect 1524 530 1684 649
rect 1737 482 1787 596
rect 1894 516 1960 649
rect 2118 516 2184 649
rect 1737 476 2190 482
rect 1524 448 2190 476
rect 1524 416 1877 448
rect 1737 394 1877 416
rect 1388 280 1614 314
rect 1388 119 1435 280
rect 1580 260 1614 280
rect 1756 260 1809 310
rect 1469 85 1534 246
rect 1580 226 1809 260
rect 1843 192 1877 394
rect 1942 364 2081 414
rect 1942 238 2013 364
rect 2156 330 2190 448
rect 1320 51 1534 85
rect 1617 17 1683 192
rect 1717 85 1783 192
rect 1817 119 1877 192
rect 1911 85 1945 204
rect 1717 51 1945 85
rect 1979 162 2013 238
rect 2156 264 2224 330
rect 1979 70 2077 162
rect 2113 17 2179 162
rect 2328 406 2378 582
rect 2328 317 2362 406
rect 2415 364 2465 649
rect 2328 251 2471 317
rect 2328 70 2375 251
rect 2411 17 2461 162
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2592 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
<< metal1 >>
rect 0 683 2592 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2592 683
rect 0 617 2592 649
rect 0 17 2592 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2592 17
rect 0 -49 2592 -17
<< obsm1 >>
rect 1075 273 1133 282
rect 1939 273 1997 282
rect 1075 245 1997 273
rect 1075 236 1133 245
rect 1939 236 1997 245
<< labels >>
rlabel locali s 392 365 458 431 6 D
port 1 nsew signal input
rlabel locali s 2505 70 2572 596 6 Q
port 2 nsew signal output
rlabel locali s 2258 226 2292 364 6 Q_N
port 3 nsew signal output
rlabel locali s 2224 364 2292 596 6 Q_N
port 3 nsew signal output
rlabel locali s 2213 70 2292 226 6 Q_N
port 3 nsew signal output
rlabel locali s 2047 196 2116 330 6 RESET_B
port 4 nsew signal input
rlabel locali s 1648 294 1714 348 6 SET_B
port 5 nsew signal input
rlabel locali s 1456 382 1490 581 6 SET_B
port 5 nsew signal input
rlabel locali s 1456 360 1703 382 6 SET_B
port 5 nsew signal input
rlabel locali s 1456 348 1714 360 6 SET_B
port 5 nsew signal input
rlabel locali s 1208 581 1490 615 6 SET_B
port 5 nsew signal input
rlabel locali s 1208 467 1242 581 6 SET_B
port 5 nsew signal input
rlabel locali s 1032 467 1066 581 6 SET_B
port 5 nsew signal input
rlabel locali s 1032 433 1242 467 6 SET_B
port 5 nsew signal input
rlabel locali s 872 581 1066 615 6 SET_B
port 5 nsew signal input
rlabel locali s 872 331 906 581 6 SET_B
port 5 nsew signal input
rlabel locali s 846 282 912 331 6 SET_B
port 5 nsew signal input
rlabel locali s 85 236 161 310 6 CLK
port 6 nsew clock input
rlabel metal1 s 0 -49 2592 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 617 2592 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2592 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 2660358
string GDS_START 2641094
<< end >>
