magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 101 236 167 302
rect 409 270 551 356
rect 601 270 712 356
rect 914 394 980 596
rect 1114 394 1180 596
rect 914 360 1319 394
rect 1187 226 1221 360
rect 1273 310 1319 360
rect 993 192 1221 226
rect 993 70 1043 192
rect 1185 70 1221 192
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 95 370 161 572
rect 195 404 261 649
rect 295 424 361 572
rect 395 458 461 649
rect 495 424 561 572
rect 595 458 661 649
rect 707 424 780 572
rect 295 390 780 424
rect 23 336 261 370
rect 295 364 373 390
rect 23 202 57 336
rect 227 330 261 336
rect 227 264 305 330
rect 339 230 373 364
rect 746 326 780 390
rect 814 364 880 649
rect 1014 428 1080 649
rect 1214 428 1280 649
rect 746 292 1153 326
rect 951 260 1153 292
rect 23 70 89 202
rect 123 17 175 202
rect 235 85 301 230
rect 337 119 373 230
rect 407 144 473 230
rect 507 202 857 236
rect 507 178 573 202
rect 407 94 659 144
rect 407 85 473 94
rect 235 51 473 85
rect 705 17 771 168
rect 807 90 857 202
rect 893 17 959 226
rect 1079 17 1145 158
rect 1255 17 1321 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
<< metal1 >>
rect 0 683 1344 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 0 617 1344 649
rect 0 17 1344 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
rect 0 -49 1344 -17
<< labels >>
rlabel locali s 101 236 167 302 6 A_N
port 1 nsew signal input
rlabel locali s 409 270 551 356 6 B
port 2 nsew signal input
rlabel locali s 601 270 712 356 6 C
port 3 nsew signal input
rlabel locali s 1273 310 1319 360 6 X
port 4 nsew signal output
rlabel locali s 1187 226 1221 360 6 X
port 4 nsew signal output
rlabel locali s 1185 70 1221 192 6 X
port 4 nsew signal output
rlabel locali s 1114 394 1180 596 6 X
port 4 nsew signal output
rlabel locali s 993 192 1221 226 6 X
port 4 nsew signal output
rlabel locali s 993 70 1043 192 6 X
port 4 nsew signal output
rlabel locali s 914 394 980 596 6 X
port 4 nsew signal output
rlabel locali s 914 360 1319 394 6 X
port 4 nsew signal output
rlabel metal1 s 0 -49 1344 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 617 1344 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1344 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3261000
string GDS_START 3250274
<< end >>
