magic
tech sky130A
magscale 1 2
timestamp 1604502697
<< nwell >>
rect -38 261 2338 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 89 47 119 177
rect 183 47 213 177
rect 277 47 307 177
rect 371 47 401 177
rect 455 47 485 177
rect 549 47 579 177
rect 643 47 673 177
rect 747 47 777 177
rect 955 47 985 177
rect 1049 47 1079 177
rect 1143 47 1173 177
rect 1237 47 1267 177
rect 1349 47 1379 177
rect 1443 47 1473 177
rect 1537 47 1567 177
rect 1641 47 1671 177
rect 1829 47 1859 177
rect 1923 47 1953 177
rect 2017 47 2047 177
rect 2121 47 2151 177
<< pmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 457 297 493 497
rect 551 297 587 497
rect 645 297 681 497
rect 739 297 775 497
rect 837 297 873 497
rect 931 297 967 497
rect 1025 297 1061 497
rect 1210 297 1246 497
rect 1351 297 1387 497
rect 1445 297 1481 497
rect 1539 297 1575 497
rect 1633 297 1669 497
rect 1831 297 1867 497
rect 1925 297 1961 497
rect 2019 297 2055 497
rect 2113 297 2149 497
<< ndiff >>
rect 27 101 89 177
rect 27 67 35 101
rect 69 67 89 101
rect 27 47 89 67
rect 119 93 183 177
rect 119 59 129 93
rect 163 59 183 93
rect 119 47 183 59
rect 213 101 277 177
rect 213 67 223 101
rect 257 67 277 101
rect 213 47 277 67
rect 307 93 371 177
rect 307 59 317 93
rect 351 59 371 93
rect 307 47 371 59
rect 401 109 455 177
rect 401 75 411 109
rect 445 75 455 109
rect 401 47 455 75
rect 485 161 549 177
rect 485 127 505 161
rect 539 127 549 161
rect 485 47 549 127
rect 579 93 643 177
rect 579 59 599 93
rect 633 59 643 93
rect 579 47 643 59
rect 673 161 747 177
rect 673 127 693 161
rect 727 127 747 161
rect 673 47 747 127
rect 777 93 829 177
rect 777 59 787 93
rect 821 59 829 93
rect 777 47 829 59
rect 893 93 955 177
rect 893 59 901 93
rect 935 59 955 93
rect 893 47 955 59
rect 985 161 1049 177
rect 985 127 995 161
rect 1029 127 1049 161
rect 985 47 1049 127
rect 1079 93 1143 177
rect 1079 59 1089 93
rect 1123 59 1143 93
rect 1079 47 1143 59
rect 1173 161 1237 177
rect 1173 127 1183 161
rect 1217 127 1237 161
rect 1173 47 1237 127
rect 1267 93 1349 177
rect 1267 59 1277 93
rect 1311 59 1349 93
rect 1267 47 1349 59
rect 1379 161 1443 177
rect 1379 127 1399 161
rect 1433 127 1443 161
rect 1379 47 1443 127
rect 1473 93 1537 177
rect 1473 59 1493 93
rect 1527 59 1537 93
rect 1473 47 1537 59
rect 1567 161 1641 177
rect 1567 127 1587 161
rect 1621 127 1641 161
rect 1567 47 1641 127
rect 1671 93 1723 177
rect 1671 59 1681 93
rect 1715 59 1723 93
rect 1671 47 1723 59
rect 1777 93 1829 177
rect 1777 59 1785 93
rect 1819 59 1829 93
rect 1777 47 1829 59
rect 1859 101 1923 177
rect 1859 67 1879 101
rect 1913 67 1923 101
rect 1859 47 1923 67
rect 1953 93 2017 177
rect 1953 59 1973 93
rect 2007 59 2017 93
rect 1953 47 2017 59
rect 2047 101 2121 177
rect 2047 67 2067 101
rect 2101 67 2121 101
rect 2047 47 2121 67
rect 2151 93 2207 177
rect 2151 59 2163 93
rect 2197 59 2207 93
rect 2151 47 2207 59
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 297 81 451
rect 117 417 175 497
rect 117 383 129 417
rect 163 383 175 417
rect 117 349 175 383
rect 117 315 129 349
rect 163 315 175 349
rect 117 297 175 315
rect 211 485 269 497
rect 211 451 223 485
rect 257 451 269 485
rect 211 297 269 451
rect 305 417 363 497
rect 305 383 317 417
rect 351 383 363 417
rect 305 349 363 383
rect 305 315 317 349
rect 351 315 363 349
rect 305 297 363 315
rect 399 485 457 497
rect 399 451 411 485
rect 445 451 457 485
rect 399 297 457 451
rect 493 417 551 497
rect 493 383 505 417
rect 539 383 551 417
rect 493 349 551 383
rect 493 315 505 349
rect 539 315 551 349
rect 493 297 551 315
rect 587 485 645 497
rect 587 451 599 485
rect 633 451 645 485
rect 587 297 645 451
rect 681 417 739 497
rect 681 383 693 417
rect 727 383 739 417
rect 681 349 739 383
rect 681 315 693 349
rect 727 315 739 349
rect 681 297 739 315
rect 775 469 837 497
rect 775 435 787 469
rect 821 435 837 469
rect 775 297 837 435
rect 873 485 931 497
rect 873 451 885 485
rect 919 451 931 485
rect 873 417 931 451
rect 873 383 885 417
rect 919 383 931 417
rect 873 297 931 383
rect 967 477 1025 497
rect 967 443 979 477
rect 1013 443 1025 477
rect 967 409 1025 443
rect 967 375 979 409
rect 1013 375 1025 409
rect 967 297 1025 375
rect 1061 485 1210 497
rect 1061 383 1080 485
rect 1182 383 1210 485
rect 1061 297 1210 383
rect 1246 477 1351 497
rect 1246 443 1258 477
rect 1292 443 1351 477
rect 1246 409 1351 443
rect 1246 375 1258 409
rect 1292 375 1351 409
rect 1246 297 1351 375
rect 1387 485 1445 497
rect 1387 451 1399 485
rect 1433 451 1445 485
rect 1387 417 1445 451
rect 1387 383 1399 417
rect 1433 383 1445 417
rect 1387 297 1445 383
rect 1481 477 1539 497
rect 1481 443 1493 477
rect 1527 443 1539 477
rect 1481 409 1539 443
rect 1481 375 1493 409
rect 1527 375 1539 409
rect 1481 297 1539 375
rect 1575 485 1633 497
rect 1575 451 1587 485
rect 1621 451 1633 485
rect 1575 297 1633 451
rect 1669 477 1831 497
rect 1669 443 1681 477
rect 1715 443 1831 477
rect 1669 409 1831 443
rect 1669 375 1681 409
rect 1715 375 1831 409
rect 1669 297 1831 375
rect 1867 485 1925 497
rect 1867 451 1879 485
rect 1913 451 1925 485
rect 1867 417 1925 451
rect 1867 383 1879 417
rect 1913 383 1925 417
rect 1867 297 1925 383
rect 1961 477 2019 497
rect 1961 443 1973 477
rect 2007 443 2019 477
rect 1961 409 2019 443
rect 1961 375 1973 409
rect 2007 375 2019 409
rect 1961 297 2019 375
rect 2055 485 2113 497
rect 2055 451 2067 485
rect 2101 451 2113 485
rect 2055 417 2113 451
rect 2055 383 2067 417
rect 2101 383 2113 417
rect 2055 297 2113 383
rect 2149 477 2203 497
rect 2149 443 2161 477
rect 2195 443 2203 477
rect 2149 409 2203 443
rect 2149 375 2161 409
rect 2195 375 2203 409
rect 2149 297 2203 375
<< ndiffc >>
rect 35 67 69 101
rect 129 59 163 93
rect 223 67 257 101
rect 317 59 351 93
rect 411 75 445 109
rect 505 127 539 161
rect 599 59 633 93
rect 693 127 727 161
rect 787 59 821 93
rect 901 59 935 93
rect 995 127 1029 161
rect 1089 59 1123 93
rect 1183 127 1217 161
rect 1277 59 1311 93
rect 1399 127 1433 161
rect 1493 59 1527 93
rect 1587 127 1621 161
rect 1681 59 1715 93
rect 1785 59 1819 93
rect 1879 67 1913 101
rect 1973 59 2007 93
rect 2067 67 2101 101
rect 2163 59 2197 93
<< pdiffc >>
rect 35 451 69 485
rect 129 383 163 417
rect 129 315 163 349
rect 223 451 257 485
rect 317 383 351 417
rect 317 315 351 349
rect 411 451 445 485
rect 505 383 539 417
rect 505 315 539 349
rect 599 451 633 485
rect 693 383 727 417
rect 693 315 727 349
rect 787 435 821 469
rect 885 451 919 485
rect 885 383 919 417
rect 979 443 1013 477
rect 979 375 1013 409
rect 1080 383 1182 485
rect 1258 443 1292 477
rect 1258 375 1292 409
rect 1399 451 1433 485
rect 1399 383 1433 417
rect 1493 443 1527 477
rect 1493 375 1527 409
rect 1587 451 1621 485
rect 1681 443 1715 477
rect 1681 375 1715 409
rect 1879 451 1913 485
rect 1879 383 1913 417
rect 1973 443 2007 477
rect 1973 375 2007 409
rect 2067 451 2101 485
rect 2067 383 2101 417
rect 2161 443 2195 477
rect 2161 375 2195 409
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 457 497 493 523
rect 551 497 587 523
rect 645 497 681 523
rect 739 497 775 523
rect 837 497 873 523
rect 931 497 967 523
rect 1025 497 1061 523
rect 1210 497 1246 523
rect 1351 497 1387 523
rect 1445 497 1481 523
rect 1539 497 1575 523
rect 1633 497 1669 523
rect 1831 497 1867 523
rect 1925 497 1961 523
rect 2019 497 2055 523
rect 2113 497 2149 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 457 282 493 297
rect 551 282 587 297
rect 645 282 681 297
rect 739 282 775 297
rect 837 282 873 297
rect 931 282 967 297
rect 1025 282 1061 297
rect 1210 282 1246 297
rect 1351 282 1387 297
rect 1445 282 1481 297
rect 1539 282 1575 297
rect 1633 282 1669 297
rect 1831 282 1867 297
rect 1925 282 1961 297
rect 2019 282 2055 297
rect 2113 282 2149 297
rect 79 265 119 282
rect 173 265 213 282
rect 267 265 307 282
rect 361 265 401 282
rect 79 261 401 265
rect 22 249 401 261
rect 22 215 38 249
rect 72 215 106 249
rect 140 215 184 249
rect 218 215 262 249
rect 296 215 401 249
rect 22 205 401 215
rect 89 199 401 205
rect 89 177 119 199
rect 183 177 213 199
rect 277 177 307 199
rect 371 177 401 199
rect 455 265 495 282
rect 549 265 589 282
rect 643 265 683 282
rect 737 265 777 282
rect 455 249 777 265
rect 455 215 567 249
rect 601 215 645 249
rect 679 215 723 249
rect 757 215 777 249
rect 455 199 777 215
rect 835 269 875 282
rect 929 269 969 282
rect 1023 269 1063 282
rect 1208 269 1248 282
rect 835 265 1248 269
rect 1349 269 1389 282
rect 1443 269 1483 282
rect 1537 269 1577 282
rect 1631 269 1671 282
rect 835 249 1267 265
rect 835 215 851 249
rect 885 215 929 249
rect 963 215 1007 249
rect 1041 215 1085 249
rect 1119 215 1153 249
rect 1187 215 1267 249
rect 835 202 1267 215
rect 835 199 1173 202
rect 455 177 485 199
rect 549 177 579 199
rect 643 177 673 199
rect 747 177 777 199
rect 955 177 985 199
rect 1049 177 1079 199
rect 1143 177 1173 199
rect 1237 177 1267 202
rect 1349 249 1671 269
rect 1349 215 1365 249
rect 1399 215 1443 249
rect 1477 215 1521 249
rect 1555 215 1599 249
rect 1633 215 1671 249
rect 1349 202 1671 215
rect 1349 199 1567 202
rect 1349 177 1379 199
rect 1443 177 1473 199
rect 1537 177 1567 199
rect 1641 177 1671 202
rect 1829 265 1869 282
rect 1923 265 1963 282
rect 2017 265 2057 282
rect 2111 265 2151 282
rect 1829 261 2151 265
rect 1829 249 2207 261
rect 1829 215 1845 249
rect 1879 215 1923 249
rect 1957 215 2001 249
rect 2035 215 2079 249
rect 2113 215 2157 249
rect 2191 215 2207 249
rect 1829 203 2207 215
rect 1829 199 2151 203
rect 1829 177 1859 199
rect 1923 177 1953 199
rect 2017 177 2047 199
rect 2121 177 2151 199
rect 89 21 119 47
rect 183 21 213 47
rect 277 21 307 47
rect 371 21 401 47
rect 455 21 485 47
rect 549 21 579 47
rect 643 21 673 47
rect 747 21 777 47
rect 955 21 985 47
rect 1049 21 1079 47
rect 1143 21 1173 47
rect 1237 21 1267 47
rect 1349 21 1379 47
rect 1443 21 1473 47
rect 1537 21 1567 47
rect 1641 21 1671 47
rect 1829 21 1859 47
rect 1923 21 1953 47
rect 2017 21 2047 47
rect 2121 21 2151 47
<< polycont >>
rect 38 215 72 249
rect 106 215 140 249
rect 184 215 218 249
rect 262 215 296 249
rect 567 215 601 249
rect 645 215 679 249
rect 723 215 757 249
rect 851 215 885 249
rect 929 215 963 249
rect 1007 215 1041 249
rect 1085 215 1119 249
rect 1153 215 1187 249
rect 1365 215 1399 249
rect 1443 215 1477 249
rect 1521 215 1555 249
rect 1599 215 1633 249
rect 1845 215 1879 249
rect 1923 215 1957 249
rect 2001 215 2035 249
rect 2079 215 2113 249
rect 2157 215 2191 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2300 561
rect 859 485 935 527
rect 19 451 35 485
rect 69 451 223 485
rect 257 451 411 485
rect 445 451 599 485
rect 633 469 821 485
rect 633 451 787 469
rect 22 261 66 393
rect 103 383 129 417
rect 163 383 179 417
rect 103 349 179 383
rect 291 383 317 417
rect 351 383 367 417
rect 291 349 367 383
rect 435 383 505 417
rect 539 383 555 417
rect 435 349 555 383
rect 667 383 693 417
rect 727 383 743 417
rect 667 349 743 383
rect 103 315 129 349
rect 163 315 317 349
rect 351 315 505 349
rect 539 315 693 349
rect 727 315 743 349
rect 787 349 821 435
rect 859 451 885 485
rect 919 451 935 485
rect 859 417 935 451
rect 859 383 885 417
rect 919 383 935 417
rect 979 477 1013 493
rect 979 409 1013 443
rect 1064 485 1208 527
rect 1064 383 1080 485
rect 1182 383 1208 485
rect 1258 477 1292 493
rect 1258 409 1292 443
rect 979 349 1013 375
rect 1373 485 1449 527
rect 1373 451 1399 485
rect 1433 451 1449 485
rect 1373 417 1449 451
rect 1373 383 1399 417
rect 1433 383 1449 417
rect 1493 477 1527 493
rect 1493 409 1527 443
rect 1258 349 1292 375
rect 1561 485 1637 527
rect 1561 451 1587 485
rect 1621 451 1637 485
rect 1561 383 1637 451
rect 1681 477 1715 493
rect 1681 409 1715 443
rect 1493 349 1527 375
rect 1853 485 1929 527
rect 1853 451 1879 485
rect 1913 451 1929 485
rect 1853 417 1929 451
rect 1853 383 1879 417
rect 1913 383 1929 417
rect 1973 477 2007 493
rect 1973 409 2007 443
rect 1681 349 1715 375
rect 2041 485 2117 527
rect 2041 451 2067 485
rect 2101 451 2117 485
rect 2041 417 2117 451
rect 2041 383 2067 417
rect 2101 383 2117 417
rect 2161 477 2195 493
rect 2161 409 2195 443
rect 1973 349 2007 375
rect 2161 349 2195 375
rect 787 315 2195 349
rect 22 249 380 261
rect 22 215 38 249
rect 72 215 106 249
rect 140 215 184 249
rect 218 215 262 249
rect 296 215 380 249
rect 435 198 523 315
rect 567 249 791 265
rect 601 215 645 249
rect 679 215 723 249
rect 757 215 791 249
rect 835 249 1213 257
rect 835 215 851 249
rect 885 215 929 249
rect 963 215 1007 249
rect 1041 215 1085 249
rect 1119 215 1153 249
rect 1187 215 1213 249
rect 1349 249 1709 260
rect 1349 215 1365 249
rect 1399 215 1443 249
rect 1477 215 1521 249
rect 1555 215 1599 249
rect 1633 215 1709 249
rect 1829 249 2207 256
rect 1829 215 1845 249
rect 1879 215 1923 249
rect 1957 215 2001 249
rect 2035 215 2079 249
rect 2113 215 2157 249
rect 2191 215 2207 249
rect 567 199 791 215
rect 479 161 523 198
rect 35 127 445 161
rect 479 127 505 161
rect 539 127 693 161
rect 727 127 995 161
rect 1029 127 1183 161
rect 1217 127 1233 161
rect 1373 127 1399 161
rect 1433 127 1587 161
rect 1621 127 2101 161
rect 2151 151 2207 215
rect 35 101 69 127
rect 223 101 257 127
rect 35 51 69 67
rect 103 59 129 93
rect 163 59 179 93
rect 103 17 179 59
rect 411 109 445 127
rect 223 51 257 67
rect 291 59 317 93
rect 351 59 367 93
rect 1879 101 1913 127
rect 445 75 599 93
rect 411 59 599 75
rect 633 59 787 93
rect 821 59 837 93
rect 885 59 901 93
rect 935 59 1089 93
rect 1123 59 1277 93
rect 1311 59 1493 93
rect 1527 59 1681 93
rect 1715 59 1731 93
rect 1769 59 1785 93
rect 1819 59 1835 93
rect 291 17 367 59
rect 1769 17 1835 59
rect 2067 101 2101 127
rect 1879 51 1913 67
rect 1947 59 1973 93
rect 2007 59 2023 93
rect 1947 17 2023 59
rect 2067 51 2101 67
rect 2137 59 2163 93
rect 2197 59 2215 93
rect 2137 17 2215 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2300 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
<< metal1 >>
rect 0 561 2300 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2300 561
rect 0 496 2300 527
rect 0 17 2300 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2300 17
rect 0 -48 2300 -17
<< labels >>
flabel corelocali s 1968 221 2002 255 0 FreeSans 200 0 0 0 A3
port 3 nsew
flabel corelocali s 1864 221 1908 255 0 FreeSans 200 0 0 0 A3
port 3 nsew
flabel corelocali s 1673 221 1707 255 0 FreeSans 200 0 0 0 A2
port 2 nsew
flabel corelocali s 1498 221 1532 255 0 FreeSans 200 0 0 0 A2
port 2 nsew
flabel corelocali s 1402 221 1446 255 0 FreeSans 200 0 0 0 A2
port 2 nsew
flabel corelocali s 1596 221 1630 255 0 FreeSans 200 0 0 0 A2
port 2 nsew
flabel corelocali s 947 221 981 255 0 FreeSans 200 0 0 0 A1
port 1 nsew
flabel corelocali s 859 221 893 255 0 FreeSans 200 0 0 0 A1
port 1 nsew
flabel corelocali s 1138 221 1172 255 0 FreeSans 200 0 0 0 A1
port 1 nsew
flabel corelocali s 2153 153 2187 187 0 FreeSans 200 0 0 0 A3
port 3 nsew
flabel corelocali s 673 221 707 255 0 FreeSans 200 0 0 0 B1
port 4 nsew
flabel corelocali s 459 374 459 374 0 FreeSans 200 0 0 0 Y
port 10 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 200 0 0 0 B2
port 5 nsew
flabel corelocali s 214 221 248 255 0 FreeSans 200 0 0 0 B2
port 5 nsew
flabel corelocali s 123 221 157 255 0 FreeSans 200 0 0 0 B2
port 5 nsew
flabel corelocali s 30 289 64 323 0 FreeSans 200 0 0 0 B2
port 5 nsew
flabel corelocali s 30 357 64 391 0 FreeSans 200 0 0 0 B2
port 5 nsew
flabel corelocali s 305 221 339 255 0 FreeSans 200 0 0 0 B2
port 5 nsew
flabel corelocali s 459 238 459 238 0 FreeSans 200 0 0 0 Y
port 10 nsew
flabel corelocali s 459 306 459 306 0 FreeSans 200 0 0 0 Y
port 10 nsew
flabel corelocali s 581 221 615 255 0 FreeSans 200 0 0 0 B1
port 4 nsew
flabel corelocali s 1041 221 1075 255 0 FreeSans 200 0 0 0 A1
port 1 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel pwell s 47 0 47 0 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel nbase s 47 544 47 544 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew
flabel metal1 s 46 0 46 0 0 FreeSans 200 0 0 0 VGND
port 6 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew
flabel metal1 s 46 544 46 544 0 FreeSans 200 0 0 0 VPWR
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 2300 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1478552
string GDS_START 1461808
<< end >>
