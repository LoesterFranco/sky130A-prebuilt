magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 2918 704
rect 989 330 1209 332
rect 2374 329 2588 332
<< pwell >>
rect 0 0 2880 49
<< scnmos >>
rect 115 74 145 158
rect 193 74 223 158
rect 395 74 425 158
rect 497 74 527 158
rect 575 74 605 158
rect 788 74 818 222
rect 978 74 1008 222
rect 1168 97 1198 181
rect 1304 97 1334 181
rect 1419 97 1449 181
rect 1555 74 1585 202
rect 1777 74 1807 222
rect 1849 74 1879 222
rect 2197 118 2227 202
rect 2275 118 2305 202
rect 2406 74 2436 202
rect 2614 78 2644 226
rect 2766 78 2796 226
<< pmoshvt >>
rect 86 508 116 592
rect 164 508 194 592
rect 390 460 420 588
rect 526 504 556 588
rect 604 504 634 588
rect 806 368 836 592
rect 1084 366 1114 590
rect 1303 508 1333 592
rect 1393 508 1423 592
rect 1495 508 1525 592
rect 1619 424 1649 592
rect 1978 392 2008 592
rect 2062 392 2092 592
rect 2176 443 2206 527
rect 2272 443 2302 527
rect 2463 365 2493 565
rect 2665 368 2695 592
rect 2755 368 2785 592
<< ndiff >>
rect 731 186 788 222
rect 27 134 115 158
rect 27 100 70 134
rect 104 100 115 134
rect 27 74 115 100
rect 145 74 193 158
rect 223 133 280 158
rect 223 99 234 133
rect 268 99 280 133
rect 223 74 280 99
rect 334 146 395 158
rect 334 112 348 146
rect 382 112 395 146
rect 334 74 395 112
rect 425 133 497 158
rect 425 99 450 133
rect 484 99 497 133
rect 425 74 497 99
rect 527 74 575 158
rect 605 133 662 158
rect 605 99 616 133
rect 650 99 662 133
rect 605 74 662 99
rect 731 152 743 186
rect 777 152 788 186
rect 731 118 788 152
rect 731 84 743 118
rect 777 84 788 118
rect 731 74 788 84
rect 818 196 871 222
rect 818 162 829 196
rect 863 162 871 196
rect 818 120 871 162
rect 818 86 829 120
rect 863 86 871 120
rect 818 74 871 86
rect 925 127 978 222
rect 925 93 933 127
rect 967 93 978 127
rect 925 74 978 93
rect 1008 210 1061 222
rect 1008 176 1019 210
rect 1053 176 1061 210
rect 1505 181 1555 202
rect 1008 120 1061 176
rect 1008 86 1019 120
rect 1053 86 1061 120
rect 1115 169 1168 181
rect 1115 135 1123 169
rect 1157 135 1168 169
rect 1115 97 1168 135
rect 1198 169 1304 181
rect 1198 135 1259 169
rect 1293 135 1304 169
rect 1198 97 1304 135
rect 1334 97 1419 181
rect 1449 143 1555 181
rect 1449 109 1460 143
rect 1494 109 1555 143
rect 1449 97 1555 109
rect 1008 74 1061 86
rect 1505 74 1555 97
rect 1585 179 1642 202
rect 1585 145 1596 179
rect 1630 145 1642 179
rect 1585 74 1642 145
rect 1720 136 1777 222
rect 1720 102 1732 136
rect 1766 102 1777 136
rect 1720 74 1777 102
rect 1807 74 1849 222
rect 1879 202 1929 222
rect 1879 174 2197 202
rect 1879 140 1908 174
rect 1942 140 1991 174
rect 2025 140 2074 174
rect 2108 140 2152 174
rect 2186 140 2197 174
rect 1879 118 2197 140
rect 2227 118 2275 202
rect 2305 190 2406 202
rect 2305 156 2347 190
rect 2381 156 2406 190
rect 2305 120 2406 156
rect 2305 118 2347 120
rect 1879 74 1929 118
rect 2335 86 2347 118
rect 2381 86 2406 120
rect 2335 74 2406 86
rect 2436 190 2493 202
rect 2436 156 2447 190
rect 2481 156 2493 190
rect 2436 120 2493 156
rect 2436 86 2447 120
rect 2481 86 2493 120
rect 2436 74 2493 86
rect 2557 179 2614 226
rect 2557 145 2569 179
rect 2603 145 2614 179
rect 2557 78 2614 145
rect 2644 214 2766 226
rect 2644 180 2721 214
rect 2755 180 2766 214
rect 2644 124 2766 180
rect 2644 90 2721 124
rect 2755 90 2766 124
rect 2644 78 2766 90
rect 2796 214 2853 226
rect 2796 180 2807 214
rect 2841 180 2853 214
rect 2796 124 2853 180
rect 2796 90 2807 124
rect 2841 90 2853 124
rect 2796 78 2853 90
<< pdiff >>
rect 1543 627 1601 639
rect 27 567 86 592
rect 27 533 39 567
rect 73 533 86 567
rect 27 508 86 533
rect 116 508 164 592
rect 194 578 253 592
rect 194 544 207 578
rect 241 544 253 578
rect 194 508 253 544
rect 331 518 390 588
rect 331 484 343 518
rect 377 484 390 518
rect 331 460 390 484
rect 420 576 526 588
rect 420 542 479 576
rect 513 542 526 576
rect 420 504 526 542
rect 556 504 604 588
rect 634 563 693 588
rect 634 529 647 563
rect 681 529 693 563
rect 634 504 693 529
rect 747 580 806 592
rect 747 546 759 580
rect 793 546 806 580
rect 420 460 473 504
rect 747 368 806 546
rect 836 421 895 592
rect 1227 612 1285 624
rect 1025 571 1084 590
rect 1025 537 1037 571
rect 1071 537 1084 571
rect 836 387 849 421
rect 883 387 895 421
rect 836 368 895 387
rect 1025 366 1084 537
rect 1114 412 1173 590
rect 1227 578 1239 612
rect 1273 592 1285 612
rect 1543 593 1555 627
rect 1589 593 1601 627
rect 1543 592 1601 593
rect 1273 578 1303 592
rect 1227 508 1303 578
rect 1333 570 1393 592
rect 1333 536 1346 570
rect 1380 536 1393 570
rect 1333 508 1393 536
rect 1423 508 1495 592
rect 1525 508 1619 592
rect 1114 378 1127 412
rect 1161 378 1173 412
rect 1114 366 1173 378
rect 1566 424 1619 508
rect 1649 475 1708 592
rect 1919 580 1978 592
rect 1919 546 1931 580
rect 1965 546 1978 580
rect 1649 441 1662 475
rect 1696 441 1708 475
rect 1649 424 1708 441
rect 1919 511 1978 546
rect 1919 477 1931 511
rect 1965 477 1978 511
rect 1919 442 1978 477
rect 1919 408 1931 442
rect 1965 408 1978 442
rect 1919 392 1978 408
rect 2008 392 2062 592
rect 2092 580 2151 592
rect 2092 546 2105 580
rect 2139 546 2151 580
rect 2606 580 2665 592
rect 2092 527 2151 546
rect 2410 527 2463 565
rect 2092 511 2176 527
rect 2092 477 2105 511
rect 2139 477 2176 511
rect 2092 443 2176 477
rect 2206 443 2272 527
rect 2302 515 2463 527
rect 2302 481 2315 515
rect 2349 481 2406 515
rect 2440 481 2463 515
rect 2302 443 2463 481
rect 2092 442 2151 443
rect 2092 408 2105 442
rect 2139 408 2151 442
rect 2092 392 2151 408
rect 2410 365 2463 443
rect 2493 553 2552 565
rect 2493 519 2506 553
rect 2540 519 2552 553
rect 2493 482 2552 519
rect 2493 448 2506 482
rect 2540 448 2552 482
rect 2493 411 2552 448
rect 2493 377 2506 411
rect 2540 377 2552 411
rect 2493 365 2552 377
rect 2606 546 2618 580
rect 2652 546 2665 580
rect 2606 497 2665 546
rect 2606 463 2618 497
rect 2652 463 2665 497
rect 2606 414 2665 463
rect 2606 380 2618 414
rect 2652 380 2665 414
rect 2606 368 2665 380
rect 2695 580 2755 592
rect 2695 546 2708 580
rect 2742 546 2755 580
rect 2695 497 2755 546
rect 2695 463 2708 497
rect 2742 463 2755 497
rect 2695 414 2755 463
rect 2695 380 2708 414
rect 2742 380 2755 414
rect 2695 368 2755 380
rect 2785 580 2844 592
rect 2785 546 2798 580
rect 2832 546 2844 580
rect 2785 497 2844 546
rect 2785 463 2798 497
rect 2832 463 2844 497
rect 2785 414 2844 463
rect 2785 380 2798 414
rect 2832 380 2844 414
rect 2785 368 2844 380
<< ndiffc >>
rect 70 100 104 134
rect 234 99 268 133
rect 348 112 382 146
rect 450 99 484 133
rect 616 99 650 133
rect 743 152 777 186
rect 743 84 777 118
rect 829 162 863 196
rect 829 86 863 120
rect 933 93 967 127
rect 1019 176 1053 210
rect 1019 86 1053 120
rect 1123 135 1157 169
rect 1259 135 1293 169
rect 1460 109 1494 143
rect 1596 145 1630 179
rect 1732 102 1766 136
rect 1908 140 1942 174
rect 1991 140 2025 174
rect 2074 140 2108 174
rect 2152 140 2186 174
rect 2347 156 2381 190
rect 2347 86 2381 120
rect 2447 156 2481 190
rect 2447 86 2481 120
rect 2569 145 2603 179
rect 2721 180 2755 214
rect 2721 90 2755 124
rect 2807 180 2841 214
rect 2807 90 2841 124
<< pdiffc >>
rect 39 533 73 567
rect 207 544 241 578
rect 343 484 377 518
rect 479 542 513 576
rect 647 529 681 563
rect 759 546 793 580
rect 1037 537 1071 571
rect 849 387 883 421
rect 1239 578 1273 612
rect 1555 593 1589 627
rect 1346 536 1380 570
rect 1127 378 1161 412
rect 1931 546 1965 580
rect 1662 441 1696 475
rect 1931 477 1965 511
rect 1931 408 1965 442
rect 2105 546 2139 580
rect 2105 477 2139 511
rect 2315 481 2349 515
rect 2406 481 2440 515
rect 2105 408 2139 442
rect 2506 519 2540 553
rect 2506 448 2540 482
rect 2506 377 2540 411
rect 2618 546 2652 580
rect 2618 463 2652 497
rect 2618 380 2652 414
rect 2708 546 2742 580
rect 2708 463 2742 497
rect 2708 380 2742 414
rect 2798 546 2832 580
rect 2798 463 2832 497
rect 2798 380 2832 414
<< poly >>
rect 86 592 116 618
rect 164 592 194 618
rect 390 588 420 614
rect 526 588 556 614
rect 604 588 634 614
rect 806 592 836 618
rect 86 493 116 508
rect 164 493 194 508
rect 83 398 119 493
rect 161 476 197 493
rect 161 446 231 476
rect 526 489 556 504
rect 604 489 634 504
rect 523 476 559 489
rect 201 424 231 446
rect 390 445 420 460
rect 488 446 559 476
rect 201 408 267 424
rect 387 408 423 445
rect 488 408 518 446
rect 83 382 151 398
rect 83 348 101 382
rect 135 348 151 382
rect 83 314 151 348
rect 83 280 101 314
rect 135 280 151 314
rect 201 374 217 408
rect 251 374 267 408
rect 201 340 267 374
rect 201 306 217 340
rect 251 306 267 340
rect 201 290 267 306
rect 315 378 518 408
rect 601 398 637 489
rect 575 382 641 398
rect 315 340 423 378
rect 315 306 331 340
rect 365 306 423 340
rect 575 348 591 382
rect 625 348 641 382
rect 1084 590 1114 616
rect 927 412 1008 428
rect 927 378 943 412
rect 977 378 1008 412
rect 806 353 836 368
rect 315 290 423 306
rect 467 314 533 330
rect 83 246 151 280
rect 83 212 101 246
rect 135 212 151 246
rect 83 196 151 212
rect 315 203 345 290
rect 467 280 483 314
rect 517 280 533 314
rect 467 246 533 280
rect 467 212 483 246
rect 517 212 533 246
rect 115 158 145 196
rect 193 173 425 203
rect 467 196 533 212
rect 575 314 641 348
rect 575 280 591 314
rect 625 280 641 314
rect 803 310 839 353
rect 927 351 1008 378
rect 1303 592 1333 618
rect 1393 592 1423 618
rect 1495 592 1525 618
rect 1619 592 1649 618
rect 1978 592 2008 618
rect 2062 592 2092 618
rect 2665 592 2695 618
rect 2755 592 2785 618
rect 1303 493 1333 508
rect 1393 493 1423 508
rect 1495 493 1525 508
rect 1300 481 1336 493
rect 1205 460 1336 481
rect 1390 476 1426 493
rect 1205 426 1221 460
rect 1255 451 1336 460
rect 1378 460 1444 476
rect 1255 426 1271 451
rect 1205 410 1271 426
rect 1378 426 1394 460
rect 1428 426 1444 460
rect 1378 403 1444 426
rect 1319 373 1444 403
rect 1084 351 1114 366
rect 1319 351 1349 373
rect 927 321 1349 351
rect 1492 325 1528 493
rect 1740 501 1807 517
rect 1740 467 1756 501
rect 1790 467 1807 501
rect 1740 433 1807 467
rect 1619 409 1649 424
rect 1616 391 1652 409
rect 575 246 641 280
rect 575 212 591 246
rect 625 212 641 246
rect 743 294 877 310
rect 743 260 759 294
rect 793 260 827 294
rect 861 260 877 294
rect 743 244 877 260
rect 788 222 818 244
rect 978 222 1008 321
rect 575 196 641 212
rect 193 158 223 173
rect 395 158 425 173
rect 497 158 527 196
rect 575 158 605 196
rect 1168 181 1198 321
rect 1441 304 1528 325
rect 1441 273 1457 304
rect 1419 270 1457 273
rect 1491 295 1528 304
rect 1586 375 1652 391
rect 1586 341 1602 375
rect 1636 341 1652 375
rect 1586 325 1652 341
rect 1740 399 1756 433
rect 1790 399 1807 433
rect 1740 377 1807 399
rect 2463 565 2493 591
rect 2176 527 2206 553
rect 2272 527 2302 553
rect 2176 428 2206 443
rect 2272 428 2302 443
rect 1978 377 2008 392
rect 2062 377 2092 392
rect 1740 365 2011 377
rect 1740 331 1756 365
rect 1790 347 2011 365
rect 2059 358 2095 377
rect 2173 360 2209 428
rect 2272 411 2305 428
rect 2272 408 2378 411
rect 2275 395 2378 408
rect 2275 361 2328 395
rect 2362 361 2378 395
rect 1790 331 1807 347
rect 1491 270 1507 295
rect 1304 253 1377 269
rect 1304 219 1327 253
rect 1361 219 1377 253
rect 1304 203 1377 219
rect 1419 254 1507 270
rect 1419 243 1471 254
rect 1586 247 1616 325
rect 1740 315 1807 331
rect 1304 181 1334 203
rect 1419 181 1449 243
rect 1555 217 1616 247
rect 1777 222 1807 315
rect 2059 342 2125 358
rect 2059 308 2075 342
rect 2109 308 2125 342
rect 2059 292 2125 308
rect 2167 344 2233 360
rect 2167 310 2183 344
rect 2217 310 2233 344
rect 2167 294 2233 310
rect 2275 345 2378 361
rect 2463 350 2493 365
rect 2665 353 2695 368
rect 2755 353 2785 368
rect 2460 349 2496 350
rect 1951 274 2017 290
rect 1951 267 1967 274
rect 1849 240 1967 267
rect 2001 240 2017 274
rect 1849 237 2017 240
rect 1849 222 1879 237
rect 1951 224 2017 237
rect 2095 252 2125 292
rect 2095 222 2227 252
rect 1555 202 1585 217
rect 115 48 145 74
rect 193 48 223 74
rect 395 48 425 74
rect 497 48 527 74
rect 575 48 605 74
rect 788 48 818 74
rect 978 48 1008 74
rect 1168 71 1198 97
rect 1304 71 1334 97
rect 1419 71 1449 97
rect 2197 202 2227 222
rect 2275 202 2305 345
rect 2426 303 2496 349
rect 2662 303 2698 353
rect 2752 330 2788 353
rect 2426 297 2698 303
rect 2347 281 2698 297
rect 2347 247 2363 281
rect 2397 247 2698 281
rect 2740 314 2806 330
rect 2740 280 2756 314
rect 2790 280 2806 314
rect 2740 264 2806 280
rect 2347 241 2698 247
rect 2347 231 2456 241
rect 2406 202 2436 231
rect 2614 226 2644 241
rect 2766 226 2796 264
rect 2197 92 2227 118
rect 2275 92 2305 118
rect 1555 48 1585 74
rect 1777 48 1807 74
rect 1849 48 1879 74
rect 2406 48 2436 74
rect 2614 52 2644 78
rect 2766 52 2796 78
<< polycont >>
rect 101 348 135 382
rect 101 280 135 314
rect 217 374 251 408
rect 217 306 251 340
rect 331 306 365 340
rect 591 348 625 382
rect 943 378 977 412
rect 101 212 135 246
rect 483 280 517 314
rect 483 212 517 246
rect 591 280 625 314
rect 1221 426 1255 460
rect 1394 426 1428 460
rect 1756 467 1790 501
rect 591 212 625 246
rect 759 260 793 294
rect 827 260 861 294
rect 1457 270 1491 304
rect 1602 341 1636 375
rect 1756 399 1790 433
rect 1756 331 1790 365
rect 2328 361 2362 395
rect 1327 219 1361 253
rect 2075 308 2109 342
rect 2183 310 2217 344
rect 1967 240 2001 274
rect 2363 247 2397 281
rect 2756 280 2790 314
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2880 683
rect 17 567 89 596
rect 17 533 39 567
rect 73 533 89 567
rect 17 492 89 533
rect 191 578 241 649
rect 191 544 207 578
rect 191 526 241 544
rect 275 581 445 615
rect 275 492 309 581
rect 17 458 309 492
rect 343 518 377 547
rect 17 150 51 458
rect 343 424 377 484
rect 411 492 445 581
rect 479 576 529 649
rect 513 542 529 576
rect 479 526 529 542
rect 631 563 709 592
rect 631 529 647 563
rect 681 529 709 563
rect 743 580 809 649
rect 743 546 759 580
rect 793 546 809 580
rect 743 530 809 546
rect 1021 571 1087 649
rect 1539 627 1605 649
rect 1021 537 1037 571
rect 1071 537 1087 571
rect 1021 530 1087 537
rect 1121 578 1239 612
rect 1273 578 1289 612
rect 631 496 709 529
rect 1121 496 1155 578
rect 1330 570 1396 596
rect 1539 593 1555 627
rect 1589 593 1605 627
rect 1539 577 1605 593
rect 1330 544 1346 570
rect 631 492 1155 496
rect 411 462 1155 492
rect 1310 536 1346 544
rect 1380 536 1396 570
rect 1639 551 1881 585
rect 1639 543 1673 551
rect 1310 510 1396 536
rect 411 458 709 462
rect 201 408 533 424
rect 85 382 167 398
rect 85 348 101 382
rect 135 348 167 382
rect 85 314 167 348
rect 85 280 101 314
rect 135 280 167 314
rect 85 246 167 280
rect 85 212 101 246
rect 135 212 167 246
rect 201 374 217 408
rect 251 390 533 408
rect 251 374 267 390
rect 201 340 267 374
rect 201 306 217 340
rect 251 306 267 340
rect 201 256 267 306
rect 313 340 381 356
rect 313 306 331 340
rect 365 306 381 340
rect 313 290 381 306
rect 467 314 533 390
rect 467 280 483 314
rect 517 280 533 314
rect 201 222 400 256
rect 85 196 167 212
rect 17 134 120 150
rect 17 100 70 134
rect 104 100 120 134
rect 17 84 120 100
rect 218 133 284 162
rect 218 99 234 133
rect 268 99 284 133
rect 218 17 284 99
rect 330 146 400 222
rect 467 246 533 280
rect 467 212 483 246
rect 517 212 533 246
rect 467 196 533 212
rect 575 382 641 398
rect 575 348 591 382
rect 625 350 641 382
rect 575 316 607 348
rect 575 314 641 316
rect 575 280 591 314
rect 625 280 641 314
rect 575 246 641 280
rect 575 212 591 246
rect 625 212 641 246
rect 575 196 641 212
rect 675 162 709 458
rect 833 421 993 428
rect 833 387 849 421
rect 883 412 993 421
rect 883 387 943 412
rect 833 378 943 387
rect 977 378 993 412
rect 833 362 993 378
rect 743 294 877 310
rect 743 260 759 294
rect 793 260 827 294
rect 861 260 877 294
rect 743 236 877 260
rect 911 202 945 362
rect 1043 294 1077 462
rect 1191 460 1271 476
rect 1191 428 1221 460
rect 1111 426 1221 428
rect 1255 426 1271 460
rect 1111 412 1271 426
rect 1111 378 1127 412
rect 1161 394 1271 412
rect 1161 378 1225 394
rect 1111 362 1225 378
rect 1043 260 1157 294
rect 330 112 348 146
rect 382 112 400 146
rect 330 96 400 112
rect 434 133 500 162
rect 434 99 450 133
rect 484 99 500 133
rect 434 17 500 99
rect 600 133 709 162
rect 600 99 616 133
rect 650 99 709 133
rect 600 70 709 99
rect 743 186 777 202
rect 743 118 777 152
rect 743 17 777 84
rect 813 196 945 202
rect 813 162 829 196
rect 863 168 945 196
rect 1019 210 1069 226
rect 1053 176 1069 210
rect 863 162 879 168
rect 813 120 879 162
rect 813 86 829 120
rect 863 86 879 120
rect 813 70 879 86
rect 917 127 983 134
rect 917 93 933 127
rect 967 93 983 127
rect 917 17 983 93
rect 1019 120 1069 176
rect 1053 86 1069 120
rect 1107 169 1157 260
rect 1107 135 1123 169
rect 1107 119 1157 135
rect 1019 85 1069 86
rect 1191 85 1225 362
rect 1310 382 1344 510
rect 1430 509 1673 543
rect 1430 476 1464 509
rect 1378 460 1464 476
rect 1740 501 1806 517
rect 1740 475 1756 501
rect 1378 426 1394 460
rect 1428 426 1464 460
rect 1378 416 1464 426
rect 1646 441 1662 475
rect 1696 467 1756 475
rect 1790 467 1806 501
rect 1696 441 1806 467
rect 1646 433 1806 441
rect 1646 425 1756 433
rect 1740 399 1756 425
rect 1790 399 1806 433
rect 1586 382 1652 391
rect 1310 375 1652 382
rect 1310 348 1602 375
rect 1310 337 1344 348
rect 1259 303 1344 337
rect 1586 341 1602 348
rect 1636 341 1652 375
rect 1586 329 1652 341
rect 1740 365 1806 399
rect 1740 331 1756 365
rect 1790 331 1806 365
rect 1441 304 1507 314
rect 1259 169 1293 303
rect 1441 270 1457 304
rect 1491 295 1507 304
rect 1740 295 1806 331
rect 1847 358 1881 551
rect 1915 580 1981 649
rect 1915 546 1931 580
rect 1965 546 1981 580
rect 1915 511 1981 546
rect 1915 477 1931 511
rect 1965 477 1981 511
rect 1915 442 1981 477
rect 1915 408 1931 442
rect 1965 408 1981 442
rect 1915 392 1981 408
rect 2089 580 2155 596
rect 2089 546 2105 580
rect 2139 546 2155 580
rect 2089 511 2155 546
rect 2089 477 2105 511
rect 2139 477 2155 511
rect 2089 442 2155 477
rect 2299 515 2456 649
rect 2585 580 2668 596
rect 2299 481 2315 515
rect 2349 481 2406 515
rect 2440 481 2456 515
rect 2299 465 2456 481
rect 2490 553 2540 569
rect 2490 519 2506 553
rect 2490 482 2540 519
rect 2089 408 2105 442
rect 2139 431 2155 442
rect 2490 448 2506 482
rect 2139 408 2289 431
rect 2490 424 2540 448
rect 2089 397 2289 408
rect 1847 342 2125 358
rect 1847 324 2075 342
rect 1491 270 1806 295
rect 2059 308 2075 324
rect 2109 308 2125 342
rect 2059 292 2125 308
rect 2167 344 2221 360
rect 2167 310 2183 344
rect 2217 310 2221 344
rect 1259 119 1293 135
rect 1327 253 1377 269
rect 1441 261 1806 270
rect 1840 274 2017 290
rect 1361 227 1377 253
rect 1361 219 1562 227
rect 1327 193 1562 219
rect 1327 85 1377 193
rect 1019 51 1377 85
rect 1444 143 1494 159
rect 1444 109 1460 143
rect 1444 17 1494 109
rect 1528 85 1562 193
rect 1596 179 1630 261
rect 1840 240 1967 274
rect 2001 258 2017 274
rect 2167 258 2221 310
rect 2001 240 2221 258
rect 1840 227 2221 240
rect 1596 119 1630 145
rect 1664 224 2221 227
rect 2255 297 2289 397
rect 2323 411 2540 424
rect 2323 395 2506 411
rect 2323 361 2328 395
rect 2362 377 2506 395
rect 2362 361 2540 377
rect 2585 546 2618 580
rect 2652 546 2668 580
rect 2585 497 2668 546
rect 2585 463 2618 497
rect 2652 463 2668 497
rect 2585 414 2668 463
rect 2585 380 2618 414
rect 2652 380 2668 414
rect 2585 364 2668 380
rect 2708 580 2758 649
rect 2742 546 2758 580
rect 2708 497 2758 546
rect 2742 463 2758 497
rect 2708 414 2758 463
rect 2742 380 2758 414
rect 2708 364 2758 380
rect 2798 580 2863 596
rect 2832 546 2863 580
rect 2798 497 2863 546
rect 2832 463 2863 497
rect 2798 414 2863 463
rect 2832 380 2863 414
rect 2798 364 2863 380
rect 2323 350 2497 361
rect 2323 345 2431 350
rect 2465 316 2497 350
rect 2255 281 2397 297
rect 2255 247 2363 281
rect 2255 231 2397 247
rect 1664 193 1874 224
rect 1664 85 1698 193
rect 2255 190 2289 231
rect 1908 174 2289 190
rect 1528 51 1698 85
rect 1732 136 1782 154
rect 1766 102 1782 136
rect 1942 140 1991 174
rect 2025 140 2074 174
rect 2108 140 2152 174
rect 2186 140 2289 174
rect 1908 124 2289 140
rect 2331 190 2397 197
rect 2331 156 2347 190
rect 2381 156 2397 190
rect 1732 17 1782 102
rect 2331 120 2397 156
rect 2331 86 2347 120
rect 2381 86 2397 120
rect 2331 17 2397 86
rect 2431 190 2497 316
rect 2585 200 2619 364
rect 2431 156 2447 190
rect 2481 156 2497 190
rect 2431 120 2497 156
rect 2553 179 2619 200
rect 2553 145 2569 179
rect 2603 145 2619 179
rect 2553 124 2619 145
rect 2653 314 2795 330
rect 2653 280 2756 314
rect 2790 280 2795 314
rect 2653 264 2795 280
rect 2431 86 2447 120
rect 2481 86 2497 120
rect 2431 85 2497 86
rect 2653 85 2687 264
rect 2829 230 2863 364
rect 2431 51 2687 85
rect 2721 214 2755 230
rect 2721 124 2755 180
rect 2721 17 2755 90
rect 2791 214 2863 230
rect 2791 180 2807 214
rect 2841 180 2863 214
rect 2791 124 2863 180
rect 2791 90 2807 124
rect 2841 90 2863 124
rect 2791 74 2863 90
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2880 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 607 348 625 350
rect 625 348 641 350
rect 607 316 641 348
rect 2431 316 2465 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
<< metal1 >>
rect 0 683 2880 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2880 683
rect 0 617 2880 649
rect 595 350 653 356
rect 595 316 607 350
rect 641 347 653 350
rect 2419 350 2477 356
rect 2419 347 2431 350
rect 641 319 2431 347
rect 641 316 653 319
rect 595 310 653 316
rect 2419 316 2431 319
rect 2465 316 2477 350
rect 2419 310 2477 316
rect 0 17 2880 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2880 17
rect 0 -49 2880 -17
<< labels >>
flabel comment s 1137 335 1137 335 0 FreeSans 200 0 0 0 no_jumper_check
rlabel comment s 0 0 0 0 4 edfxbp_1
flabel pwell s 0 0 2880 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 2880 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 2880 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 2880 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 799 242 833 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 2623 390 2657 424 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 2623 464 2657 498 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 2623 538 2657 572 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 127 242 161 276 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 DE
port 3 nsew
flabel corelocali s 2815 94 2849 128 0 FreeSans 340 0 0 0 Q_N
port 9 nsew
flabel corelocali s 2815 168 2849 202 0 FreeSans 340 0 0 0 Q_N
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 2880 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2170224
string GDS_START 2149858
<< end >>
