magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1288 561
rect 44 365 94 527
rect 128 323 178 493
rect 212 359 262 527
rect 296 323 346 493
rect 380 425 534 527
rect 820 425 886 527
rect 17 289 346 323
rect 17 181 74 289
rect 484 289 836 323
rect 484 215 591 289
rect 625 215 736 255
rect 770 215 836 289
rect 870 289 1147 323
rect 1181 291 1222 527
rect 870 215 936 289
rect 1113 255 1147 289
rect 980 215 1079 255
rect 1113 215 1271 255
rect 17 145 354 181
rect 52 17 86 111
rect 120 53 186 145
rect 220 17 254 111
rect 288 51 354 145
rect 388 17 422 111
rect 928 17 962 111
rect 1096 17 1130 111
rect 0 -17 1288 17
<< obsli1 >>
rect 568 459 786 493
rect 568 425 618 459
rect 736 425 786 459
rect 920 459 1138 493
rect 920 425 970 459
rect 652 391 702 425
rect 1004 391 1054 425
rect 380 357 1054 391
rect 1088 357 1138 459
rect 380 255 446 357
rect 108 215 446 255
rect 388 181 446 215
rect 388 147 794 181
rect 483 129 794 147
rect 828 147 1230 181
rect 828 95 894 147
rect 996 145 1230 147
rect 476 51 894 95
rect 996 51 1062 145
rect 1164 51 1230 145
<< metal1 >>
rect 0 496 1288 592
rect 0 -48 1288 48
<< labels >>
rlabel locali s 1113 255 1147 289 6 A1
port 1 nsew signal input
rlabel locali s 1113 215 1271 255 6 A1
port 1 nsew signal input
rlabel locali s 870 289 1147 323 6 A1
port 1 nsew signal input
rlabel locali s 870 215 936 289 6 A1
port 1 nsew signal input
rlabel locali s 980 215 1079 255 6 A2
port 2 nsew signal input
rlabel locali s 770 215 836 289 6 B1
port 3 nsew signal input
rlabel locali s 484 289 836 323 6 B1
port 3 nsew signal input
rlabel locali s 484 215 591 289 6 B1
port 3 nsew signal input
rlabel locali s 625 215 736 255 6 B2
port 4 nsew signal input
rlabel locali s 296 323 346 493 6 X
port 5 nsew signal output
rlabel locali s 288 51 354 145 6 X
port 5 nsew signal output
rlabel locali s 128 323 178 493 6 X
port 5 nsew signal output
rlabel locali s 120 53 186 145 6 X
port 5 nsew signal output
rlabel locali s 17 289 346 323 6 X
port 5 nsew signal output
rlabel locali s 17 181 74 289 6 X
port 5 nsew signal output
rlabel locali s 17 145 354 181 6 X
port 5 nsew signal output
rlabel locali s 1096 17 1130 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 928 17 962 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 388 17 422 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 220 17 254 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 52 17 86 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 1288 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1288 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1181 291 1222 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 820 425 886 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 380 425 534 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 212 359 262 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 44 365 94 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 1288 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 1288 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1288 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1489128
string GDS_START 1479502
<< end >>
