magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1472 561
rect 40 297 82 527
rect 116 333 182 493
rect 216 367 250 527
rect 284 333 350 493
rect 384 367 418 527
rect 452 333 518 493
rect 552 367 586 527
rect 620 333 686 493
rect 720 367 754 527
rect 788 333 854 493
rect 888 367 922 527
rect 956 333 1022 493
rect 1056 367 1090 527
rect 1124 333 1190 493
rect 1224 367 1258 527
rect 1292 333 1358 493
rect 1392 367 1434 527
rect 116 299 1358 333
rect 17 215 1105 263
rect 1292 181 1358 299
rect 36 17 82 177
rect 116 143 1358 181
rect 116 51 182 143
rect 216 17 250 109
rect 284 51 350 143
rect 384 17 418 109
rect 452 51 518 143
rect 552 17 586 109
rect 620 51 686 143
rect 720 17 754 109
rect 788 51 854 143
rect 888 17 922 109
rect 956 51 1022 143
rect 1056 17 1090 109
rect 1124 51 1190 143
rect 1224 17 1258 109
rect 1292 51 1358 143
rect 1392 17 1434 177
rect 0 -17 1472 17
<< metal1 >>
rect 0 496 1472 592
rect 0 -48 1472 48
<< labels >>
rlabel locali s 17 215 1105 263 6 A
port 1 nsew signal input
rlabel locali s 1292 333 1358 493 6 Y
port 2 nsew signal output
rlabel locali s 1292 181 1358 299 6 Y
port 2 nsew signal output
rlabel locali s 1292 51 1358 143 6 Y
port 2 nsew signal output
rlabel locali s 1124 333 1190 493 6 Y
port 2 nsew signal output
rlabel locali s 1124 51 1190 143 6 Y
port 2 nsew signal output
rlabel locali s 956 333 1022 493 6 Y
port 2 nsew signal output
rlabel locali s 956 51 1022 143 6 Y
port 2 nsew signal output
rlabel locali s 788 333 854 493 6 Y
port 2 nsew signal output
rlabel locali s 788 51 854 143 6 Y
port 2 nsew signal output
rlabel locali s 620 333 686 493 6 Y
port 2 nsew signal output
rlabel locali s 620 51 686 143 6 Y
port 2 nsew signal output
rlabel locali s 452 333 518 493 6 Y
port 2 nsew signal output
rlabel locali s 452 51 518 143 6 Y
port 2 nsew signal output
rlabel locali s 284 333 350 493 6 Y
port 2 nsew signal output
rlabel locali s 284 51 350 143 6 Y
port 2 nsew signal output
rlabel locali s 116 333 182 493 6 Y
port 2 nsew signal output
rlabel locali s 116 299 1358 333 6 Y
port 2 nsew signal output
rlabel locali s 116 143 1358 181 6 Y
port 2 nsew signal output
rlabel locali s 116 51 182 143 6 Y
port 2 nsew signal output
rlabel locali s 1392 17 1434 177 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1224 17 1258 109 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1056 17 1090 109 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 888 17 922 109 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 720 17 754 109 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 552 17 586 109 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 384 17 418 109 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 216 17 250 109 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 36 17 82 177 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 0 -17 1472 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1472 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1392 367 1434 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1224 367 1258 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1056 367 1090 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 888 367 922 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 720 367 754 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 552 367 586 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 384 367 418 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 216 367 250 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 40 297 82 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 0 527 1472 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 496 1472 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1472 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2170790
string GDS_START 2159302
<< end >>
