magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 109 403 163 596
rect 293 403 343 596
rect 109 369 343 403
rect 109 310 167 369
rect 109 235 159 310
rect 451 269 551 356
rect 585 290 651 356
rect 109 201 345 235
rect 109 95 159 201
rect 295 95 345 201
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 23 364 73 649
rect 203 437 253 649
rect 387 458 453 649
rect 494 424 560 581
rect 594 458 660 649
rect 700 424 734 581
rect 377 390 734 424
rect 774 405 840 649
rect 377 335 411 390
rect 23 17 73 251
rect 201 269 411 335
rect 700 256 734 390
rect 195 17 261 167
rect 397 17 463 235
rect 499 85 565 235
rect 599 222 734 256
rect 599 119 665 222
rect 701 85 735 188
rect 499 51 735 85
rect 775 17 841 251
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel locali s 585 290 651 356 6 A
port 1 nsew signal input
rlabel locali s 451 269 551 356 6 B
port 2 nsew signal input
rlabel locali s 295 95 345 201 6 X
port 3 nsew signal output
rlabel locali s 293 403 343 596 6 X
port 3 nsew signal output
rlabel locali s 109 403 163 596 6 X
port 3 nsew signal output
rlabel locali s 109 369 343 403 6 X
port 3 nsew signal output
rlabel locali s 109 310 167 369 6 X
port 3 nsew signal output
rlabel locali s 109 235 159 310 6 X
port 3 nsew signal output
rlabel locali s 109 201 345 235 6 X
port 3 nsew signal output
rlabel locali s 109 95 159 201 6 X
port 3 nsew signal output
rlabel metal1 s 0 -49 864 49 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 617 864 715 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3204348
string GDS_START 3196774
<< end >>
