magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 103 333 179 417
rect 291 333 370 417
rect 972 333 1038 417
rect 1150 333 1226 417
rect 103 299 1226 333
rect 22 215 367 255
rect 411 181 447 299
rect 481 215 788 255
rect 834 215 1196 255
rect 1304 215 1602 255
rect 1818 215 2185 255
rect 103 131 746 181
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 18 451 448 493
rect 18 299 69 451
rect 223 367 257 451
rect 414 401 448 451
rect 482 435 558 527
rect 602 401 636 485
rect 670 435 746 527
rect 790 401 840 493
rect 414 367 840 401
rect 878 451 1696 493
rect 878 367 928 451
rect 1082 367 1116 451
rect 1270 367 1304 451
rect 1338 333 1414 417
rect 1458 367 1492 451
rect 1526 333 1602 417
rect 1646 367 1696 451
rect 1734 367 1784 527
rect 1818 333 1894 493
rect 1938 367 1972 527
rect 2006 333 2082 493
rect 1338 299 2082 333
rect 2135 299 2185 527
rect 18 93 69 181
rect 790 147 2185 181
rect 790 93 840 147
rect 18 51 840 93
rect 884 17 918 109
rect 952 51 1028 147
rect 1072 17 1138 109
rect 1182 51 1316 147
rect 1364 17 1398 109
rect 1432 51 1508 147
rect 1552 17 1586 109
rect 1620 51 1768 147
rect 1844 17 1878 109
rect 1912 51 1988 147
rect 2032 17 2075 109
rect 2109 51 2185 147
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
<< metal1 >>
rect 0 561 2208 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 0 496 2208 527
rect 0 17 2208 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
rect 0 -48 2208 -17
<< labels >>
rlabel locali s 1818 215 2185 255 6 A1
port 1 nsew signal input
rlabel locali s 1304 215 1602 255 6 A2
port 2 nsew signal input
rlabel locali s 834 215 1196 255 6 A3
port 3 nsew signal input
rlabel locali s 481 215 788 255 6 B1
port 4 nsew signal input
rlabel locali s 22 215 367 255 6 B2
port 5 nsew signal input
rlabel locali s 1150 333 1226 417 6 Y
port 6 nsew signal output
rlabel locali s 972 333 1038 417 6 Y
port 6 nsew signal output
rlabel locali s 411 181 447 299 6 Y
port 6 nsew signal output
rlabel locali s 291 333 370 417 6 Y
port 6 nsew signal output
rlabel locali s 103 333 179 417 6 Y
port 6 nsew signal output
rlabel locali s 103 299 1226 333 6 Y
port 6 nsew signal output
rlabel locali s 103 131 746 181 6 Y
port 6 nsew signal output
rlabel metal1 s 0 -48 2208 48 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 496 2208 592 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2208 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 608194
string GDS_START 591224
<< end >>
