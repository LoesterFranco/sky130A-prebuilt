magic
tech sky130A
magscale 1 2
timestamp 1601050047
<< nwell >>
rect -38 332 1862 704
<< pwell >>
rect 0 0 1824 49
<< scpmos >>
rect 117 392 147 592
rect 247 392 277 592
rect 354 392 384 560
rect 455 392 485 520
rect 549 392 579 520
rect 656 379 686 547
rect 963 368 993 592
rect 1185 396 1215 564
rect 1336 396 1366 564
rect 1570 373 1600 501
rect 1708 368 1738 592
<< nmoslvt >>
rect 84 134 114 262
rect 250 134 280 262
rect 386 86 416 214
rect 486 130 516 214
rect 620 86 650 214
rect 738 125 768 253
rect 972 74 1002 222
rect 1216 121 1246 249
rect 1352 121 1382 249
rect 1608 84 1638 168
rect 1710 84 1740 232
<< ndiff >>
rect 27 248 84 262
rect 27 214 39 248
rect 73 214 84 248
rect 27 180 84 214
rect 27 146 39 180
rect 73 146 84 180
rect 27 134 84 146
rect 114 134 250 262
rect 280 250 337 262
rect 280 216 291 250
rect 325 216 337 250
rect 280 214 337 216
rect 665 241 738 253
rect 665 214 677 241
rect 280 134 386 214
rect 129 82 235 134
rect 336 86 386 134
rect 416 202 486 214
rect 416 168 427 202
rect 461 168 486 202
rect 416 132 486 168
rect 416 98 427 132
rect 461 130 486 132
rect 516 189 620 214
rect 516 155 536 189
rect 570 155 620 189
rect 516 130 620 155
rect 461 98 471 130
rect 416 86 471 98
rect 531 86 620 130
rect 650 207 677 214
rect 711 207 738 241
rect 650 132 738 207
rect 650 98 677 132
rect 711 125 738 132
rect 768 237 857 253
rect 768 203 813 237
rect 847 203 857 237
rect 768 125 857 203
rect 711 98 723 125
rect 650 86 723 98
rect 129 48 165 82
rect 199 48 235 82
rect 129 36 235 48
rect 917 189 972 222
rect 917 155 927 189
rect 961 155 972 189
rect 917 74 972 155
rect 1002 120 1107 222
rect 1161 177 1216 249
rect 1161 143 1171 177
rect 1205 143 1216 177
rect 1161 121 1216 143
rect 1246 237 1352 249
rect 1246 203 1307 237
rect 1341 203 1352 237
rect 1246 121 1352 203
rect 1382 169 1457 249
rect 1653 220 1710 232
rect 1382 135 1402 169
rect 1436 135 1457 169
rect 1653 186 1665 220
rect 1699 186 1710 220
rect 1653 168 1710 186
rect 1382 121 1457 135
rect 1551 143 1608 168
rect 1002 86 1063 120
rect 1097 86 1107 120
rect 1551 109 1563 143
rect 1597 109 1608 143
rect 1002 74 1107 86
rect 1551 84 1608 109
rect 1638 130 1710 168
rect 1638 96 1665 130
rect 1699 96 1710 130
rect 1638 84 1710 96
rect 1740 220 1797 232
rect 1740 186 1751 220
rect 1785 186 1797 220
rect 1740 130 1797 186
rect 1740 96 1751 130
rect 1785 96 1797 130
rect 1740 84 1797 96
<< pdiff >>
rect 58 580 117 592
rect 58 546 70 580
rect 104 546 117 580
rect 58 502 117 546
rect 58 468 70 502
rect 104 468 117 502
rect 58 392 117 468
rect 147 580 247 592
rect 147 546 170 580
rect 204 546 247 580
rect 147 502 247 546
rect 147 468 170 502
rect 204 468 247 502
rect 147 392 247 468
rect 277 580 332 592
rect 277 546 290 580
rect 324 560 332 580
rect 324 546 354 560
rect 277 510 354 546
rect 277 476 290 510
rect 324 476 354 510
rect 277 438 354 476
rect 277 404 290 438
rect 324 404 354 438
rect 277 392 354 404
rect 384 520 437 560
rect 603 520 656 547
rect 384 508 455 520
rect 384 474 402 508
rect 436 474 455 508
rect 384 438 455 474
rect 384 404 402 438
rect 436 404 455 438
rect 384 392 455 404
rect 485 458 549 520
rect 485 424 502 458
rect 536 424 549 458
rect 485 392 549 424
rect 579 444 656 520
rect 579 410 609 444
rect 643 410 656 444
rect 579 392 656 410
rect 597 379 656 392
rect 686 535 807 547
rect 686 501 745 535
rect 779 501 807 535
rect 686 431 807 501
rect 686 397 745 431
rect 779 397 807 431
rect 686 379 807 397
rect 904 580 963 592
rect 904 546 916 580
rect 950 546 963 580
rect 904 497 963 546
rect 904 463 916 497
rect 950 463 963 497
rect 904 414 963 463
rect 904 380 916 414
rect 950 380 963 414
rect 904 368 963 380
rect 993 580 1052 592
rect 993 546 1006 580
rect 1040 546 1052 580
rect 1649 580 1708 592
rect 993 510 1052 546
rect 993 476 1006 510
rect 1040 476 1052 510
rect 993 440 1052 476
rect 993 406 1006 440
rect 1040 406 1052 440
rect 993 368 1052 406
rect 1109 552 1185 564
rect 1109 518 1121 552
rect 1155 518 1185 552
rect 1109 442 1185 518
rect 1109 408 1121 442
rect 1155 408 1185 442
rect 1109 396 1185 408
rect 1215 531 1336 564
rect 1215 497 1289 531
rect 1323 497 1336 531
rect 1215 442 1336 497
rect 1215 408 1289 442
rect 1323 408 1336 442
rect 1215 396 1336 408
rect 1366 531 1437 564
rect 1366 497 1391 531
rect 1425 497 1437 531
rect 1649 546 1661 580
rect 1695 546 1708 580
rect 1649 510 1708 546
rect 1649 501 1661 510
rect 1366 442 1437 497
rect 1366 408 1391 442
rect 1425 408 1437 442
rect 1366 396 1437 408
rect 1491 489 1570 501
rect 1491 455 1513 489
rect 1547 455 1570 489
rect 1491 373 1570 455
rect 1600 476 1661 501
rect 1695 476 1708 510
rect 1600 440 1708 476
rect 1600 406 1661 440
rect 1695 406 1708 440
rect 1600 373 1708 406
rect 1649 368 1708 373
rect 1738 580 1797 592
rect 1738 546 1751 580
rect 1785 546 1797 580
rect 1738 497 1797 546
rect 1738 463 1751 497
rect 1785 463 1797 497
rect 1738 414 1797 463
rect 1738 380 1751 414
rect 1785 380 1797 414
rect 1738 368 1797 380
<< ndiffc >>
rect 39 214 73 248
rect 39 146 73 180
rect 291 216 325 250
rect 427 168 461 202
rect 427 98 461 132
rect 536 155 570 189
rect 677 207 711 241
rect 677 98 711 132
rect 813 203 847 237
rect 165 48 199 82
rect 927 155 961 189
rect 1171 143 1205 177
rect 1307 203 1341 237
rect 1402 135 1436 169
rect 1665 186 1699 220
rect 1063 86 1097 120
rect 1563 109 1597 143
rect 1665 96 1699 130
rect 1751 186 1785 220
rect 1751 96 1785 130
<< pdiffc >>
rect 70 546 104 580
rect 70 468 104 502
rect 170 546 204 580
rect 170 468 204 502
rect 290 546 324 580
rect 290 476 324 510
rect 290 404 324 438
rect 402 474 436 508
rect 402 404 436 438
rect 502 424 536 458
rect 609 410 643 444
rect 745 501 779 535
rect 745 397 779 431
rect 916 546 950 580
rect 916 463 950 497
rect 916 380 950 414
rect 1006 546 1040 580
rect 1006 476 1040 510
rect 1006 406 1040 440
rect 1121 518 1155 552
rect 1121 408 1155 442
rect 1289 497 1323 531
rect 1289 408 1323 442
rect 1391 497 1425 531
rect 1661 546 1695 580
rect 1391 408 1425 442
rect 1513 455 1547 489
rect 1661 476 1695 510
rect 1661 406 1695 440
rect 1751 546 1785 580
rect 1751 463 1785 497
rect 1751 380 1785 414
<< poly >>
rect 117 592 147 618
rect 247 592 277 618
rect 351 615 889 645
rect 351 575 387 615
rect 354 560 384 575
rect 455 520 485 546
rect 546 535 582 615
rect 656 547 686 573
rect 549 520 579 535
rect 117 377 147 392
rect 247 377 277 392
rect 114 360 150 377
rect 84 344 150 360
rect 244 350 280 377
rect 354 366 384 392
rect 455 377 485 392
rect 84 310 100 344
rect 134 310 150 344
rect 84 294 150 310
rect 192 334 280 350
rect 192 300 208 334
rect 242 300 280 334
rect 84 262 114 294
rect 192 284 280 300
rect 452 318 488 377
rect 549 366 579 392
rect 656 364 686 379
rect 653 318 689 364
rect 738 331 811 347
rect 738 318 761 331
rect 452 297 761 318
rect 795 297 811 331
rect 452 288 811 297
rect 250 262 280 284
rect 386 214 416 240
rect 486 214 516 288
rect 738 281 811 288
rect 859 300 889 615
rect 963 592 993 618
rect 1708 592 1738 618
rect 1185 564 1215 590
rect 1336 564 1366 590
rect 1570 501 1600 527
rect 1185 381 1215 396
rect 1336 381 1366 396
rect 963 353 993 368
rect 1182 364 1218 381
rect 960 336 996 353
rect 1157 348 1246 364
rect 960 320 1050 336
rect 960 300 1000 320
rect 859 286 1000 300
rect 1034 286 1050 320
rect 1157 314 1177 348
rect 1211 314 1246 348
rect 1157 298 1246 314
rect 1333 337 1369 381
rect 1570 358 1600 373
rect 1333 321 1441 337
rect 1333 307 1391 321
rect 738 253 768 281
rect 859 270 1050 286
rect 620 214 650 240
rect 84 108 114 134
rect 250 108 280 134
rect 486 104 516 130
rect 738 99 768 125
rect 386 51 416 86
rect 620 51 650 86
rect 872 51 902 270
rect 972 222 1002 270
rect 1216 249 1246 298
rect 1352 287 1391 307
rect 1425 301 1441 321
rect 1567 301 1603 358
rect 1708 353 1738 368
rect 1705 336 1741 353
rect 1651 320 1741 336
rect 1425 287 1597 301
rect 1352 271 1597 287
rect 1352 249 1382 271
rect 1567 213 1597 271
rect 1651 286 1667 320
rect 1701 306 1741 320
rect 1701 286 1740 306
rect 1651 270 1740 286
rect 1710 232 1740 270
rect 1567 183 1638 213
rect 1608 168 1638 183
rect 1216 95 1246 121
rect 1352 95 1382 121
rect 386 21 902 51
rect 972 48 1002 74
rect 1608 58 1638 84
rect 1710 58 1740 84
<< polycont >>
rect 100 310 134 344
rect 208 300 242 334
rect 761 297 795 331
rect 1000 286 1034 320
rect 1177 314 1211 348
rect 1391 287 1425 321
rect 1667 286 1701 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 17 580 120 596
rect 17 546 70 580
rect 104 546 120 580
rect 17 502 120 546
rect 17 468 70 502
rect 104 468 120 502
rect 17 452 120 468
rect 154 580 220 649
rect 154 546 170 580
rect 204 546 220 580
rect 154 502 220 546
rect 154 468 170 502
rect 204 468 220 502
rect 154 452 220 468
rect 274 581 779 615
rect 274 580 340 581
rect 274 546 290 580
rect 324 546 340 580
rect 745 551 779 581
rect 916 580 950 596
rect 274 510 340 546
rect 274 476 290 510
rect 324 476 340 510
rect 17 260 51 452
rect 274 438 340 476
rect 274 418 290 438
rect 85 404 290 418
rect 324 404 340 438
rect 85 388 340 404
rect 386 513 711 547
rect 386 508 452 513
rect 386 474 402 508
rect 436 474 452 508
rect 386 438 452 474
rect 386 404 402 438
rect 436 404 452 438
rect 386 388 452 404
rect 486 458 552 479
rect 486 424 502 458
rect 536 424 552 458
rect 85 384 325 388
rect 85 344 150 384
rect 85 310 100 344
rect 134 310 150 344
rect 85 294 150 310
rect 192 334 257 350
rect 192 300 208 334
rect 242 300 257 334
rect 17 248 89 260
rect 17 214 39 248
rect 73 214 89 248
rect 192 236 257 300
rect 291 250 325 384
rect 486 286 552 424
rect 593 444 643 479
rect 593 410 609 444
rect 593 375 643 410
rect 17 180 89 214
rect 291 200 325 216
rect 359 252 552 286
rect 17 146 39 180
rect 73 166 89 180
rect 359 166 393 252
rect 518 218 552 252
rect 604 350 643 375
rect 604 316 607 350
rect 641 316 643 350
rect 73 146 393 166
rect 17 132 393 146
rect 427 202 477 218
rect 461 168 477 202
rect 427 132 477 168
rect 17 130 89 132
rect 461 98 477 132
rect 518 189 570 218
rect 518 155 536 189
rect 518 126 570 155
rect 125 82 239 98
rect 125 48 165 82
rect 199 48 239 82
rect 427 92 477 98
rect 604 92 643 316
rect 427 58 643 92
rect 677 241 711 513
rect 745 535 879 551
rect 779 501 879 535
rect 745 431 879 501
rect 779 397 879 431
rect 745 381 879 397
rect 677 132 711 207
rect 745 331 811 347
rect 745 297 761 331
rect 795 297 811 331
rect 745 287 811 297
rect 745 153 779 287
rect 845 253 879 381
rect 813 237 879 253
rect 847 203 879 237
rect 813 187 879 203
rect 916 497 950 546
rect 916 414 950 463
rect 990 580 1040 649
rect 990 546 1006 580
rect 1205 581 1521 615
rect 990 510 1040 546
rect 990 476 1006 510
rect 990 440 1040 476
rect 990 406 1006 440
rect 990 390 1040 406
rect 1081 552 1171 568
rect 1081 518 1121 552
rect 1155 518 1171 552
rect 1081 442 1171 518
rect 1081 408 1121 442
rect 1155 408 1171 442
rect 1081 398 1171 408
rect 1081 390 1125 398
rect 916 226 950 380
rect 984 320 1050 356
rect 984 286 1000 320
rect 1034 286 1050 320
rect 984 270 1050 286
rect 1084 350 1125 390
rect 1205 364 1239 581
rect 1084 316 1087 350
rect 1121 316 1125 350
rect 1084 272 1125 316
rect 1161 348 1239 364
rect 1161 314 1177 348
rect 1211 314 1239 348
rect 1161 306 1239 314
rect 1273 531 1341 547
rect 1273 497 1289 531
rect 1323 497 1341 531
rect 1273 442 1341 497
rect 1273 408 1289 442
rect 1323 408 1341 442
rect 1273 350 1341 408
rect 1375 531 1441 547
rect 1375 497 1391 531
rect 1425 497 1441 531
rect 1375 442 1441 497
rect 1375 408 1391 442
rect 1425 408 1441 442
rect 1487 505 1521 581
rect 1645 580 1711 649
rect 1645 546 1661 580
rect 1695 546 1711 580
rect 1645 510 1711 546
rect 1487 489 1597 505
rect 1487 455 1513 489
rect 1547 455 1597 489
rect 1487 439 1597 455
rect 1375 405 1441 408
rect 1375 371 1529 405
rect 1273 316 1279 350
rect 1313 316 1341 350
rect 1273 310 1341 316
rect 1084 238 1273 272
rect 916 189 961 226
rect 916 155 927 189
rect 916 153 961 155
rect 745 119 961 153
rect 995 177 1205 204
rect 995 170 1171 177
rect 677 85 711 98
rect 995 85 1029 170
rect 1155 143 1171 170
rect 677 51 1029 85
rect 1063 120 1113 136
rect 1097 86 1113 120
rect 125 17 239 48
rect 1063 17 1113 86
rect 1155 85 1205 143
rect 1239 153 1273 238
rect 1307 237 1341 310
rect 1375 321 1441 337
rect 1375 287 1391 321
rect 1425 287 1441 321
rect 1375 236 1441 287
rect 1307 187 1341 203
rect 1377 169 1461 185
rect 1377 153 1402 169
rect 1239 135 1402 153
rect 1436 135 1461 169
rect 1239 119 1461 135
rect 1495 85 1529 371
rect 1155 51 1529 85
rect 1563 172 1597 439
rect 1645 476 1661 510
rect 1695 476 1711 510
rect 1645 440 1711 476
rect 1645 406 1661 440
rect 1695 406 1711 440
rect 1645 390 1711 406
rect 1751 580 1801 596
rect 1785 546 1801 580
rect 1751 497 1801 546
rect 1785 463 1801 497
rect 1751 414 1801 463
rect 1785 380 1801 414
rect 1651 350 1717 356
rect 1651 316 1663 350
rect 1697 320 1717 350
rect 1651 286 1667 316
rect 1701 286 1717 320
rect 1651 270 1717 286
rect 1649 220 1715 236
rect 1649 186 1665 220
rect 1699 186 1715 220
rect 1563 143 1613 172
rect 1597 109 1613 143
rect 1563 80 1613 109
rect 1649 130 1715 186
rect 1649 96 1665 130
rect 1699 96 1715 130
rect 1649 17 1715 96
rect 1751 220 1801 380
rect 1785 186 1801 220
rect 1751 130 1801 186
rect 1785 96 1801 130
rect 1751 80 1801 96
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 607 316 641 350
rect 1087 316 1121 350
rect 1279 316 1313 350
rect 1663 320 1697 350
rect 1663 316 1667 320
rect 1667 316 1697 320
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
<< metal1 >>
rect 0 683 1824 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 0 617 1824 649
rect 595 350 653 356
rect 595 316 607 350
rect 641 347 653 350
rect 1075 350 1133 356
rect 1075 347 1087 350
rect 641 319 1087 347
rect 641 316 653 319
rect 595 310 653 316
rect 1075 316 1087 319
rect 1121 316 1133 350
rect 1075 310 1133 316
rect 1267 350 1325 356
rect 1267 316 1279 350
rect 1313 347 1325 350
rect 1651 350 1709 356
rect 1651 347 1663 350
rect 1313 319 1663 347
rect 1313 316 1325 319
rect 1267 310 1325 316
rect 1651 316 1663 319
rect 1697 316 1709 350
rect 1651 310 1709 316
rect 0 17 1824 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
rect 0 -49 1824 -17
<< labels >>
rlabel comment s 0 0 0 0 4 xor3_1
flabel pwell s 0 0 1824 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 1824 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 1824 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 1824 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 1375 242 1409 276 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 223 242 257 276 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 1759 94 1793 128 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 1759 168 1793 202 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 1759 242 1793 276 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 1759 316 1793 350 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 1759 390 1793 424 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 1759 464 1793 498 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 1759 538 1793 572 0 FreeSans 340 0 0 0 X
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 1824 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 585532
string GDS_START 571620
<< end >>
