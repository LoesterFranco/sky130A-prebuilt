magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 2154 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 89 47 119 177
rect 176 47 206 177
rect 457 47 487 177
rect 551 47 581 177
rect 645 47 675 177
rect 739 47 769 177
rect 823 47 853 177
rect 917 47 947 177
rect 1011 47 1041 177
rect 1115 47 1145 177
rect 1319 47 1349 177
rect 1413 47 1443 177
rect 1507 47 1537 177
rect 1601 47 1631 177
rect 1685 47 1715 177
rect 1779 47 1809 177
rect 1873 47 1903 177
rect 1967 47 1997 177
<< pmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 449 297 485 497
rect 543 297 579 497
rect 637 297 673 497
rect 731 297 767 497
rect 825 297 861 497
rect 919 297 955 497
rect 1013 297 1049 497
rect 1107 297 1143 497
rect 1311 297 1347 497
rect 1405 297 1441 497
rect 1499 297 1535 497
rect 1593 297 1629 497
rect 1687 297 1723 497
rect 1781 297 1817 497
rect 1875 297 1911 497
rect 1969 297 2005 497
<< ndiff >>
rect 27 109 89 177
rect 27 75 35 109
rect 69 75 89 109
rect 27 47 89 75
rect 119 93 176 177
rect 119 59 129 93
rect 163 59 176 93
rect 119 47 176 59
rect 206 93 302 177
rect 206 59 239 93
rect 273 59 302 93
rect 206 47 302 59
rect 395 165 457 177
rect 395 131 403 165
rect 437 131 457 165
rect 395 47 457 131
rect 487 165 551 177
rect 487 131 497 165
rect 531 131 551 165
rect 487 47 551 131
rect 581 97 645 177
rect 581 63 591 97
rect 625 63 645 97
rect 581 47 645 63
rect 675 165 739 177
rect 675 131 685 165
rect 719 131 739 165
rect 675 47 739 131
rect 769 97 823 177
rect 769 63 779 97
rect 813 63 823 97
rect 769 47 823 63
rect 853 165 917 177
rect 853 131 873 165
rect 907 131 917 165
rect 853 47 917 131
rect 947 97 1011 177
rect 947 63 967 97
rect 1001 63 1011 97
rect 947 47 1011 63
rect 1041 165 1115 177
rect 1041 131 1061 165
rect 1095 131 1115 165
rect 1041 47 1115 131
rect 1145 97 1197 177
rect 1145 63 1155 97
rect 1189 63 1197 97
rect 1145 47 1197 63
rect 1251 97 1319 177
rect 1251 63 1269 97
rect 1303 63 1319 97
rect 1251 47 1319 63
rect 1349 165 1413 177
rect 1349 131 1364 165
rect 1398 131 1413 165
rect 1349 47 1413 131
rect 1443 97 1507 177
rect 1443 63 1457 97
rect 1491 63 1507 97
rect 1443 47 1507 63
rect 1537 165 1601 177
rect 1537 131 1552 165
rect 1586 131 1601 165
rect 1537 47 1601 131
rect 1631 124 1685 177
rect 1631 90 1641 124
rect 1675 90 1685 124
rect 1631 47 1685 90
rect 1715 97 1779 177
rect 1715 63 1735 97
rect 1769 63 1779 97
rect 1715 47 1779 63
rect 1809 165 1873 177
rect 1809 131 1826 165
rect 1860 131 1873 165
rect 1809 47 1873 131
rect 1903 97 1967 177
rect 1903 63 1923 97
rect 1957 63 1967 97
rect 1903 47 1967 63
rect 1997 165 2062 177
rect 1997 131 2007 165
rect 2041 131 2062 165
rect 1997 47 2062 131
<< pdiff >>
rect 27 472 81 497
rect 27 438 35 472
rect 69 438 81 472
rect 27 297 81 438
rect 117 489 175 497
rect 117 455 129 489
rect 163 455 175 489
rect 117 297 175 455
rect 211 483 302 497
rect 211 449 223 483
rect 257 449 302 483
rect 211 297 302 449
rect 395 485 449 497
rect 395 451 403 485
rect 437 451 449 485
rect 395 417 449 451
rect 395 383 403 417
rect 437 383 449 417
rect 395 349 449 383
rect 395 315 403 349
rect 437 315 449 349
rect 395 297 449 315
rect 485 477 543 497
rect 485 443 497 477
rect 531 443 543 477
rect 485 374 543 443
rect 485 340 497 374
rect 531 340 543 374
rect 485 297 543 340
rect 579 485 637 497
rect 579 451 591 485
rect 625 451 637 485
rect 579 417 637 451
rect 579 383 591 417
rect 625 383 637 417
rect 579 297 637 383
rect 673 485 731 497
rect 673 451 685 485
rect 719 451 731 485
rect 673 417 731 451
rect 673 383 685 417
rect 719 383 731 417
rect 673 349 731 383
rect 673 315 685 349
rect 719 315 731 349
rect 673 297 731 315
rect 767 485 825 497
rect 767 451 779 485
rect 813 451 825 485
rect 767 417 825 451
rect 767 383 779 417
rect 813 383 825 417
rect 767 297 825 383
rect 861 485 919 497
rect 861 451 873 485
rect 907 451 919 485
rect 861 417 919 451
rect 861 383 873 417
rect 907 383 919 417
rect 861 349 919 383
rect 861 315 873 349
rect 907 315 919 349
rect 861 297 919 315
rect 955 485 1013 497
rect 955 451 967 485
rect 1001 451 1013 485
rect 955 417 1013 451
rect 955 383 967 417
rect 1001 383 1013 417
rect 955 297 1013 383
rect 1049 485 1107 497
rect 1049 451 1061 485
rect 1095 451 1107 485
rect 1049 417 1107 451
rect 1049 383 1061 417
rect 1095 383 1107 417
rect 1049 349 1107 383
rect 1049 315 1061 349
rect 1095 315 1107 349
rect 1049 297 1107 315
rect 1143 485 1311 497
rect 1143 451 1165 485
rect 1199 451 1234 485
rect 1268 451 1311 485
rect 1143 417 1311 451
rect 1143 383 1165 417
rect 1199 383 1234 417
rect 1268 383 1311 417
rect 1143 297 1311 383
rect 1347 485 1405 497
rect 1347 451 1359 485
rect 1393 451 1405 485
rect 1347 417 1405 451
rect 1347 383 1359 417
rect 1393 383 1405 417
rect 1347 349 1405 383
rect 1347 315 1359 349
rect 1393 315 1405 349
rect 1347 297 1405 315
rect 1441 485 1499 497
rect 1441 451 1453 485
rect 1487 451 1499 485
rect 1441 417 1499 451
rect 1441 383 1453 417
rect 1487 383 1499 417
rect 1441 297 1499 383
rect 1535 485 1593 497
rect 1535 451 1547 485
rect 1581 451 1593 485
rect 1535 417 1593 451
rect 1535 383 1547 417
rect 1581 383 1593 417
rect 1535 349 1593 383
rect 1535 315 1547 349
rect 1581 315 1593 349
rect 1535 297 1593 315
rect 1629 485 1687 497
rect 1629 451 1641 485
rect 1675 451 1687 485
rect 1629 417 1687 451
rect 1629 383 1641 417
rect 1675 383 1687 417
rect 1629 297 1687 383
rect 1723 485 1781 497
rect 1723 451 1735 485
rect 1769 451 1781 485
rect 1723 417 1781 451
rect 1723 383 1735 417
rect 1769 383 1781 417
rect 1723 349 1781 383
rect 1723 315 1735 349
rect 1769 315 1781 349
rect 1723 297 1781 315
rect 1817 485 1875 497
rect 1817 451 1829 485
rect 1863 451 1875 485
rect 1817 417 1875 451
rect 1817 383 1829 417
rect 1863 383 1875 417
rect 1817 297 1875 383
rect 1911 485 1969 497
rect 1911 451 1923 485
rect 1957 451 1969 485
rect 1911 417 1969 451
rect 1911 383 1923 417
rect 1957 383 1969 417
rect 1911 349 1969 383
rect 1911 315 1923 349
rect 1957 315 1969 349
rect 1911 297 1969 315
rect 2005 485 2062 497
rect 2005 451 2017 485
rect 2051 451 2062 485
rect 2005 417 2062 451
rect 2005 383 2017 417
rect 2051 383 2062 417
rect 2005 349 2062 383
rect 2005 315 2017 349
rect 2051 315 2062 349
rect 2005 297 2062 315
<< ndiffc >>
rect 35 75 69 109
rect 129 59 163 93
rect 239 59 273 93
rect 403 131 437 165
rect 497 131 531 165
rect 591 63 625 97
rect 685 131 719 165
rect 779 63 813 97
rect 873 131 907 165
rect 967 63 1001 97
rect 1061 131 1095 165
rect 1155 63 1189 97
rect 1269 63 1303 97
rect 1364 131 1398 165
rect 1457 63 1491 97
rect 1552 131 1586 165
rect 1641 90 1675 124
rect 1735 63 1769 97
rect 1826 131 1860 165
rect 1923 63 1957 97
rect 2007 131 2041 165
<< pdiffc >>
rect 35 438 69 472
rect 129 455 163 489
rect 223 449 257 483
rect 403 451 437 485
rect 403 383 437 417
rect 403 315 437 349
rect 497 443 531 477
rect 497 340 531 374
rect 591 451 625 485
rect 591 383 625 417
rect 685 451 719 485
rect 685 383 719 417
rect 685 315 719 349
rect 779 451 813 485
rect 779 383 813 417
rect 873 451 907 485
rect 873 383 907 417
rect 873 315 907 349
rect 967 451 1001 485
rect 967 383 1001 417
rect 1061 451 1095 485
rect 1061 383 1095 417
rect 1061 315 1095 349
rect 1165 451 1199 485
rect 1234 451 1268 485
rect 1165 383 1199 417
rect 1234 383 1268 417
rect 1359 451 1393 485
rect 1359 383 1393 417
rect 1359 315 1393 349
rect 1453 451 1487 485
rect 1453 383 1487 417
rect 1547 451 1581 485
rect 1547 383 1581 417
rect 1547 315 1581 349
rect 1641 451 1675 485
rect 1641 383 1675 417
rect 1735 451 1769 485
rect 1735 383 1769 417
rect 1735 315 1769 349
rect 1829 451 1863 485
rect 1829 383 1863 417
rect 1923 451 1957 485
rect 1923 383 1957 417
rect 1923 315 1957 349
rect 2017 451 2051 485
rect 2017 383 2051 417
rect 2017 315 2051 349
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 449 497 485 523
rect 543 497 579 523
rect 637 497 673 523
rect 731 497 767 523
rect 825 497 861 523
rect 919 497 955 523
rect 1013 497 1049 523
rect 1107 497 1143 523
rect 1311 497 1347 523
rect 1405 497 1441 523
rect 1499 497 1535 523
rect 1593 497 1629 523
rect 1687 497 1723 523
rect 1781 497 1817 523
rect 1875 497 1911 523
rect 1969 497 2005 523
rect 81 282 117 297
rect 175 282 211 297
rect 449 282 485 297
rect 543 282 579 297
rect 637 282 673 297
rect 731 282 767 297
rect 825 282 861 297
rect 919 282 955 297
rect 1013 282 1049 297
rect 1107 282 1143 297
rect 1311 282 1347 297
rect 1405 282 1441 297
rect 1499 282 1535 297
rect 1593 282 1629 297
rect 1687 282 1723 297
rect 1781 282 1817 297
rect 1875 282 1911 297
rect 1969 282 2005 297
rect 79 265 119 282
rect 173 265 213 282
rect 447 265 487 282
rect 21 249 119 265
rect 21 215 32 249
rect 66 215 119 249
rect 21 199 119 215
rect 161 249 215 265
rect 161 215 171 249
rect 205 215 215 249
rect 161 199 215 215
rect 257 259 487 265
rect 541 259 581 282
rect 635 259 675 282
rect 729 259 769 282
rect 257 249 769 259
rect 257 215 267 249
rect 301 215 497 249
rect 531 215 590 249
rect 624 215 769 249
rect 257 205 769 215
rect 257 199 487 205
rect 89 177 119 199
rect 176 177 206 199
rect 457 177 487 199
rect 551 177 581 205
rect 645 177 675 205
rect 739 177 769 205
rect 823 259 863 282
rect 917 259 957 282
rect 1011 259 1051 282
rect 1105 259 1145 282
rect 1309 259 1349 282
rect 1403 259 1443 282
rect 1497 259 1537 282
rect 1591 259 1631 282
rect 823 249 1145 259
rect 823 215 874 249
rect 908 215 966 249
rect 1000 215 1061 249
rect 1095 215 1145 249
rect 823 205 1145 215
rect 1243 249 1631 259
rect 1243 215 1259 249
rect 1293 215 1359 249
rect 1393 215 1453 249
rect 1487 215 1547 249
rect 1581 215 1631 249
rect 1243 205 1631 215
rect 823 177 853 205
rect 917 177 947 205
rect 1011 177 1041 205
rect 1115 177 1145 205
rect 1319 177 1349 205
rect 1413 177 1443 205
rect 1507 177 1537 205
rect 1601 177 1631 205
rect 1685 259 1725 282
rect 1779 259 1819 282
rect 1873 259 1913 282
rect 1967 261 2007 282
rect 1967 259 2068 261
rect 1685 249 2068 259
rect 1685 215 1735 249
rect 1769 215 1829 249
rect 1863 215 1923 249
rect 1957 215 2017 249
rect 2051 215 2068 249
rect 1685 205 2068 215
rect 1685 177 1715 205
rect 1779 177 1809 205
rect 1873 177 1903 205
rect 1967 177 1997 205
rect 89 21 119 47
rect 176 21 206 47
rect 457 21 487 47
rect 551 21 581 47
rect 645 21 675 47
rect 739 21 769 47
rect 823 21 853 47
rect 917 21 947 47
rect 1011 21 1041 47
rect 1115 21 1145 47
rect 1319 21 1349 47
rect 1413 21 1443 47
rect 1507 21 1537 47
rect 1601 21 1631 47
rect 1685 21 1715 47
rect 1779 21 1809 47
rect 1873 21 1903 47
rect 1967 21 1997 47
<< polycont >>
rect 32 215 66 249
rect 171 215 205 249
rect 267 215 301 249
rect 497 215 531 249
rect 590 215 624 249
rect 874 215 908 249
rect 966 215 1000 249
rect 1061 215 1095 249
rect 1259 215 1293 249
rect 1359 215 1393 249
rect 1453 215 1487 249
rect 1547 215 1581 249
rect 1735 215 1769 249
rect 1829 215 1863 249
rect 1923 215 1957 249
rect 2017 215 2051 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 108 489 163 527
rect 17 472 74 488
rect 17 438 35 472
rect 69 438 74 472
rect 108 455 129 489
rect 108 439 163 455
rect 197 483 369 493
rect 197 449 223 483
rect 257 449 369 483
rect 17 396 74 438
rect 197 430 369 449
rect 17 357 301 396
rect 20 249 66 323
rect 20 215 32 249
rect 20 199 66 215
rect 117 249 205 323
rect 117 215 171 249
rect 117 199 205 215
rect 239 249 301 357
rect 239 215 267 249
rect 239 161 301 215
rect 17 127 301 161
rect 335 261 369 430
rect 403 485 437 527
rect 403 417 437 451
rect 403 349 437 383
rect 403 299 437 315
rect 471 477 531 493
rect 471 443 497 477
rect 471 374 531 443
rect 471 340 497 374
rect 565 485 625 527
rect 565 451 591 485
rect 565 417 625 451
rect 565 383 591 417
rect 565 367 625 383
rect 659 485 735 493
rect 659 451 685 485
rect 719 451 735 485
rect 659 417 735 451
rect 659 383 685 417
rect 719 383 735 417
rect 471 333 531 340
rect 659 349 735 383
rect 779 485 813 527
rect 779 417 813 451
rect 779 367 813 383
rect 847 485 923 493
rect 847 451 873 485
rect 907 451 923 485
rect 847 417 923 451
rect 847 383 873 417
rect 907 383 923 417
rect 659 333 685 349
rect 471 315 685 333
rect 719 333 735 349
rect 847 349 923 383
rect 967 485 1001 527
rect 967 417 1001 451
rect 967 367 1001 383
rect 1035 485 1111 493
rect 1035 451 1061 485
rect 1095 451 1111 485
rect 1035 417 1111 451
rect 1035 383 1061 417
rect 1095 383 1111 417
rect 847 333 873 349
rect 719 315 873 333
rect 907 333 923 349
rect 1035 349 1111 383
rect 1165 485 1293 527
rect 1199 451 1234 485
rect 1268 451 1293 485
rect 1165 417 1293 451
rect 1199 383 1234 417
rect 1268 383 1293 417
rect 1165 367 1293 383
rect 1333 485 1409 493
rect 1333 451 1359 485
rect 1393 451 1409 485
rect 1333 417 1409 451
rect 1333 383 1359 417
rect 1393 383 1409 417
rect 1035 333 1061 349
rect 907 315 1061 333
rect 1095 333 1111 349
rect 1333 349 1409 383
rect 1453 485 1487 527
rect 1453 417 1487 451
rect 1453 367 1487 383
rect 1521 485 1597 493
rect 1521 451 1547 485
rect 1581 451 1597 485
rect 1521 417 1597 451
rect 1521 383 1547 417
rect 1581 383 1597 417
rect 1333 333 1359 349
rect 1095 315 1359 333
rect 1393 333 1409 349
rect 1521 349 1597 383
rect 1641 485 1675 527
rect 1641 417 1675 451
rect 1641 367 1675 383
rect 1709 485 1785 493
rect 1709 451 1735 485
rect 1769 451 1785 485
rect 1709 417 1785 451
rect 1709 383 1735 417
rect 1769 383 1785 417
rect 1521 333 1547 349
rect 1393 315 1547 333
rect 1581 333 1597 349
rect 1709 349 1785 383
rect 1829 485 1863 527
rect 1829 417 1863 451
rect 1829 367 1863 383
rect 1897 485 1973 493
rect 1897 451 1923 485
rect 1957 451 1973 485
rect 1897 417 1973 451
rect 1897 383 1923 417
rect 1957 383 1973 417
rect 1709 333 1735 349
rect 1581 315 1735 333
rect 1769 333 1785 349
rect 1897 349 1973 383
rect 1897 333 1923 349
rect 1769 315 1923 333
rect 1957 315 1973 349
rect 471 289 1973 315
rect 2017 485 2072 527
rect 2051 451 2072 485
rect 2017 417 2072 451
rect 2051 383 2072 417
rect 2017 349 2072 383
rect 2051 315 2072 349
rect 2017 289 2072 315
rect 335 255 405 261
rect 335 221 359 255
rect 393 221 405 255
rect 335 215 405 221
rect 471 215 497 249
rect 531 215 590 249
rect 624 215 640 249
rect 17 109 69 127
rect 17 75 35 109
rect 335 93 369 215
rect 733 181 803 289
rect 837 221 866 255
rect 900 249 1111 255
rect 837 215 874 221
rect 908 215 966 249
rect 1000 215 1061 249
rect 1095 215 1111 249
rect 1209 249 1597 255
rect 1209 215 1259 249
rect 1293 215 1359 249
rect 1393 215 1453 249
rect 1487 215 1547 249
rect 1581 215 1597 249
rect 1679 249 2068 255
rect 1679 215 1735 249
rect 1769 215 1829 249
rect 1863 215 1923 249
rect 1957 215 2017 249
rect 2051 215 2068 249
rect 17 51 69 75
rect 103 59 129 93
rect 163 59 179 93
rect 103 17 179 59
rect 223 59 239 93
rect 273 59 369 93
rect 223 51 369 59
rect 403 165 437 181
rect 471 165 803 181
rect 471 131 497 165
rect 531 131 685 165
rect 719 131 803 165
rect 847 165 1602 181
rect 847 131 873 165
rect 907 131 1061 165
rect 1095 131 1364 165
rect 1398 131 1552 165
rect 1586 131 1602 165
rect 1641 131 1826 165
rect 1860 131 2007 165
rect 2041 131 2057 165
rect 403 97 437 131
rect 1641 124 1675 131
rect 403 63 591 97
rect 625 63 779 97
rect 813 63 967 97
rect 1001 63 1155 97
rect 1189 63 1205 97
rect 403 51 1205 63
rect 1253 63 1269 97
rect 1303 63 1457 97
rect 1491 90 1641 97
rect 1491 63 1675 90
rect 1253 51 1675 63
rect 1719 63 1735 97
rect 1769 63 1785 97
rect 1719 17 1785 63
rect 1907 63 1923 97
rect 1957 63 1973 97
rect 1907 17 1973 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 359 221 393 255
rect 866 249 900 255
rect 866 221 874 249
rect 874 221 900 249
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
<< metal1 >>
rect 0 561 2116 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 0 496 2116 527
rect 347 255 405 261
rect 347 221 359 255
rect 393 252 405 255
rect 847 255 915 261
rect 847 252 866 255
rect 393 224 866 252
rect 393 221 405 224
rect 347 215 405 221
rect 847 221 866 224
rect 900 221 915 255
rect 847 215 915 221
rect 0 17 2116 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
rect 0 -48 2116 -17
<< labels >>
flabel corelocali s 132 221 166 255 0 FreeSans 200 0 0 0 B_N
port 2 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 200 0 0 0 A_N
port 1 nsew
flabel corelocali s 1209 221 1243 255 0 FreeSans 200 0 0 0 C
port 3 nsew
flabel corelocali s 757 153 791 187 0 FreeSans 200 0 0 0 Y
port 9 nsew
flabel corelocali s 757 289 791 323 0 FreeSans 200 0 0 0 Y
port 9 nsew
flabel corelocali s 1301 221 1335 255 0 FreeSans 200 0 0 0 C
port 3 nsew
flabel corelocali s 1403 221 1437 255 0 FreeSans 200 0 0 0 C
port 3 nsew
flabel corelocali s 1505 221 1539 255 0 FreeSans 200 0 0 0 C
port 3 nsew
flabel corelocali s 1719 221 1753 255 0 FreeSans 200 0 0 0 D
port 4 nsew
flabel corelocali s 1923 221 1957 255 0 FreeSans 200 0 0 0 D
port 4 nsew
flabel corelocali s 2025 221 2059 255 0 FreeSans 200 0 0 0 D
port 4 nsew
flabel corelocali s 1821 221 1855 255 0 FreeSans 200 0 0 0 D
port 4 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
rlabel comment s 0 0 0 0 4 nand4bb_4
<< properties >>
string FIXED_BBOX 0 0 2116 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2380958
string GDS_START 2365442
<< end >>
