magic
tech sky130A
magscale 1 2
timestamp 1604502729
<< locali >>
rect 21 236 87 310
rect 189 270 263 356
rect 297 270 363 356
rect 405 270 471 578
rect 666 378 732 596
rect 505 270 585 356
rect 666 344 839 378
rect 793 210 839 344
rect 687 162 839 210
rect 687 70 737 162
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 45 424 121 572
rect 155 458 221 649
rect 267 424 333 596
rect 45 390 333 424
rect 45 364 155 390
rect 121 236 155 364
rect 549 390 615 649
rect 766 412 832 649
rect 619 244 702 310
rect 619 236 653 244
rect 121 202 653 236
rect 41 70 155 202
rect 236 134 532 168
rect 236 70 302 134
rect 338 17 430 100
rect 466 70 532 134
rect 566 17 632 168
rect 771 17 841 120
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel locali s 505 270 585 356 6 A1
port 1 nsew signal input
rlabel locali s 405 270 471 578 6 A2
port 2 nsew signal input
rlabel locali s 297 270 363 356 6 A3
port 3 nsew signal input
rlabel locali s 189 270 263 356 6 B1
port 4 nsew signal input
rlabel locali s 21 236 87 310 6 C1
port 5 nsew signal input
rlabel locali s 793 210 839 344 6 X
port 6 nsew signal output
rlabel locali s 687 162 839 210 6 X
port 6 nsew signal output
rlabel locali s 687 70 737 162 6 X
port 6 nsew signal output
rlabel locali s 666 378 732 596 6 X
port 6 nsew signal output
rlabel locali s 666 344 839 378 6 X
port 6 nsew signal output
rlabel metal1 s 0 -49 864 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 617 864 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1332132
string GDS_START 1324156
<< end >>
