magic
tech sky130A
magscale 1 2
timestamp 1604502741
<< locali >>
rect 123 424 189 547
rect 313 424 379 547
rect 25 390 379 424
rect 25 236 71 390
rect 105 270 375 356
rect 487 270 757 356
rect 793 270 1319 356
rect 1409 260 1703 326
rect 1561 236 1703 260
rect 25 226 918 236
rect 25 202 1514 226
rect 123 70 348 202
rect 482 70 718 202
rect 852 192 1572 202
rect 852 70 918 192
rect 1448 68 1572 192
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 23 581 453 615
rect 23 458 89 581
rect 229 458 279 581
rect 419 424 453 581
rect 493 581 1215 615
rect 493 458 559 581
rect 594 424 638 547
rect 673 458 739 581
rect 779 424 829 547
rect 419 390 829 424
rect 875 424 925 547
rect 965 460 1031 581
rect 1068 424 1112 547
rect 1149 460 1215 581
rect 1251 424 1305 596
rect 1339 458 1405 649
rect 1439 424 1505 596
rect 1539 458 1605 649
rect 1639 424 1705 596
rect 875 390 1705 424
rect 419 364 453 390
rect 1639 364 1705 390
rect 23 17 89 168
rect 382 17 448 168
rect 752 17 818 168
rect 952 17 1414 158
rect 1606 17 1672 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
<< metal1 >>
rect 0 683 1728 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 0 617 1728 649
rect 0 17 1728 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
rect 0 -49 1728 -17
<< labels >>
rlabel locali s 1561 236 1703 260 6 A
port 1 nsew signal input
rlabel locali s 1409 260 1703 326 6 A
port 1 nsew signal input
rlabel locali s 793 270 1319 356 6 B
port 2 nsew signal input
rlabel locali s 487 270 757 356 6 C
port 3 nsew signal input
rlabel locali s 105 270 375 356 6 D
port 4 nsew signal input
rlabel locali s 1448 68 1572 192 6 Y
port 5 nsew signal output
rlabel locali s 852 192 1572 202 6 Y
port 5 nsew signal output
rlabel locali s 852 70 918 192 6 Y
port 5 nsew signal output
rlabel locali s 482 70 718 202 6 Y
port 5 nsew signal output
rlabel locali s 313 424 379 547 6 Y
port 5 nsew signal output
rlabel locali s 123 424 189 547 6 Y
port 5 nsew signal output
rlabel locali s 123 70 348 202 6 Y
port 5 nsew signal output
rlabel locali s 25 390 379 424 6 Y
port 5 nsew signal output
rlabel locali s 25 236 71 390 6 Y
port 5 nsew signal output
rlabel locali s 25 226 918 236 6 Y
port 5 nsew signal output
rlabel locali s 25 202 1514 226 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -49 1728 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 1728 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1728 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1626040
string GDS_START 1612554
<< end >>
