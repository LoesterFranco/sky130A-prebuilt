magic
tech sky130A
magscale 1 2
timestamp 1601050058
<< locali >>
rect 28 195 98 325
rect 293 397 346 493
rect 297 214 346 397
rect 573 357 624 493
rect 547 271 624 357
rect 804 142 879 340
rect 804 57 855 142
rect 1301 187 1407 209
rect 1301 153 1373 187
rect 2505 416 2565 493
rect 1905 221 1938 255
rect 1972 221 2023 255
rect 1905 213 2023 221
rect 1965 187 2023 213
rect 1965 153 1989 187
rect 1965 127 2023 153
rect 2315 53 2385 339
rect 2487 307 2565 416
rect 2531 165 2565 307
rect 2489 62 2565 165
<< viali >>
rect 1373 153 1407 187
rect 1938 221 1972 255
rect 1989 153 2023 187
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2668 561
rect 18 393 69 493
rect 106 427 172 527
rect 18 359 173 393
rect 132 265 173 359
rect 207 380 241 493
rect 380 411 430 480
rect 207 346 263 380
rect 132 199 195 265
rect 132 161 167 199
rect 19 127 167 161
rect 229 135 263 346
rect 396 291 430 411
rect 464 408 498 527
rect 692 421 726 493
rect 860 455 926 527
rect 981 437 1055 487
rect 981 421 1015 437
rect 1094 427 1167 493
rect 396 252 494 291
rect 658 387 1015 421
rect 411 237 494 252
rect 658 237 692 387
rect 411 199 617 237
rect 411 180 445 199
rect 19 69 69 127
rect 103 17 169 93
rect 203 69 263 135
rect 307 146 445 180
rect 307 79 341 146
rect 375 17 441 112
rect 479 17 545 165
rect 583 85 617 199
rect 651 203 692 237
rect 651 135 685 203
rect 736 85 770 337
rect 583 51 770 85
rect 913 179 947 387
rect 1049 315 1099 391
rect 981 213 1015 279
rect 1065 207 1099 315
rect 1133 277 1167 427
rect 1201 421 1235 475
rect 1282 471 1348 527
rect 1399 421 1433 475
rect 1475 435 1549 527
rect 1201 387 1433 421
rect 1594 401 1628 493
rect 1664 425 1838 493
rect 1872 439 1922 527
rect 1803 423 1838 425
rect 1803 407 1842 423
rect 1491 367 1628 401
rect 1662 387 1768 391
rect 1491 353 1543 367
rect 1257 319 1543 353
rect 1662 333 1774 387
rect 1133 243 1475 277
rect 913 143 1029 179
rect 889 17 955 108
rect 995 101 1029 143
rect 1065 141 1195 207
rect 995 67 1063 101
rect 1233 95 1267 243
rect 1441 201 1475 243
rect 1509 167 1543 319
rect 1097 61 1267 95
rect 1383 17 1449 109
rect 1491 89 1543 167
rect 1577 331 1774 333
rect 1808 349 1842 407
rect 1956 417 1990 475
rect 2024 451 2090 527
rect 1956 383 2109 417
rect 1577 299 1704 331
rect 1808 315 2041 349
rect 1577 141 1619 299
rect 1808 297 1842 315
rect 1681 184 1715 265
rect 1749 263 1842 297
rect 2075 265 2109 383
rect 2143 407 2178 493
rect 2218 441 2284 527
rect 2405 451 2471 527
rect 2310 407 2453 417
rect 2143 373 2453 407
rect 2143 359 2281 373
rect 1749 107 1783 263
rect 2075 259 2212 265
rect 1825 173 1859 229
rect 1825 139 1931 173
rect 1491 55 1557 89
rect 1601 51 1783 107
rect 1817 17 1851 105
rect 1897 93 1931 139
rect 2069 211 2212 259
rect 2069 93 2103 211
rect 2246 177 2281 359
rect 1897 59 2103 93
rect 2143 143 2281 177
rect 2143 69 2177 143
rect 2218 17 2273 109
rect 2419 265 2453 373
rect 2419 199 2497 265
rect 2599 299 2649 527
rect 2421 17 2455 165
rect 2599 17 2633 186
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2668 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
<< metal1 >>
rect 0 561 2668 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2668 561
rect 0 496 2668 527
rect 1926 255 1984 261
rect 1926 221 1938 255
rect 1972 221 1984 255
rect 1926 193 1984 221
rect 1289 187 1419 193
rect 1289 153 1373 187
rect 1407 184 1419 187
rect 1926 187 2035 193
rect 1926 184 1989 187
rect 1407 156 1989 184
rect 1407 153 1419 156
rect 1289 147 1419 153
rect 1977 153 1989 156
rect 2023 153 2035 187
rect 1977 147 2035 153
rect 0 17 2668 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2668 17
rect 0 -48 2668 -17
<< obsm1 >>
rect 194 388 254 397
rect 1053 388 1111 397
rect 1677 388 1735 397
rect 194 360 1735 388
rect 194 351 254 360
rect 1053 351 1111 360
rect 1677 351 1735 360
rect 149 252 207 261
rect 969 252 1027 261
rect 1669 252 1727 261
rect 149 224 1727 252
rect 149 215 207 224
rect 969 215 1027 224
rect 1669 215 1727 224
<< labels >>
rlabel locali s 573 357 624 493 6 D
port 1 nsew signal input
rlabel locali s 547 271 624 357 6 D
port 1 nsew signal input
rlabel locali s 2315 53 2385 339 6 Q
port 2 nsew signal output
rlabel locali s 2531 165 2565 307 6 Q_N
port 3 nsew signal output
rlabel locali s 2505 416 2565 493 6 Q_N
port 3 nsew signal output
rlabel locali s 2489 62 2565 165 6 Q_N
port 3 nsew signal output
rlabel locali s 2487 307 2565 416 6 Q_N
port 3 nsew signal output
rlabel viali s 1373 153 1407 187 6 RESET_B
port 4 nsew signal input
rlabel locali s 1301 153 1407 209 6 RESET_B
port 4 nsew signal input
rlabel viali s 1989 153 2023 187 6 RESET_B
port 4 nsew signal input
rlabel viali s 1938 221 1972 255 6 RESET_B
port 4 nsew signal input
rlabel locali s 1965 127 2023 213 6 RESET_B
port 4 nsew signal input
rlabel locali s 1905 213 2023 255 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 1977 147 2035 156 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 1926 193 1984 261 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 1926 184 2035 193 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 1289 184 1419 193 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 1289 156 2035 184 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 1289 147 1419 156 6 RESET_B
port 4 nsew signal input
rlabel locali s 804 142 879 340 6 SCD
port 5 nsew signal input
rlabel locali s 804 57 855 142 6 SCD
port 5 nsew signal input
rlabel locali s 297 214 346 397 6 SCE
port 6 nsew signal input
rlabel locali s 293 397 346 493 6 SCE
port 6 nsew signal input
rlabel locali s 28 195 98 325 6 CLK
port 7 nsew clock input
rlabel metal1 s 0 -48 2668 48 8 VGND
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 496 2668 592 6 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2668 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 197554
string GDS_START 176912
<< end >>
