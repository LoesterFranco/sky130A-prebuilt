magic
tech sky130A
magscale 1 2
timestamp 1601050056
<< nwell >>
rect -38 332 1478 704
<< pwell >>
rect 0 0 1440 49
<< scpmos >>
rect 84 368 120 592
rect 174 368 210 592
rect 264 368 300 592
rect 354 368 390 592
rect 444 368 480 592
rect 534 368 570 592
rect 624 368 660 592
rect 724 368 760 592
rect 936 368 972 592
rect 1029 368 1065 592
rect 1231 424 1267 592
rect 1321 424 1357 592
<< nmoslvt >>
rect 84 74 114 222
rect 180 74 210 222
rect 266 74 296 222
rect 352 74 382 222
rect 438 74 468 222
rect 524 74 554 222
rect 610 74 640 222
rect 728 74 758 222
rect 828 74 858 222
rect 914 74 944 222
rect 1014 74 1044 222
rect 1114 74 1144 222
rect 1326 104 1356 252
<< ndiff >>
rect 1269 240 1326 252
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 152 180 222
rect 114 118 125 152
rect 159 118 180 152
rect 114 74 180 118
rect 210 210 266 222
rect 210 176 221 210
rect 255 176 266 210
rect 210 120 266 176
rect 210 86 221 120
rect 255 86 266 120
rect 210 74 266 86
rect 296 152 352 222
rect 296 118 307 152
rect 341 118 352 152
rect 296 74 352 118
rect 382 210 438 222
rect 382 176 393 210
rect 427 176 438 210
rect 382 120 438 176
rect 382 86 393 120
rect 427 86 438 120
rect 382 74 438 86
rect 468 152 524 222
rect 468 118 479 152
rect 513 118 524 152
rect 468 74 524 118
rect 554 210 610 222
rect 554 176 565 210
rect 599 176 610 210
rect 554 120 610 176
rect 554 86 565 120
rect 599 86 610 120
rect 554 74 610 86
rect 640 84 728 222
rect 640 74 667 84
rect 655 50 667 74
rect 701 74 728 84
rect 758 136 828 222
rect 758 102 769 136
rect 803 102 828 136
rect 758 74 828 102
rect 858 181 914 222
rect 858 147 869 181
rect 903 147 914 181
rect 858 74 914 147
rect 944 144 1014 222
rect 944 110 969 144
rect 1003 110 1014 144
rect 944 74 1014 110
rect 1044 189 1114 222
rect 1044 155 1069 189
rect 1103 155 1114 189
rect 1044 74 1114 155
rect 1144 188 1215 222
rect 1144 154 1169 188
rect 1203 154 1215 188
rect 1144 120 1215 154
rect 1144 86 1169 120
rect 1203 86 1215 120
rect 1269 206 1281 240
rect 1315 206 1326 240
rect 1269 150 1326 206
rect 1269 116 1281 150
rect 1315 116 1326 150
rect 1269 104 1326 116
rect 1356 240 1413 252
rect 1356 206 1367 240
rect 1401 206 1413 240
rect 1356 150 1413 206
rect 1356 116 1367 150
rect 1401 116 1413 150
rect 1356 104 1413 116
rect 1144 74 1215 86
rect 701 50 713 74
rect 655 38 713 50
<< pdiff >>
rect 28 580 84 592
rect 28 546 40 580
rect 74 546 84 580
rect 28 505 84 546
rect 28 471 40 505
rect 74 471 84 505
rect 28 424 84 471
rect 28 390 40 424
rect 74 390 84 424
rect 28 368 84 390
rect 120 580 174 592
rect 120 546 130 580
rect 164 546 174 580
rect 120 508 174 546
rect 120 474 130 508
rect 164 474 174 508
rect 120 368 174 474
rect 210 580 264 592
rect 210 546 220 580
rect 254 546 264 580
rect 210 505 264 546
rect 210 471 220 505
rect 254 471 264 505
rect 210 424 264 471
rect 210 390 220 424
rect 254 390 264 424
rect 210 368 264 390
rect 300 580 354 592
rect 300 546 310 580
rect 344 546 354 580
rect 300 508 354 546
rect 300 474 310 508
rect 344 474 354 508
rect 300 368 354 474
rect 390 580 444 592
rect 390 546 400 580
rect 434 546 444 580
rect 390 497 444 546
rect 390 463 400 497
rect 434 463 444 497
rect 390 414 444 463
rect 390 380 400 414
rect 434 380 444 414
rect 390 368 444 380
rect 480 531 534 592
rect 480 497 490 531
rect 524 497 534 531
rect 480 424 534 497
rect 480 390 490 424
rect 524 390 534 424
rect 480 368 534 390
rect 570 580 624 592
rect 570 546 580 580
rect 614 546 624 580
rect 570 508 624 546
rect 570 474 580 508
rect 614 474 624 508
rect 570 368 624 474
rect 660 531 724 592
rect 660 497 680 531
rect 714 497 724 531
rect 660 424 724 497
rect 660 390 680 424
rect 714 390 724 424
rect 660 368 724 390
rect 760 580 826 592
rect 760 546 780 580
rect 814 546 826 580
rect 760 492 826 546
rect 760 458 780 492
rect 814 458 826 492
rect 760 368 826 458
rect 880 580 936 592
rect 880 546 892 580
rect 926 546 936 580
rect 880 500 936 546
rect 880 466 892 500
rect 926 466 936 500
rect 880 420 936 466
rect 880 386 892 420
rect 926 386 936 420
rect 880 368 936 386
rect 972 580 1029 592
rect 972 546 982 580
rect 1016 546 1029 580
rect 972 488 1029 546
rect 972 454 982 488
rect 1016 454 1029 488
rect 972 368 1029 454
rect 1065 580 1121 592
rect 1065 546 1075 580
rect 1109 546 1121 580
rect 1065 500 1121 546
rect 1065 466 1075 500
rect 1109 466 1121 500
rect 1065 420 1121 466
rect 1175 580 1231 592
rect 1175 546 1187 580
rect 1221 546 1231 580
rect 1175 508 1231 546
rect 1175 474 1187 508
rect 1221 474 1231 508
rect 1175 424 1231 474
rect 1267 580 1321 592
rect 1267 546 1277 580
rect 1311 546 1321 580
rect 1267 470 1321 546
rect 1267 436 1277 470
rect 1311 436 1321 470
rect 1267 424 1321 436
rect 1357 580 1413 592
rect 1357 546 1367 580
rect 1401 546 1413 580
rect 1357 470 1413 546
rect 1357 436 1367 470
rect 1401 436 1413 470
rect 1357 424 1413 436
rect 1065 386 1075 420
rect 1109 386 1121 420
rect 1065 368 1121 386
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 125 118 159 152
rect 221 176 255 210
rect 221 86 255 120
rect 307 118 341 152
rect 393 176 427 210
rect 393 86 427 120
rect 479 118 513 152
rect 565 176 599 210
rect 565 86 599 120
rect 667 50 701 84
rect 769 102 803 136
rect 869 147 903 181
rect 969 110 1003 144
rect 1069 155 1103 189
rect 1169 154 1203 188
rect 1169 86 1203 120
rect 1281 206 1315 240
rect 1281 116 1315 150
rect 1367 206 1401 240
rect 1367 116 1401 150
<< pdiffc >>
rect 40 546 74 580
rect 40 471 74 505
rect 40 390 74 424
rect 130 546 164 580
rect 130 474 164 508
rect 220 546 254 580
rect 220 471 254 505
rect 220 390 254 424
rect 310 546 344 580
rect 310 474 344 508
rect 400 546 434 580
rect 400 463 434 497
rect 400 380 434 414
rect 490 497 524 531
rect 490 390 524 424
rect 580 546 614 580
rect 580 474 614 508
rect 680 497 714 531
rect 680 390 714 424
rect 780 546 814 580
rect 780 458 814 492
rect 892 546 926 580
rect 892 466 926 500
rect 892 386 926 420
rect 982 546 1016 580
rect 982 454 1016 488
rect 1075 546 1109 580
rect 1075 466 1109 500
rect 1187 546 1221 580
rect 1187 474 1221 508
rect 1277 546 1311 580
rect 1277 436 1311 470
rect 1367 546 1401 580
rect 1367 436 1401 470
rect 1075 386 1109 420
<< poly >>
rect 84 592 120 618
rect 174 592 210 618
rect 264 592 300 618
rect 354 592 390 618
rect 444 592 480 618
rect 534 592 570 618
rect 624 592 660 618
rect 724 592 760 618
rect 936 592 972 618
rect 1029 592 1065 618
rect 1231 592 1267 618
rect 1321 592 1357 618
rect 84 336 120 368
rect 174 336 210 368
rect 264 336 300 368
rect 84 320 300 336
rect 84 286 100 320
rect 134 286 168 320
rect 202 286 236 320
rect 270 300 300 320
rect 354 300 390 368
rect 444 300 480 368
rect 534 336 570 368
rect 624 336 660 368
rect 724 336 760 368
rect 936 336 972 368
rect 1029 336 1065 368
rect 1231 356 1267 424
rect 1321 356 1357 424
rect 1237 340 1357 356
rect 524 320 760 336
rect 524 300 540 320
rect 270 286 390 300
rect 84 270 390 286
rect 438 286 540 300
rect 574 286 608 320
rect 642 286 676 320
rect 710 300 760 320
rect 828 320 1144 336
rect 710 286 758 300
rect 438 270 758 286
rect 84 222 114 270
rect 180 222 210 270
rect 266 222 296 270
rect 352 222 382 270
rect 438 222 468 270
rect 524 222 554 270
rect 610 222 640 270
rect 728 222 758 270
rect 828 286 890 320
rect 924 286 958 320
rect 992 286 1026 320
rect 1060 286 1094 320
rect 1128 286 1144 320
rect 1237 306 1289 340
rect 1323 306 1357 340
rect 1237 290 1357 306
rect 828 270 1144 286
rect 828 222 858 270
rect 914 222 944 270
rect 1014 222 1044 270
rect 1114 222 1144 270
rect 1326 252 1356 290
rect 84 48 114 74
rect 180 48 210 74
rect 266 48 296 74
rect 352 48 382 74
rect 438 48 468 74
rect 524 48 554 74
rect 610 48 640 74
rect 1326 78 1356 104
rect 728 48 758 74
rect 828 48 858 74
rect 914 48 944 74
rect 1014 48 1044 74
rect 1114 48 1144 74
<< polycont >>
rect 100 286 134 320
rect 168 286 202 320
rect 236 286 270 320
rect 540 286 574 320
rect 608 286 642 320
rect 676 286 710 320
rect 890 286 924 320
rect 958 286 992 320
rect 1026 286 1060 320
rect 1094 286 1128 320
rect 1289 306 1323 340
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 24 580 74 596
rect 24 546 40 580
rect 24 505 74 546
rect 24 471 40 505
rect 24 424 74 471
rect 114 580 164 649
rect 114 546 130 580
rect 114 508 164 546
rect 114 474 130 508
rect 114 458 164 474
rect 204 580 254 596
rect 204 546 220 580
rect 204 505 254 546
rect 204 471 220 505
rect 204 424 254 471
rect 294 580 360 649
rect 294 546 310 580
rect 344 546 360 580
rect 294 508 360 546
rect 294 474 310 508
rect 344 474 360 508
rect 294 458 360 474
rect 400 581 830 615
rect 400 580 434 581
rect 564 580 630 581
rect 400 497 434 546
rect 400 424 434 463
rect 24 390 40 424
rect 74 390 220 424
rect 254 414 434 424
rect 254 390 400 414
rect 474 531 524 547
rect 474 497 490 531
rect 474 424 524 497
rect 564 546 580 580
rect 614 546 630 580
rect 764 580 830 581
rect 564 508 630 546
rect 564 474 580 508
rect 614 474 630 508
rect 564 458 630 474
rect 664 531 730 547
rect 664 497 680 531
rect 714 497 730 531
rect 664 424 730 497
rect 764 546 780 580
rect 814 546 830 580
rect 764 492 830 546
rect 764 458 780 492
rect 814 458 830 492
rect 876 580 942 596
rect 876 546 892 580
rect 926 546 942 580
rect 876 500 942 546
rect 876 466 892 500
rect 926 466 942 500
rect 876 424 942 466
rect 982 580 1016 649
rect 982 488 1016 546
rect 982 438 1016 454
rect 1059 580 1125 596
rect 1059 546 1075 580
rect 1109 546 1125 580
rect 1059 500 1125 546
rect 1059 466 1075 500
rect 1109 466 1125 500
rect 474 390 490 424
rect 524 390 680 424
rect 714 420 942 424
rect 714 390 892 420
rect 400 364 434 380
rect 25 320 359 356
rect 25 286 100 320
rect 134 286 168 320
rect 202 286 236 320
rect 270 286 359 320
rect 25 270 359 286
rect 505 320 743 356
rect 505 286 540 320
rect 574 286 608 320
rect 642 286 676 320
rect 710 286 743 320
rect 505 270 743 286
rect 793 236 839 390
rect 876 386 892 390
rect 926 404 942 420
rect 1059 420 1125 466
rect 1171 580 1221 649
rect 1171 546 1187 580
rect 1171 508 1221 546
rect 1171 474 1187 508
rect 1171 458 1221 474
rect 1261 580 1311 596
rect 1261 546 1277 580
rect 1261 470 1311 546
rect 1261 436 1277 470
rect 1261 424 1311 436
rect 1059 404 1075 420
rect 926 386 1075 404
rect 1109 386 1125 420
rect 876 370 1125 386
rect 1159 390 1311 424
rect 1351 580 1417 649
rect 1351 546 1367 580
rect 1401 546 1417 580
rect 1351 470 1417 546
rect 1351 436 1367 470
rect 1401 436 1417 470
rect 1351 420 1417 436
rect 1159 336 1193 390
rect 874 320 1193 336
rect 874 286 890 320
rect 924 286 958 320
rect 992 286 1026 320
rect 1060 286 1094 320
rect 1128 286 1193 320
rect 1273 340 1415 356
rect 1273 306 1289 340
rect 1323 306 1415 340
rect 1273 290 1415 306
rect 874 270 1193 286
rect 1159 256 1193 270
rect 1159 240 1315 256
rect 23 210 615 236
rect 23 176 39 210
rect 73 202 221 210
rect 23 120 73 176
rect 255 202 393 210
rect 23 86 39 120
rect 23 70 73 86
rect 109 152 175 168
rect 109 118 125 152
rect 159 118 175 152
rect 109 17 175 118
rect 221 120 255 176
rect 427 202 565 210
rect 221 70 255 86
rect 291 152 357 168
rect 291 118 307 152
rect 341 118 357 152
rect 291 17 357 118
rect 393 120 427 176
rect 599 176 615 210
rect 793 202 1119 236
rect 1159 222 1281 240
rect 565 168 615 176
rect 853 181 919 202
rect 393 70 427 86
rect 463 152 529 168
rect 463 118 479 152
rect 513 118 529 152
rect 463 17 529 118
rect 565 136 819 168
rect 565 134 769 136
rect 565 120 615 134
rect 599 86 615 120
rect 753 102 769 134
rect 803 102 819 136
rect 853 147 869 181
rect 903 147 919 181
rect 1053 189 1119 202
rect 853 119 919 147
rect 953 144 1019 168
rect 565 70 615 86
rect 651 84 717 100
rect 651 50 667 84
rect 701 50 717 84
rect 753 85 819 102
rect 953 110 969 144
rect 1003 110 1019 144
rect 1053 155 1069 189
rect 1103 155 1119 189
rect 1265 206 1281 222
rect 1053 119 1119 155
rect 1153 154 1169 188
rect 1203 154 1219 188
rect 1153 120 1219 154
rect 953 85 1019 110
rect 1153 86 1169 120
rect 1203 86 1219 120
rect 1265 150 1315 206
rect 1265 116 1281 150
rect 1265 100 1315 116
rect 1351 240 1417 256
rect 1351 206 1367 240
rect 1401 206 1417 240
rect 1351 150 1417 206
rect 1351 116 1367 150
rect 1401 116 1417 150
rect 1153 85 1219 86
rect 753 51 1219 85
rect 651 17 717 50
rect 1351 17 1417 116
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 683 1440 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 0 617 1440 649
rect 0 17 1440 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -49 1440 -17
<< labels >>
flabel pwell s 0 0 1440 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 1440 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
rlabel comment s 0 0 0 0 4 o21bai_4
flabel metal1 s 0 617 1440 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 1440 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 799 242 833 276 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 1279 316 1313 350 0 FreeSans 340 0 0 0 B1_N
port 3 nsew
flabel corelocali s 1375 316 1409 350 0 FreeSans 340 0 0 0 B1_N
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 1440 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1134832
string GDS_START 1122932
<< end >>
