magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 17 191 66 333
rect 171 191 247 391
rect 1397 51 1447 493
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 17 367 69 527
rect 103 425 256 493
rect 322 425 460 493
rect 103 157 137 425
rect 293 241 392 391
rect 426 275 460 425
rect 504 415 621 527
rect 665 417 709 493
rect 777 451 1147 527
rect 1191 417 1225 493
rect 1277 451 1343 527
rect 665 383 1147 417
rect 665 381 709 383
rect 494 327 709 381
rect 494 315 533 327
rect 426 241 641 275
rect 17 123 259 157
rect 293 141 360 241
rect 394 141 461 207
rect 495 199 641 241
rect 17 51 69 123
rect 103 17 179 89
rect 223 51 259 123
rect 495 107 529 199
rect 293 51 529 107
rect 582 17 616 165
rect 675 51 709 327
rect 747 315 829 349
rect 747 187 781 315
rect 873 299 1043 349
rect 873 255 910 299
rect 815 221 910 255
rect 747 51 813 187
rect 876 157 910 221
rect 949 255 1012 265
rect 949 221 961 255
rect 995 221 1012 255
rect 949 199 1012 221
rect 1077 199 1147 383
rect 1191 299 1363 417
rect 1191 255 1279 265
rect 1191 221 1200 255
rect 1234 221 1279 255
rect 1191 199 1279 221
rect 1329 157 1363 299
rect 876 123 1043 157
rect 857 17 923 89
rect 993 51 1043 123
rect 1107 123 1363 157
rect 1107 51 1141 123
rect 1265 17 1337 89
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 961 221 995 255
rect 1200 221 1234 255
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 949 255 1007 261
rect 949 221 961 255
rect 995 252 1007 255
rect 1188 255 1246 261
rect 1188 252 1200 255
rect 995 224 1200 252
rect 995 221 1007 224
rect 949 215 1007 221
rect 1188 221 1200 224
rect 1234 221 1246 255
rect 1188 215 1246 221
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< obsm1 >>
rect 313 320 371 329
rect 861 320 919 329
rect 313 292 919 320
rect 313 283 371 292
rect 861 283 919 292
rect 415 184 473 193
rect 748 184 806 193
rect 415 156 806 184
rect 415 147 473 156
rect 748 147 806 156
<< labels >>
rlabel metal1 s 1188 252 1246 261 6 CLK
port 1 nsew signal input
rlabel metal1 s 1188 215 1246 224 6 CLK
port 1 nsew signal input
rlabel metal1 s 949 252 1007 261 6 CLK
port 1 nsew signal input
rlabel metal1 s 949 224 1246 252 6 CLK
port 1 nsew signal input
rlabel metal1 s 949 215 1007 224 6 CLK
port 1 nsew signal input
rlabel locali s 171 191 247 391 6 GATE
port 2 nsew signal input
rlabel locali s 1397 51 1447 493 6 GCLK
port 3 nsew signal output
rlabel locali s 17 191 66 333 6 SCE
port 4 nsew signal input
rlabel metal1 s 0 -48 1472 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 1472 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1472 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 381274
string GDS_START 369770
<< end >>
