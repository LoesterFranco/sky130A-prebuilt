magic
tech sky130A
magscale 1 2
timestamp 1599588232
<< locali >>
rect 107 316 173 416
rect 217 356 396 424
rect 107 282 409 316
rect 560 305 647 430
rect 375 191 510 282
rect 855 242 935 310
rect 2695 70 2761 596
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 23 492 73 596
rect 113 526 179 649
rect 563 594 629 649
rect 281 560 444 592
rect 686 560 736 596
rect 281 526 736 560
rect 23 458 509 492
rect 23 248 73 458
rect 443 316 509 458
rect 686 479 736 526
rect 956 500 1022 649
rect 686 470 929 479
rect 686 468 940 470
rect 686 466 944 468
rect 1171 466 1223 547
rect 686 439 1223 466
rect 1257 489 1314 547
rect 1257 447 1411 489
rect 1445 476 1479 649
rect 781 434 1223 439
rect 681 350 747 405
rect 681 316 703 350
rect 737 316 747 350
rect 23 210 324 248
rect 23 84 89 210
rect 258 187 324 210
rect 681 271 747 316
rect 781 237 815 434
rect 932 432 1223 434
rect 1377 442 1411 447
rect 1515 442 1590 547
rect 1659 462 1725 649
rect 1377 428 1590 442
rect 1759 428 1913 596
rect 851 398 920 400
rect 1299 398 1343 413
rect 851 364 1006 398
rect 969 321 1006 364
rect 1046 355 1343 398
rect 1085 347 1343 355
rect 1377 408 1704 428
rect 969 247 1051 321
rect 1085 293 1135 347
rect 1085 253 1299 293
rect 544 203 815 237
rect 969 208 1033 247
rect 1085 217 1135 253
rect 123 17 189 176
rect 544 153 578 203
rect 233 85 299 153
rect 391 119 578 153
rect 612 85 678 169
rect 781 140 815 203
rect 849 174 1033 208
rect 1069 174 1135 217
rect 1181 140 1231 219
rect 781 106 1231 140
rect 1265 109 1299 253
rect 1377 219 1411 408
rect 1529 394 1704 408
rect 1445 260 1495 374
rect 1537 350 1607 360
rect 1537 316 1567 350
rect 1601 316 1607 350
rect 1537 294 1607 316
rect 1645 294 1704 394
rect 1738 394 1913 428
rect 1738 260 1772 394
rect 1947 376 2013 596
rect 2121 530 2242 649
rect 2276 492 2342 596
rect 2376 526 2442 649
rect 2087 458 2447 492
rect 2087 410 2137 458
rect 2171 390 2379 424
rect 2171 376 2205 390
rect 1806 308 1870 360
rect 1947 342 2205 376
rect 2239 350 2279 356
rect 2273 316 2279 350
rect 2239 308 2279 316
rect 1806 294 2079 308
rect 1836 274 2079 294
rect 1445 226 1802 260
rect 2013 245 2079 274
rect 2199 242 2279 308
rect 1333 145 1411 219
rect 1899 192 1965 240
rect 2313 208 2379 390
rect 1499 158 1965 192
rect 1999 174 2379 208
rect 1499 109 1544 158
rect 1999 124 2033 174
rect 2413 140 2447 458
rect 233 51 678 85
rect 715 17 813 72
rect 961 17 1033 72
rect 1265 51 1544 109
rect 1578 17 1644 124
rect 1838 58 2033 124
rect 2146 17 2240 136
rect 2338 90 2447 140
rect 2488 337 2559 596
rect 2595 364 2661 649
rect 2488 271 2562 337
rect 2488 70 2559 271
rect 2595 17 2661 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 703 316 737 350
rect 1567 316 1601 350
rect 2239 316 2273 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
<< metal1 >>
rect 0 683 2784 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 0 617 2784 649
rect 0 616 50 617
rect 691 350 749 356
rect 691 316 703 350
rect 737 347 749 350
rect 1555 350 1613 356
rect 1555 347 1567 350
rect 737 319 1567 347
rect 737 316 749 319
rect 691 310 749 316
rect 1555 316 1567 319
rect 1601 347 1613 350
rect 2227 350 2285 356
rect 2227 347 2239 350
rect 1601 319 2239 347
rect 1601 316 1613 319
rect 1555 310 1613 316
rect 2227 316 2239 319
rect 2273 316 2285 350
rect 2227 310 2285 316
rect 0 49 50 50
rect 0 17 2784 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
rect 0 -49 2784 -17
<< labels >>
rlabel locali s 217 356 396 424 6 D
port 1 nsew signal input
rlabel locali s 2695 70 2761 596 6 Q
port 2 nsew signal output
rlabel metal1 s 2227 347 2285 356 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 2227 310 2285 319 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 1555 347 1613 356 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 1555 310 1613 319 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 691 347 749 356 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 691 319 2285 347 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 691 310 749 319 6 RESET_B
port 3 nsew signal input
rlabel locali s 560 305 647 430 6 SCD
port 4 nsew signal input
rlabel locali s 375 191 510 282 6 SCE
port 5 nsew signal input
rlabel locali s 107 316 173 416 6 SCE
port 5 nsew signal input
rlabel locali s 107 282 409 316 6 SCE
port 5 nsew signal input
rlabel locali s 855 242 935 310 6 CLK_N
port 6 nsew clock input
rlabel metal1 s 0 -49 2784 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 8 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 9 nsew power bidirectional
rlabel metal1 s 0 617 2784 715 6 VPWR
port 10 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2784 666
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 256034
string GDS_START 235588
<< end >>
