magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 2438 704
<< pwell >>
rect 0 0 2400 49
<< scnmos >>
rect 93 74 123 158
rect 193 74 223 158
rect 271 74 301 158
rect 412 74 442 158
rect 490 74 520 158
rect 604 74 634 222
rect 816 74 846 222
rect 1014 100 1044 184
rect 1189 100 1219 184
rect 1303 100 1333 184
rect 1487 74 1517 184
rect 1655 74 1685 184
rect 1757 74 1787 158
rect 1835 74 1865 158
rect 1935 74 1965 222
rect 2186 74 2216 222
rect 2281 74 2311 222
<< pmoshvt >>
rect 86 453 116 581
rect 186 453 216 581
rect 270 453 300 581
rect 409 453 439 581
rect 493 453 523 581
rect 641 368 671 592
rect 888 368 918 592
rect 1090 508 1120 592
rect 1180 508 1210 592
rect 1290 508 1320 592
rect 1426 424 1456 592
rect 1562 424 1592 592
rect 1674 496 1704 580
rect 1832 496 1862 580
rect 1992 380 2022 580
rect 2194 368 2224 592
rect 2284 368 2314 592
<< ndiff >>
rect 547 158 604 222
rect 27 128 93 158
rect 27 94 43 128
rect 77 94 93 128
rect 27 74 93 94
rect 123 124 193 158
rect 123 90 148 124
rect 182 90 193 124
rect 123 74 193 90
rect 223 74 271 158
rect 301 120 412 158
rect 301 86 339 120
rect 373 86 412 120
rect 301 74 412 86
rect 442 74 490 158
rect 520 133 604 158
rect 520 99 554 133
rect 588 99 604 133
rect 520 74 604 99
rect 634 184 691 222
rect 634 150 645 184
rect 679 150 691 184
rect 634 116 691 150
rect 634 82 645 116
rect 679 82 691 116
rect 634 74 691 82
rect 745 136 816 222
rect 745 102 757 136
rect 791 102 816 136
rect 745 74 816 102
rect 846 210 903 222
rect 846 176 857 210
rect 891 176 903 210
rect 846 120 903 176
rect 846 86 857 120
rect 891 86 903 120
rect 957 170 1014 184
rect 957 136 969 170
rect 1003 136 1014 170
rect 957 100 1014 136
rect 1044 170 1189 184
rect 1044 136 1105 170
rect 1139 136 1189 170
rect 1044 100 1189 136
rect 1219 100 1303 184
rect 1333 100 1487 184
rect 846 74 903 86
rect 1348 94 1487 100
rect 1348 60 1360 94
rect 1394 74 1487 94
rect 1517 170 1655 184
rect 1517 136 1528 170
rect 1562 136 1655 170
rect 1517 74 1655 136
rect 1685 158 1742 184
rect 1885 158 1935 222
rect 1685 133 1757 158
rect 1685 99 1696 133
rect 1730 99 1757 133
rect 1685 74 1757 99
rect 1787 74 1835 158
rect 1865 133 1935 158
rect 1865 99 1876 133
rect 1910 99 1935 133
rect 1865 74 1935 99
rect 1965 210 2022 222
rect 1965 176 1976 210
rect 2010 176 2022 210
rect 1965 120 2022 176
rect 1965 86 1976 120
rect 2010 86 2022 120
rect 1965 74 2022 86
rect 2115 194 2186 222
rect 2115 160 2141 194
rect 2175 160 2186 194
rect 2115 120 2186 160
rect 2115 86 2141 120
rect 2175 86 2186 120
rect 2115 74 2186 86
rect 2216 210 2281 222
rect 2216 176 2227 210
rect 2261 176 2281 210
rect 2216 120 2281 176
rect 2216 86 2227 120
rect 2261 86 2281 120
rect 2216 74 2281 86
rect 2311 210 2373 222
rect 2311 176 2327 210
rect 2361 176 2373 210
rect 2311 120 2373 176
rect 2311 86 2327 120
rect 2361 86 2373 120
rect 2311 74 2373 86
rect 1394 60 1406 74
rect 1348 48 1406 60
<< pdiff >>
rect 541 608 623 620
rect 541 581 565 608
rect 27 569 86 581
rect 27 535 39 569
rect 73 535 86 569
rect 27 499 86 535
rect 27 465 39 499
rect 73 465 86 499
rect 27 453 86 465
rect 116 573 186 581
rect 116 539 139 573
rect 173 539 186 573
rect 116 505 186 539
rect 116 471 139 505
rect 173 471 186 505
rect 116 453 186 471
rect 216 453 270 581
rect 300 573 409 581
rect 300 539 337 573
rect 371 539 409 573
rect 300 505 409 539
rect 300 471 337 505
rect 371 471 409 505
rect 300 453 409 471
rect 439 453 493 581
rect 523 574 565 581
rect 599 592 623 608
rect 784 608 870 620
rect 599 574 641 592
rect 523 453 641 574
rect 588 368 641 453
rect 671 440 730 592
rect 671 406 684 440
rect 718 406 730 440
rect 671 368 730 406
rect 784 574 810 608
rect 844 592 870 608
rect 844 574 888 592
rect 784 368 888 574
rect 918 427 977 592
rect 1031 567 1090 592
rect 1031 533 1043 567
rect 1077 533 1090 567
rect 1031 508 1090 533
rect 1120 567 1180 592
rect 1120 533 1133 567
rect 1167 533 1180 567
rect 1120 508 1180 533
rect 1210 508 1290 592
rect 1320 567 1426 592
rect 1320 533 1333 567
rect 1367 533 1426 567
rect 1320 508 1426 533
rect 918 393 931 427
rect 965 393 977 427
rect 918 368 977 393
rect 1373 424 1426 508
rect 1456 499 1562 592
rect 1456 465 1469 499
rect 1503 465 1562 499
rect 1456 424 1562 465
rect 1592 580 1645 592
rect 2135 580 2194 592
rect 1592 558 1674 580
rect 1592 524 1605 558
rect 1639 524 1674 558
rect 1592 496 1674 524
rect 1704 496 1832 580
rect 1862 568 1992 580
rect 1862 534 1875 568
rect 1909 534 1945 568
rect 1979 534 1992 568
rect 1862 496 1992 534
rect 1592 424 1651 496
rect 1939 380 1992 496
rect 2022 550 2081 580
rect 2022 516 2035 550
rect 2069 516 2081 550
rect 2022 380 2081 516
rect 2135 546 2147 580
rect 2181 546 2194 580
rect 2135 497 2194 546
rect 2135 463 2147 497
rect 2181 463 2194 497
rect 2135 414 2194 463
rect 2135 380 2147 414
rect 2181 380 2194 414
rect 2135 368 2194 380
rect 2224 580 2284 592
rect 2224 546 2237 580
rect 2271 546 2284 580
rect 2224 497 2284 546
rect 2224 463 2237 497
rect 2271 463 2284 497
rect 2224 414 2284 463
rect 2224 380 2237 414
rect 2271 380 2284 414
rect 2224 368 2284 380
rect 2314 580 2373 592
rect 2314 546 2327 580
rect 2361 546 2373 580
rect 2314 497 2373 546
rect 2314 463 2327 497
rect 2361 463 2373 497
rect 2314 414 2373 463
rect 2314 380 2327 414
rect 2361 380 2373 414
rect 2314 368 2373 380
<< ndiffc >>
rect 43 94 77 128
rect 148 90 182 124
rect 339 86 373 120
rect 554 99 588 133
rect 645 150 679 184
rect 645 82 679 116
rect 757 102 791 136
rect 857 176 891 210
rect 857 86 891 120
rect 969 136 1003 170
rect 1105 136 1139 170
rect 1360 60 1394 94
rect 1528 136 1562 170
rect 1696 99 1730 133
rect 1876 99 1910 133
rect 1976 176 2010 210
rect 1976 86 2010 120
rect 2141 160 2175 194
rect 2141 86 2175 120
rect 2227 176 2261 210
rect 2227 86 2261 120
rect 2327 176 2361 210
rect 2327 86 2361 120
<< pdiffc >>
rect 39 535 73 569
rect 39 465 73 499
rect 139 539 173 573
rect 139 471 173 505
rect 337 539 371 573
rect 337 471 371 505
rect 565 574 599 608
rect 684 406 718 440
rect 810 574 844 608
rect 1043 533 1077 567
rect 1133 533 1167 567
rect 1333 533 1367 567
rect 931 393 965 427
rect 1469 465 1503 499
rect 1605 524 1639 558
rect 1875 534 1909 568
rect 1945 534 1979 568
rect 2035 516 2069 550
rect 2147 546 2181 580
rect 2147 463 2181 497
rect 2147 380 2181 414
rect 2237 546 2271 580
rect 2237 463 2271 497
rect 2237 380 2271 414
rect 2327 546 2361 580
rect 2327 463 2361 497
rect 2327 380 2361 414
<< poly >>
rect 86 581 116 607
rect 186 581 216 607
rect 270 581 300 607
rect 409 581 439 607
rect 493 581 523 607
rect 641 592 671 618
rect 86 438 116 453
rect 186 438 216 453
rect 270 438 300 453
rect 409 438 439 453
rect 493 438 523 453
rect 39 408 219 438
rect 39 246 69 408
rect 267 372 303 438
rect 406 421 442 438
rect 376 405 442 421
rect 117 344 223 360
rect 117 310 133 344
rect 167 310 223 344
rect 117 294 223 310
rect 39 230 151 246
rect 39 216 101 230
rect 85 196 101 216
rect 135 196 151 230
rect 85 180 151 196
rect 93 158 123 180
rect 193 158 223 294
rect 267 356 333 372
rect 267 322 283 356
rect 317 322 333 356
rect 376 371 392 405
rect 426 371 442 405
rect 376 355 442 371
rect 490 421 526 438
rect 490 405 556 421
rect 490 371 506 405
rect 540 371 556 405
rect 267 288 333 322
rect 267 254 283 288
rect 317 254 333 288
rect 267 238 333 254
rect 490 337 556 371
rect 888 592 918 618
rect 1090 592 1120 618
rect 1180 592 1210 618
rect 1290 592 1320 618
rect 1426 592 1456 618
rect 1562 592 1592 618
rect 1090 493 1120 508
rect 1180 493 1210 508
rect 1290 493 1320 508
rect 1087 456 1123 493
rect 1009 440 1123 456
rect 1009 406 1025 440
rect 1059 426 1123 440
rect 1177 460 1213 493
rect 1177 444 1245 460
rect 1059 406 1075 426
rect 1009 372 1075 406
rect 1177 410 1195 444
rect 1229 410 1245 444
rect 1177 378 1245 410
rect 641 353 671 368
rect 888 353 918 368
rect 490 303 506 337
rect 540 303 556 337
rect 638 336 674 353
rect 490 287 556 303
rect 604 320 724 336
rect 885 326 921 353
rect 271 158 301 238
rect 375 230 442 246
rect 375 196 391 230
rect 425 196 442 230
rect 375 180 442 196
rect 412 158 442 180
rect 490 158 520 287
rect 604 286 674 320
rect 708 286 724 320
rect 604 270 724 286
rect 767 310 921 326
rect 1009 338 1025 372
rect 1059 338 1075 372
rect 1009 322 1075 338
rect 1117 348 1245 378
rect 1287 350 1323 493
rect 1674 580 1704 606
rect 1832 580 1862 606
rect 1992 580 2022 606
rect 2194 592 2224 618
rect 2284 592 2314 618
rect 1674 481 1704 496
rect 1832 481 1862 496
rect 1671 464 1707 481
rect 1671 448 1749 464
rect 1426 409 1456 424
rect 1562 409 1592 424
rect 1671 414 1699 448
rect 1733 414 1749 448
rect 1423 392 1459 409
rect 1369 376 1509 392
rect 1559 386 1595 409
rect 1671 398 1749 414
rect 1829 398 1865 481
rect 767 276 783 310
rect 817 276 921 310
rect 767 274 921 276
rect 1117 274 1147 348
rect 1287 320 1327 350
rect 1369 342 1385 376
rect 1419 342 1509 376
rect 1369 326 1509 342
rect 604 222 634 270
rect 767 244 1147 274
rect 1297 278 1327 320
rect 1189 256 1255 272
rect 816 222 846 244
rect 1014 184 1044 244
rect 1189 222 1205 256
rect 1239 222 1255 256
rect 1189 206 1255 222
rect 1297 262 1431 278
rect 1297 228 1313 262
rect 1347 228 1381 262
rect 1415 228 1431 262
rect 1297 212 1431 228
rect 1479 229 1509 326
rect 1557 370 1623 386
rect 1557 336 1573 370
rect 1607 350 1623 370
rect 1835 381 1865 398
rect 1835 365 1907 381
rect 1992 365 2022 380
rect 1607 336 1787 350
rect 1557 320 1787 336
rect 1619 256 1685 272
rect 1189 184 1219 206
rect 1303 184 1333 212
rect 1479 199 1517 229
rect 1619 222 1635 256
rect 1669 222 1685 256
rect 1619 206 1685 222
rect 1487 184 1517 199
rect 1655 184 1685 206
rect 1014 74 1044 100
rect 1189 74 1219 100
rect 1303 74 1333 100
rect 93 48 123 74
rect 193 48 223 74
rect 271 48 301 74
rect 412 48 442 74
rect 490 48 520 74
rect 604 48 634 74
rect 816 48 846 74
rect 1757 158 1787 320
rect 1835 331 1857 365
rect 1891 331 1907 365
rect 1989 348 2025 365
rect 2194 353 2224 368
rect 2284 353 2314 368
rect 1835 315 1907 331
rect 1955 332 2025 348
rect 1835 158 1865 315
rect 1955 298 1971 332
rect 2005 298 2025 332
rect 2191 310 2227 353
rect 2281 310 2317 353
rect 1955 282 2025 298
rect 2075 294 2317 310
rect 1955 267 1985 282
rect 1935 237 1985 267
rect 2075 260 2091 294
rect 2125 260 2159 294
rect 2193 260 2317 294
rect 2075 244 2317 260
rect 1935 222 1965 237
rect 2186 222 2216 244
rect 2281 222 2311 244
rect 1487 48 1517 74
rect 1655 48 1685 74
rect 1757 48 1787 74
rect 1835 48 1865 74
rect 1935 48 1965 74
rect 2186 48 2216 74
rect 2281 48 2311 74
<< polycont >>
rect 133 310 167 344
rect 101 196 135 230
rect 283 322 317 356
rect 392 371 426 405
rect 506 371 540 405
rect 283 254 317 288
rect 1025 406 1059 440
rect 1195 410 1229 444
rect 506 303 540 337
rect 391 196 425 230
rect 674 286 708 320
rect 1025 338 1059 372
rect 1699 414 1733 448
rect 783 276 817 310
rect 1385 342 1419 376
rect 1205 222 1239 256
rect 1313 228 1347 262
rect 1381 228 1415 262
rect 1573 336 1607 370
rect 1635 222 1669 256
rect 1857 331 1891 365
rect 1971 298 2005 332
rect 2091 260 2125 294
rect 2159 260 2193 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2400 683
rect 17 569 89 585
rect 17 535 39 569
rect 73 535 89 569
rect 17 499 89 535
rect 17 465 39 499
rect 73 465 89 499
rect 123 573 189 649
rect 537 608 627 649
rect 123 539 139 573
rect 173 539 189 573
rect 123 505 189 539
rect 123 471 139 505
rect 173 471 189 505
rect 297 573 412 589
rect 297 539 337 573
rect 371 539 412 573
rect 537 574 565 608
rect 599 574 627 608
rect 537 558 627 574
rect 780 608 874 649
rect 780 574 810 608
rect 844 574 874 608
rect 780 558 874 574
rect 1027 567 1077 596
rect 297 524 412 539
rect 1027 533 1043 567
rect 1027 524 1077 533
rect 297 505 1077 524
rect 297 471 337 505
rect 371 490 1077 505
rect 1111 567 1183 596
rect 1111 533 1133 567
rect 1167 533 1183 567
rect 1111 504 1183 533
rect 1317 567 1367 649
rect 1317 533 1333 567
rect 1317 504 1367 533
rect 1401 581 1571 615
rect 371 471 624 490
rect 17 437 89 465
rect 17 405 442 437
rect 17 403 392 405
rect 17 344 183 403
rect 376 371 392 403
rect 426 371 442 405
rect 17 310 133 344
rect 167 310 183 344
rect 17 294 183 310
rect 217 356 333 369
rect 217 322 283 356
rect 317 322 333 356
rect 376 355 442 371
rect 490 405 556 430
rect 490 371 506 405
rect 540 371 556 405
rect 17 128 51 294
rect 217 288 333 322
rect 217 254 283 288
rect 317 254 333 288
rect 490 337 556 371
rect 490 303 506 337
rect 540 303 556 337
rect 490 287 556 303
rect 85 230 167 246
rect 217 238 333 254
rect 590 253 624 471
rect 668 440 829 456
rect 668 406 684 440
rect 718 406 829 440
rect 668 390 829 406
rect 658 320 737 356
rect 658 286 674 320
rect 708 286 737 320
rect 658 270 737 286
rect 771 310 829 390
rect 771 276 783 310
rect 817 276 829 310
rect 85 196 101 230
rect 135 204 167 230
rect 375 230 441 246
rect 375 204 391 230
rect 135 196 391 204
rect 425 196 441 230
rect 85 170 441 196
rect 475 219 624 253
rect 771 260 829 276
rect 863 294 897 490
rect 931 440 1075 456
rect 931 427 1025 440
rect 965 406 1025 427
rect 1059 406 1075 440
rect 965 393 1075 406
rect 931 372 1075 393
rect 931 364 1025 372
rect 1009 338 1025 364
rect 1059 338 1075 372
rect 1009 322 1075 338
rect 1111 360 1145 504
rect 1401 460 1435 581
rect 1179 444 1435 460
rect 1179 410 1195 444
rect 1229 426 1435 444
rect 1469 499 1503 522
rect 1229 410 1245 426
rect 1179 394 1245 410
rect 1369 376 1435 392
rect 1369 360 1385 376
rect 1111 342 1385 360
rect 1419 342 1435 376
rect 1111 326 1435 342
rect 863 260 975 294
rect 771 236 805 260
rect 85 162 167 170
rect 475 136 509 219
rect 661 202 805 236
rect 841 210 907 226
rect 661 184 695 202
rect 17 94 43 128
rect 77 94 98 128
rect 17 78 98 94
rect 132 124 198 128
rect 132 90 148 124
rect 182 90 198 124
rect 132 17 198 90
rect 296 120 509 136
rect 296 86 339 120
rect 373 86 509 120
rect 296 70 509 86
rect 543 133 595 162
rect 543 99 554 133
rect 588 99 595 133
rect 543 17 595 99
rect 629 150 645 184
rect 679 150 695 184
rect 841 176 857 210
rect 891 176 907 210
rect 629 116 695 150
rect 629 82 645 116
rect 679 82 695 116
rect 629 66 695 82
rect 741 136 807 168
rect 741 102 757 136
rect 791 102 807 136
rect 741 17 807 102
rect 841 120 907 176
rect 841 86 857 120
rect 891 86 907 120
rect 941 188 975 260
rect 941 170 1003 188
rect 941 136 969 170
rect 941 119 1003 136
rect 841 85 907 86
rect 1037 85 1071 322
rect 1111 188 1155 326
rect 1469 278 1503 465
rect 1537 386 1571 581
rect 1605 558 1655 584
rect 1639 532 1655 558
rect 1859 568 1985 649
rect 1859 534 1875 568
rect 1909 534 1945 568
rect 1979 534 1985 568
rect 1639 524 1812 532
rect 1605 498 1812 524
rect 1859 518 1985 534
rect 2019 550 2089 584
rect 1657 448 1744 464
rect 1657 414 1699 448
rect 1733 414 1744 448
rect 1657 398 1744 414
rect 1778 449 1812 498
rect 2019 516 2035 550
rect 2069 516 2089 550
rect 2019 483 2089 516
rect 1778 415 2021 449
rect 1537 370 1623 386
rect 1537 336 1573 370
rect 1607 336 1623 370
rect 1537 320 1623 336
rect 1105 170 1155 188
rect 1139 136 1155 170
rect 1105 119 1155 136
rect 1189 256 1255 272
rect 1189 222 1205 256
rect 1239 222 1255 256
rect 1189 178 1255 222
rect 1297 262 1503 278
rect 1657 272 1691 398
rect 1297 228 1313 262
rect 1347 228 1381 262
rect 1415 246 1503 262
rect 1612 256 1691 272
rect 1415 228 1578 246
rect 1297 212 1578 228
rect 1189 144 1478 178
rect 1189 85 1223 144
rect 841 51 1223 85
rect 1344 94 1410 110
rect 1344 60 1360 94
rect 1394 60 1410 94
rect 1344 17 1410 60
rect 1444 85 1478 144
rect 1512 170 1578 212
rect 1512 136 1528 170
rect 1562 136 1578 170
rect 1512 119 1578 136
rect 1612 222 1635 256
rect 1669 222 1691 256
rect 1612 206 1691 222
rect 1612 85 1646 206
rect 1778 162 1812 415
rect 1846 365 1907 381
rect 1846 331 1857 365
rect 1891 331 1907 365
rect 1846 248 1907 331
rect 1955 332 2021 415
rect 1955 298 1971 332
rect 2005 298 2021 332
rect 1955 282 2021 298
rect 2055 310 2089 483
rect 2131 580 2181 649
rect 2131 546 2147 580
rect 2131 497 2181 546
rect 2131 463 2147 497
rect 2131 414 2181 463
rect 2131 380 2147 414
rect 2131 364 2181 380
rect 2221 580 2287 596
rect 2221 546 2237 580
rect 2271 546 2287 580
rect 2221 497 2287 546
rect 2221 463 2237 497
rect 2271 463 2287 497
rect 2221 414 2287 463
rect 2221 380 2237 414
rect 2271 380 2287 414
rect 2221 364 2287 380
rect 2327 580 2377 649
rect 2361 546 2377 580
rect 2327 497 2377 546
rect 2361 463 2377 497
rect 2327 414 2377 463
rect 2361 380 2377 414
rect 2327 364 2377 380
rect 2055 294 2209 310
rect 2055 260 2091 294
rect 2125 260 2159 294
rect 2193 260 2209 294
rect 2055 248 2209 260
rect 1846 244 2209 248
rect 1846 214 2089 244
rect 1960 210 2026 214
rect 2243 210 2277 364
rect 1960 176 1976 210
rect 2010 176 2026 210
rect 1444 51 1646 85
rect 1680 133 1812 162
rect 1680 99 1696 133
rect 1730 128 1812 133
rect 1860 133 1926 162
rect 1730 99 1759 128
rect 1680 70 1759 99
rect 1860 99 1876 133
rect 1910 99 1926 133
rect 1860 17 1926 99
rect 1960 120 2026 176
rect 1960 86 1976 120
rect 2010 86 2026 120
rect 1960 70 2026 86
rect 2123 194 2177 210
rect 2123 160 2141 194
rect 2175 160 2177 194
rect 2123 120 2177 160
rect 2123 86 2141 120
rect 2175 86 2177 120
rect 2123 17 2177 86
rect 2211 176 2227 210
rect 2261 176 2277 210
rect 2211 120 2277 176
rect 2211 86 2227 120
rect 2261 86 2277 120
rect 2211 70 2277 86
rect 2311 210 2377 226
rect 2311 176 2327 210
rect 2361 176 2377 210
rect 2311 120 2377 176
rect 2311 86 2327 120
rect 2361 86 2377 120
rect 2311 17 2377 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2400 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
<< metal1 >>
rect 0 683 2400 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2400 683
rect 0 617 2400 649
rect 0 17 2400 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2400 17
rect 0 -49 2400 -17
<< labels >>
rlabel comment s 0 0 0 0 4 sdfxtp_2
flabel comment s 993 260 993 260 0 FreeSans 200 0 0 0 no_jumper_check
flabel pwell s 0 0 2400 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 2400 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 2400 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 2400 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 127 168 161 202 0 FreeSans 340 0 0 0 SCE
port 4 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 SCD
port 3 nsew
flabel corelocali s 511 390 545 424 0 FreeSans 340 0 0 0 SCD
port 3 nsew
flabel corelocali s 2239 390 2273 424 0 FreeSans 340 0 0 0 Q
port 9 nsew
flabel corelocali s 2239 464 2273 498 0 FreeSans 340 0 0 0 Q
port 9 nsew
flabel corelocali s 2239 538 2273 572 0 FreeSans 340 0 0 0 Q
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 2400 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 241456
string GDS_START 224414
<< end >>
