magic
tech sky130A
magscale 1 2
timestamp 1601050056
<< nwell >>
rect -38 351 2246 704
rect -38 332 230 351
rect 1064 332 2246 351
rect 1064 311 1280 332
<< pwell >>
rect 0 0 2208 49
<< scpmos >>
rect 81 523 117 607
rect 171 523 207 607
rect 367 387 403 611
rect 457 387 493 611
rect 665 463 701 547
rect 755 463 791 547
rect 833 463 869 547
rect 954 463 990 547
rect 1158 347 1194 547
rect 1259 377 1295 577
rect 1435 493 1471 577
rect 1519 493 1555 577
rect 1634 493 1670 577
rect 1724 493 1760 577
rect 1831 409 1867 577
rect 2088 368 2124 592
<< nmoslvt >>
rect 87 78 117 162
rect 165 78 195 162
rect 376 119 406 267
rect 480 119 510 267
rect 694 138 724 222
rect 791 138 821 222
rect 864 138 894 222
rect 942 138 972 222
rect 1073 74 1103 222
rect 1236 74 1266 222
rect 1446 81 1476 165
rect 1524 81 1554 165
rect 1626 81 1656 165
rect 1698 81 1728 165
rect 1896 74 1926 184
rect 2094 74 2124 222
<< ndiff >>
rect 310 228 376 267
rect 310 194 322 228
rect 356 194 376 228
rect 30 137 87 162
rect 30 103 42 137
rect 76 103 87 137
rect 30 78 87 103
rect 117 78 165 162
rect 195 137 252 162
rect 195 103 206 137
rect 240 103 252 137
rect 310 160 376 194
rect 310 126 322 160
rect 356 126 376 160
rect 310 119 376 126
rect 406 160 480 267
rect 406 126 426 160
rect 460 126 480 160
rect 406 119 480 126
rect 510 222 560 267
rect 510 161 576 222
rect 510 127 526 161
rect 560 127 576 161
rect 630 197 694 222
rect 630 163 641 197
rect 675 163 694 197
rect 630 138 694 163
rect 724 189 791 222
rect 724 155 741 189
rect 775 155 791 189
rect 724 138 791 155
rect 821 138 864 222
rect 894 138 942 222
rect 972 138 1073 222
rect 510 119 576 127
rect 310 118 361 119
rect 195 78 252 103
rect 421 118 465 119
rect 987 79 1073 138
rect 987 45 1005 79
rect 1039 74 1073 79
rect 1103 188 1236 222
rect 1103 154 1180 188
rect 1214 154 1236 188
rect 1103 74 1236 154
rect 1266 165 1316 222
rect 2037 210 2094 222
rect 1266 153 1446 165
rect 1266 119 1280 153
rect 1314 119 1366 153
rect 1400 119 1446 153
rect 1266 81 1446 119
rect 1476 81 1524 165
rect 1554 140 1626 165
rect 1554 106 1565 140
rect 1599 106 1626 140
rect 1554 81 1626 106
rect 1656 81 1698 165
rect 1728 140 1785 165
rect 1728 106 1739 140
rect 1773 106 1785 140
rect 1728 81 1785 106
rect 1839 136 1896 184
rect 1839 102 1851 136
rect 1885 102 1896 136
rect 1266 74 1316 81
rect 1039 45 1058 74
rect 1839 74 1896 102
rect 1926 146 1983 184
rect 1926 112 1937 146
rect 1971 112 1983 146
rect 1926 74 1983 112
rect 2037 176 2049 210
rect 2083 176 2094 210
rect 2037 120 2094 176
rect 2037 86 2049 120
rect 2083 86 2094 120
rect 2037 74 2094 86
rect 2124 210 2181 222
rect 2124 176 2135 210
rect 2169 176 2181 210
rect 2124 120 2181 176
rect 2124 86 2135 120
rect 2169 86 2181 120
rect 2124 74 2181 86
rect 987 33 1058 45
<< pdiff >>
rect 27 581 81 607
rect 27 547 37 581
rect 71 547 81 581
rect 27 523 81 547
rect 117 581 171 607
rect 117 547 127 581
rect 161 547 171 581
rect 117 523 171 547
rect 207 595 263 607
rect 207 561 217 595
rect 251 561 263 595
rect 207 523 263 561
rect 317 462 367 611
rect 299 437 367 462
rect 299 403 307 437
rect 341 403 367 437
rect 299 387 367 403
rect 403 591 457 611
rect 403 557 413 591
rect 447 557 457 591
rect 403 387 457 557
rect 493 439 547 611
rect 493 405 503 439
rect 537 405 547 439
rect 493 387 547 405
rect 884 582 939 597
rect 884 548 894 582
rect 928 548 939 582
rect 2023 580 2088 592
rect 884 547 939 548
rect 1209 547 1259 577
rect 609 524 665 547
rect 609 490 621 524
rect 655 490 665 524
rect 609 463 665 490
rect 701 539 755 547
rect 701 505 711 539
rect 745 505 755 539
rect 701 463 755 505
rect 791 463 833 547
rect 869 463 954 547
rect 990 514 1046 547
rect 990 480 1000 514
rect 1034 480 1046 514
rect 990 463 1046 480
rect 1100 535 1158 547
rect 1100 501 1112 535
rect 1146 501 1158 535
rect 1100 467 1158 501
rect 1100 433 1112 467
rect 1146 433 1158 467
rect 1100 399 1158 433
rect 1100 365 1112 399
rect 1146 365 1158 399
rect 1100 347 1158 365
rect 1194 535 1259 547
rect 1194 501 1212 535
rect 1246 501 1259 535
rect 1194 423 1259 501
rect 1194 389 1212 423
rect 1246 389 1259 423
rect 1194 377 1259 389
rect 1295 545 1435 577
rect 1295 511 1312 545
rect 1346 511 1391 545
rect 1425 511 1435 545
rect 1295 493 1435 511
rect 1471 493 1519 577
rect 1555 552 1634 577
rect 1555 518 1577 552
rect 1611 518 1634 552
rect 1555 493 1634 518
rect 1670 552 1724 577
rect 1670 518 1680 552
rect 1714 518 1724 552
rect 1670 493 1724 518
rect 1760 565 1831 577
rect 1760 531 1787 565
rect 1821 531 1831 565
rect 1760 493 1831 531
rect 1295 377 1345 493
rect 1194 347 1244 377
rect 1775 489 1831 493
rect 1775 455 1787 489
rect 1821 455 1831 489
rect 1775 409 1831 455
rect 1867 565 1923 577
rect 1867 531 1877 565
rect 1911 531 1923 565
rect 1867 455 1923 531
rect 1867 421 1877 455
rect 1911 421 1923 455
rect 1867 409 1923 421
rect 2023 546 2035 580
rect 2069 546 2088 580
rect 2023 503 2088 546
rect 2023 469 2035 503
rect 2069 469 2088 503
rect 2023 427 2088 469
rect 2023 393 2035 427
rect 2069 393 2088 427
rect 2023 368 2088 393
rect 2124 580 2181 592
rect 2124 546 2135 580
rect 2169 546 2181 580
rect 2124 497 2181 546
rect 2124 463 2135 497
rect 2169 463 2181 497
rect 2124 414 2181 463
rect 2124 380 2135 414
rect 2169 380 2181 414
rect 2124 368 2181 380
<< ndiffc >>
rect 322 194 356 228
rect 42 103 76 137
rect 206 103 240 137
rect 322 126 356 160
rect 426 126 460 160
rect 526 127 560 161
rect 641 163 675 197
rect 741 155 775 189
rect 1005 45 1039 79
rect 1180 154 1214 188
rect 1280 119 1314 153
rect 1366 119 1400 153
rect 1565 106 1599 140
rect 1739 106 1773 140
rect 1851 102 1885 136
rect 1937 112 1971 146
rect 2049 176 2083 210
rect 2049 86 2083 120
rect 2135 176 2169 210
rect 2135 86 2169 120
<< pdiffc >>
rect 37 547 71 581
rect 127 547 161 581
rect 217 561 251 595
rect 307 403 341 437
rect 413 557 447 591
rect 503 405 537 439
rect 894 548 928 582
rect 621 490 655 524
rect 711 505 745 539
rect 1000 480 1034 514
rect 1112 501 1146 535
rect 1112 433 1146 467
rect 1112 365 1146 399
rect 1212 501 1246 535
rect 1212 389 1246 423
rect 1312 511 1346 545
rect 1391 511 1425 545
rect 1577 518 1611 552
rect 1680 518 1714 552
rect 1787 531 1821 565
rect 1787 455 1821 489
rect 1877 531 1911 565
rect 1877 421 1911 455
rect 2035 546 2069 580
rect 2035 469 2069 503
rect 2035 393 2069 427
rect 2135 546 2169 580
rect 2135 463 2169 497
rect 2135 380 2169 414
<< poly >>
rect 81 607 117 633
rect 171 607 207 633
rect 367 611 403 637
rect 457 611 493 637
rect 562 615 1295 645
rect 81 402 117 523
rect 171 428 207 523
rect 44 386 117 402
rect 44 352 60 386
rect 94 352 117 386
rect 44 318 117 352
rect 44 284 60 318
rect 94 284 117 318
rect 44 250 117 284
rect 44 216 60 250
rect 94 216 117 250
rect 44 200 117 216
rect 87 162 117 200
rect 165 412 264 428
rect 165 378 214 412
rect 248 378 264 412
rect 165 344 264 378
rect 367 355 403 387
rect 457 355 493 387
rect 562 355 592 615
rect 665 547 701 573
rect 755 547 791 615
rect 833 547 869 573
rect 1259 577 1295 615
rect 1435 577 1471 603
rect 1519 577 1555 603
rect 1634 577 1670 603
rect 1724 577 1760 603
rect 1831 577 1867 603
rect 2088 592 2124 618
rect 954 547 990 573
rect 1158 547 1194 573
rect 665 403 701 463
rect 755 437 791 463
rect 165 310 214 344
rect 248 310 264 344
rect 165 276 264 310
rect 349 339 415 355
rect 349 305 365 339
rect 399 305 415 339
rect 349 289 415 305
rect 457 339 592 355
rect 457 305 503 339
rect 537 318 592 339
rect 634 387 701 403
rect 833 425 869 463
rect 954 437 990 463
rect 955 425 990 437
rect 833 409 905 425
rect 833 400 855 409
rect 634 353 650 387
rect 684 367 701 387
rect 839 375 855 400
rect 889 375 905 409
rect 684 353 796 367
rect 839 359 905 375
rect 955 409 1057 425
rect 955 375 1007 409
rect 1041 375 1057 409
rect 955 359 1057 375
rect 634 337 796 353
rect 537 313 596 318
rect 766 317 796 337
rect 537 307 599 313
rect 537 305 604 307
rect 457 304 604 305
rect 457 295 608 304
rect 165 242 214 276
rect 248 242 264 276
rect 376 267 406 289
rect 457 282 724 295
rect 766 287 821 317
rect 480 267 510 282
rect 571 278 724 282
rect 165 226 264 242
rect 165 162 195 226
rect 575 265 724 278
rect 694 222 724 265
rect 791 222 821 287
rect 864 222 894 359
rect 960 267 990 359
rect 1435 461 1471 493
rect 1393 445 1471 461
rect 1393 411 1409 445
rect 1443 411 1471 445
rect 1393 395 1471 411
rect 1259 347 1295 377
rect 1519 349 1555 493
rect 1634 451 1670 493
rect 1603 435 1670 451
rect 1603 401 1619 435
rect 1653 401 1670 435
rect 1603 385 1670 401
rect 1158 315 1194 347
rect 1259 317 1476 347
rect 942 237 990 267
rect 1064 299 1194 315
rect 1064 265 1080 299
rect 1114 285 1194 299
rect 1114 265 1130 285
rect 1064 249 1130 265
rect 1236 253 1404 269
rect 942 222 972 237
rect 1073 222 1103 249
rect 1236 239 1354 253
rect 1236 222 1266 239
rect 376 93 406 119
rect 480 93 510 119
rect 694 112 724 138
rect 791 112 821 138
rect 864 112 894 138
rect 87 52 117 78
rect 165 51 195 78
rect 942 51 972 138
rect 165 21 972 51
rect 1338 219 1354 239
rect 1388 219 1404 253
rect 1338 203 1404 219
rect 1446 165 1476 317
rect 1519 269 1549 349
rect 1518 253 1584 269
rect 1518 219 1534 253
rect 1568 219 1584 253
rect 1518 203 1584 219
rect 1524 165 1554 203
rect 1626 165 1656 385
rect 1724 337 1760 493
rect 1831 337 1867 409
rect 2088 343 2124 368
rect 1704 321 1867 337
rect 1704 301 1720 321
rect 1698 287 1720 301
rect 1754 287 1867 321
rect 1698 271 1867 287
rect 1921 327 2124 343
rect 1921 293 1937 327
rect 1971 293 2124 327
rect 1921 277 2124 293
rect 1698 165 1728 271
rect 1831 229 1861 271
rect 1831 199 1926 229
rect 2094 222 2124 277
rect 1896 184 1926 199
rect 1073 48 1103 74
rect 1236 48 1266 74
rect 1446 55 1476 81
rect 1524 55 1554 81
rect 1626 55 1656 81
rect 1698 55 1728 81
rect 1896 48 1926 74
rect 2094 48 2124 74
<< polycont >>
rect 60 352 94 386
rect 60 284 94 318
rect 60 216 94 250
rect 214 378 248 412
rect 214 310 248 344
rect 365 305 399 339
rect 503 305 537 339
rect 650 353 684 387
rect 855 375 889 409
rect 1007 375 1041 409
rect 214 242 248 276
rect 1409 411 1443 445
rect 1619 401 1653 435
rect 1080 265 1114 299
rect 1354 219 1388 253
rect 1534 219 1568 253
rect 1720 287 1754 321
rect 1937 293 1971 327
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 21 581 71 649
rect 21 547 37 581
rect 21 531 71 547
rect 105 581 167 607
rect 105 547 127 581
rect 161 547 167 581
rect 201 595 267 649
rect 201 561 217 595
rect 251 561 267 595
rect 201 557 267 561
rect 397 591 463 649
rect 397 557 413 591
rect 447 557 463 591
rect 878 582 944 649
rect 105 530 167 547
rect 105 525 173 530
rect 105 523 177 525
rect 605 524 661 551
rect 605 523 621 524
rect 105 504 621 523
rect 137 490 621 504
rect 655 490 661 524
rect 695 539 843 551
rect 878 548 894 582
rect 928 548 944 582
rect 695 505 711 539
rect 745 512 843 539
rect 990 514 1050 536
rect 990 512 1000 514
rect 745 505 1000 512
rect 137 489 661 490
rect 25 386 103 434
rect 25 352 60 386
rect 94 352 103 386
rect 25 318 103 352
rect 25 284 60 318
rect 94 284 103 318
rect 25 250 103 284
rect 25 216 60 250
rect 94 216 103 250
rect 25 200 103 216
rect 137 166 171 489
rect 621 471 661 489
rect 787 480 1000 505
rect 1034 480 1050 514
rect 787 472 1050 480
rect 291 437 357 455
rect 205 424 257 428
rect 205 412 223 424
rect 205 378 214 412
rect 248 378 257 390
rect 205 344 257 378
rect 205 310 214 344
rect 248 310 257 344
rect 205 276 257 310
rect 205 242 214 276
rect 248 242 257 276
rect 205 226 257 242
rect 291 403 307 437
rect 341 403 357 437
rect 291 389 357 403
rect 503 439 587 455
rect 621 447 753 471
rect 537 426 587 439
rect 634 437 753 447
rect 537 422 592 426
rect 537 418 596 422
rect 537 412 603 418
rect 537 407 606 412
rect 537 405 610 407
rect 503 403 610 405
rect 503 389 685 403
rect 291 228 325 389
rect 561 387 685 389
rect 561 380 650 387
rect 409 355 455 356
rect 359 339 455 355
rect 359 305 365 339
rect 399 305 455 339
rect 503 339 537 355
rect 359 262 455 305
rect 489 305 503 310
rect 489 228 537 305
rect 291 194 322 228
rect 356 195 537 228
rect 571 353 650 380
rect 684 353 685 387
rect 571 315 685 353
rect 356 194 500 195
rect 26 137 171 166
rect 26 103 42 137
rect 76 132 171 137
rect 206 137 256 166
rect 76 103 92 132
rect 26 74 92 103
rect 240 103 256 137
rect 291 160 374 194
rect 571 161 607 315
rect 719 274 753 437
rect 291 126 322 160
rect 356 126 374 160
rect 291 110 374 126
rect 410 126 426 160
rect 460 126 476 160
rect 206 17 256 103
rect 410 17 476 126
rect 510 127 526 161
rect 560 127 607 161
rect 510 85 607 127
rect 641 240 753 274
rect 641 197 699 240
rect 787 206 821 472
rect 923 464 1050 472
rect 1096 535 1162 649
rect 1096 501 1112 535
rect 1146 501 1162 535
rect 1096 467 1162 501
rect 675 163 699 197
rect 641 119 699 163
rect 733 189 821 206
rect 733 155 741 189
rect 775 155 821 189
rect 855 409 889 425
rect 855 215 889 375
rect 923 315 957 464
rect 1096 433 1112 467
rect 1146 433 1162 467
rect 991 424 1057 430
rect 1025 409 1057 424
rect 991 375 1007 390
rect 1041 375 1057 409
rect 991 359 1057 375
rect 1096 399 1162 433
rect 1096 365 1112 399
rect 1146 365 1162 399
rect 1096 349 1162 365
rect 1196 535 1262 551
rect 1196 501 1212 535
rect 1246 501 1262 535
rect 1196 423 1262 501
rect 1196 389 1212 423
rect 1246 389 1262 423
rect 1196 373 1262 389
rect 1296 545 1527 561
rect 1296 511 1312 545
rect 1346 511 1391 545
rect 1425 511 1527 545
rect 1296 495 1527 511
rect 923 299 1130 315
rect 923 281 1080 299
rect 1038 265 1080 281
rect 1114 265 1130 299
rect 1038 257 1130 265
rect 1196 226 1230 373
rect 1296 337 1330 495
rect 1164 215 1230 226
rect 855 188 1230 215
rect 855 181 1180 188
rect 733 119 821 155
rect 1164 154 1180 181
rect 1214 154 1230 188
rect 862 113 1130 147
rect 1164 133 1230 154
rect 1264 303 1330 337
rect 1393 445 1459 461
rect 1393 411 1409 445
rect 1443 411 1459 445
rect 1264 169 1298 303
rect 1393 269 1459 411
rect 1493 337 1527 495
rect 1561 552 1627 649
rect 1561 518 1577 552
rect 1611 518 1627 552
rect 1561 489 1627 518
rect 1664 552 1737 581
rect 1664 518 1680 552
rect 1714 518 1737 552
rect 1664 489 1737 518
rect 1561 435 1669 451
rect 1561 424 1619 435
rect 1561 390 1567 424
rect 1601 401 1619 424
rect 1653 401 1669 435
rect 1601 390 1669 401
rect 1561 384 1669 390
rect 1703 405 1737 489
rect 1771 565 1837 649
rect 1771 531 1787 565
rect 1821 531 1837 565
rect 1771 489 1837 531
rect 1771 455 1787 489
rect 1821 455 1837 489
rect 1771 439 1837 455
rect 1877 565 1911 581
rect 1877 455 1911 531
rect 1703 371 1838 405
rect 1493 321 1770 337
rect 1493 303 1720 321
rect 1704 287 1720 303
rect 1754 287 1770 321
rect 1704 271 1770 287
rect 1338 253 1484 269
rect 1338 219 1354 253
rect 1388 219 1484 253
rect 1338 203 1484 219
rect 1518 253 1584 269
rect 1518 219 1534 253
rect 1568 237 1584 253
rect 1804 237 1838 371
rect 1877 343 1911 421
rect 1945 580 2085 596
rect 1945 546 2035 580
rect 2069 546 2085 580
rect 1945 503 2085 546
rect 1945 469 2035 503
rect 2069 469 2085 503
rect 1945 427 2085 469
rect 1945 393 2035 427
rect 2069 393 2085 427
rect 1945 377 2085 393
rect 1877 327 1987 343
rect 1877 293 1937 327
rect 1971 293 1987 327
rect 1877 277 1987 293
rect 1568 219 1838 237
rect 1518 203 1838 219
rect 1264 153 1416 169
rect 1264 119 1280 153
rect 1314 119 1366 153
rect 1400 119 1416 153
rect 862 85 896 113
rect 510 51 896 85
rect 1096 85 1130 113
rect 1450 85 1484 203
rect 983 45 1005 79
rect 1039 45 1062 79
rect 1096 51 1484 85
rect 1549 140 1615 169
rect 1549 106 1565 140
rect 1599 106 1615 140
rect 983 17 1062 45
rect 1549 17 1615 106
rect 1723 140 1789 203
rect 1723 106 1739 140
rect 1773 106 1789 140
rect 1723 77 1789 106
rect 1835 136 1885 169
rect 1835 102 1851 136
rect 1835 17 1885 102
rect 1921 146 1987 277
rect 1921 112 1937 146
rect 1971 112 1987 146
rect 1921 70 1987 112
rect 2033 226 2085 377
rect 2119 580 2185 649
rect 2119 546 2135 580
rect 2169 546 2185 580
rect 2119 497 2185 546
rect 2119 463 2135 497
rect 2169 463 2185 497
rect 2119 414 2185 463
rect 2119 380 2135 414
rect 2169 380 2185 414
rect 2119 364 2185 380
rect 2033 210 2099 226
rect 2033 176 2049 210
rect 2083 176 2099 210
rect 2033 120 2099 176
rect 2033 86 2049 120
rect 2083 86 2099 120
rect 2033 70 2099 86
rect 2135 210 2185 226
rect 2169 176 2185 210
rect 2135 120 2185 176
rect 2169 86 2185 120
rect 2135 17 2185 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 223 412 257 424
rect 223 390 248 412
rect 248 390 257 412
rect 991 409 1025 424
rect 991 390 1007 409
rect 1007 390 1025 409
rect 1567 390 1601 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
<< metal1 >>
rect 0 683 2208 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 0 617 2208 649
rect 211 424 269 430
rect 211 390 223 424
rect 257 421 269 424
rect 979 424 1037 430
rect 979 421 991 424
rect 257 393 991 421
rect 257 390 269 393
rect 211 384 269 390
rect 979 390 991 393
rect 1025 421 1037 424
rect 1555 424 1613 430
rect 1555 421 1567 424
rect 1025 393 1567 421
rect 1025 390 1037 393
rect 979 384 1037 390
rect 1555 390 1567 393
rect 1601 390 1613 424
rect 1555 384 1613 390
rect 0 17 2208 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
rect 0 -49 2208 -17
<< labels >>
flabel pwell s 0 0 2208 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 2208 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel comment s 940 630 940 630 0 FreeSans 300 0 0 0 no_jumper_check
flabel comment s 540 36 540 36 0 FreeSans 300 0 0 0 no_jumper_check
rlabel comment s 0 0 0 0 4 dfrtp_1
flabel metal1 s 223 390 257 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew
flabel metal1 s 0 617 2208 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 2208 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 1951 390 1985 424 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 1951 464 1985 498 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 1951 538 1985 572 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 31 390 65 424 0 FreeSans 340 0 0 0 D
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 2208 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 2884472
string GDS_START 2867466
<< end >>
