magic
tech sky130A
magscale 1 2
timestamp 1599588238
<< locali >>
rect 23 260 89 356
rect 191 88 263 310
rect 305 88 371 310
rect 409 236 485 310
rect 567 226 647 430
rect 558 154 647 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 23 390 89 649
rect 123 378 197 596
rect 243 412 309 649
rect 353 498 419 596
rect 460 532 526 649
rect 674 532 745 649
rect 353 464 747 498
rect 353 378 419 464
rect 123 344 419 378
rect 123 226 157 344
rect 52 192 157 226
rect 52 70 118 192
rect 681 260 747 464
rect 453 17 519 202
rect 681 120 731 216
rect 644 17 731 120
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel locali s 23 260 89 356 6 A
port 1 nsew signal input
rlabel locali s 191 88 263 310 6 B
port 2 nsew signal input
rlabel locali s 305 88 371 310 6 C
port 3 nsew signal input
rlabel locali s 409 236 485 310 6 D
port 4 nsew signal input
rlabel locali s 567 226 647 430 6 X
port 5 nsew signal output
rlabel locali s 558 154 647 226 6 X
port 5 nsew signal output
rlabel metal1 s 0 -49 768 49 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 617 768 715 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3220954
string GDS_START 3213750
<< end >>
