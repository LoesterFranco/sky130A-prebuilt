magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 23 426 89 596
rect 223 426 331 547
rect 23 392 331 426
rect 25 224 119 358
rect 197 224 263 358
rect 297 356 331 392
rect 297 190 359 356
rect 395 224 461 358
rect 505 224 575 358
rect 631 224 743 358
rect 777 236 843 356
rect 28 156 672 190
rect 28 70 94 156
rect 505 66 672 156
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 123 581 531 615
rect 123 460 189 581
rect 365 426 431 547
rect 465 460 531 581
rect 565 426 631 596
rect 665 460 731 649
rect 775 426 841 596
rect 365 392 841 426
rect 192 17 436 120
rect 770 17 836 190
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel locali s 631 224 743 358 6 A1
port 1 nsew signal input
rlabel locali s 777 236 843 356 6 A2
port 2 nsew signal input
rlabel locali s 505 224 575 358 6 B1
port 3 nsew signal input
rlabel locali s 395 224 461 358 6 B2
port 4 nsew signal input
rlabel locali s 25 224 119 358 6 C1
port 5 nsew signal input
rlabel locali s 197 224 263 358 6 C2
port 6 nsew signal input
rlabel locali s 505 66 672 156 6 Y
port 7 nsew signal output
rlabel locali s 297 356 331 392 6 Y
port 7 nsew signal output
rlabel locali s 297 190 359 356 6 Y
port 7 nsew signal output
rlabel locali s 223 426 331 547 6 Y
port 7 nsew signal output
rlabel locali s 28 156 672 190 6 Y
port 7 nsew signal output
rlabel locali s 28 70 94 156 6 Y
port 7 nsew signal output
rlabel locali s 23 426 89 596 6 Y
port 7 nsew signal output
rlabel locali s 23 392 331 426 6 Y
port 7 nsew signal output
rlabel metal1 s 0 -49 864 49 8 VGND
port 8 nsew ground bidirectional
rlabel metal1 s 0 617 864 715 6 VPWR
port 9 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3664144
string GDS_START 3655310
<< end >>
