magic
tech sky130A
magscale 1 2
timestamp 1599588238
<< locali >>
rect 121 394 161 596
rect 291 394 357 596
rect 121 360 357 394
rect 121 282 155 360
rect 25 236 155 282
rect 505 290 647 356
rect 109 226 155 236
rect 109 192 361 226
rect 109 70 159 192
rect 295 70 361 192
rect 981 224 1047 358
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 21 364 87 649
rect 201 428 251 649
rect 397 388 447 649
rect 486 424 552 596
rect 592 458 642 649
rect 685 581 931 615
rect 685 424 735 581
rect 486 390 735 424
rect 685 383 735 390
rect 189 260 429 326
rect 775 290 825 547
rect 865 389 931 581
rect 975 392 1041 649
rect 395 256 429 260
rect 701 256 825 290
rect 859 289 925 355
rect 23 17 73 202
rect 395 222 751 256
rect 195 17 261 153
rect 395 17 461 188
rect 495 70 561 222
rect 601 17 667 188
rect 701 70 751 222
rect 787 17 853 206
rect 887 190 925 289
rect 1081 190 1131 596
rect 887 70 1131 190
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
rlabel locali s 505 290 647 356 6 A
port 1 nsew signal input
rlabel locali s 981 224 1047 358 6 B_N
port 2 nsew signal input
rlabel locali s 295 70 361 192 6 X
port 3 nsew signal output
rlabel locali s 291 394 357 596 6 X
port 3 nsew signal output
rlabel locali s 121 394 161 596 6 X
port 3 nsew signal output
rlabel locali s 121 360 357 394 6 X
port 3 nsew signal output
rlabel locali s 121 282 155 360 6 X
port 3 nsew signal output
rlabel locali s 109 226 155 236 6 X
port 3 nsew signal output
rlabel locali s 109 192 361 226 6 X
port 3 nsew signal output
rlabel locali s 109 70 159 192 6 X
port 3 nsew signal output
rlabel locali s 25 236 155 282 6 X
port 3 nsew signal output
rlabel metal1 s 0 -49 1152 49 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1152 715 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 997636
string GDS_START 987470
<< end >>
