magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 210 401 286 493
rect 210 367 438 401
rect 18 215 84 263
rect 118 215 237 263
rect 364 109 438 367
rect 272 51 438 109
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 126 367 176 527
rect 330 435 373 527
rect 18 333 74 365
rect 18 299 324 333
rect 290 181 324 299
rect 18 147 324 181
rect 18 105 72 147
rect 126 17 192 109
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
rlabel locali s 18 215 84 263 6 A_N
port 1 nsew signal input
rlabel locali s 118 215 237 263 6 B
port 2 nsew signal input
rlabel locali s 364 109 438 367 6 Y
port 3 nsew signal output
rlabel locali s 272 51 438 109 6 Y
port 3 nsew signal output
rlabel locali s 210 401 286 493 6 Y
port 3 nsew signal output
rlabel locali s 210 367 438 401 6 Y
port 3 nsew signal output
rlabel metal1 s 0 -48 460 48 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 496 460 592 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 460 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2222346
string GDS_START 2217752
<< end >>
