magic
tech sky130A
magscale 1 2
timestamp 1601050088
<< locali >>
rect 21 236 155 310
rect 209 270 275 356
rect 391 364 462 596
rect 428 226 462 364
rect 391 70 462 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 59 424 125 540
rect 233 458 357 649
rect 59 390 357 424
rect 59 364 125 390
rect 323 326 357 390
rect 323 260 394 326
rect 323 236 357 260
rect 189 202 357 236
rect 59 17 130 199
rect 189 108 248 202
rect 291 17 357 168
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< metal1 >>
rect 0 683 480 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 0 617 480 649
rect 0 17 480 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
rect 0 -49 480 -17
<< labels >>
rlabel locali s 209 270 275 356 6 A
port 1 nsew signal input
rlabel locali s 21 236 155 310 6 B
port 2 nsew signal input
rlabel locali s 428 226 462 364 6 X
port 3 nsew signal output
rlabel locali s 391 364 462 596 6 X
port 3 nsew signal output
rlabel locali s 391 70 462 226 6 X
port 3 nsew signal output
rlabel metal1 s 0 -49 480 49 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 617 480 715 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 480 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 743660
string GDS_START 738986
<< end >>
