magic
tech sky130A
magscale 1 2
timestamp 1601050088
<< locali >>
rect 105 294 263 360
rect 299 294 365 360
rect 595 404 645 547
rect 595 370 857 404
rect 823 356 857 370
rect 823 310 935 356
rect 1081 327 1223 356
rect 823 236 857 310
rect 972 270 1223 327
rect 1262 270 1415 356
rect 791 202 1315 236
rect 791 168 857 202
rect 578 134 857 168
rect 578 70 644 134
rect 791 70 857 134
rect 993 70 1043 202
rect 1265 70 1315 202
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 23 394 89 596
rect 123 394 343 649
rect 377 428 443 596
rect 499 581 745 615
rect 377 394 465 428
rect 23 260 57 394
rect 431 336 465 394
rect 499 370 555 581
rect 679 472 745 581
rect 779 581 1137 615
rect 779 506 835 581
rect 869 472 935 547
rect 679 438 935 472
rect 981 424 1031 547
rect 1071 458 1137 581
rect 1171 424 1237 596
rect 1277 458 1311 649
rect 1351 424 1417 596
rect 981 390 1417 424
rect 981 364 1031 390
rect 431 270 633 336
rect 723 270 789 336
rect 431 260 465 270
rect 23 226 163 260
rect 97 176 163 226
rect 324 210 465 260
rect 723 236 757 270
rect 499 202 757 236
rect 499 176 533 202
rect 97 142 533 176
rect 97 72 163 142
rect 198 17 303 108
rect 439 17 542 108
rect 680 17 755 100
rect 891 17 957 168
rect 1077 17 1231 168
rect 1351 17 1417 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 683 1440 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 0 617 1440 649
rect 0 17 1440 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -49 1440 -17
<< labels >>
rlabel locali s 1262 270 1415 356 6 A
port 1 nsew signal input
rlabel locali s 1081 327 1223 356 6 B
port 2 nsew signal input
rlabel locali s 972 270 1223 327 6 B
port 2 nsew signal input
rlabel locali s 105 294 263 360 6 C_N
port 3 nsew signal input
rlabel locali s 299 294 365 360 6 D_N
port 4 nsew signal input
rlabel locali s 1265 70 1315 202 6 Y
port 5 nsew signal output
rlabel locali s 993 70 1043 202 6 Y
port 5 nsew signal output
rlabel locali s 823 356 857 370 6 Y
port 5 nsew signal output
rlabel locali s 823 310 935 356 6 Y
port 5 nsew signal output
rlabel locali s 823 236 857 310 6 Y
port 5 nsew signal output
rlabel locali s 791 202 1315 236 6 Y
port 5 nsew signal output
rlabel locali s 791 168 857 202 6 Y
port 5 nsew signal output
rlabel locali s 791 70 857 134 6 Y
port 5 nsew signal output
rlabel locali s 595 404 645 547 6 Y
port 5 nsew signal output
rlabel locali s 595 370 857 404 6 Y
port 5 nsew signal output
rlabel locali s 578 134 857 168 6 Y
port 5 nsew signal output
rlabel locali s 578 70 644 134 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -49 1440 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 1440 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1440 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1573848
string GDS_START 1562212
<< end >>
