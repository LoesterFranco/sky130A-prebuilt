magic
tech sky130A
magscale 1 2
timestamp 1604502697
<< nwell >>
rect -38 261 2154 582
<< pwell >>
rect 47 -17 81 17
<< scnmos >>
rect 89 47 119 177
rect 183 47 213 177
rect 277 47 307 177
rect 371 47 401 177
rect 518 93 548 177
rect 722 49 752 177
rect 842 49 872 177
rect 1124 47 1154 177
rect 1320 49 1350 177
rect 1482 49 1512 133
rect 1641 49 1671 177
rect 1781 47 1811 167
rect 1891 47 1921 175
rect 1993 47 2023 175
<< pmoshvt >>
rect 101 297 137 497
rect 195 297 231 497
rect 289 297 325 497
rect 383 297 419 497
rect 492 297 528 425
rect 706 325 742 493
rect 822 325 858 493
rect 1073 297 1109 497
rect 1312 297 1348 465
rect 1474 297 1510 425
rect 1659 329 1695 457
rect 1772 329 1808 497
rect 1883 297 1919 497
rect 1985 297 2021 497
<< ndiff >>
rect 27 93 89 177
rect 27 59 35 93
rect 69 59 89 93
rect 27 47 89 59
rect 119 129 183 177
rect 119 95 129 129
rect 163 95 183 129
rect 119 47 183 95
rect 213 93 277 177
rect 213 59 223 93
rect 257 59 277 93
rect 213 47 277 59
rect 307 129 371 177
rect 307 95 317 129
rect 351 95 371 129
rect 307 47 371 95
rect 401 93 518 177
rect 548 169 604 177
rect 548 135 558 169
rect 592 135 604 169
rect 548 93 604 135
rect 658 165 722 177
rect 658 131 668 165
rect 702 131 722 165
rect 401 89 493 93
rect 401 55 411 89
rect 445 55 493 89
rect 401 47 493 55
rect 658 49 722 131
rect 752 91 842 177
rect 752 57 762 91
rect 796 57 842 91
rect 752 49 842 57
rect 872 169 971 177
rect 872 135 924 169
rect 958 135 971 169
rect 872 49 971 135
rect 1052 161 1124 177
rect 1052 127 1060 161
rect 1094 127 1124 161
rect 1052 93 1124 127
rect 1052 59 1060 93
rect 1094 59 1124 93
rect 1052 47 1124 59
rect 1154 161 1206 177
rect 1154 127 1164 161
rect 1198 127 1206 161
rect 1154 121 1206 127
rect 1154 47 1204 121
rect 1260 105 1320 177
rect 1258 97 1320 105
rect 1258 63 1266 97
rect 1300 63 1320 97
rect 1258 49 1320 63
rect 1350 133 1451 177
rect 1537 169 1641 177
rect 1537 135 1583 169
rect 1617 135 1641 169
rect 1537 133 1641 135
rect 1350 126 1482 133
rect 1350 92 1360 126
rect 1394 92 1482 126
rect 1350 49 1482 92
rect 1512 49 1641 133
rect 1671 167 1731 177
rect 1831 167 1891 175
rect 1671 93 1781 167
rect 1671 59 1693 93
rect 1727 59 1781 93
rect 1671 49 1781 59
rect 1698 47 1781 49
rect 1811 142 1891 167
rect 1811 108 1837 142
rect 1871 108 1891 142
rect 1811 47 1891 108
rect 1921 97 1993 175
rect 1921 63 1939 97
rect 1973 63 1993 97
rect 1921 47 1993 63
rect 2023 101 2075 175
rect 2023 67 2033 101
rect 2067 67 2075 101
rect 2023 47 2075 67
<< pdiff >>
rect 47 477 101 497
rect 47 443 55 477
rect 89 443 101 477
rect 47 297 101 443
rect 137 477 195 497
rect 137 443 149 477
rect 183 443 195 477
rect 137 409 195 443
rect 137 375 149 409
rect 183 375 195 409
rect 137 341 195 375
rect 137 307 149 341
rect 183 307 195 341
rect 137 297 195 307
rect 231 477 289 497
rect 231 443 243 477
rect 277 443 289 477
rect 231 297 289 443
rect 325 477 383 497
rect 325 443 337 477
rect 371 443 383 477
rect 325 409 383 443
rect 325 375 337 409
rect 371 375 383 409
rect 325 341 383 375
rect 325 307 337 341
rect 371 307 383 341
rect 325 297 383 307
rect 419 477 473 497
rect 419 443 431 477
rect 465 443 473 477
rect 419 425 473 443
rect 419 297 492 425
rect 528 341 594 425
rect 528 307 548 341
rect 582 307 594 341
rect 652 413 706 493
rect 652 379 660 413
rect 694 379 706 413
rect 652 325 706 379
rect 742 481 822 493
rect 742 447 763 481
rect 797 447 822 481
rect 742 325 822 447
rect 858 481 965 493
rect 858 447 920 481
rect 954 447 965 481
rect 858 325 965 447
rect 1019 481 1073 497
rect 1019 447 1027 481
rect 1061 447 1073 481
rect 528 297 594 307
rect 1019 297 1073 447
rect 1109 349 1171 497
rect 1712 489 1772 497
rect 1225 405 1312 465
rect 1225 371 1233 405
rect 1267 371 1312 405
rect 1225 365 1312 371
rect 1109 343 1173 349
rect 1109 309 1121 343
rect 1155 309 1173 343
rect 1109 297 1173 309
rect 1227 297 1312 365
rect 1348 425 1450 465
rect 1712 457 1724 489
rect 1572 425 1659 457
rect 1348 409 1474 425
rect 1348 375 1401 409
rect 1435 375 1474 409
rect 1348 341 1474 375
rect 1348 307 1401 341
rect 1435 307 1474 341
rect 1348 297 1474 307
rect 1510 421 1659 425
rect 1510 387 1613 421
rect 1647 387 1659 421
rect 1510 329 1659 387
rect 1695 455 1724 457
rect 1758 455 1772 489
rect 1695 329 1772 455
rect 1808 341 1883 497
rect 1808 329 1837 341
rect 1510 297 1607 329
rect 1825 307 1837 329
rect 1871 307 1883 341
rect 1825 297 1883 307
rect 1919 489 1985 497
rect 1919 455 1939 489
rect 1973 455 1985 489
rect 1919 297 1985 455
rect 2021 477 2075 497
rect 2021 443 2033 477
rect 2067 443 2075 477
rect 2021 409 2075 443
rect 2021 375 2033 409
rect 2067 375 2075 409
rect 2021 297 2075 375
<< ndiffc >>
rect 35 59 69 93
rect 129 95 163 129
rect 223 59 257 93
rect 317 95 351 129
rect 558 135 592 169
rect 668 131 702 165
rect 411 55 445 89
rect 762 57 796 91
rect 924 135 958 169
rect 1060 127 1094 161
rect 1060 59 1094 93
rect 1164 127 1198 161
rect 1266 63 1300 97
rect 1583 135 1617 169
rect 1360 92 1394 126
rect 1693 59 1727 93
rect 1837 108 1871 142
rect 1939 63 1973 97
rect 2033 67 2067 101
<< pdiffc >>
rect 55 443 89 477
rect 149 443 183 477
rect 149 375 183 409
rect 149 307 183 341
rect 243 443 277 477
rect 337 443 371 477
rect 337 375 371 409
rect 337 307 371 341
rect 431 443 465 477
rect 548 307 582 341
rect 660 379 694 413
rect 763 447 797 481
rect 920 447 954 481
rect 1027 447 1061 481
rect 1233 371 1267 405
rect 1121 309 1155 343
rect 1401 375 1435 409
rect 1401 307 1435 341
rect 1613 387 1647 421
rect 1724 455 1758 489
rect 1837 307 1871 341
rect 1939 455 1973 489
rect 2033 443 2067 477
rect 2033 375 2067 409
<< poly >>
rect 101 497 137 523
rect 195 497 231 523
rect 289 497 325 523
rect 383 497 419 523
rect 706 493 742 519
rect 822 493 858 519
rect 1073 497 1109 523
rect 490 451 530 483
rect 492 425 528 451
rect 706 310 742 325
rect 822 310 858 325
rect 101 282 137 297
rect 195 282 231 297
rect 289 282 325 297
rect 383 282 419 297
rect 492 282 528 297
rect 99 265 139 282
rect 193 265 233 282
rect 287 265 327 282
rect 381 265 421 282
rect 490 265 530 282
rect 704 271 744 310
rect 704 265 753 271
rect 820 265 860 310
rect 1310 493 1697 523
rect 1772 497 1808 523
rect 1883 497 1919 523
rect 1985 497 2021 523
rect 1310 491 1350 493
rect 1312 465 1348 491
rect 1657 483 1697 493
rect 1659 457 1695 483
rect 1474 425 1510 451
rect 1659 314 1695 329
rect 1772 314 1808 329
rect 1073 282 1109 297
rect 1312 282 1348 297
rect 1474 282 1510 297
rect 80 249 448 265
rect 80 215 404 249
rect 438 215 448 249
rect 80 207 448 215
rect 89 199 448 207
rect 490 249 753 265
rect 490 215 631 249
rect 665 215 699 249
rect 733 215 753 249
rect 490 199 753 215
rect 808 249 872 265
rect 808 215 818 249
rect 852 215 872 249
rect 1071 247 1111 282
rect 1310 247 1350 282
rect 1472 265 1512 282
rect 1657 265 1697 314
rect 1071 217 1350 247
rect 808 199 872 215
rect 89 177 119 199
rect 183 177 213 199
rect 277 177 307 199
rect 371 177 401 199
rect 518 177 548 199
rect 722 197 753 199
rect 722 177 752 197
rect 842 177 872 199
rect 1124 177 1154 217
rect 1320 177 1350 217
rect 1392 249 1512 265
rect 1392 215 1402 249
rect 1436 215 1512 249
rect 1392 199 1512 215
rect 518 67 548 93
rect 89 21 119 47
rect 183 21 213 47
rect 277 21 307 47
rect 371 21 401 47
rect 722 21 752 49
rect 842 21 872 49
rect 1482 133 1512 199
rect 1641 249 1705 265
rect 1770 256 1810 314
rect 1883 282 1919 297
rect 1985 282 2021 297
rect 1881 265 1921 282
rect 1983 265 2023 282
rect 1770 255 1811 256
rect 1641 215 1651 249
rect 1685 215 1705 249
rect 1641 199 1705 215
rect 1747 239 1811 255
rect 1747 205 1757 239
rect 1791 205 1811 239
rect 1641 177 1671 199
rect 1747 189 1811 205
rect 1853 249 1921 265
rect 1853 215 1863 249
rect 1897 215 1921 249
rect 1853 199 1921 215
rect 1963 249 2027 265
rect 1963 215 1973 249
rect 2007 215 2027 249
rect 1963 199 2027 215
rect 1781 167 1811 189
rect 1891 175 1921 199
rect 1993 175 2023 199
rect 1124 21 1154 47
rect 1320 21 1350 49
rect 1482 23 1512 49
rect 1641 21 1671 49
rect 1781 21 1811 47
rect 1891 21 1921 47
rect 1993 21 2023 47
<< polycont >>
rect 404 215 438 249
rect 631 215 665 249
rect 699 215 733 249
rect 818 215 852 249
rect 1402 215 1436 249
rect 1651 215 1685 249
rect 1757 205 1791 239
rect 1863 215 1897 249
rect 1973 215 2007 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 55 477 89 527
rect 55 427 89 443
rect 149 477 183 493
rect 227 477 293 527
rect 227 443 243 477
rect 277 443 293 477
rect 337 477 371 493
rect 415 477 481 527
rect 1011 481 1077 527
rect 1923 489 1989 527
rect 415 443 431 477
rect 465 443 481 477
rect 515 447 763 481
rect 797 447 843 481
rect 896 447 920 481
rect 954 447 977 481
rect 1011 447 1027 481
rect 1061 447 1077 481
rect 1164 455 1724 489
rect 1758 455 1823 489
rect 1923 455 1939 489
rect 1973 455 1989 489
rect 2033 477 2085 493
rect 149 409 183 443
rect 337 409 371 443
rect 515 409 559 447
rect 943 413 977 447
rect 1164 413 1198 455
rect 183 375 337 409
rect 149 341 371 375
rect 183 307 337 341
rect 149 291 371 307
rect 415 375 559 409
rect 628 379 660 413
rect 694 379 909 413
rect 943 379 1198 413
rect 1233 405 1267 421
rect 149 288 314 291
rect 241 185 314 288
rect 415 265 449 375
rect 514 307 548 341
rect 582 307 831 341
rect 404 249 449 265
rect 438 215 449 249
rect 404 193 449 215
rect 129 132 351 185
rect 415 173 449 193
rect 415 139 513 173
rect 129 129 163 132
rect 35 93 69 109
rect 129 70 163 95
rect 317 129 351 132
rect 35 17 69 59
rect 197 59 223 93
rect 257 59 273 93
rect 317 70 351 95
rect 411 89 445 105
rect 197 17 273 59
rect 411 17 445 55
rect 479 85 513 139
rect 558 169 592 307
rect 797 265 831 307
rect 875 339 909 379
rect 875 323 981 339
rect 875 305 947 323
rect 924 289 947 305
rect 924 275 981 289
rect 626 249 763 265
rect 626 215 631 249
rect 665 215 699 249
rect 733 215 763 249
rect 626 199 763 215
rect 797 249 881 265
rect 797 215 818 249
rect 852 215 881 249
rect 797 199 881 215
rect 924 169 958 275
rect 1015 241 1049 379
rect 1095 309 1121 343
rect 1155 309 1198 343
rect 1095 289 1198 309
rect 558 119 592 135
rect 648 131 668 165
rect 702 131 890 165
rect 732 85 762 91
rect 479 57 762 85
rect 796 57 812 91
rect 479 51 812 57
rect 846 85 890 131
rect 924 119 958 135
rect 992 210 1049 241
rect 992 209 1048 210
rect 992 208 1046 209
rect 992 207 1043 208
rect 992 85 1026 207
rect 1140 187 1198 289
rect 846 51 1026 85
rect 1060 161 1094 177
rect 1060 93 1094 127
rect 1140 153 1141 187
rect 1175 161 1198 187
rect 1140 127 1164 153
rect 1140 83 1198 127
rect 1233 119 1267 371
rect 1305 178 1339 455
rect 2067 443 2085 477
rect 2033 421 2085 443
rect 1383 375 1401 409
rect 1435 375 1466 409
rect 1383 341 1466 375
rect 1383 307 1401 341
rect 1435 323 1466 341
rect 1583 387 1613 421
rect 1647 409 2085 421
rect 1647 387 2033 409
rect 1435 307 1437 323
rect 1383 289 1437 307
rect 1471 289 1549 323
rect 1386 249 1471 254
rect 1386 215 1402 249
rect 1436 215 1471 249
rect 1386 199 1471 215
rect 1428 187 1471 199
rect 1305 165 1355 178
rect 1305 144 1394 165
rect 1311 131 1394 144
rect 1360 126 1394 131
rect 1428 153 1437 187
rect 1428 126 1471 153
rect 1233 85 1243 119
rect 1060 17 1094 59
rect 1233 63 1266 85
rect 1300 63 1316 97
rect 1360 64 1394 92
rect 1515 85 1549 289
rect 1583 169 1617 387
rect 1978 375 2033 387
rect 2067 375 2085 409
rect 1651 289 1728 323
rect 1821 307 1837 341
rect 1871 307 1995 341
rect 1821 299 1995 307
rect 1651 249 1695 289
rect 1961 265 1995 299
rect 1685 215 1695 249
rect 1651 199 1695 215
rect 1729 239 1791 255
rect 1729 205 1757 239
rect 1835 249 1927 265
rect 1835 215 1863 249
rect 1897 215 1927 249
rect 1961 249 2007 265
rect 1961 215 1973 249
rect 1729 189 1791 205
rect 1961 199 2007 215
rect 1729 187 1770 189
rect 1729 153 1733 187
rect 1767 153 1770 187
rect 1961 181 1995 199
rect 1729 146 1770 153
rect 1837 150 1995 181
rect 1829 147 1995 150
rect 1583 119 1617 135
rect 1829 142 1887 147
rect 1829 119 1837 142
rect 1651 85 1693 93
rect 1233 53 1316 63
rect 1515 59 1693 85
rect 1727 59 1754 93
rect 1829 85 1835 119
rect 1871 108 1887 142
rect 2051 117 2085 375
rect 1869 85 1887 108
rect 1829 59 1887 85
rect 1939 97 1973 113
rect 1515 51 1754 59
rect 1939 17 1973 63
rect 2033 101 2085 117
rect 2067 67 2085 101
rect 2033 51 2085 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 947 289 981 323
rect 1141 161 1175 187
rect 1141 153 1164 161
rect 1164 153 1175 161
rect 1437 289 1471 323
rect 1437 153 1471 187
rect 1243 97 1277 119
rect 1243 85 1266 97
rect 1266 85 1277 97
rect 1733 153 1767 187
rect 1835 108 1837 119
rect 1837 108 1869 119
rect 1835 85 1869 108
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
<< metal1 >>
rect 0 561 2116 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 0 496 2116 527
rect 935 323 993 329
rect 935 289 947 323
rect 981 320 993 323
rect 1425 323 1483 329
rect 1425 320 1437 323
rect 981 292 1437 320
rect 981 289 993 292
rect 935 283 993 289
rect 1425 289 1437 292
rect 1471 289 1483 323
rect 1425 283 1483 289
rect 1129 187 1197 193
rect 1129 153 1141 187
rect 1175 184 1197 187
rect 1425 187 1483 193
rect 1425 184 1437 187
rect 1175 156 1437 184
rect 1175 153 1197 156
rect 1129 147 1197 153
rect 1425 153 1437 156
rect 1471 184 1483 187
rect 1721 187 1779 193
rect 1721 184 1733 187
rect 1471 156 1733 184
rect 1471 153 1483 156
rect 1425 147 1483 153
rect 1721 153 1733 156
rect 1767 153 1779 187
rect 1721 147 1779 153
rect 1231 119 1289 125
rect 1231 85 1243 119
rect 1277 116 1289 119
rect 1823 119 1881 125
rect 1823 116 1835 119
rect 1277 88 1835 116
rect 1277 85 1289 88
rect 1231 79 1289 85
rect 1823 85 1835 88
rect 1869 85 1881 119
rect 1823 79 1881 85
rect 0 17 2116 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
rect 0 -48 2116 -17
<< labels >>
flabel corelocali s 209 374 209 374 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 673 221 707 255 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 1684 289 1718 323 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 1870 221 1904 255 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel pwell s 47 -17 81 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 47 527 81 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 44 0 44 0 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 46 544 46 544 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
rlabel comment s 0 0 0 0 4 hkscl5hdv1_xor3_1
flabel comment s 0 544 0 544 3 FreeSans 200 0 0 0 HHNEC
<< properties >>
string FIXED_BBOX 0 0 2116 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 820024
string GDS_START 806038
<< end >>
