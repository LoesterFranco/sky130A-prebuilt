magic
tech sky130A
magscale 1 2
timestamp 1601050047
<< nwell >>
rect -38 332 2054 704
<< pwell >>
rect 0 0 2016 49
<< scpmos >>
rect 84 368 114 592
rect 174 368 204 592
rect 264 368 294 592
rect 354 368 384 592
rect 444 368 474 592
rect 534 368 564 592
rect 624 368 654 592
rect 714 368 744 592
rect 804 368 834 592
rect 894 368 924 592
rect 984 368 1014 592
rect 1074 368 1104 592
rect 1272 368 1302 592
rect 1362 368 1392 592
rect 1452 368 1482 592
rect 1542 368 1572 592
rect 1632 368 1662 592
rect 1722 368 1752 592
rect 1812 368 1842 592
rect 1902 368 1932 592
<< nmoslvt >>
rect 84 74 114 222
rect 170 74 200 222
rect 258 74 288 222
rect 344 74 374 222
rect 430 74 460 222
rect 516 74 546 222
rect 621 74 651 222
rect 716 74 746 222
rect 914 74 944 222
rect 1000 74 1030 222
rect 1086 74 1116 222
rect 1172 74 1202 222
rect 1258 74 1288 222
rect 1358 74 1388 222
rect 1444 74 1474 222
rect 1544 74 1574 222
rect 1630 74 1660 222
rect 1716 74 1746 222
rect 1802 74 1832 222
rect 1902 74 1932 222
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 136 170 222
rect 114 102 125 136
rect 159 102 170 136
rect 114 74 170 102
rect 200 210 258 222
rect 200 176 212 210
rect 246 176 258 210
rect 200 120 258 176
rect 200 86 212 120
rect 246 86 258 120
rect 200 74 258 86
rect 288 136 344 222
rect 288 102 299 136
rect 333 102 344 136
rect 288 74 344 102
rect 374 210 430 222
rect 374 176 385 210
rect 419 176 430 210
rect 374 120 430 176
rect 374 86 385 120
rect 419 86 430 120
rect 374 74 430 86
rect 460 181 516 222
rect 460 147 471 181
rect 505 147 516 181
rect 460 74 516 147
rect 546 136 621 222
rect 546 102 571 136
rect 605 102 621 136
rect 546 74 621 102
rect 651 189 716 222
rect 651 155 671 189
rect 705 155 716 189
rect 651 74 716 155
rect 746 210 803 222
rect 746 176 757 210
rect 791 176 803 210
rect 746 120 803 176
rect 746 86 757 120
rect 791 86 803 120
rect 746 74 803 86
rect 857 210 914 222
rect 857 176 869 210
rect 903 176 914 210
rect 857 120 914 176
rect 857 86 869 120
rect 903 86 914 120
rect 857 74 914 86
rect 944 189 1000 222
rect 944 155 955 189
rect 989 155 1000 189
rect 944 74 1000 155
rect 1030 131 1086 222
rect 1030 97 1041 131
rect 1075 97 1086 131
rect 1030 74 1086 97
rect 1116 189 1172 222
rect 1116 155 1127 189
rect 1161 155 1172 189
rect 1116 74 1172 155
rect 1202 210 1258 222
rect 1202 176 1213 210
rect 1247 176 1258 210
rect 1202 120 1258 176
rect 1202 86 1213 120
rect 1247 86 1258 120
rect 1202 74 1258 86
rect 1288 147 1358 222
rect 1288 113 1299 147
rect 1333 113 1358 147
rect 1288 74 1358 113
rect 1388 210 1444 222
rect 1388 176 1399 210
rect 1433 176 1444 210
rect 1388 120 1444 176
rect 1388 86 1399 120
rect 1433 86 1444 120
rect 1388 74 1444 86
rect 1474 147 1544 222
rect 1474 113 1485 147
rect 1519 113 1544 147
rect 1474 74 1544 113
rect 1574 210 1630 222
rect 1574 176 1585 210
rect 1619 176 1630 210
rect 1574 120 1630 176
rect 1574 86 1585 120
rect 1619 86 1630 120
rect 1574 74 1630 86
rect 1660 147 1716 222
rect 1660 113 1671 147
rect 1705 113 1716 147
rect 1660 74 1716 113
rect 1746 210 1802 222
rect 1746 176 1757 210
rect 1791 176 1802 210
rect 1746 120 1802 176
rect 1746 86 1757 120
rect 1791 86 1802 120
rect 1746 74 1802 86
rect 1832 147 1902 222
rect 1832 113 1857 147
rect 1891 113 1902 147
rect 1832 74 1902 113
rect 1932 210 1989 222
rect 1932 176 1943 210
rect 1977 176 1989 210
rect 1932 120 1989 176
rect 1932 86 1943 120
rect 1977 86 1989 120
rect 1932 74 1989 86
<< pdiff >>
rect 27 580 84 592
rect 27 546 37 580
rect 71 546 84 580
rect 27 510 84 546
rect 27 476 37 510
rect 71 476 84 510
rect 27 440 84 476
rect 27 406 37 440
rect 71 406 84 440
rect 27 368 84 406
rect 114 580 174 592
rect 114 546 127 580
rect 161 546 174 580
rect 114 505 174 546
rect 114 471 127 505
rect 161 471 174 505
rect 114 424 174 471
rect 114 390 127 424
rect 161 390 174 424
rect 114 368 174 390
rect 204 580 264 592
rect 204 546 217 580
rect 251 546 264 580
rect 204 508 264 546
rect 204 474 217 508
rect 251 474 264 508
rect 204 368 264 474
rect 294 580 354 592
rect 294 546 307 580
rect 341 546 354 580
rect 294 505 354 546
rect 294 471 307 505
rect 341 471 354 505
rect 294 424 354 471
rect 294 390 307 424
rect 341 390 354 424
rect 294 368 354 390
rect 384 580 444 592
rect 384 546 397 580
rect 431 546 444 580
rect 384 508 444 546
rect 384 474 397 508
rect 431 474 444 508
rect 384 368 444 474
rect 474 580 534 592
rect 474 546 487 580
rect 521 546 534 580
rect 474 505 534 546
rect 474 471 487 505
rect 521 471 534 505
rect 474 424 534 471
rect 474 390 487 424
rect 521 390 534 424
rect 474 368 534 390
rect 564 580 624 592
rect 564 546 577 580
rect 611 546 624 580
rect 564 508 624 546
rect 564 474 577 508
rect 611 474 624 508
rect 564 368 624 474
rect 654 580 714 592
rect 654 546 667 580
rect 701 546 714 580
rect 654 505 714 546
rect 654 471 667 505
rect 701 471 714 505
rect 654 424 714 471
rect 654 390 667 424
rect 701 390 714 424
rect 654 368 714 390
rect 744 580 804 592
rect 744 546 757 580
rect 791 546 804 580
rect 744 497 804 546
rect 744 463 757 497
rect 791 463 804 497
rect 744 414 804 463
rect 744 380 757 414
rect 791 380 804 414
rect 744 368 804 380
rect 834 580 894 592
rect 834 546 847 580
rect 881 546 894 580
rect 834 497 894 546
rect 834 463 847 497
rect 881 463 894 497
rect 834 414 894 463
rect 834 380 847 414
rect 881 380 894 414
rect 834 368 894 380
rect 924 580 984 592
rect 924 546 937 580
rect 971 546 984 580
rect 924 478 984 546
rect 924 444 937 478
rect 971 444 984 478
rect 924 368 984 444
rect 1014 580 1074 592
rect 1014 546 1027 580
rect 1061 546 1074 580
rect 1014 497 1074 546
rect 1014 463 1027 497
rect 1061 463 1074 497
rect 1014 414 1074 463
rect 1014 380 1027 414
rect 1061 380 1074 414
rect 1014 368 1074 380
rect 1104 580 1161 592
rect 1104 546 1117 580
rect 1151 546 1161 580
rect 1104 498 1161 546
rect 1104 464 1117 498
rect 1151 464 1161 498
rect 1104 368 1161 464
rect 1215 580 1272 592
rect 1215 546 1225 580
rect 1259 546 1272 580
rect 1215 508 1272 546
rect 1215 474 1225 508
rect 1259 474 1272 508
rect 1215 368 1272 474
rect 1302 537 1362 592
rect 1302 503 1315 537
rect 1349 503 1362 537
rect 1302 428 1362 503
rect 1302 394 1315 428
rect 1349 394 1362 428
rect 1302 368 1362 394
rect 1392 580 1452 592
rect 1392 546 1405 580
rect 1439 546 1452 580
rect 1392 508 1452 546
rect 1392 474 1405 508
rect 1439 474 1452 508
rect 1392 368 1452 474
rect 1482 537 1542 592
rect 1482 503 1495 537
rect 1529 503 1542 537
rect 1482 428 1542 503
rect 1482 394 1495 428
rect 1529 394 1542 428
rect 1482 368 1542 394
rect 1572 580 1632 592
rect 1572 546 1585 580
rect 1619 546 1632 580
rect 1572 510 1632 546
rect 1572 476 1585 510
rect 1619 476 1632 510
rect 1572 440 1632 476
rect 1572 406 1585 440
rect 1619 406 1632 440
rect 1572 368 1632 406
rect 1662 580 1722 592
rect 1662 546 1675 580
rect 1709 546 1722 580
rect 1662 508 1722 546
rect 1662 474 1675 508
rect 1709 474 1722 508
rect 1662 368 1722 474
rect 1752 580 1812 592
rect 1752 546 1765 580
rect 1799 546 1812 580
rect 1752 504 1812 546
rect 1752 470 1765 504
rect 1799 470 1812 504
rect 1752 424 1812 470
rect 1752 390 1765 424
rect 1799 390 1812 424
rect 1752 368 1812 390
rect 1842 580 1902 592
rect 1842 546 1855 580
rect 1889 546 1902 580
rect 1842 508 1902 546
rect 1842 474 1855 508
rect 1889 474 1902 508
rect 1842 368 1902 474
rect 1932 580 1989 592
rect 1932 546 1945 580
rect 1979 546 1989 580
rect 1932 504 1989 546
rect 1932 470 1945 504
rect 1979 470 1989 504
rect 1932 424 1989 470
rect 1932 390 1945 424
rect 1979 390 1989 424
rect 1932 368 1989 390
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 125 102 159 136
rect 212 176 246 210
rect 212 86 246 120
rect 299 102 333 136
rect 385 176 419 210
rect 385 86 419 120
rect 471 147 505 181
rect 571 102 605 136
rect 671 155 705 189
rect 757 176 791 210
rect 757 86 791 120
rect 869 176 903 210
rect 869 86 903 120
rect 955 155 989 189
rect 1041 97 1075 131
rect 1127 155 1161 189
rect 1213 176 1247 210
rect 1213 86 1247 120
rect 1299 113 1333 147
rect 1399 176 1433 210
rect 1399 86 1433 120
rect 1485 113 1519 147
rect 1585 176 1619 210
rect 1585 86 1619 120
rect 1671 113 1705 147
rect 1757 176 1791 210
rect 1757 86 1791 120
rect 1857 113 1891 147
rect 1943 176 1977 210
rect 1943 86 1977 120
<< pdiffc >>
rect 37 546 71 580
rect 37 476 71 510
rect 37 406 71 440
rect 127 546 161 580
rect 127 471 161 505
rect 127 390 161 424
rect 217 546 251 580
rect 217 474 251 508
rect 307 546 341 580
rect 307 471 341 505
rect 307 390 341 424
rect 397 546 431 580
rect 397 474 431 508
rect 487 546 521 580
rect 487 471 521 505
rect 487 390 521 424
rect 577 546 611 580
rect 577 474 611 508
rect 667 546 701 580
rect 667 471 701 505
rect 667 390 701 424
rect 757 546 791 580
rect 757 463 791 497
rect 757 380 791 414
rect 847 546 881 580
rect 847 463 881 497
rect 847 380 881 414
rect 937 546 971 580
rect 937 444 971 478
rect 1027 546 1061 580
rect 1027 463 1061 497
rect 1027 380 1061 414
rect 1117 546 1151 580
rect 1117 464 1151 498
rect 1225 546 1259 580
rect 1225 474 1259 508
rect 1315 503 1349 537
rect 1315 394 1349 428
rect 1405 546 1439 580
rect 1405 474 1439 508
rect 1495 503 1529 537
rect 1495 394 1529 428
rect 1585 546 1619 580
rect 1585 476 1619 510
rect 1585 406 1619 440
rect 1675 546 1709 580
rect 1675 474 1709 508
rect 1765 546 1799 580
rect 1765 470 1799 504
rect 1765 390 1799 424
rect 1855 546 1889 580
rect 1855 474 1889 508
rect 1945 546 1979 580
rect 1945 470 1979 504
rect 1945 390 1979 424
<< poly >>
rect 84 592 114 618
rect 174 592 204 618
rect 264 592 294 618
rect 354 592 384 618
rect 444 592 474 618
rect 534 592 564 618
rect 624 592 654 618
rect 714 592 744 618
rect 804 592 834 618
rect 894 592 924 618
rect 984 592 1014 618
rect 1074 592 1104 618
rect 1272 592 1302 618
rect 1362 592 1392 618
rect 1452 592 1482 618
rect 1542 592 1572 618
rect 1632 592 1662 618
rect 1722 592 1752 618
rect 1812 592 1842 618
rect 1902 592 1932 618
rect 84 353 114 368
rect 174 353 204 368
rect 264 353 294 368
rect 354 353 384 368
rect 444 353 474 368
rect 534 353 564 368
rect 624 353 654 368
rect 714 353 744 368
rect 804 353 834 368
rect 894 353 924 368
rect 984 353 1014 368
rect 1074 353 1104 368
rect 1272 353 1302 368
rect 1362 353 1392 368
rect 1452 353 1482 368
rect 1542 353 1572 368
rect 1632 353 1662 368
rect 1722 353 1752 368
rect 1812 353 1842 368
rect 1902 353 1932 368
rect 81 336 117 353
rect 171 336 207 353
rect 261 336 297 353
rect 351 336 387 353
rect 441 336 477 353
rect 531 336 567 353
rect 621 336 657 353
rect 49 320 387 336
rect 49 286 65 320
rect 99 286 133 320
rect 167 286 201 320
rect 235 286 269 320
rect 303 286 337 320
rect 371 286 387 320
rect 49 270 387 286
rect 430 320 657 336
rect 430 286 461 320
rect 495 286 529 320
rect 563 286 597 320
rect 631 294 657 320
rect 711 294 747 353
rect 801 326 837 353
rect 891 326 927 353
rect 981 326 1017 353
rect 1071 326 1107 353
rect 1269 336 1305 353
rect 1359 336 1395 353
rect 1449 336 1485 353
rect 1539 336 1575 353
rect 801 320 1107 326
rect 1258 320 1575 336
rect 801 310 1116 320
rect 801 296 831 310
rect 631 286 746 294
rect 84 222 114 270
rect 170 222 200 270
rect 258 222 288 270
rect 344 222 374 270
rect 430 264 746 286
rect 430 222 460 264
rect 516 222 546 264
rect 621 222 651 264
rect 716 222 746 264
rect 815 276 831 296
rect 865 276 899 310
rect 933 276 967 310
rect 1001 276 1035 310
rect 1069 290 1116 310
rect 1069 276 1202 290
rect 815 260 1202 276
rect 914 222 944 260
rect 1000 222 1030 260
rect 1086 222 1116 260
rect 1172 222 1202 260
rect 1258 286 1274 320
rect 1308 286 1342 320
rect 1376 286 1410 320
rect 1444 286 1478 320
rect 1512 286 1575 320
rect 1629 336 1665 353
rect 1719 336 1755 353
rect 1809 336 1845 353
rect 1899 336 1935 353
rect 1629 320 1968 336
rect 1629 306 1646 320
rect 1258 270 1575 286
rect 1630 286 1646 306
rect 1680 286 1714 320
rect 1748 286 1782 320
rect 1816 286 1850 320
rect 1884 286 1918 320
rect 1952 286 1968 320
rect 1630 270 1968 286
rect 1258 222 1288 270
rect 1358 222 1388 270
rect 1444 222 1474 270
rect 1544 222 1574 270
rect 1630 222 1660 270
rect 1716 222 1746 270
rect 1802 222 1832 270
rect 1902 222 1932 270
rect 84 48 114 74
rect 170 48 200 74
rect 258 48 288 74
rect 344 48 374 74
rect 430 48 460 74
rect 516 48 546 74
rect 621 48 651 74
rect 716 48 746 74
rect 914 48 944 74
rect 1000 48 1030 74
rect 1086 48 1116 74
rect 1172 48 1202 74
rect 1258 48 1288 74
rect 1358 48 1388 74
rect 1444 48 1474 74
rect 1544 48 1574 74
rect 1630 48 1660 74
rect 1716 48 1746 74
rect 1802 48 1832 74
rect 1902 48 1932 74
<< polycont >>
rect 65 286 99 320
rect 133 286 167 320
rect 201 286 235 320
rect 269 286 303 320
rect 337 286 371 320
rect 461 286 495 320
rect 529 286 563 320
rect 597 286 631 320
rect 831 276 865 310
rect 899 276 933 310
rect 967 276 1001 310
rect 1035 276 1069 310
rect 1274 286 1308 320
rect 1342 286 1376 320
rect 1410 286 1444 320
rect 1478 286 1512 320
rect 1646 286 1680 320
rect 1714 286 1748 320
rect 1782 286 1816 320
rect 1850 286 1884 320
rect 1918 286 1952 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 21 580 71 649
rect 21 546 37 580
rect 21 510 71 546
rect 21 476 37 510
rect 21 440 71 476
rect 21 406 37 440
rect 21 390 71 406
rect 111 580 177 596
rect 111 546 127 580
rect 161 546 177 580
rect 111 505 177 546
rect 111 471 127 505
rect 161 471 177 505
rect 111 424 177 471
rect 217 580 251 649
rect 217 508 251 546
rect 217 458 251 474
rect 291 580 357 596
rect 291 546 307 580
rect 341 546 357 580
rect 291 505 357 546
rect 291 471 307 505
rect 341 471 357 505
rect 291 424 357 471
rect 397 580 431 649
rect 397 508 431 546
rect 397 458 431 474
rect 471 580 537 596
rect 471 546 487 580
rect 521 546 537 580
rect 471 505 537 546
rect 471 471 487 505
rect 521 471 537 505
rect 471 424 537 471
rect 577 580 611 649
rect 577 508 611 546
rect 577 458 611 474
rect 651 580 717 596
rect 651 546 667 580
rect 701 546 717 580
rect 651 505 717 546
rect 651 471 667 505
rect 701 471 717 505
rect 651 424 717 471
rect 111 390 127 424
rect 161 390 307 424
rect 341 390 487 424
rect 521 390 667 424
rect 701 390 717 424
rect 25 320 387 356
rect 25 286 65 320
rect 99 286 133 320
rect 167 286 201 320
rect 235 286 269 320
rect 303 286 337 320
rect 371 286 387 320
rect 25 270 387 286
rect 445 320 647 356
rect 445 286 461 320
rect 495 286 529 320
rect 563 286 597 320
rect 631 286 647 320
rect 445 270 647 286
rect 683 326 717 390
rect 757 580 791 649
rect 757 497 791 546
rect 757 414 791 463
rect 757 364 791 380
rect 831 580 897 596
rect 831 546 847 580
rect 881 546 897 580
rect 831 497 897 546
rect 831 463 847 497
rect 881 463 897 497
rect 831 414 897 463
rect 937 580 971 649
rect 937 478 971 546
rect 937 428 971 444
rect 1011 580 1061 596
rect 1011 546 1027 580
rect 1011 497 1061 546
rect 1011 463 1027 497
rect 1101 580 1167 649
rect 1101 546 1117 580
rect 1151 546 1167 580
rect 1101 498 1167 546
rect 1101 464 1117 498
rect 1151 464 1167 498
rect 1209 581 1622 615
rect 1209 580 1262 581
rect 1209 546 1225 580
rect 1259 546 1262 580
rect 1402 580 1442 581
rect 1209 508 1262 546
rect 1209 474 1225 508
rect 1259 474 1262 508
rect 1011 430 1061 463
rect 1209 458 1262 474
rect 1299 537 1365 547
rect 1299 503 1315 537
rect 1349 503 1365 537
rect 831 380 847 414
rect 881 394 897 414
rect 1011 424 1127 430
rect 1299 428 1365 503
rect 1402 546 1405 580
rect 1439 546 1442 580
rect 1582 580 1622 581
rect 1402 508 1442 546
rect 1402 474 1405 508
rect 1439 474 1442 508
rect 1402 458 1442 474
rect 1479 537 1545 547
rect 1479 503 1495 537
rect 1529 503 1545 537
rect 1299 424 1315 428
rect 1011 414 1315 424
rect 1011 394 1027 414
rect 881 380 1027 394
rect 1061 394 1315 414
rect 1349 424 1365 428
rect 1479 428 1545 503
rect 1479 424 1495 428
rect 1349 394 1495 424
rect 1529 394 1545 428
rect 1061 390 1545 394
rect 1582 546 1585 580
rect 1619 546 1622 580
rect 1582 510 1622 546
rect 1582 476 1585 510
rect 1619 476 1622 510
rect 1582 440 1622 476
rect 1659 580 1712 649
rect 1659 546 1675 580
rect 1709 546 1712 580
rect 1659 508 1712 546
rect 1659 474 1675 508
rect 1709 474 1712 508
rect 1659 458 1712 474
rect 1749 580 1815 596
rect 1749 546 1765 580
rect 1799 546 1815 580
rect 1749 504 1815 546
rect 1749 470 1765 504
rect 1799 470 1815 504
rect 1582 406 1585 440
rect 1619 424 1622 440
rect 1749 424 1815 470
rect 1852 580 1893 649
rect 1852 546 1855 580
rect 1889 546 1893 580
rect 1852 508 1893 546
rect 1852 474 1855 508
rect 1889 474 1893 508
rect 1852 458 1893 474
rect 1929 580 1995 596
rect 1929 546 1945 580
rect 1979 546 1995 580
rect 1929 504 1995 546
rect 1929 470 1945 504
rect 1979 470 1995 504
rect 1929 424 1995 470
rect 1619 406 1765 424
rect 1582 390 1765 406
rect 1799 390 1945 424
rect 1979 390 1995 424
rect 1061 380 1143 390
rect 831 360 1143 380
rect 683 310 1075 326
rect 683 276 831 310
rect 865 276 899 310
rect 933 276 967 310
rect 1001 276 1035 310
rect 1069 276 1075 310
rect 683 260 1075 276
rect 683 236 721 260
rect 23 210 419 236
rect 23 176 39 210
rect 73 202 212 210
rect 23 120 73 176
rect 211 176 212 202
rect 246 202 385 210
rect 246 176 247 202
rect 23 86 39 120
rect 23 70 73 86
rect 109 136 175 168
rect 109 102 125 136
rect 159 102 175 136
rect 109 17 175 102
rect 211 120 247 176
rect 211 86 212 120
rect 246 86 247 120
rect 211 70 247 86
rect 283 136 349 168
rect 283 102 299 136
rect 333 102 349 136
rect 283 17 349 102
rect 385 120 419 176
rect 455 202 721 236
rect 1109 226 1143 360
rect 1177 320 1528 356
rect 1177 286 1274 320
rect 1308 286 1342 320
rect 1376 286 1410 320
rect 1444 286 1478 320
rect 1512 286 1528 320
rect 1177 270 1528 286
rect 1630 320 1991 356
rect 1630 286 1646 320
rect 1680 286 1714 320
rect 1748 286 1782 320
rect 1816 286 1850 320
rect 1884 286 1918 320
rect 1952 286 1991 320
rect 1630 270 1991 286
rect 455 181 521 202
rect 455 147 471 181
rect 505 147 521 181
rect 655 189 721 202
rect 455 119 521 147
rect 555 136 621 168
rect 385 85 419 86
rect 555 102 571 136
rect 605 102 621 136
rect 655 155 671 189
rect 705 155 721 189
rect 655 119 721 155
rect 757 210 807 226
rect 791 176 807 210
rect 757 120 807 176
rect 555 85 621 102
rect 791 86 807 120
rect 757 85 807 86
rect 385 51 807 85
rect 853 210 903 226
rect 853 176 869 210
rect 853 120 903 176
rect 853 86 869 120
rect 939 192 1177 226
rect 939 189 1005 192
rect 939 155 955 189
rect 989 155 1005 189
rect 1109 189 1177 192
rect 939 119 1005 155
rect 1041 131 1075 158
rect 853 85 903 86
rect 1109 155 1127 189
rect 1161 155 1177 189
rect 1109 119 1177 155
rect 1213 210 1993 236
rect 1247 202 1399 210
rect 1213 120 1247 176
rect 1383 176 1399 202
rect 1433 202 1585 210
rect 1041 85 1075 97
rect 1213 85 1247 86
rect 853 51 1247 85
rect 1283 147 1349 166
rect 1283 113 1299 147
rect 1333 113 1349 147
rect 1283 17 1349 113
rect 1383 120 1433 176
rect 1569 176 1585 202
rect 1619 202 1757 210
rect 1383 86 1399 120
rect 1383 70 1433 86
rect 1469 147 1535 166
rect 1469 113 1485 147
rect 1519 113 1535 147
rect 1469 17 1535 113
rect 1569 120 1619 176
rect 1791 202 1943 210
rect 1791 176 1807 202
rect 1569 86 1585 120
rect 1569 70 1619 86
rect 1655 147 1721 166
rect 1655 113 1671 147
rect 1705 113 1721 147
rect 1655 17 1721 113
rect 1757 120 1807 176
rect 1977 176 1993 210
rect 1791 86 1807 120
rect 1757 70 1807 86
rect 1841 147 1907 166
rect 1841 113 1857 147
rect 1891 113 1907 147
rect 1841 17 1907 113
rect 1943 120 1993 176
rect 1977 86 1993 120
rect 1943 70 1993 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o2bb2ai_4
flabel pwell s 0 0 2016 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 2016 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 2016 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 2016 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 1087 390 1121 424 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 A2_N
port 2 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 A2_N
port 2 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 A1_N
port 1 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 A1_N
port 1 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A1_N
port 1 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A1_N
port 1 nsew
flabel corelocali s 1663 316 1697 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 1759 316 1793 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 1855 316 1889 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 1951 316 1985 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 1183 316 1217 350 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 1279 316 1313 350 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 1375 316 1409 350 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 1471 316 1505 350 0 FreeSans 340 0 0 0 B2
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 2016 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1406338
string GDS_START 1389172
<< end >>
