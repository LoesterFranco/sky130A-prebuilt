magic
tech sky130A
magscale 1 2
timestamp 1599588238
<< locali >>
rect 25 260 91 356
rect 197 290 263 356
rect 1252 384 1327 578
rect 1283 225 1317 384
rect 1264 70 1317 225
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 53 424 119 596
rect 153 458 219 649
rect 253 522 331 596
rect 472 556 541 649
rect 575 581 838 615
rect 575 522 609 581
rect 253 488 609 522
rect 53 390 159 424
rect 253 420 331 488
rect 125 226 159 390
rect 297 354 331 420
rect 365 394 445 454
rect 666 428 770 547
rect 365 388 702 394
rect 411 360 702 388
rect 297 234 377 354
rect 23 150 159 226
rect 227 184 377 234
rect 297 152 377 184
rect 23 116 263 150
rect 411 119 461 360
rect 495 260 594 326
rect 636 294 702 360
rect 229 85 263 116
rect 495 85 529 260
rect 125 17 191 82
rect 229 51 529 85
rect 563 17 629 211
rect 663 117 697 294
rect 736 211 770 428
rect 804 363 838 581
rect 872 525 1016 649
rect 1050 471 1116 591
rect 872 405 1116 471
rect 1050 393 1116 405
rect 804 297 870 363
rect 1050 359 1135 393
rect 1169 364 1212 649
rect 1101 325 1135 359
rect 998 263 1067 325
rect 816 259 1067 263
rect 1101 259 1249 325
rect 816 229 1032 259
rect 816 211 850 229
rect 1101 225 1135 259
rect 1367 364 1417 649
rect 731 161 850 211
rect 663 51 875 117
rect 964 17 1030 195
rect 1066 191 1135 225
rect 1066 71 1116 191
rect 1169 17 1228 225
rect 1351 17 1417 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 683 1440 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 0 617 1440 649
rect 0 17 1440 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -49 1440 -17
<< labels >>
rlabel locali s 25 260 91 356 6 D
port 1 nsew signal input
rlabel locali s 1283 225 1317 384 6 Q
port 2 nsew signal output
rlabel locali s 1264 70 1317 225 6 Q
port 2 nsew signal output
rlabel locali s 1252 384 1327 578 6 Q
port 2 nsew signal output
rlabel locali s 197 290 263 356 6 GATE_N
port 3 nsew clock input
rlabel metal1 s 0 -49 1440 49 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1440 715 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1440 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2993948
string GDS_START 2982644
<< end >>
