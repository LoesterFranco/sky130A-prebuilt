magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 644 561
rect 17 425 69 527
rect 17 215 85 391
rect 201 426 324 527
rect 285 391 324 426
rect 358 425 453 493
rect 487 418 530 527
rect 285 353 351 391
rect 572 353 627 493
rect 17 17 69 181
rect 397 145 479 249
rect 593 147 627 353
rect 397 61 437 145
rect 475 17 541 109
rect 575 51 627 147
rect 0 -17 644 17
<< obsli1 >>
rect 119 249 153 493
rect 201 319 251 392
rect 395 319 538 378
rect 201 285 559 319
rect 119 199 278 249
rect 119 181 169 199
rect 103 97 169 181
rect 312 114 363 285
rect 205 61 363 114
rect 513 199 559 285
<< metal1 >>
rect 0 496 644 592
rect 0 -48 644 48
<< labels >>
rlabel locali s 17 215 85 391 6 A_N
port 1 nsew signal input
rlabel locali s 358 425 453 493 6 B
port 2 nsew signal input
rlabel locali s 397 145 479 249 6 C
port 3 nsew signal input
rlabel locali s 397 61 437 145 6 C
port 3 nsew signal input
rlabel locali s 593 147 627 353 6 X
port 4 nsew signal output
rlabel locali s 575 51 627 147 6 X
port 4 nsew signal output
rlabel locali s 572 353 627 493 6 X
port 4 nsew signal output
rlabel locali s 475 17 541 109 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 17 17 69 181 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 644 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 644 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 487 418 530 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 285 391 324 426 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 285 353 351 391 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 201 426 324 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 17 425 69 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 644 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 644 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3800670
string GDS_START 3794328
<< end >>
