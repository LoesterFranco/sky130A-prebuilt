magic
tech sky130A
magscale 1 2
timestamp 1604502711
<< locali >>
rect 17 459 85 493
rect 17 425 31 459
rect 65 425 85 459
rect 17 333 85 425
rect 17 75 65 265
rect 119 258 153 493
rect 187 459 259 493
rect 187 425 211 459
rect 245 425 259 459
rect 187 333 259 425
rect 119 189 259 258
rect 118 152 259 189
rect 118 51 168 152
<< viali >>
rect 31 425 65 459
rect 211 425 245 459
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 276 561
rect 202 17 259 118
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 276 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
<< metal1 >>
rect 0 561 276 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 276 561
rect 0 496 276 527
rect 14 459 262 468
rect 14 428 31 459
rect 19 425 31 428
rect 65 428 211 459
rect 65 425 77 428
rect 19 416 77 425
rect 199 425 211 428
rect 245 428 262 459
rect 245 425 257 428
rect 199 416 257 425
rect 0 17 276 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 276 17
rect 0 -48 276 -17
<< labels >>
rlabel locali s 17 75 65 265 6 A
port 1 nsew signal input
rlabel locali s 119 258 153 493 6 Y
port 2 nsew signal output
rlabel locali s 119 189 259 258 6 Y
port 2 nsew signal output
rlabel locali s 118 152 259 189 6 Y
port 2 nsew signal output
rlabel locali s 118 51 168 152 6 Y
port 2 nsew signal output
rlabel viali s 31 425 65 459 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 17 333 85 493 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel viali s 211 425 245 459 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 187 333 259 493 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 199 416 257 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 19 416 77 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 14 428 262 468 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 0 -48 276 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 276 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 276 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2174986
string GDS_START 2170860
<< end >>
