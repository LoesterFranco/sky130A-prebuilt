magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 1050 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 97 93 127 177
rect 186 93 216 177
rect 398 47 428 131
rect 495 47 525 131
rect 586 47 616 131
rect 683 47 713 131
rect 791 47 821 177
rect 885 47 915 177
<< pmoshvt >>
rect 81 410 117 494
rect 390 413 426 497
rect 188 297 224 381
rect 496 297 532 381
rect 578 297 614 381
rect 675 297 711 381
rect 783 297 819 497
rect 877 297 913 497
<< ndiff >>
rect 35 149 97 177
rect 35 115 43 149
rect 77 115 97 149
rect 35 93 97 115
rect 127 149 186 177
rect 127 115 142 149
rect 176 115 186 149
rect 127 93 186 115
rect 216 149 278 177
rect 216 115 236 149
rect 270 115 278 149
rect 728 131 791 177
rect 216 93 278 115
rect 332 97 398 131
rect 332 63 340 97
rect 374 63 398 97
rect 332 47 398 63
rect 428 111 495 131
rect 428 77 438 111
rect 472 77 495 111
rect 428 47 495 77
rect 525 97 586 131
rect 525 63 535 97
rect 569 63 586 97
rect 525 47 586 63
rect 616 111 683 131
rect 616 77 629 111
rect 663 77 683 111
rect 616 47 683 77
rect 713 97 791 131
rect 713 63 733 97
rect 767 63 791 97
rect 713 47 791 63
rect 821 135 885 177
rect 821 101 831 135
rect 865 101 885 135
rect 821 47 885 101
rect 915 163 972 177
rect 915 129 930 163
rect 964 129 972 163
rect 915 95 972 129
rect 915 61 930 95
rect 964 61 972 95
rect 915 47 972 61
<< pdiff >>
rect 27 475 81 494
rect 27 441 35 475
rect 69 441 81 475
rect 27 410 81 441
rect 117 475 171 494
rect 117 441 129 475
rect 163 441 171 475
rect 117 410 171 441
rect 336 475 390 497
rect 336 441 344 475
rect 378 441 390 475
rect 336 413 390 441
rect 426 413 479 497
rect 134 381 171 410
rect 134 297 188 381
rect 224 339 282 381
rect 224 305 236 339
rect 270 305 282 339
rect 224 297 282 305
rect 443 381 479 413
rect 728 485 783 497
rect 728 451 736 485
rect 770 451 783 485
rect 728 417 783 451
rect 728 383 736 417
rect 770 383 783 417
rect 728 381 783 383
rect 443 297 496 381
rect 532 297 578 381
rect 614 297 675 381
rect 711 297 783 381
rect 819 454 877 497
rect 819 420 831 454
rect 865 420 877 454
rect 819 386 877 420
rect 819 352 831 386
rect 865 352 877 386
rect 819 297 877 352
rect 913 485 972 497
rect 913 451 930 485
rect 964 451 972 485
rect 913 417 972 451
rect 913 383 930 417
rect 964 383 972 417
rect 913 349 972 383
rect 913 315 930 349
rect 964 315 972 349
rect 913 297 972 315
<< ndiffc >>
rect 43 115 77 149
rect 142 115 176 149
rect 236 115 270 149
rect 340 63 374 97
rect 438 77 472 111
rect 535 63 569 97
rect 629 77 663 111
rect 733 63 767 97
rect 831 101 865 135
rect 930 129 964 163
rect 930 61 964 95
<< pdiffc >>
rect 35 441 69 475
rect 129 441 163 475
rect 344 441 378 475
rect 236 305 270 339
rect 736 451 770 485
rect 736 383 770 417
rect 831 420 865 454
rect 831 352 865 386
rect 930 451 964 485
rect 930 383 964 417
rect 930 315 964 349
<< poly >>
rect 81 494 117 520
rect 390 497 426 523
rect 783 497 819 523
rect 877 497 913 523
rect 81 395 117 410
rect 79 265 119 395
rect 188 381 224 407
rect 390 398 426 413
rect 188 282 224 297
rect 186 265 226 282
rect 388 265 428 398
rect 576 484 646 494
rect 576 450 592 484
rect 626 450 646 484
rect 576 440 646 450
rect 576 407 616 440
rect 496 381 532 407
rect 578 381 614 407
rect 675 381 711 407
rect 496 282 532 297
rect 578 282 614 297
rect 675 282 711 297
rect 783 282 819 297
rect 877 282 913 297
rect 494 265 534 282
rect 79 249 140 265
rect 79 215 89 249
rect 123 215 140 249
rect 79 199 140 215
rect 186 249 260 265
rect 186 215 200 249
rect 234 215 260 249
rect 186 199 260 215
rect 327 249 428 265
rect 327 215 337 249
rect 371 215 428 249
rect 327 199 428 215
rect 470 249 534 265
rect 470 215 480 249
rect 514 215 534 249
rect 470 199 534 215
rect 97 177 127 199
rect 186 177 216 199
rect 398 131 428 199
rect 495 131 525 199
rect 576 152 616 282
rect 673 265 713 282
rect 781 265 821 282
rect 875 265 915 282
rect 658 249 722 265
rect 658 215 668 249
rect 702 215 722 249
rect 658 199 722 215
rect 764 249 915 265
rect 764 215 774 249
rect 808 215 915 249
rect 764 199 915 215
rect 586 131 616 152
rect 683 131 713 199
rect 791 177 821 199
rect 885 177 915 199
rect 97 67 127 93
rect 186 67 216 93
rect 398 21 428 47
rect 495 21 525 47
rect 586 21 616 47
rect 683 21 713 47
rect 791 21 821 47
rect 885 21 915 47
<< polycont >>
rect 592 450 626 484
rect 89 215 123 249
rect 200 215 234 249
rect 337 215 371 249
rect 480 215 514 249
rect 668 215 702 249
rect 774 215 808 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 17 475 69 491
rect 17 441 35 475
rect 103 475 179 527
rect 541 484 679 491
rect 103 441 129 475
rect 163 441 179 475
rect 327 441 344 475
rect 378 441 486 475
rect 17 407 69 441
rect 17 373 408 407
rect 17 165 52 373
rect 86 249 166 339
rect 209 305 236 339
rect 270 305 340 339
rect 86 215 89 249
rect 123 215 166 249
rect 86 199 166 215
rect 200 249 268 265
rect 234 215 268 249
rect 200 199 268 215
rect 302 249 340 305
rect 374 317 408 373
rect 452 391 486 441
rect 541 450 592 484
rect 626 450 679 484
rect 541 425 679 450
rect 723 485 779 527
rect 723 451 736 485
rect 770 451 779 485
rect 723 417 779 451
rect 452 357 679 391
rect 723 383 736 417
rect 770 383 779 417
rect 723 367 779 383
rect 831 454 891 493
rect 865 420 891 454
rect 831 386 891 420
rect 645 333 679 357
rect 865 352 891 386
rect 374 283 514 317
rect 645 299 787 333
rect 831 299 891 352
rect 480 249 514 283
rect 753 265 787 299
rect 302 215 337 249
rect 371 215 391 249
rect 302 165 340 215
rect 480 199 514 215
rect 568 249 719 265
rect 568 215 668 249
rect 702 215 719 249
rect 568 199 719 215
rect 753 249 808 265
rect 753 215 774 249
rect 753 199 808 215
rect 753 165 787 199
rect 17 149 81 165
rect 17 115 43 149
rect 77 115 81 149
rect 17 90 81 115
rect 142 149 176 165
rect 142 17 176 115
rect 236 149 340 165
rect 270 131 340 149
rect 438 131 787 165
rect 852 152 891 299
rect 930 485 964 527
rect 930 417 964 451
rect 930 349 964 383
rect 930 288 964 315
rect 831 135 891 152
rect 236 90 270 115
rect 438 111 472 131
rect 319 63 340 97
rect 374 63 394 97
rect 319 17 394 63
rect 629 111 663 131
rect 438 61 472 77
rect 509 63 535 97
rect 569 63 585 97
rect 509 17 585 63
rect 865 101 891 135
rect 629 61 663 77
rect 697 63 733 97
rect 767 63 783 97
rect 831 83 891 101
rect 930 163 964 183
rect 930 95 964 129
rect 697 17 783 63
rect 930 17 964 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
flabel corelocali s 603 238 603 238 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 840 357 874 391 0 FreeSans 400 0 0 0 X
port 9 nsew
flabel corelocali s 603 442 603 442 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel corelocali s 231 238 231 238 0 FreeSans 400 0 0 0 D_N
port 4 nsew
flabel corelocali s 132 221 166 255 0 FreeSans 400 0 0 0 C_N
port 3 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
rlabel comment s 0 0 0 0 4 or4bb_2
<< properties >>
string FIXED_BBOX 0 0 1012 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 8094
string GDS_START 134
<< end >>
