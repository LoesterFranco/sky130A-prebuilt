magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 2852 561
rect 103 455 169 527
rect 541 428 620 527
rect 17 153 68 335
rect 108 153 164 335
rect 210 153 267 335
rect 729 455 795 527
rect 581 323 620 394
rect 481 215 547 318
rect 581 211 713 323
rect 581 145 620 211
rect 17 17 140 119
rect 368 17 418 109
rect 1200 455 1266 527
rect 540 17 620 111
rect 1412 425 1603 527
rect 1832 447 1898 527
rect 2020 447 2086 527
rect 1328 289 1413 353
rect 728 17 788 109
rect 1776 305 1987 345
rect 1776 287 1823 305
rect 2216 297 2258 527
rect 1133 17 1233 93
rect 1344 17 1541 161
rect 2007 17 2057 109
rect 2224 17 2258 177
rect 2292 51 2371 493
rect 2405 297 2463 527
rect 2577 327 2648 527
rect 2682 299 2748 490
rect 2405 17 2463 177
rect 2703 165 2748 299
rect 2782 297 2835 527
rect 2577 17 2648 165
rect 2682 55 2748 165
rect 2782 17 2835 177
rect 0 -17 2852 17
<< obsli1 >>
rect 17 415 69 493
rect 203 451 421 493
rect 203 415 237 451
rect 455 417 507 493
rect 17 369 237 415
rect 271 369 339 417
rect 301 323 339 369
rect 301 289 305 323
rect 301 144 339 289
rect 300 141 339 144
rect 396 352 507 417
rect 654 400 695 465
rect 829 427 888 493
rect 396 181 447 352
rect 654 391 799 400
rect 654 366 765 391
rect 747 357 765 366
rect 396 143 506 181
rect 747 177 799 357
rect 299 129 339 141
rect 299 119 334 129
rect 174 51 334 119
rect 452 51 506 143
rect 654 143 799 177
rect 833 284 888 427
rect 933 323 978 493
rect 1012 427 1161 493
rect 1041 357 1052 391
rect 1086 357 1093 391
rect 933 318 960 323
rect 943 289 960 318
rect 1041 315 1093 357
rect 833 255 898 284
rect 833 221 857 255
rect 891 221 898 255
rect 833 218 898 221
rect 654 51 694 143
rect 833 117 867 218
rect 943 184 977 289
rect 1127 279 1161 427
rect 1321 421 1364 490
rect 1637 425 1798 492
rect 1195 387 1364 421
rect 1764 413 1798 425
rect 1932 413 1986 490
rect 1195 315 1229 387
rect 1477 357 1512 391
rect 1546 357 1611 391
rect 1477 341 1611 357
rect 1028 255 1295 279
rect 1471 255 1541 265
rect 822 51 867 117
rect 901 51 977 184
rect 1011 245 1541 255
rect 1011 51 1090 245
rect 1124 161 1203 203
rect 1261 195 1541 245
rect 1577 179 1611 341
rect 1684 255 1730 381
rect 1764 379 2086 413
rect 2021 305 2086 379
rect 2120 271 2169 493
rect 1684 221 1696 255
rect 1684 215 1730 221
rect 1766 179 1817 253
rect 1124 127 1310 161
rect 1267 51 1310 127
rect 1577 139 1817 179
rect 1857 237 2182 271
rect 1857 171 1903 237
rect 1937 169 2112 203
rect 1937 103 1971 169
rect 2146 117 2182 237
rect 1693 55 1971 103
rect 2093 51 2182 117
rect 2506 265 2543 493
rect 2506 199 2669 265
rect 2506 51 2543 199
<< obsli1c >>
rect 305 289 339 323
rect 765 357 799 391
rect 1052 357 1086 391
rect 960 289 994 323
rect 857 221 891 255
rect 1512 357 1546 391
rect 1696 221 1730 255
<< metal1 >>
rect 0 496 2852 592
rect 1316 320 1374 329
rect 1776 320 1834 329
rect 1316 292 1834 320
rect 1316 283 1374 292
rect 1776 283 1834 292
rect 109 252 167 261
rect 477 252 535 261
rect 109 224 535 252
rect 109 215 167 224
rect 477 215 535 224
rect 0 -48 2852 48
<< obsm1 >>
rect 753 391 811 397
rect 753 357 765 391
rect 799 388 811 391
rect 1040 391 1098 397
rect 1040 388 1052 391
rect 799 360 1052 388
rect 799 357 811 360
rect 753 351 811 357
rect 1040 357 1052 360
rect 1086 388 1098 391
rect 1500 391 1558 397
rect 1500 388 1512 391
rect 1086 360 1512 388
rect 1086 357 1098 360
rect 1040 351 1098 357
rect 1500 357 1512 360
rect 1546 357 1558 391
rect 1500 351 1558 357
rect 293 323 351 329
rect 293 289 305 323
rect 339 320 351 323
rect 948 323 1006 329
rect 948 320 960 323
rect 339 292 960 320
rect 339 289 351 292
rect 293 283 351 289
rect 948 289 960 292
rect 994 289 1006 323
rect 948 283 1006 289
rect 845 255 903 261
rect 845 221 857 255
rect 891 252 903 255
rect 1684 255 1742 261
rect 1684 252 1696 255
rect 891 224 1696 252
rect 891 221 903 224
rect 845 215 903 221
rect 1684 221 1696 224
rect 1730 221 1742 255
rect 1684 215 1742 221
<< labels >>
rlabel locali s 210 153 267 335 6 D
port 1 nsew signal input
rlabel locali s 2703 165 2748 299 6 Q
port 2 nsew signal output
rlabel locali s 2682 299 2748 490 6 Q
port 2 nsew signal output
rlabel locali s 2682 55 2748 165 6 Q
port 2 nsew signal output
rlabel locali s 2292 51 2371 493 6 Q_N
port 3 nsew signal output
rlabel locali s 17 153 68 335 6 SCD
port 4 nsew signal input
rlabel locali s 108 153 164 335 6 SCE
port 5 nsew signal input
rlabel locali s 481 215 547 318 6 SCE
port 5 nsew signal input
rlabel metal1 s 477 252 535 261 6 SCE
port 5 nsew signal input
rlabel metal1 s 477 215 535 224 6 SCE
port 5 nsew signal input
rlabel metal1 s 109 252 167 261 6 SCE
port 5 nsew signal input
rlabel metal1 s 109 224 535 252 6 SCE
port 5 nsew signal input
rlabel metal1 s 109 215 167 224 6 SCE
port 5 nsew signal input
rlabel locali s 1328 289 1413 353 6 SET_B
port 6 nsew signal input
rlabel locali s 1776 305 1987 345 6 SET_B
port 6 nsew signal input
rlabel locali s 1776 287 1823 305 6 SET_B
port 6 nsew signal input
rlabel metal1 s 1776 320 1834 329 6 SET_B
port 6 nsew signal input
rlabel metal1 s 1776 283 1834 292 6 SET_B
port 6 nsew signal input
rlabel metal1 s 1316 320 1374 329 6 SET_B
port 6 nsew signal input
rlabel metal1 s 1316 292 1834 320 6 SET_B
port 6 nsew signal input
rlabel metal1 s 1316 283 1374 292 6 SET_B
port 6 nsew signal input
rlabel locali s 581 323 620 394 6 CLK
port 7 nsew clock input
rlabel locali s 581 211 713 323 6 CLK
port 7 nsew clock input
rlabel locali s 581 145 620 211 6 CLK
port 7 nsew clock input
rlabel locali s 2782 17 2835 177 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 2577 17 2648 165 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 2405 17 2463 177 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 2224 17 2258 177 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 2007 17 2057 109 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 1344 17 1541 161 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 1133 17 1233 93 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 728 17 788 109 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 540 17 620 111 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 368 17 418 109 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 17 17 140 119 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 0 -17 2852 17 8 VGND
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 2852 48 8 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 2782 297 2835 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 2577 327 2648 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 2405 297 2463 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 2216 297 2258 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 2020 447 2086 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 1832 447 1898 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 1412 425 1603 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 1200 455 1266 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 729 455 795 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 541 428 620 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 103 455 169 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 0 527 2852 561 6 VPWR
port 9 nsew power bidirectional abutment
rlabel metal1 s 0 496 2852 592 6 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2852 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 77464
string GDS_START 54832
<< end >>
