magic
tech sky130A
magscale 1 2
timestamp 1604502711
<< locali >>
rect 105 459 171 493
rect 105 425 122 459
rect 156 425 171 459
rect 105 367 171 425
rect 205 401 253 493
rect 287 462 353 493
rect 287 428 299 462
rect 333 428 353 462
rect 205 400 265 401
rect 205 396 266 400
rect 205 395 274 396
rect 205 394 277 395
rect 205 393 278 394
rect 387 393 433 493
rect 205 367 433 393
rect 237 365 433 367
rect 239 364 433 365
rect 241 363 433 364
rect 243 361 433 363
rect 249 357 433 361
rect 254 350 433 357
rect 467 459 524 493
rect 467 425 475 459
rect 509 425 524 459
rect 467 353 524 425
rect 85 151 155 265
rect 381 317 433 350
rect 381 283 532 317
rect 451 181 532 283
rect 202 147 532 181
rect 202 69 261 147
rect 381 69 433 147
<< viali >>
rect 122 425 156 459
rect 299 428 333 462
rect 475 425 509 459
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 17 333 71 493
rect 17 299 223 333
rect 17 117 51 299
rect 189 249 223 299
rect 189 215 417 249
rect 17 51 77 117
rect 111 17 166 113
rect 295 17 346 113
rect 467 17 523 113
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 14 462 538 468
rect 14 459 299 462
rect 14 428 122 459
rect 110 425 122 428
rect 156 428 299 459
rect 333 459 538 462
rect 333 428 475 459
rect 156 425 168 428
rect 110 416 168 425
rect 287 416 345 428
rect 463 425 475 428
rect 509 428 538 459
rect 509 425 521 428
rect 463 416 521 425
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
rlabel locali s 85 151 155 265 6 A
port 1 nsew signal input
rlabel locali s 451 181 532 283 6 X
port 2 nsew signal output
rlabel locali s 387 393 433 493 6 X
port 2 nsew signal output
rlabel locali s 381 317 433 350 6 X
port 2 nsew signal output
rlabel locali s 381 283 532 317 6 X
port 2 nsew signal output
rlabel locali s 381 69 433 147 6 X
port 2 nsew signal output
rlabel locali s 254 350 433 357 6 X
port 2 nsew signal output
rlabel locali s 249 357 433 361 6 X
port 2 nsew signal output
rlabel locali s 243 361 433 363 6 X
port 2 nsew signal output
rlabel locali s 241 363 433 364 6 X
port 2 nsew signal output
rlabel locali s 239 364 433 365 6 X
port 2 nsew signal output
rlabel locali s 237 365 433 367 6 X
port 2 nsew signal output
rlabel locali s 205 401 253 493 6 X
port 2 nsew signal output
rlabel locali s 205 400 265 401 6 X
port 2 nsew signal output
rlabel locali s 205 396 266 400 6 X
port 2 nsew signal output
rlabel locali s 205 395 274 396 6 X
port 2 nsew signal output
rlabel locali s 205 394 277 395 6 X
port 2 nsew signal output
rlabel locali s 205 393 278 394 6 X
port 2 nsew signal output
rlabel locali s 205 367 433 393 6 X
port 2 nsew signal output
rlabel locali s 202 147 532 181 6 X
port 2 nsew signal output
rlabel locali s 202 69 261 147 6 X
port 2 nsew signal output
rlabel viali s 122 425 156 459 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 105 367 171 493 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel viali s 475 425 509 459 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel viali s 299 428 333 462 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 467 353 524 493 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 287 428 353 493 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 463 416 521 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 287 416 345 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 110 416 168 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 14 428 538 468 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 0 -48 552 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 552 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 552 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2189892
string GDS_START 2183970
<< end >>
