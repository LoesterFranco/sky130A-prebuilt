magic
tech sky130A
magscale 1 2
timestamp 1601050056
<< nwell >>
rect -38 332 902 704
<< pwell >>
rect 0 0 864 49
<< scpmos >>
rect 83 368 119 592
rect 173 368 209 592
rect 263 368 299 592
rect 353 368 389 592
rect 460 388 496 588
rect 550 388 586 588
rect 640 388 676 588
rect 740 388 776 588
<< nmoslvt >>
rect 84 74 114 222
rect 170 74 200 222
rect 256 74 286 222
rect 359 74 389 222
rect 459 74 489 222
rect 556 74 586 222
<< ndiff >>
rect 27 131 84 222
rect 27 97 39 131
rect 73 97 84 131
rect 27 74 84 97
rect 114 210 170 222
rect 114 176 125 210
rect 159 176 170 210
rect 114 120 170 176
rect 114 86 125 120
rect 159 86 170 120
rect 114 74 170 86
rect 200 131 256 222
rect 200 97 211 131
rect 245 97 256 131
rect 200 74 256 97
rect 286 210 359 222
rect 286 176 301 210
rect 335 176 359 210
rect 286 120 359 176
rect 286 86 301 120
rect 335 86 359 120
rect 286 74 359 86
rect 389 152 459 222
rect 389 118 400 152
rect 434 118 459 152
rect 389 74 459 118
rect 489 210 556 222
rect 489 176 500 210
rect 534 176 556 210
rect 489 120 556 176
rect 489 86 500 120
rect 534 86 556 120
rect 489 74 556 86
rect 586 152 837 222
rect 586 118 597 152
rect 631 118 692 152
rect 726 118 788 152
rect 822 118 837 152
rect 586 74 837 118
<< pdiff >>
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 478 83 546
rect 27 444 39 478
rect 73 444 83 478
rect 27 368 83 444
rect 119 580 173 592
rect 119 546 129 580
rect 163 546 173 580
rect 119 497 173 546
rect 119 463 129 497
rect 163 463 173 497
rect 119 414 173 463
rect 119 380 129 414
rect 163 380 173 414
rect 119 368 173 380
rect 209 580 263 592
rect 209 546 219 580
rect 253 546 263 580
rect 209 478 263 546
rect 209 444 219 478
rect 253 444 263 478
rect 209 368 263 444
rect 299 580 353 592
rect 299 546 309 580
rect 343 546 353 580
rect 299 497 353 546
rect 299 463 309 497
rect 343 463 353 497
rect 299 414 353 463
rect 299 380 309 414
rect 343 380 353 414
rect 299 368 353 380
rect 389 588 445 592
rect 389 580 460 588
rect 389 546 399 580
rect 433 546 460 580
rect 389 474 460 546
rect 389 440 399 474
rect 433 440 460 474
rect 389 388 460 440
rect 496 576 550 588
rect 496 542 506 576
rect 540 542 550 576
rect 496 508 550 542
rect 496 474 506 508
rect 540 474 550 508
rect 496 388 550 474
rect 586 519 640 588
rect 586 485 596 519
rect 630 485 640 519
rect 586 388 640 485
rect 676 576 740 588
rect 676 542 696 576
rect 730 542 740 576
rect 676 388 740 542
rect 776 576 837 588
rect 776 542 788 576
rect 822 542 837 576
rect 776 388 837 542
rect 389 368 445 388
<< ndiffc >>
rect 39 97 73 131
rect 125 176 159 210
rect 125 86 159 120
rect 211 97 245 131
rect 301 176 335 210
rect 301 86 335 120
rect 400 118 434 152
rect 500 176 534 210
rect 500 86 534 120
rect 597 118 631 152
rect 692 118 726 152
rect 788 118 822 152
<< pdiffc >>
rect 39 546 73 580
rect 39 444 73 478
rect 129 546 163 580
rect 129 463 163 497
rect 129 380 163 414
rect 219 546 253 580
rect 219 444 253 478
rect 309 546 343 580
rect 309 463 343 497
rect 309 380 343 414
rect 399 546 433 580
rect 399 440 433 474
rect 506 542 540 576
rect 506 474 540 508
rect 596 485 630 519
rect 696 542 730 576
rect 788 542 822 576
<< poly >>
rect 83 592 119 618
rect 173 592 209 618
rect 263 592 299 618
rect 353 592 389 618
rect 460 588 496 614
rect 550 588 586 614
rect 640 588 676 614
rect 740 588 776 614
rect 83 326 119 368
rect 173 326 209 368
rect 263 326 299 368
rect 353 326 389 368
rect 460 336 496 388
rect 550 356 586 388
rect 640 356 676 388
rect 740 356 776 388
rect 550 340 676 356
rect 83 310 389 326
rect 83 276 135 310
rect 169 276 203 310
rect 237 276 271 310
rect 305 276 339 310
rect 373 276 389 310
rect 83 260 389 276
rect 442 320 508 336
rect 550 326 601 340
rect 442 286 458 320
rect 492 286 508 320
rect 442 270 508 286
rect 556 306 601 326
rect 635 326 676 340
rect 718 340 784 356
rect 635 306 651 326
rect 556 290 651 306
rect 718 306 734 340
rect 768 306 784 340
rect 718 290 784 306
rect 84 222 114 260
rect 170 222 200 260
rect 256 222 286 260
rect 359 222 389 260
rect 459 222 489 270
rect 556 222 586 290
rect 84 48 114 74
rect 170 48 200 74
rect 256 48 286 74
rect 359 48 389 74
rect 459 48 489 74
rect 556 48 586 74
<< polycont >>
rect 135 276 169 310
rect 203 276 237 310
rect 271 276 305 310
rect 339 276 373 310
rect 458 286 492 320
rect 601 306 635 340
rect 734 306 768 340
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 23 580 73 649
rect 23 546 39 580
rect 23 478 73 546
rect 23 444 39 478
rect 23 428 73 444
rect 113 580 179 596
rect 113 546 129 580
rect 163 546 179 580
rect 113 497 179 546
rect 113 463 129 497
rect 163 463 179 497
rect 113 414 179 463
rect 219 580 253 649
rect 219 478 253 546
rect 219 428 253 444
rect 293 580 359 596
rect 293 546 309 580
rect 343 546 359 580
rect 293 497 359 546
rect 293 463 309 497
rect 343 463 359 497
rect 113 394 129 414
rect 25 380 129 394
rect 163 394 179 414
rect 293 414 359 463
rect 399 580 449 649
rect 433 546 449 580
rect 399 474 449 546
rect 433 440 449 474
rect 490 581 746 615
rect 490 576 556 581
rect 490 542 506 576
rect 540 542 556 576
rect 680 576 746 581
rect 490 508 556 542
rect 490 474 506 508
rect 540 474 556 508
rect 490 458 556 474
rect 596 519 646 547
rect 680 542 696 576
rect 730 542 746 576
rect 680 526 746 542
rect 786 576 841 649
rect 786 542 788 576
rect 822 542 841 576
rect 786 526 841 542
rect 630 492 646 519
rect 630 485 847 492
rect 596 458 847 485
rect 399 424 449 440
rect 293 394 309 414
rect 163 380 309 394
rect 343 380 359 414
rect 504 390 779 424
rect 25 360 359 380
rect 25 226 71 360
rect 119 310 408 326
rect 119 276 135 310
rect 169 276 203 310
rect 237 276 271 310
rect 305 276 339 310
rect 373 276 408 310
rect 119 260 408 276
rect 442 320 551 390
rect 442 286 458 320
rect 492 286 551 320
rect 585 340 651 356
rect 585 306 601 340
rect 635 306 651 340
rect 585 290 651 306
rect 718 340 779 390
rect 718 306 734 340
rect 768 306 779 340
rect 718 290 779 306
rect 442 270 551 286
rect 374 236 408 260
rect 813 236 847 458
rect 25 210 340 226
rect 25 192 125 210
rect 109 176 125 192
rect 159 192 301 210
rect 23 131 73 158
rect 23 97 39 131
rect 23 17 73 97
rect 109 120 159 176
rect 281 176 301 192
rect 335 176 340 210
rect 374 210 847 236
rect 374 202 500 210
rect 109 86 125 120
rect 109 70 159 86
rect 195 131 245 158
rect 195 97 211 131
rect 195 17 245 97
rect 281 120 340 176
rect 484 176 500 202
rect 534 202 847 210
rect 534 176 550 202
rect 281 86 301 120
rect 335 86 340 120
rect 281 70 340 86
rect 384 152 450 168
rect 384 118 400 152
rect 434 118 450 152
rect 384 17 450 118
rect 484 120 550 176
rect 484 86 500 120
rect 534 86 550 120
rect 484 70 550 86
rect 584 152 841 168
rect 584 118 597 152
rect 631 118 692 152
rect 726 118 788 152
rect 822 118 841 152
rect 584 17 841 118
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
rlabel comment s 0 0 0 0 4 or2_4
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 7 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 7 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 A
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 864 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 756024
string GDS_START 748964
<< end >>
