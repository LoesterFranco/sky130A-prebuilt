magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 871 424 937 547
rect 1051 424 1117 547
rect 505 390 1117 424
rect 157 270 455 356
rect 505 236 551 390
rect 585 270 787 356
rect 847 270 1049 356
rect 505 202 1118 236
rect 505 176 930 202
rect 505 119 556 176
rect 880 70 930 176
rect 1068 70 1118 202
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 61 424 111 596
rect 151 458 201 649
rect 241 424 307 596
rect 347 458 381 649
rect 421 492 471 596
rect 511 526 561 649
rect 601 492 667 596
rect 707 526 741 649
rect 781 581 1207 615
rect 781 492 831 581
rect 421 458 831 492
rect 421 424 471 458
rect 977 458 1011 581
rect 61 390 471 424
rect 61 364 111 390
rect 1157 364 1207 581
rect 76 202 470 236
rect 76 70 126 202
rect 162 17 228 168
rect 264 70 298 202
rect 334 17 400 168
rect 436 85 470 202
rect 592 85 658 142
rect 764 85 830 142
rect 436 51 830 85
rect 966 17 1032 168
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
<< metal1 >>
rect 0 683 1248 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 0 617 1248 649
rect 0 17 1248 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
rect 0 -49 1248 -17
<< labels >>
rlabel locali s 585 270 787 356 6 A1
port 1 nsew signal input
rlabel locali s 157 270 455 356 6 A2
port 2 nsew signal input
rlabel locali s 847 270 1049 356 6 B1
port 3 nsew signal input
rlabel locali s 1068 70 1118 202 6 Y
port 4 nsew signal output
rlabel locali s 1051 424 1117 547 6 Y
port 4 nsew signal output
rlabel locali s 880 70 930 176 6 Y
port 4 nsew signal output
rlabel locali s 871 424 937 547 6 Y
port 4 nsew signal output
rlabel locali s 505 390 1117 424 6 Y
port 4 nsew signal output
rlabel locali s 505 236 551 390 6 Y
port 4 nsew signal output
rlabel locali s 505 202 1118 236 6 Y
port 4 nsew signal output
rlabel locali s 505 176 930 202 6 Y
port 4 nsew signal output
rlabel locali s 505 119 556 176 6 Y
port 4 nsew signal output
rlabel metal1 s 0 -49 1248 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 617 1248 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1248 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 4128258
string GDS_START 4117992
<< end >>
