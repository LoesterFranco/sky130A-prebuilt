magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 828 561
rect 110 442 182 527
rect 284 442 350 527
rect 451 442 519 527
rect 17 215 85 328
rect 187 283 444 340
rect 480 283 544 340
rect 187 181 221 283
rect 187 147 405 181
rect 124 17 158 113
rect 200 57 266 147
rect 371 117 405 147
rect 507 199 544 283
rect 578 199 640 340
rect 300 17 334 113
rect 371 51 418 117
rect 452 17 518 97
rect 620 17 698 97
rect 0 -17 828 17
<< obsli1 >>
rect 17 408 69 444
rect 704 442 811 485
rect 17 374 724 408
rect 17 362 153 374
rect 119 181 153 362
rect 17 147 153 181
rect 255 215 473 249
rect 17 58 69 147
rect 439 178 473 215
rect 678 265 724 374
rect 678 199 736 265
rect 439 165 480 178
rect 770 165 811 442
rect 439 144 811 165
rect 450 131 811 144
rect 552 61 586 131
rect 732 121 811 131
rect 732 61 783 121
<< metal1 >>
rect 0 496 828 592
rect 0 -48 828 48
<< labels >>
rlabel locali s 507 199 544 283 6 A
port 1 nsew signal input
rlabel locali s 480 283 544 340 6 A
port 1 nsew signal input
rlabel locali s 578 199 640 340 6 B
port 2 nsew signal input
rlabel locali s 17 215 85 328 6 C_N
port 3 nsew signal input
rlabel locali s 371 117 405 147 6 X
port 4 nsew signal output
rlabel locali s 371 51 418 117 6 X
port 4 nsew signal output
rlabel locali s 200 57 266 147 6 X
port 4 nsew signal output
rlabel locali s 187 283 444 340 6 X
port 4 nsew signal output
rlabel locali s 187 181 221 283 6 X
port 4 nsew signal output
rlabel locali s 187 147 405 181 6 X
port 4 nsew signal output
rlabel locali s 620 17 698 97 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 452 17 518 97 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 300 17 334 113 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 124 17 158 113 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 828 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 828 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 451 442 519 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 284 442 350 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 110 442 182 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 828 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 828 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1062984
string GDS_START 1056550
<< end >>
