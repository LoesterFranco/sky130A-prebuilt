magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 356 998 704
rect -38 332 349 356
rect 622 332 998 356
<< pwell >>
rect 0 0 960 49
<< scnmos >>
rect 84 74 114 222
rect 275 130 305 258
rect 361 130 391 258
rect 467 139 497 267
rect 665 119 695 247
rect 737 119 767 247
rect 837 99 867 247
<< pmoshvt >>
rect 86 368 116 592
rect 255 392 285 560
rect 356 392 386 592
rect 470 392 500 592
rect 635 424 665 592
rect 725 424 755 592
rect 835 368 865 592
<< ndiff >>
rect 417 258 467 267
rect 218 238 275 258
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 132 164 222
rect 218 204 230 238
rect 264 204 275 238
rect 218 186 275 204
rect 114 120 171 132
rect 225 130 275 186
rect 305 244 361 258
rect 305 210 316 244
rect 350 210 361 244
rect 305 176 361 210
rect 305 142 316 176
rect 350 142 361 176
rect 305 130 361 142
rect 391 176 467 258
rect 391 142 404 176
rect 438 142 467 176
rect 391 139 467 142
rect 497 236 554 267
rect 497 202 508 236
rect 542 202 554 236
rect 497 139 554 202
rect 608 235 665 247
rect 608 201 620 235
rect 654 201 665 235
rect 608 165 665 201
rect 391 130 452 139
rect 114 86 125 120
rect 159 86 171 120
rect 608 131 620 165
rect 654 131 665 165
rect 608 119 665 131
rect 695 119 737 247
rect 767 229 837 247
rect 767 195 778 229
rect 812 195 837 229
rect 767 161 837 195
rect 767 127 778 161
rect 812 127 837 161
rect 767 119 837 127
rect 114 74 171 86
rect 787 99 837 119
rect 867 220 924 247
rect 867 186 878 220
rect 912 186 924 220
rect 867 145 924 186
rect 867 111 878 145
rect 912 111 924 145
rect 867 99 924 111
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 497 86 546
rect 27 463 39 497
rect 73 463 86 497
rect 27 414 86 463
rect 27 380 39 414
rect 73 380 86 414
rect 27 368 86 380
rect 116 572 237 592
rect 116 538 167 572
rect 201 560 237 572
rect 303 560 356 592
rect 201 538 255 560
rect 116 392 255 538
rect 285 528 356 560
rect 285 494 298 528
rect 332 494 356 528
rect 285 392 356 494
rect 386 392 470 592
rect 500 580 635 592
rect 500 546 513 580
rect 547 546 588 580
rect 622 546 635 580
rect 500 496 635 546
rect 500 462 513 496
rect 547 462 588 496
rect 622 462 635 496
rect 500 424 635 462
rect 665 580 725 592
rect 665 546 678 580
rect 712 546 725 580
rect 665 470 725 546
rect 665 436 678 470
rect 712 436 725 470
rect 665 424 725 436
rect 755 580 835 592
rect 755 546 778 580
rect 812 546 835 580
rect 755 470 835 546
rect 755 436 778 470
rect 812 436 835 470
rect 755 424 835 436
rect 500 392 553 424
rect 116 368 169 392
rect 782 368 835 424
rect 865 580 924 592
rect 865 546 878 580
rect 912 546 924 580
rect 865 500 924 546
rect 865 466 878 500
rect 912 466 924 500
rect 865 420 924 466
rect 865 386 878 420
rect 912 386 924 420
rect 865 368 924 386
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 230 204 264 238
rect 316 210 350 244
rect 316 142 350 176
rect 404 142 438 176
rect 508 202 542 236
rect 620 201 654 235
rect 125 86 159 120
rect 620 131 654 165
rect 778 195 812 229
rect 778 127 812 161
rect 878 186 912 220
rect 878 111 912 145
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 167 538 201 572
rect 298 494 332 528
rect 513 546 547 580
rect 588 546 622 580
rect 513 462 547 496
rect 588 462 622 496
rect 678 546 712 580
rect 678 436 712 470
rect 778 546 812 580
rect 778 436 812 470
rect 878 546 912 580
rect 878 466 912 500
rect 878 386 912 420
<< poly >>
rect 86 592 116 618
rect 356 592 386 618
rect 470 592 500 618
rect 635 592 665 618
rect 725 592 755 618
rect 835 592 865 618
rect 255 560 285 586
rect 635 409 665 424
rect 725 409 755 424
rect 255 377 285 392
rect 356 377 386 392
rect 470 377 500 392
rect 86 353 116 368
rect 252 360 288 377
rect 353 360 389 377
rect 83 326 119 353
rect 239 344 305 360
rect 83 310 171 326
rect 83 276 121 310
rect 155 276 171 310
rect 239 310 255 344
rect 289 310 305 344
rect 239 294 305 310
rect 353 344 419 360
rect 353 310 369 344
rect 403 310 419 344
rect 353 294 419 310
rect 83 260 171 276
rect 84 222 114 260
rect 275 258 305 294
rect 361 258 391 294
rect 467 282 503 377
rect 632 360 668 409
rect 722 402 758 409
rect 722 372 767 402
rect 594 344 668 360
rect 594 310 610 344
rect 644 324 668 344
rect 644 310 695 324
rect 594 294 695 310
rect 467 267 497 282
rect 665 247 695 294
rect 737 247 767 372
rect 835 353 865 368
rect 832 336 868 353
rect 809 320 875 336
rect 809 286 825 320
rect 859 286 875 320
rect 809 270 875 286
rect 837 247 867 270
rect 275 104 305 130
rect 361 104 391 130
rect 467 117 497 139
rect 467 101 556 117
rect 84 48 114 74
rect 467 67 506 101
rect 540 67 556 101
rect 665 93 695 119
rect 467 51 556 67
rect 737 51 767 119
rect 837 73 867 99
rect 467 21 767 51
<< polycont >>
rect 121 276 155 310
rect 255 310 289 344
rect 369 310 403 344
rect 610 310 644 344
rect 825 286 859 320
rect 506 67 540 101
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 23 580 89 596
rect 23 546 39 580
rect 73 546 89 580
rect 23 497 89 546
rect 123 572 241 649
rect 123 538 167 572
rect 201 538 241 572
rect 497 580 638 649
rect 123 530 241 538
rect 23 463 39 497
rect 73 463 89 497
rect 282 528 348 560
rect 282 496 298 528
rect 23 414 89 463
rect 23 380 39 414
rect 73 380 89 414
rect 23 364 89 380
rect 137 494 298 496
rect 332 494 348 528
rect 137 462 348 494
rect 497 546 513 580
rect 547 546 588 580
rect 622 546 638 580
rect 497 496 638 546
rect 497 462 513 496
rect 547 462 588 496
rect 622 462 638 496
rect 672 580 728 596
rect 672 546 678 580
rect 712 546 728 580
rect 672 470 728 546
rect 23 226 71 364
rect 137 326 171 462
rect 672 436 678 470
rect 712 436 728 470
rect 672 428 728 436
rect 105 310 171 326
rect 105 276 121 310
rect 155 276 171 310
rect 239 394 728 428
rect 762 580 828 649
rect 762 546 778 580
rect 812 546 828 580
rect 762 470 828 546
rect 762 436 778 470
rect 812 436 828 470
rect 762 420 828 436
rect 862 580 943 596
rect 862 546 878 580
rect 912 546 943 580
rect 862 500 943 546
rect 862 466 878 500
rect 912 466 943 500
rect 862 420 943 466
rect 239 344 305 394
rect 239 310 255 344
rect 289 310 305 344
rect 239 294 305 310
rect 353 344 660 360
rect 353 310 369 344
rect 403 310 610 344
rect 644 310 660 344
rect 353 294 419 310
rect 594 294 660 310
rect 694 336 728 394
rect 862 386 878 420
rect 912 386 943 420
rect 862 370 943 386
rect 694 320 875 336
rect 105 260 171 276
rect 694 286 825 320
rect 859 286 875 320
rect 492 260 558 271
rect 137 238 280 260
rect 137 226 230 238
rect 23 210 89 226
rect 23 176 39 210
rect 73 176 89 210
rect 214 204 230 226
rect 264 204 280 238
rect 214 182 280 204
rect 316 244 558 260
rect 694 270 875 286
rect 694 251 728 270
rect 350 236 558 244
rect 350 226 508 236
rect 23 120 89 176
rect 316 176 350 210
rect 492 202 508 226
rect 542 202 558 236
rect 23 86 39 120
rect 73 86 89 120
rect 23 70 89 86
rect 125 120 175 159
rect 316 126 350 142
rect 386 176 456 192
rect 386 142 404 176
rect 438 142 456 176
rect 492 168 558 202
rect 604 235 728 251
rect 909 236 943 370
rect 604 201 620 235
rect 654 217 728 235
rect 762 229 828 236
rect 654 201 670 217
rect 159 86 175 120
rect 125 17 175 86
rect 386 17 456 142
rect 604 165 670 201
rect 490 101 556 134
rect 604 131 620 165
rect 654 131 670 165
rect 604 115 670 131
rect 762 195 778 229
rect 812 195 828 229
rect 762 161 828 195
rect 762 127 778 161
rect 812 127 828 161
rect 490 67 506 101
rect 540 67 556 101
rect 490 51 556 67
rect 762 17 828 127
rect 862 220 943 236
rect 862 186 878 220
rect 912 186 943 220
rect 862 145 943 186
rect 862 111 878 145
rect 912 111 943 145
rect 862 95 943 111
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
rlabel comment s 0 0 0 0 4 ha_1
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 31 94 65 128 0 FreeSans 340 0 0 0 SUM
port 8 nsew
flabel corelocali s 31 168 65 202 0 FreeSans 340 0 0 0 SUM
port 8 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 SUM
port 8 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 SUM
port 8 nsew
flabel corelocali s 31 390 65 424 0 FreeSans 340 0 0 0 SUM
port 8 nsew
flabel corelocali s 31 464 65 498 0 FreeSans 340 0 0 0 SUM
port 8 nsew
flabel corelocali s 31 538 65 572 0 FreeSans 340 0 0 0 SUM
port 8 nsew
flabel corelocali s 895 390 929 424 0 FreeSans 340 0 0 0 COUT
port 7 nsew
flabel corelocali s 895 464 929 498 0 FreeSans 340 0 0 0 COUT
port 7 nsew
flabel corelocali s 895 538 929 572 0 FreeSans 340 0 0 0 COUT
port 7 nsew
flabel corelocali s 511 94 545 128 0 FreeSans 340 0 0 0 A
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 960 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2383768
string GDS_START 2374626
<< end >>
