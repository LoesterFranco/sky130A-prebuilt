magic
tech sky130A
magscale 1 2
timestamp 1604502729
<< locali >>
rect 123 394 189 596
rect 323 394 389 596
rect 25 360 389 394
rect 25 226 71 360
rect 501 287 567 356
rect 690 290 756 356
rect 25 192 352 226
rect 116 70 166 192
rect 302 70 352 192
rect 985 290 1167 356
rect 1215 290 1319 356
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 23 428 89 649
rect 223 428 289 649
rect 423 458 489 649
rect 555 424 621 563
rect 655 458 721 649
rect 758 424 824 563
rect 865 458 931 649
rect 965 581 1221 615
rect 965 458 1031 581
rect 1065 424 1131 547
rect 423 390 1131 424
rect 1171 390 1221 581
rect 1255 390 1321 649
rect 423 326 457 390
rect 123 260 457 326
rect 30 17 80 158
rect 202 17 268 158
rect 388 17 454 226
rect 506 85 556 253
rect 608 153 642 257
rect 790 256 824 390
rect 678 222 824 256
rect 880 256 930 257
rect 880 222 1321 256
rect 678 187 744 222
rect 778 153 844 188
rect 608 119 844 153
rect 880 85 930 222
rect 506 51 930 85
rect 966 17 1035 187
rect 1069 121 1119 222
rect 1155 17 1221 188
rect 1255 121 1321 222
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
<< metal1 >>
rect 0 683 1344 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 0 617 1344 649
rect 0 17 1344 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
rect 0 -49 1344 -17
<< labels >>
rlabel locali s 1215 290 1319 356 6 A1
port 1 nsew signal input
rlabel locali s 985 290 1167 356 6 A2
port 2 nsew signal input
rlabel locali s 501 287 567 356 6 B1
port 3 nsew signal input
rlabel locali s 690 290 756 356 6 C1
port 4 nsew signal input
rlabel locali s 323 394 389 596 6 X
port 5 nsew signal output
rlabel locali s 302 70 352 192 6 X
port 5 nsew signal output
rlabel locali s 123 394 189 596 6 X
port 5 nsew signal output
rlabel locali s 116 70 166 192 6 X
port 5 nsew signal output
rlabel locali s 25 360 389 394 6 X
port 5 nsew signal output
rlabel locali s 25 226 71 360 6 X
port 5 nsew signal output
rlabel locali s 25 192 352 226 6 X
port 5 nsew signal output
rlabel metal1 s 0 -49 1344 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 1344 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1344 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1777828
string GDS_START 1766756
<< end >>
