magic
tech sky130A
magscale 1 2
timestamp 1601050082
<< locali >>
rect 165 497 271 615
rect 17 169 79 467
rect 211 199 271 497
rect 17 51 123 169
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 288 683
rect 57 501 123 649
rect 165 17 231 165
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 288 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
<< metal1 >>
rect 0 683 288 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 288 683
rect 0 617 288 649
rect 0 17 288 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 288 17
rect 0 -49 288 -17
<< labels >>
rlabel locali s 17 169 79 467 6 HI
port 1 nsew signal output
rlabel locali s 17 51 123 169 6 HI
port 1 nsew signal output
rlabel locali s 211 199 271 497 6 LO
port 2 nsew signal output
rlabel locali s 165 497 271 615 6 LO
port 2 nsew signal output
rlabel metal1 s 0 -49 288 49 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 617 288 715 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 288 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3431206
string GDS_START 3426798
<< end >>
