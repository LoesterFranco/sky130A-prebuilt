magic
tech sky130A
magscale 1 2
timestamp 1601050088
<< locali >>
rect 17 364 89 596
rect 17 226 51 364
rect 191 270 263 356
rect 299 270 365 356
rect 407 270 473 356
rect 507 270 579 356
rect 682 236 747 356
rect 17 70 112 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 123 458 189 649
rect 441 424 519 576
rect 664 458 730 649
rect 123 390 647 424
rect 682 394 730 458
rect 123 330 157 390
rect 85 264 157 330
rect 613 236 647 390
rect 146 17 212 206
rect 246 202 512 236
rect 246 70 312 202
rect 346 17 412 164
rect 446 104 512 202
rect 546 202 647 236
rect 546 140 645 202
rect 681 104 731 202
rect 446 68 731 104
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel locali s 191 270 263 356 6 A1
port 1 nsew signal input
rlabel locali s 299 270 365 356 6 A2
port 2 nsew signal input
rlabel locali s 407 270 473 356 6 A3
port 3 nsew signal input
rlabel locali s 682 236 747 356 6 B1
port 4 nsew signal input
rlabel locali s 507 270 579 356 6 B2
port 5 nsew signal input
rlabel locali s 17 364 89 596 6 X
port 6 nsew signal output
rlabel locali s 17 226 51 364 6 X
port 6 nsew signal output
rlabel locali s 17 70 112 226 6 X
port 6 nsew signal output
rlabel metal1 s 0 -49 768 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 617 768 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 672486
string GDS_START 665594
<< end >>
