magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 19 195 89 325
rect 372 157 406 337
rect 551 271 625 337
rect 663 157 707 223
rect 763 211 869 331
rect 372 123 707 157
rect 1996 301 2088 493
rect 2044 165 2088 301
rect 1992 61 2088 165
rect 2323 53 2374 465
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2392 561
rect 35 393 69 493
rect 103 427 179 527
rect 35 359 179 393
rect 133 194 179 359
rect 133 161 172 194
rect 35 127 172 161
rect 35 69 69 127
rect 103 17 179 93
rect 223 69 257 493
rect 304 415 361 489
rect 395 449 471 527
rect 575 449 774 483
rect 304 372 706 415
rect 304 89 338 372
rect 450 225 484 372
rect 667 337 706 372
rect 740 399 774 449
rect 818 433 852 527
rect 903 414 960 488
rect 999 438 1243 472
rect 903 399 937 414
rect 740 365 937 399
rect 667 271 711 337
rect 450 191 539 225
rect 903 177 937 365
rect 741 143 937 177
rect 741 89 775 143
rect 304 51 381 89
rect 429 17 495 89
rect 610 55 775 89
rect 819 17 859 109
rect 903 107 937 143
rect 971 207 1029 381
rect 1067 331 1165 402
rect 1199 315 1243 438
rect 1277 367 1311 527
rect 1345 427 1405 493
rect 1450 433 1657 467
rect 1199 297 1311 315
rect 1141 263 1311 297
rect 971 141 1097 207
rect 1141 107 1175 263
rect 1277 249 1311 263
rect 1219 213 1253 219
rect 1345 213 1389 427
rect 1423 249 1471 393
rect 1505 315 1579 381
rect 1219 153 1389 213
rect 1505 207 1543 315
rect 1623 281 1657 433
rect 1703 427 1764 527
rect 1822 381 1880 491
rect 1697 315 1880 381
rect 1924 325 1958 527
rect 903 73 973 107
rect 1017 73 1175 107
rect 1235 17 1309 117
rect 1345 107 1389 153
rect 1423 141 1543 207
rect 1587 265 1657 281
rect 1843 265 1880 315
rect 1587 199 1809 265
rect 1843 199 2010 265
rect 1587 107 1631 199
rect 1843 165 1880 199
rect 1345 73 1447 107
rect 1503 73 1631 107
rect 1676 17 1760 123
rect 1814 60 1880 165
rect 1924 17 1958 139
rect 2122 265 2172 485
rect 2218 299 2279 527
rect 2122 199 2288 265
rect 2122 69 2172 199
rect 2213 17 2279 161
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2392 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
<< metal1 >>
rect 0 561 2392 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2392 561
rect 0 496 2392 527
rect 0 17 2392 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2392 17
rect 0 -48 2392 -17
<< obsm1 >>
rect 127 388 185 397
rect 1111 388 1169 397
rect 1423 388 1481 397
rect 127 360 1481 388
rect 127 351 185 360
rect 1111 351 1169 360
rect 1423 351 1481 360
rect 1029 184 1087 193
rect 1425 184 1483 193
rect 1029 156 1483 184
rect 1029 147 1087 156
rect 1425 147 1483 156
rect 201 116 269 125
rect 1029 116 1057 147
rect 201 88 1057 116
rect 201 79 269 88
<< labels >>
rlabel locali s 19 195 89 325 6 CLK
port 1 nsew signal input
rlabel locali s 551 271 625 337 6 D
port 2 nsew signal input
rlabel locali s 2044 165 2088 301 6 Q
port 3 nsew signal output
rlabel locali s 1996 301 2088 493 6 Q
port 3 nsew signal output
rlabel locali s 1992 61 2088 165 6 Q
port 3 nsew signal output
rlabel locali s 2323 53 2374 465 6 Q_N
port 4 nsew signal output
rlabel locali s 763 211 869 331 6 SCD
port 5 nsew signal input
rlabel locali s 663 157 707 223 6 SCE
port 6 nsew signal input
rlabel locali s 372 157 406 337 6 SCE
port 6 nsew signal input
rlabel locali s 372 123 707 157 6 SCE
port 6 nsew signal input
rlabel metal1 s 0 -48 2392 48 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 496 2392 592 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2392 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 302806
string GDS_START 285468
<< end >>
