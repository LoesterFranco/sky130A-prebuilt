magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 949 323 1025 493
rect 1137 323 1213 493
rect 1325 323 1401 493
rect 1513 323 1589 493
rect 1701 323 1777 493
rect 1889 323 1965 493
rect 2077 323 2153 493
rect 2265 323 2341 493
rect 949 289 2441 323
rect 18 215 273 255
rect 2386 181 2441 289
rect 949 147 2441 181
rect 949 52 1025 147
rect 949 51 1009 52
rect 1137 52 1213 147
rect 1163 51 1197 52
rect 1325 52 1401 147
rect 1351 51 1385 52
rect 1513 52 1589 147
rect 1701 52 1777 147
rect 1889 52 1965 147
rect 2077 52 2153 147
rect 2265 52 2341 147
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2484 561
rect 19 323 85 493
rect 129 357 163 527
rect 197 323 273 493
rect 317 357 351 527
rect 385 323 461 493
rect 505 367 539 527
rect 573 323 649 493
rect 693 367 727 527
rect 761 323 837 493
rect 881 367 915 527
rect 1069 367 1103 527
rect 1257 367 1291 527
rect 1445 367 1479 527
rect 1633 367 1667 527
rect 1821 367 1855 527
rect 2009 367 2043 527
rect 2197 367 2231 527
rect 2385 367 2419 527
rect 19 289 351 323
rect 385 289 915 323
rect 317 255 351 289
rect 880 255 915 289
rect 317 215 829 255
rect 880 215 2342 255
rect 317 181 351 215
rect 880 181 915 215
rect 19 147 351 181
rect 385 147 915 181
rect 19 52 85 147
rect 129 17 163 113
rect 197 52 273 147
rect 317 17 351 113
rect 385 52 461 147
rect 505 17 539 113
rect 573 52 649 147
rect 693 17 727 113
rect 761 52 837 147
rect 881 17 915 113
rect 1069 17 1103 113
rect 1257 17 1291 113
rect 1445 17 1479 113
rect 1633 17 1667 113
rect 1821 17 1855 113
rect 2009 17 2043 113
rect 2197 17 2231 113
rect 2385 17 2419 113
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2484 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
<< metal1 >>
rect 0 561 2484 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2484 561
rect 0 496 2484 527
rect 0 17 2484 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2484 17
rect 0 -48 2484 -17
<< labels >>
rlabel locali s 18 215 273 255 6 A
port 1 nsew signal input
rlabel locali s 2386 181 2441 289 6 Y
port 2 nsew signal output
rlabel locali s 2265 323 2341 493 6 Y
port 2 nsew signal output
rlabel locali s 2265 52 2341 147 6 Y
port 2 nsew signal output
rlabel locali s 2077 323 2153 493 6 Y
port 2 nsew signal output
rlabel locali s 2077 52 2153 147 6 Y
port 2 nsew signal output
rlabel locali s 1889 323 1965 493 6 Y
port 2 nsew signal output
rlabel locali s 1889 52 1965 147 6 Y
port 2 nsew signal output
rlabel locali s 1701 323 1777 493 6 Y
port 2 nsew signal output
rlabel locali s 1701 52 1777 147 6 Y
port 2 nsew signal output
rlabel locali s 1513 323 1589 493 6 Y
port 2 nsew signal output
rlabel locali s 1513 52 1589 147 6 Y
port 2 nsew signal output
rlabel locali s 1351 51 1385 52 6 Y
port 2 nsew signal output
rlabel locali s 1325 323 1401 493 6 Y
port 2 nsew signal output
rlabel locali s 1325 52 1401 147 6 Y
port 2 nsew signal output
rlabel locali s 1163 51 1197 52 6 Y
port 2 nsew signal output
rlabel locali s 1137 323 1213 493 6 Y
port 2 nsew signal output
rlabel locali s 1137 52 1213 147 6 Y
port 2 nsew signal output
rlabel locali s 949 323 1025 493 6 Y
port 2 nsew signal output
rlabel locali s 949 289 2441 323 6 Y
port 2 nsew signal output
rlabel locali s 949 147 2441 181 6 Y
port 2 nsew signal output
rlabel locali s 949 52 1025 147 6 Y
port 2 nsew signal output
rlabel locali s 949 51 1009 52 6 Y
port 2 nsew signal output
rlabel metal1 s 0 -48 2484 48 8 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 496 2484 592 6 VPWR
port 4 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2484 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1732416
string GDS_START 1714374
<< end >>
