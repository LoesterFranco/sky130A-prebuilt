magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 1009 391 1043 493
rect 1197 391 1231 493
rect 987 357 1356 391
rect 29 289 631 323
rect 29 215 105 289
rect 155 181 251 255
rect 291 215 371 255
rect 437 215 513 255
rect 555 215 631 289
rect 437 181 474 215
rect 155 147 474 181
rect 785 215 891 257
rect 843 149 891 215
rect 1317 165 1356 357
rect 981 131 1356 165
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 35 391 69 493
rect 103 425 179 527
rect 223 391 257 493
rect 291 425 367 527
rect 411 391 445 493
rect 479 425 555 527
rect 623 459 845 493
rect 623 391 657 459
rect 35 357 657 391
rect 691 325 767 423
rect 811 359 845 459
rect 899 425 965 527
rect 1077 425 1153 527
rect 1265 425 1341 527
rect 691 291 964 325
rect 35 17 69 181
rect 691 174 739 291
rect 930 265 964 291
rect 520 161 739 174
rect 520 140 767 161
rect 930 199 1271 265
rect 520 113 554 140
rect 291 79 554 113
rect 590 17 657 106
rect 691 59 767 140
rect 827 17 933 113
rect 1077 17 1153 97
rect 1265 17 1341 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
<< metal1 >>
rect 0 561 1380 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 0 496 1380 527
rect 0 17 1380 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
rect 0 -48 1380 -17
<< labels >>
rlabel locali s 291 215 371 255 6 A1
port 1 nsew signal input
rlabel locali s 437 215 513 255 6 A2
port 2 nsew signal input
rlabel locali s 437 181 474 215 6 A2
port 2 nsew signal input
rlabel locali s 155 181 251 255 6 A2
port 2 nsew signal input
rlabel locali s 155 147 474 181 6 A2
port 2 nsew signal input
rlabel locali s 555 215 631 289 6 A3
port 3 nsew signal input
rlabel locali s 29 289 631 323 6 A3
port 3 nsew signal input
rlabel locali s 29 215 105 289 6 A3
port 3 nsew signal input
rlabel locali s 843 149 891 215 6 B1
port 4 nsew signal input
rlabel locali s 785 215 891 257 6 B1
port 4 nsew signal input
rlabel locali s 1317 165 1356 357 6 X
port 5 nsew signal output
rlabel locali s 1197 391 1231 493 6 X
port 5 nsew signal output
rlabel locali s 1009 391 1043 493 6 X
port 5 nsew signal output
rlabel locali s 987 357 1356 391 6 X
port 5 nsew signal output
rlabel locali s 981 131 1356 165 6 X
port 5 nsew signal output
rlabel metal1 s 0 -48 1380 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 1380 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1380 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1387316
string GDS_START 1377110
<< end >>
