magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 460 561
rect 18 299 84 527
rect 187 435 253 527
rect 375 333 442 489
rect 214 289 291 333
rect 17 199 73 265
rect 18 17 86 163
rect 122 67 211 255
rect 254 199 291 289
rect 325 299 442 333
rect 325 165 359 299
rect 393 199 443 265
rect 276 143 359 165
rect 276 59 357 143
rect 391 17 443 113
rect 0 -17 460 17
<< obsli1 >>
rect 118 401 153 483
rect 294 401 339 483
rect 118 367 339 401
<< metal1 >>
rect 0 496 460 592
rect 0 -48 460 48
<< labels >>
rlabel locali s 254 199 291 289 6 A1
port 1 nsew signal input
rlabel locali s 214 289 291 333 6 A1
port 1 nsew signal input
rlabel locali s 122 67 211 255 6 A2
port 2 nsew signal input
rlabel locali s 17 199 73 265 6 A3
port 3 nsew signal input
rlabel locali s 393 199 443 265 6 B1
port 4 nsew signal input
rlabel locali s 375 333 442 489 6 Y
port 5 nsew signal output
rlabel locali s 325 299 442 333 6 Y
port 5 nsew signal output
rlabel locali s 325 165 359 299 6 Y
port 5 nsew signal output
rlabel locali s 276 143 359 165 6 Y
port 5 nsew signal output
rlabel locali s 276 59 357 143 6 Y
port 5 nsew signal output
rlabel locali s 391 17 443 113 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 18 17 86 163 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 460 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 460 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 187 435 253 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 18 299 84 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 460 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 460 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 460 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3546296
string GDS_START 3541050
<< end >>
