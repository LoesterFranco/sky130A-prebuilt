magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 2154 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 79 47 109 177
rect 173 47 203 177
rect 277 47 307 177
rect 361 47 391 177
rect 455 47 485 177
rect 549 47 579 177
rect 653 47 683 177
rect 747 47 777 177
rect 831 47 861 177
rect 925 47 955 177
rect 1019 47 1049 177
rect 1123 47 1153 177
rect 1311 47 1341 177
rect 1405 47 1435 177
rect 1499 47 1529 177
rect 1603 47 1633 177
rect 1687 47 1717 177
rect 1781 47 1811 177
rect 1875 47 1905 177
rect 1979 47 2009 177
<< pmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 457 297 493 497
rect 551 297 587 497
rect 645 297 681 497
rect 739 297 775 497
rect 833 297 869 497
rect 927 297 963 497
rect 1021 297 1057 497
rect 1115 297 1151 497
rect 1313 297 1349 497
rect 1407 297 1443 497
rect 1501 297 1537 497
rect 1595 297 1631 497
rect 1689 297 1725 497
rect 1783 297 1819 497
rect 1877 297 1913 497
rect 1971 297 2007 497
<< ndiff >>
rect 27 163 79 177
rect 27 129 35 163
rect 69 129 79 163
rect 27 95 79 129
rect 27 61 35 95
rect 69 61 79 95
rect 27 47 79 61
rect 109 163 173 177
rect 109 129 129 163
rect 163 129 173 163
rect 109 95 173 129
rect 109 61 129 95
rect 163 61 173 95
rect 109 47 173 61
rect 203 95 277 177
rect 203 61 223 95
rect 257 61 277 95
rect 203 47 277 61
rect 307 163 361 177
rect 307 129 317 163
rect 351 129 361 163
rect 307 95 361 129
rect 307 61 317 95
rect 351 61 361 95
rect 307 47 361 61
rect 391 163 455 177
rect 391 129 411 163
rect 445 129 455 163
rect 391 47 455 129
rect 485 95 549 177
rect 485 61 505 95
rect 539 61 549 95
rect 485 47 549 61
rect 579 163 653 177
rect 579 129 599 163
rect 633 129 653 163
rect 579 47 653 129
rect 683 95 747 177
rect 683 61 693 95
rect 727 61 747 95
rect 683 47 747 61
rect 777 95 831 177
rect 777 61 787 95
rect 821 61 831 95
rect 777 47 831 61
rect 861 163 925 177
rect 861 129 881 163
rect 915 129 925 163
rect 861 95 925 129
rect 861 61 881 95
rect 915 61 925 95
rect 861 47 925 61
rect 955 95 1019 177
rect 955 61 975 95
rect 1009 61 1019 95
rect 955 47 1019 61
rect 1049 163 1123 177
rect 1049 129 1069 163
rect 1103 129 1123 163
rect 1049 95 1123 129
rect 1049 61 1069 95
rect 1103 61 1123 95
rect 1049 47 1123 61
rect 1153 95 1311 177
rect 1153 61 1163 95
rect 1197 61 1267 95
rect 1301 61 1311 95
rect 1153 47 1311 61
rect 1341 163 1405 177
rect 1341 129 1361 163
rect 1395 129 1405 163
rect 1341 95 1405 129
rect 1341 61 1361 95
rect 1395 61 1405 95
rect 1341 47 1405 61
rect 1435 95 1499 177
rect 1435 61 1455 95
rect 1489 61 1499 95
rect 1435 47 1499 61
rect 1529 163 1603 177
rect 1529 129 1549 163
rect 1583 129 1603 163
rect 1529 95 1603 129
rect 1529 61 1549 95
rect 1583 61 1603 95
rect 1529 47 1603 61
rect 1633 95 1687 177
rect 1633 61 1643 95
rect 1677 61 1687 95
rect 1633 47 1687 61
rect 1717 163 1781 177
rect 1717 129 1737 163
rect 1771 129 1781 163
rect 1717 95 1781 129
rect 1717 61 1737 95
rect 1771 61 1781 95
rect 1717 47 1781 61
rect 1811 95 1875 177
rect 1811 61 1831 95
rect 1865 61 1875 95
rect 1811 47 1875 61
rect 1905 163 1979 177
rect 1905 129 1925 163
rect 1959 129 1979 163
rect 1905 95 1979 129
rect 1905 61 1925 95
rect 1959 61 1979 95
rect 1905 47 1979 61
rect 2009 95 2061 177
rect 2009 61 2019 95
rect 2053 61 2061 95
rect 2009 47 2061 61
<< pdiff >>
rect 27 483 81 497
rect 27 449 35 483
rect 69 449 81 483
rect 27 415 81 449
rect 27 381 35 415
rect 69 381 81 415
rect 27 347 81 381
rect 27 313 35 347
rect 69 313 81 347
rect 27 297 81 313
rect 117 477 175 497
rect 117 443 129 477
rect 163 443 175 477
rect 117 409 175 443
rect 117 375 129 409
rect 163 375 175 409
rect 117 297 175 375
rect 211 477 269 497
rect 211 443 223 477
rect 257 443 269 477
rect 211 409 269 443
rect 211 375 223 409
rect 257 375 269 409
rect 211 341 269 375
rect 211 307 223 341
rect 257 307 269 341
rect 211 297 269 307
rect 305 477 363 497
rect 305 443 317 477
rect 351 443 363 477
rect 305 297 363 443
rect 399 477 457 497
rect 399 443 411 477
rect 445 443 457 477
rect 399 409 457 443
rect 399 375 411 409
rect 445 375 457 409
rect 399 297 457 375
rect 493 477 551 497
rect 493 443 505 477
rect 539 443 551 477
rect 493 297 551 443
rect 587 477 645 497
rect 587 443 599 477
rect 633 443 645 477
rect 587 409 645 443
rect 587 375 599 409
rect 633 375 645 409
rect 587 297 645 375
rect 681 477 739 497
rect 681 443 693 477
rect 727 443 739 477
rect 681 297 739 443
rect 775 477 833 497
rect 775 443 787 477
rect 821 443 833 477
rect 775 409 833 443
rect 775 375 787 409
rect 821 375 833 409
rect 775 297 833 375
rect 869 409 927 497
rect 869 375 881 409
rect 915 375 927 409
rect 869 341 927 375
rect 869 307 881 341
rect 915 307 927 341
rect 869 297 927 307
rect 963 477 1021 497
rect 963 443 975 477
rect 1009 443 1021 477
rect 963 409 1021 443
rect 963 375 975 409
rect 1009 375 1021 409
rect 963 297 1021 375
rect 1057 409 1115 497
rect 1057 375 1069 409
rect 1103 375 1115 409
rect 1057 341 1115 375
rect 1057 307 1069 341
rect 1103 307 1115 341
rect 1057 297 1115 307
rect 1151 483 1205 497
rect 1151 449 1163 483
rect 1197 449 1205 483
rect 1151 415 1205 449
rect 1151 381 1163 415
rect 1197 381 1205 415
rect 1151 347 1205 381
rect 1151 313 1163 347
rect 1197 313 1205 347
rect 1151 297 1205 313
rect 1259 483 1313 497
rect 1259 449 1267 483
rect 1301 449 1313 483
rect 1259 415 1313 449
rect 1259 381 1267 415
rect 1301 381 1313 415
rect 1259 347 1313 381
rect 1259 313 1267 347
rect 1301 313 1313 347
rect 1259 297 1313 313
rect 1349 477 1407 497
rect 1349 443 1361 477
rect 1395 443 1407 477
rect 1349 409 1407 443
rect 1349 375 1361 409
rect 1395 375 1407 409
rect 1349 297 1407 375
rect 1443 477 1501 497
rect 1443 443 1455 477
rect 1489 443 1501 477
rect 1443 409 1501 443
rect 1443 375 1455 409
rect 1489 375 1501 409
rect 1443 341 1501 375
rect 1443 307 1455 341
rect 1489 307 1501 341
rect 1443 297 1501 307
rect 1537 477 1595 497
rect 1537 443 1549 477
rect 1583 443 1595 477
rect 1537 409 1595 443
rect 1537 375 1549 409
rect 1583 375 1595 409
rect 1537 297 1595 375
rect 1631 477 1689 497
rect 1631 443 1643 477
rect 1677 443 1689 477
rect 1631 409 1689 443
rect 1631 375 1643 409
rect 1677 375 1689 409
rect 1631 341 1689 375
rect 1631 307 1643 341
rect 1677 307 1689 341
rect 1631 297 1689 307
rect 1725 409 1783 497
rect 1725 375 1737 409
rect 1771 375 1783 409
rect 1725 341 1783 375
rect 1725 307 1737 341
rect 1771 307 1783 341
rect 1725 297 1783 307
rect 1819 477 1877 497
rect 1819 443 1831 477
rect 1865 443 1877 477
rect 1819 297 1877 443
rect 1913 409 1971 497
rect 1913 375 1925 409
rect 1959 375 1971 409
rect 1913 341 1971 375
rect 1913 307 1925 341
rect 1959 307 1971 341
rect 1913 297 1971 307
rect 2007 477 2065 497
rect 2007 443 2019 477
rect 2053 443 2065 477
rect 2007 409 2065 443
rect 2007 375 2019 409
rect 2053 375 2065 409
rect 2007 297 2065 375
<< ndiffc >>
rect 35 129 69 163
rect 35 61 69 95
rect 129 129 163 163
rect 129 61 163 95
rect 223 61 257 95
rect 317 129 351 163
rect 317 61 351 95
rect 411 129 445 163
rect 505 61 539 95
rect 599 129 633 163
rect 693 61 727 95
rect 787 61 821 95
rect 881 129 915 163
rect 881 61 915 95
rect 975 61 1009 95
rect 1069 129 1103 163
rect 1069 61 1103 95
rect 1163 61 1197 95
rect 1267 61 1301 95
rect 1361 129 1395 163
rect 1361 61 1395 95
rect 1455 61 1489 95
rect 1549 129 1583 163
rect 1549 61 1583 95
rect 1643 61 1677 95
rect 1737 129 1771 163
rect 1737 61 1771 95
rect 1831 61 1865 95
rect 1925 129 1959 163
rect 1925 61 1959 95
rect 2019 61 2053 95
<< pdiffc >>
rect 35 449 69 483
rect 35 381 69 415
rect 35 313 69 347
rect 129 443 163 477
rect 129 375 163 409
rect 223 443 257 477
rect 223 375 257 409
rect 223 307 257 341
rect 317 443 351 477
rect 411 443 445 477
rect 411 375 445 409
rect 505 443 539 477
rect 599 443 633 477
rect 599 375 633 409
rect 693 443 727 477
rect 787 443 821 477
rect 787 375 821 409
rect 881 375 915 409
rect 881 307 915 341
rect 975 443 1009 477
rect 975 375 1009 409
rect 1069 375 1103 409
rect 1069 307 1103 341
rect 1163 449 1197 483
rect 1163 381 1197 415
rect 1163 313 1197 347
rect 1267 449 1301 483
rect 1267 381 1301 415
rect 1267 313 1301 347
rect 1361 443 1395 477
rect 1361 375 1395 409
rect 1455 443 1489 477
rect 1455 375 1489 409
rect 1455 307 1489 341
rect 1549 443 1583 477
rect 1549 375 1583 409
rect 1643 443 1677 477
rect 1643 375 1677 409
rect 1643 307 1677 341
rect 1737 375 1771 409
rect 1737 307 1771 341
rect 1831 443 1865 477
rect 1925 375 1959 409
rect 1925 307 1959 341
rect 2019 443 2053 477
rect 2019 375 2053 409
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 457 497 493 523
rect 551 497 587 523
rect 645 497 681 523
rect 739 497 775 523
rect 833 497 869 523
rect 927 497 963 523
rect 1021 497 1057 523
rect 1115 497 1151 523
rect 1313 497 1349 523
rect 1407 497 1443 523
rect 1501 497 1537 523
rect 1595 497 1631 523
rect 1689 497 1725 523
rect 1783 497 1819 523
rect 1877 497 1913 523
rect 1971 497 2007 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 457 282 493 297
rect 551 282 587 297
rect 645 282 681 297
rect 739 282 775 297
rect 833 282 869 297
rect 927 282 963 297
rect 1021 282 1057 297
rect 1115 282 1151 297
rect 1313 282 1349 297
rect 1407 282 1443 297
rect 1501 282 1537 297
rect 1595 282 1631 297
rect 1689 282 1725 297
rect 1783 282 1819 297
rect 1877 282 1913 297
rect 1971 282 2007 297
rect 79 265 119 282
rect 173 265 213 282
rect 267 265 307 282
rect 79 249 307 265
rect 79 215 94 249
rect 128 215 172 249
rect 206 215 250 249
rect 284 215 307 249
rect 79 199 307 215
rect 79 177 109 199
rect 173 177 203 199
rect 277 177 307 199
rect 361 265 401 282
rect 455 265 495 282
rect 549 265 589 282
rect 643 265 683 282
rect 737 265 777 282
rect 831 265 871 282
rect 925 265 965 282
rect 1019 265 1059 282
rect 1113 265 1153 282
rect 361 249 683 265
rect 361 215 401 249
rect 435 215 469 249
rect 503 215 547 249
rect 581 215 625 249
rect 659 215 683 249
rect 361 199 683 215
rect 725 249 789 265
rect 725 215 735 249
rect 769 215 789 249
rect 725 199 789 215
rect 831 249 1153 265
rect 831 215 926 249
rect 960 215 1004 249
rect 1038 215 1082 249
rect 1116 215 1153 249
rect 831 199 1153 215
rect 361 177 391 199
rect 455 177 485 199
rect 549 177 579 199
rect 653 177 683 199
rect 747 177 777 199
rect 831 177 861 199
rect 925 177 955 199
rect 1019 177 1049 199
rect 1123 177 1153 199
rect 1311 265 1351 282
rect 1405 265 1445 282
rect 1499 265 1539 282
rect 1593 265 1633 282
rect 1311 249 1633 265
rect 1311 215 1330 249
rect 1364 215 1408 249
rect 1442 215 1486 249
rect 1520 215 1633 249
rect 1311 199 1633 215
rect 1311 177 1341 199
rect 1405 177 1435 199
rect 1499 177 1529 199
rect 1603 177 1633 199
rect 1687 265 1727 282
rect 1781 265 1821 282
rect 1875 265 1915 282
rect 1969 265 2009 282
rect 1687 249 2009 265
rect 1687 215 1704 249
rect 1738 215 1782 249
rect 1816 215 1860 249
rect 1894 215 1938 249
rect 1972 215 2009 249
rect 1687 199 2009 215
rect 1687 177 1717 199
rect 1781 177 1811 199
rect 1875 177 1905 199
rect 1979 177 2009 199
rect 79 21 109 47
rect 173 21 203 47
rect 277 21 307 47
rect 361 21 391 47
rect 455 21 485 47
rect 549 21 579 47
rect 653 21 683 47
rect 747 21 777 47
rect 831 21 861 47
rect 925 21 955 47
rect 1019 21 1049 47
rect 1123 21 1153 47
rect 1311 21 1341 47
rect 1405 21 1435 47
rect 1499 21 1529 47
rect 1603 21 1633 47
rect 1687 21 1717 47
rect 1781 21 1811 47
rect 1875 21 1905 47
rect 1979 21 2009 47
<< polycont >>
rect 94 215 128 249
rect 172 215 206 249
rect 250 215 284 249
rect 401 215 435 249
rect 469 215 503 249
rect 547 215 581 249
rect 625 215 659 249
rect 735 215 769 249
rect 926 215 960 249
rect 1004 215 1038 249
rect 1082 215 1116 249
rect 1330 215 1364 249
rect 1408 215 1442 249
rect 1486 215 1520 249
rect 1704 215 1738 249
rect 1782 215 1816 249
rect 1860 215 1894 249
rect 1938 215 1972 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 17 483 85 493
rect 17 449 35 483
rect 69 449 85 483
rect 17 415 85 449
rect 17 381 35 415
rect 69 381 85 415
rect 17 347 85 381
rect 129 477 171 527
rect 163 443 171 477
rect 129 409 171 443
rect 163 375 171 409
rect 129 359 171 375
rect 215 477 263 493
rect 215 443 223 477
rect 257 443 263 477
rect 215 409 263 443
rect 309 477 359 527
rect 309 443 317 477
rect 351 443 359 477
rect 309 427 359 443
rect 403 477 453 493
rect 403 443 411 477
rect 445 443 453 477
rect 215 375 223 409
rect 257 393 263 409
rect 403 409 453 443
rect 497 477 547 527
rect 497 443 505 477
rect 539 443 547 477
rect 497 427 547 443
rect 591 477 641 493
rect 591 443 599 477
rect 633 443 641 477
rect 403 393 411 409
rect 257 375 411 393
rect 445 393 453 409
rect 591 409 641 443
rect 685 477 735 527
rect 685 443 693 477
rect 727 443 735 477
rect 685 427 735 443
rect 779 483 1213 493
rect 779 477 1163 483
rect 779 443 787 477
rect 821 459 975 477
rect 821 443 829 459
rect 591 393 599 409
rect 445 375 599 393
rect 633 393 641 409
rect 779 409 829 443
rect 967 443 975 459
rect 1009 459 1163 477
rect 1009 443 1015 459
rect 779 393 787 409
rect 633 375 787 393
rect 821 375 829 409
rect 215 359 829 375
rect 873 409 923 425
rect 873 375 881 409
rect 915 375 923 409
rect 17 313 35 347
rect 69 325 85 347
rect 215 341 263 359
rect 215 325 223 341
rect 69 313 223 325
rect 17 307 223 313
rect 257 307 263 341
rect 873 341 923 375
rect 967 409 1015 443
rect 1137 449 1163 459
rect 1197 449 1213 483
rect 967 375 975 409
rect 1009 375 1015 409
rect 967 359 1015 375
rect 1049 409 1103 425
rect 1049 375 1069 409
rect 873 323 881 341
rect 17 291 263 307
rect 307 289 795 323
rect 307 257 341 289
rect 20 249 341 257
rect 20 215 94 249
rect 128 215 172 249
rect 206 215 250 249
rect 284 215 341 249
rect 375 249 685 255
rect 375 215 401 249
rect 435 215 469 249
rect 503 215 547 249
rect 581 215 625 249
rect 659 215 685 249
rect 719 249 795 289
rect 719 215 735 249
rect 769 215 795 249
rect 829 307 881 323
rect 915 323 923 341
rect 1049 341 1103 375
rect 1049 323 1069 341
rect 915 307 1069 323
rect 829 283 1103 307
rect 1137 415 1213 449
rect 1137 381 1163 415
rect 1197 381 1213 415
rect 1137 347 1213 381
rect 1137 313 1163 347
rect 1197 313 1213 347
rect 1137 291 1213 313
rect 1251 483 1317 493
rect 1251 449 1267 483
rect 1301 449 1317 483
rect 1251 415 1317 449
rect 1251 381 1267 415
rect 1301 381 1317 415
rect 1251 347 1317 381
rect 1361 477 1403 527
rect 1395 443 1403 477
rect 1361 409 1403 443
rect 1395 375 1403 409
rect 1361 359 1403 375
rect 1448 477 1496 493
rect 1448 443 1455 477
rect 1489 443 1496 477
rect 1448 409 1496 443
rect 1448 375 1455 409
rect 1489 375 1496 409
rect 1251 313 1267 347
rect 1301 325 1317 347
rect 1448 341 1496 375
rect 1541 477 1591 527
rect 1541 443 1549 477
rect 1583 443 1591 477
rect 1541 409 1591 443
rect 1541 375 1549 409
rect 1583 375 1591 409
rect 1541 359 1591 375
rect 1635 477 2062 493
rect 1635 443 1643 477
rect 1677 459 1831 477
rect 1677 443 1685 459
rect 1635 409 1685 443
rect 1823 443 1831 459
rect 1865 459 2019 477
rect 1865 443 1873 459
rect 1635 375 1643 409
rect 1677 375 1685 409
rect 1448 325 1455 341
rect 1301 313 1455 325
rect 1251 307 1455 313
rect 1489 325 1496 341
rect 1635 341 1685 375
rect 1635 325 1643 341
rect 1489 307 1643 325
rect 1677 307 1685 341
rect 1251 291 1685 307
rect 1729 409 1779 425
rect 1729 375 1737 409
rect 1771 375 1779 409
rect 1729 341 1779 375
rect 1823 359 1873 443
rect 2012 443 2019 459
rect 2053 443 2062 477
rect 1917 409 1967 425
rect 1917 375 1925 409
rect 1959 375 1967 409
rect 1729 307 1737 341
rect 1771 325 1779 341
rect 1917 341 1967 375
rect 2012 409 2062 443
rect 2012 375 2019 409
rect 2053 375 2062 409
rect 2012 359 2062 375
rect 1917 325 1925 341
rect 1771 307 1925 325
rect 1959 325 1967 341
rect 1959 307 2092 325
rect 1729 291 2092 307
rect 829 181 873 283
rect 1309 249 1614 255
rect 907 215 926 249
rect 960 215 1004 249
rect 1038 215 1082 249
rect 1116 215 1265 249
rect 1309 215 1330 249
rect 1364 215 1408 249
rect 1442 215 1486 249
rect 1520 215 1614 249
rect 1688 249 1993 255
rect 1688 215 1704 249
rect 1738 215 1782 249
rect 1816 215 1860 249
rect 1894 215 1938 249
rect 1972 215 1993 249
rect 1231 181 1265 215
rect 2027 181 2092 291
rect 35 163 69 179
rect 35 95 69 129
rect 35 17 69 61
rect 103 163 351 181
rect 103 129 129 163
rect 163 145 317 163
rect 163 129 179 145
rect 103 95 179 129
rect 291 129 317 145
rect 385 163 1119 181
rect 385 129 411 163
rect 445 129 599 163
rect 633 145 881 163
rect 633 129 659 145
rect 855 129 881 145
rect 915 145 1069 163
rect 915 129 931 145
rect 103 61 129 95
rect 163 61 179 95
rect 103 51 179 61
rect 223 95 257 111
rect 223 17 257 61
rect 291 95 351 129
rect 787 95 821 111
rect 291 61 317 95
rect 351 61 505 95
rect 539 61 693 95
rect 727 61 743 95
rect 291 51 743 61
rect 787 17 821 61
rect 855 95 931 129
rect 1043 129 1069 145
rect 1103 129 1119 163
rect 1231 163 2092 181
rect 1231 147 1361 163
rect 855 61 881 95
rect 915 61 931 95
rect 855 55 931 61
rect 975 95 1009 111
rect 975 17 1009 61
rect 1043 95 1119 129
rect 1335 129 1361 147
rect 1395 145 1549 163
rect 1395 129 1411 145
rect 1043 61 1069 95
rect 1103 61 1119 95
rect 1043 55 1119 61
rect 1163 95 1301 111
rect 1197 61 1267 95
rect 1163 17 1301 61
rect 1335 95 1411 129
rect 1523 129 1549 145
rect 1583 145 1737 163
rect 1583 129 1599 145
rect 1335 61 1361 95
rect 1395 61 1411 95
rect 1335 51 1411 61
rect 1455 95 1489 111
rect 1455 17 1489 61
rect 1523 95 1599 129
rect 1711 129 1737 145
rect 1771 145 1925 163
rect 1771 129 1787 145
rect 1523 61 1549 95
rect 1583 61 1599 95
rect 1523 51 1599 61
rect 1643 95 1677 111
rect 1643 17 1677 61
rect 1711 95 1787 129
rect 1899 129 1925 145
rect 1959 147 2092 163
rect 1959 129 1975 147
rect 1711 61 1737 95
rect 1771 61 1787 95
rect 1711 51 1787 61
rect 1831 95 1865 111
rect 1831 17 1865 61
rect 1899 95 1975 129
rect 1899 61 1925 95
rect 1959 61 1975 95
rect 1899 51 1975 61
rect 2019 95 2053 111
rect 2019 17 2053 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
<< metal1 >>
rect 0 561 2116 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 0 496 2116 527
rect 0 17 2116 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
rect 0 -48 2116 -17
<< labels >>
flabel corelocali s 967 306 967 306 0 FreeSans 400 0 0 0 Y
port 9 nsew
flabel corelocali s 1745 238 1745 238 0 FreeSans 400 180 0 0 A2_N
port 2 nsew
flabel corelocali s 415 238 415 238 0 FreeSans 400 180 0 0 B2
port 4 nsew
flabel corelocali s 1339 238 1339 238 0 FreeSans 400 0 0 0 A1_N
port 1 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 400 0 0 0 B1
port 3 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 2116 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1363674
string GDS_START 1348580
<< end >>
