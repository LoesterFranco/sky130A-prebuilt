magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 85 199 166 339
rect 200 199 254 265
rect 607 289 846 341
rect 762 181 846 289
rect 880 215 1059 255
rect 1093 215 1266 255
rect 419 145 1167 181
rect 419 51 495 145
rect 607 51 683 145
rect 903 51 979 145
rect 1091 51 1167 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 17 411 69 491
rect 103 448 179 527
rect 335 445 777 493
rect 819 443 1065 493
rect 17 377 390 411
rect 17 165 51 377
rect 209 305 322 343
rect 288 249 322 305
rect 356 317 390 377
rect 429 375 979 409
rect 356 283 573 317
rect 921 291 979 375
rect 1023 325 1065 443
rect 1109 359 1151 527
rect 1185 325 1261 493
rect 1023 291 1261 325
rect 539 255 573 283
rect 288 215 495 249
rect 539 215 728 255
rect 288 165 322 215
rect 17 90 93 165
rect 137 17 171 165
rect 231 131 322 165
rect 231 90 270 131
rect 319 17 385 96
rect 539 17 573 111
rect 727 17 869 111
rect 1023 17 1057 111
rect 1211 17 1266 181
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
rlabel locali s 1093 215 1266 255 6 A
port 1 nsew signal input
rlabel locali s 880 215 1059 255 6 B
port 2 nsew signal input
rlabel locali s 200 199 254 265 6 C_N
port 3 nsew signal input
rlabel locali s 85 199 166 339 6 D_N
port 4 nsew signal input
rlabel locali s 1091 51 1167 145 6 Y
port 5 nsew signal output
rlabel locali s 903 51 979 145 6 Y
port 5 nsew signal output
rlabel locali s 762 181 846 289 6 Y
port 5 nsew signal output
rlabel locali s 607 289 846 341 6 Y
port 5 nsew signal output
rlabel locali s 607 51 683 145 6 Y
port 5 nsew signal output
rlabel locali s 419 145 1167 181 6 Y
port 5 nsew signal output
rlabel locali s 419 51 495 145 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -48 1288 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 1288 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1288 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2546740
string GDS_START 2537208
<< end >>
