magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 1958 704
<< pwell >>
rect 0 0 1920 49
<< scnmos >>
rect 84 74 114 222
rect 212 74 242 222
rect 502 119 532 203
rect 588 119 618 203
rect 683 102 713 186
rect 755 102 785 186
rect 873 76 903 186
rect 975 120 1005 230
rect 1113 146 1143 230
rect 1191 146 1221 230
rect 1389 74 1419 184
rect 1503 74 1533 222
rect 1701 112 1731 222
rect 1803 74 1833 222
<< pmoshvt >>
rect 85 368 115 592
rect 175 368 205 592
rect 390 503 420 587
rect 513 447 543 531
rect 620 508 650 592
rect 704 508 734 592
rect 870 424 900 592
rect 1021 424 1051 592
rect 1128 482 1158 566
rect 1206 482 1236 566
rect 1405 368 1435 568
rect 1506 368 1536 592
rect 1704 368 1734 536
rect 1805 368 1835 592
<< ndiff >>
rect 257 248 315 260
rect 257 222 269 248
rect 27 153 84 222
rect 27 119 39 153
rect 73 119 84 153
rect 27 74 84 119
rect 114 96 212 222
rect 114 74 146 96
rect 129 62 146 74
rect 180 74 212 96
rect 242 214 269 222
rect 303 214 315 248
rect 242 74 315 214
rect 180 62 197 74
rect 129 50 197 62
rect 375 119 502 203
rect 532 180 588 203
rect 532 146 543 180
rect 577 146 588 180
rect 532 119 588 146
rect 618 186 668 203
rect 918 218 975 230
rect 918 186 930 218
rect 618 171 683 186
rect 618 137 629 171
rect 663 137 683 171
rect 618 119 683 137
rect 375 112 452 119
rect 375 78 389 112
rect 423 78 452 112
rect 633 102 683 119
rect 713 102 755 186
rect 785 102 873 186
rect 375 66 452 78
rect 800 82 873 102
rect 800 48 812 82
rect 846 76 873 82
rect 903 184 930 186
rect 964 184 975 218
rect 903 120 975 184
rect 1005 208 1113 230
rect 1005 174 1041 208
rect 1075 174 1113 208
rect 1005 146 1113 174
rect 1143 146 1191 230
rect 1221 192 1278 230
rect 1221 158 1232 192
rect 1266 158 1278 192
rect 1453 184 1503 222
rect 1221 146 1278 158
rect 1332 146 1389 184
rect 1005 120 1055 146
rect 903 76 953 120
rect 846 48 858 76
rect 1332 112 1344 146
rect 1378 112 1389 146
rect 1332 74 1389 112
rect 1419 120 1503 184
rect 1419 86 1444 120
rect 1478 86 1503 120
rect 1419 74 1503 86
rect 1533 210 1590 222
rect 1533 176 1544 210
rect 1578 176 1590 210
rect 1533 120 1590 176
rect 1533 86 1544 120
rect 1578 86 1590 120
rect 1644 184 1701 222
rect 1644 150 1656 184
rect 1690 150 1701 184
rect 1644 112 1701 150
rect 1731 210 1803 222
rect 1731 176 1758 210
rect 1792 176 1803 210
rect 1731 120 1803 176
rect 1731 112 1758 120
rect 1746 86 1758 112
rect 1792 86 1803 120
rect 1533 74 1590 86
rect 1746 74 1803 86
rect 1833 210 1890 222
rect 1833 176 1844 210
rect 1878 176 1890 210
rect 1833 120 1890 176
rect 1833 86 1844 120
rect 1878 86 1890 120
rect 1833 74 1890 86
rect 800 36 858 48
<< pdiff >>
rect 316 627 372 639
rect 316 593 327 627
rect 361 593 372 627
rect 752 619 822 631
rect 27 580 85 592
rect 27 546 38 580
rect 72 546 85 580
rect 27 497 85 546
rect 27 463 38 497
rect 72 463 85 497
rect 27 414 85 463
rect 27 380 38 414
rect 72 380 85 414
rect 27 368 85 380
rect 115 580 175 592
rect 115 546 128 580
rect 162 546 175 580
rect 115 462 175 546
rect 115 428 128 462
rect 162 428 175 462
rect 115 368 175 428
rect 205 580 262 592
rect 205 546 218 580
rect 252 546 262 580
rect 205 497 262 546
rect 316 587 372 593
rect 752 592 770 619
rect 316 503 390 587
rect 420 531 473 587
rect 567 531 620 592
rect 420 503 513 531
rect 205 463 218 497
rect 252 463 262 497
rect 205 414 262 463
rect 205 380 218 414
rect 252 380 262 414
rect 438 459 513 503
rect 438 425 450 459
rect 484 447 513 459
rect 543 508 620 531
rect 650 508 704 592
rect 734 585 770 592
rect 804 592 822 619
rect 804 585 870 592
rect 734 508 870 585
rect 543 493 602 508
rect 543 459 556 493
rect 590 459 602 493
rect 543 447 602 459
rect 484 425 495 447
rect 438 413 495 425
rect 205 368 262 380
rect 817 424 870 508
rect 900 501 1021 592
rect 900 467 928 501
rect 962 467 1021 501
rect 900 424 1021 467
rect 1051 566 1104 592
rect 1453 568 1506 592
rect 1051 526 1128 566
rect 1051 492 1064 526
rect 1098 492 1128 526
rect 1051 482 1128 492
rect 1158 482 1206 566
rect 1236 541 1293 566
rect 1236 507 1249 541
rect 1283 507 1293 541
rect 1236 482 1293 507
rect 1347 556 1405 568
rect 1347 522 1358 556
rect 1392 522 1405 556
rect 1347 485 1405 522
rect 1051 424 1110 482
rect 1347 451 1358 485
rect 1392 451 1405 485
rect 1347 414 1405 451
rect 1347 380 1358 414
rect 1392 380 1405 414
rect 1347 368 1405 380
rect 1435 556 1506 568
rect 1435 522 1448 556
rect 1482 522 1506 556
rect 1435 456 1506 522
rect 1435 422 1448 456
rect 1482 422 1506 456
rect 1435 368 1506 422
rect 1536 580 1593 592
rect 1536 546 1549 580
rect 1583 546 1593 580
rect 1536 456 1593 546
rect 1752 536 1805 592
rect 1536 422 1549 456
rect 1583 422 1593 456
rect 1536 368 1593 422
rect 1647 524 1704 536
rect 1647 490 1657 524
rect 1691 490 1704 524
rect 1647 414 1704 490
rect 1647 380 1657 414
rect 1691 380 1704 414
rect 1647 368 1704 380
rect 1734 524 1805 536
rect 1734 490 1747 524
rect 1781 490 1805 524
rect 1734 414 1805 490
rect 1734 380 1747 414
rect 1781 380 1805 414
rect 1734 368 1805 380
rect 1835 580 1893 592
rect 1835 546 1848 580
rect 1882 546 1893 580
rect 1835 497 1893 546
rect 1835 463 1848 497
rect 1882 463 1893 497
rect 1835 414 1893 463
rect 1835 380 1848 414
rect 1882 380 1893 414
rect 1835 368 1893 380
<< ndiffc >>
rect 39 119 73 153
rect 146 62 180 96
rect 269 214 303 248
rect 543 146 577 180
rect 629 137 663 171
rect 389 78 423 112
rect 812 48 846 82
rect 930 184 964 218
rect 1041 174 1075 208
rect 1232 158 1266 192
rect 1344 112 1378 146
rect 1444 86 1478 120
rect 1544 176 1578 210
rect 1544 86 1578 120
rect 1656 150 1690 184
rect 1758 176 1792 210
rect 1758 86 1792 120
rect 1844 176 1878 210
rect 1844 86 1878 120
<< pdiffc >>
rect 327 593 361 627
rect 38 546 72 580
rect 38 463 72 497
rect 38 380 72 414
rect 128 546 162 580
rect 128 428 162 462
rect 218 546 252 580
rect 218 463 252 497
rect 218 380 252 414
rect 450 425 484 459
rect 770 585 804 619
rect 556 459 590 493
rect 928 467 962 501
rect 1064 492 1098 526
rect 1249 507 1283 541
rect 1358 522 1392 556
rect 1358 451 1392 485
rect 1358 380 1392 414
rect 1448 522 1482 556
rect 1448 422 1482 456
rect 1549 546 1583 580
rect 1549 422 1583 456
rect 1657 490 1691 524
rect 1657 380 1691 414
rect 1747 490 1781 524
rect 1747 380 1781 414
rect 1848 546 1882 580
rect 1848 463 1882 497
rect 1848 380 1882 414
<< poly >>
rect 85 592 115 618
rect 175 592 205 618
rect 390 587 420 613
rect 620 592 650 618
rect 704 592 734 618
rect 513 531 543 557
rect 390 488 420 503
rect 387 471 423 488
rect 340 455 423 471
rect 340 421 356 455
rect 390 421 423 455
rect 340 405 423 421
rect 870 592 900 618
rect 1021 592 1051 618
rect 620 493 650 508
rect 704 493 734 508
rect 513 432 543 447
rect 85 353 115 368
rect 175 353 205 368
rect 510 363 546 432
rect 617 415 653 493
rect 701 463 762 493
rect 82 310 118 353
rect 172 310 208 353
rect 294 347 546 363
rect 294 313 310 347
rect 344 333 546 347
rect 588 399 690 415
rect 588 365 640 399
rect 674 365 690 399
rect 588 349 690 365
rect 344 313 360 333
rect 34 294 118 310
rect 34 260 50 294
rect 84 260 118 294
rect 34 244 118 260
rect 160 294 242 310
rect 294 297 360 313
rect 160 260 176 294
rect 210 260 242 294
rect 160 244 242 260
rect 84 222 114 244
rect 212 222 242 244
rect 84 48 114 74
rect 212 48 242 74
rect 330 51 360 297
rect 402 275 468 291
rect 402 241 418 275
rect 452 255 468 275
rect 452 241 532 255
rect 402 225 532 241
rect 502 203 532 225
rect 588 203 618 349
rect 732 284 762 463
rect 1128 566 1158 592
rect 1206 566 1236 592
rect 1405 568 1435 594
rect 1506 592 1536 618
rect 1805 592 1835 618
rect 1128 467 1158 482
rect 1206 467 1236 482
rect 870 409 900 424
rect 1021 409 1051 424
rect 867 392 903 409
rect 804 376 903 392
rect 1018 379 1083 409
rect 804 342 820 376
rect 854 342 903 376
rect 804 326 903 342
rect 732 258 831 284
rect 732 254 781 258
rect 755 224 781 254
rect 815 224 831 258
rect 683 186 713 212
rect 755 208 831 224
rect 755 186 785 208
rect 873 186 903 326
rect 945 321 1011 337
rect 945 287 961 321
rect 995 287 1011 321
rect 945 271 1011 287
rect 1053 275 1083 379
rect 1125 389 1161 467
rect 1203 437 1312 467
rect 1246 428 1312 437
rect 1246 394 1262 428
rect 1296 394 1312 428
rect 1125 373 1198 389
rect 1125 339 1148 373
rect 1182 339 1198 373
rect 1125 323 1198 339
rect 1246 360 1312 394
rect 1704 536 1734 562
rect 1246 326 1262 360
rect 1296 326 1312 360
rect 1405 353 1435 368
rect 1506 353 1536 368
rect 1704 353 1734 368
rect 1805 353 1835 368
rect 1246 310 1312 326
rect 1246 275 1276 310
rect 1402 304 1438 353
rect 1503 336 1539 353
rect 1701 336 1737 353
rect 1480 320 1737 336
rect 1802 326 1838 353
rect 975 230 1005 271
rect 1053 245 1143 275
rect 1113 230 1143 245
rect 1191 245 1276 275
rect 1360 288 1432 304
rect 1360 254 1376 288
rect 1410 254 1432 288
rect 1480 286 1496 320
rect 1530 306 1737 320
rect 1779 310 1845 326
rect 1530 286 1731 306
rect 1480 270 1731 286
rect 1191 230 1221 245
rect 1360 238 1432 254
rect 502 93 532 119
rect 588 93 618 119
rect 683 51 713 102
rect 755 76 785 102
rect 330 21 713 51
rect 1389 184 1419 238
rect 1503 222 1533 270
rect 1701 222 1731 270
rect 1779 276 1795 310
rect 1829 276 1845 310
rect 1779 260 1845 276
rect 1803 222 1833 260
rect 1113 124 1143 146
rect 975 94 1005 120
rect 1077 108 1143 124
rect 1191 120 1221 146
rect 873 50 903 76
rect 1077 74 1093 108
rect 1127 74 1143 108
rect 1701 86 1731 112
rect 1077 58 1143 74
rect 1389 48 1419 74
rect 1503 48 1533 74
rect 1803 48 1833 74
<< polycont >>
rect 356 421 390 455
rect 310 313 344 347
rect 640 365 674 399
rect 50 260 84 294
rect 176 260 210 294
rect 418 241 452 275
rect 820 342 854 376
rect 781 224 815 258
rect 961 287 995 321
rect 1262 394 1296 428
rect 1148 339 1182 373
rect 1262 326 1296 360
rect 1376 254 1410 288
rect 1496 286 1530 320
rect 1795 276 1829 310
rect 1093 74 1127 108
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 22 580 72 596
rect 22 546 38 580
rect 22 497 72 546
rect 22 463 38 497
rect 22 414 72 463
rect 22 380 38 414
rect 112 580 162 649
rect 311 627 377 649
rect 112 546 128 580
rect 112 462 162 546
rect 112 428 128 462
rect 112 412 162 428
rect 202 580 268 596
rect 202 546 218 580
rect 252 546 268 580
rect 311 593 327 627
rect 361 593 377 627
rect 311 577 377 593
rect 748 619 826 649
rect 748 585 770 619
rect 804 585 826 619
rect 860 581 1198 615
rect 202 543 268 546
rect 411 551 658 577
rect 860 560 1030 581
rect 860 551 894 560
rect 411 543 894 551
rect 202 509 445 543
rect 624 517 894 543
rect 202 497 287 509
rect 202 463 218 497
rect 252 463 287 497
rect 556 493 590 509
rect 202 414 287 463
rect 22 378 72 380
rect 202 380 218 414
rect 252 380 287 414
rect 340 455 416 471
rect 340 421 356 455
rect 390 421 416 455
rect 340 405 416 421
rect 450 459 522 475
rect 484 425 522 459
rect 450 409 522 425
rect 22 344 168 378
rect 202 363 287 380
rect 134 310 168 344
rect 253 347 348 363
rect 253 313 310 347
rect 344 313 348 347
rect 25 294 100 310
rect 25 260 50 294
rect 84 260 100 294
rect 25 236 100 260
rect 134 294 218 310
rect 134 260 176 294
rect 210 260 218 294
rect 23 180 89 202
rect 134 180 218 260
rect 253 297 348 313
rect 382 356 416 405
rect 253 248 319 297
rect 253 214 269 248
rect 303 214 319 248
rect 382 275 454 356
rect 382 241 418 275
rect 452 241 454 275
rect 382 225 454 241
rect 488 248 522 409
rect 928 501 962 523
rect 590 459 856 483
rect 556 449 856 459
rect 556 316 590 449
rect 624 399 731 415
rect 624 365 640 399
rect 674 365 731 399
rect 624 350 731 365
rect 556 282 663 316
rect 488 214 577 248
rect 543 180 577 214
rect 23 153 509 180
rect 23 119 39 153
rect 73 146 509 153
rect 73 119 89 146
rect 23 70 89 119
rect 125 96 201 112
rect 125 62 146 96
rect 180 62 201 96
rect 125 17 201 62
rect 371 78 389 112
rect 423 78 441 112
rect 371 17 441 78
rect 475 85 509 146
rect 543 119 577 146
rect 613 171 663 282
rect 613 137 629 171
rect 613 119 663 137
rect 697 150 731 350
rect 804 376 856 449
rect 928 405 962 467
rect 804 342 820 376
rect 854 342 856 376
rect 804 326 856 342
rect 890 371 962 405
rect 890 274 924 371
rect 996 337 1030 560
rect 765 258 924 274
rect 958 321 1030 337
rect 958 287 961 321
rect 995 287 1030 321
rect 958 271 1030 287
rect 1064 526 1114 547
rect 1098 492 1114 526
rect 1064 423 1114 492
rect 1064 276 1098 423
rect 1164 389 1198 581
rect 1233 541 1299 649
rect 1233 507 1249 541
rect 1283 507 1299 541
rect 1233 478 1299 507
rect 1342 556 1408 572
rect 1342 522 1358 556
rect 1392 522 1408 556
rect 1342 485 1408 522
rect 1342 451 1358 485
rect 1392 451 1408 485
rect 1342 444 1408 451
rect 1132 373 1198 389
rect 1132 339 1148 373
rect 1182 339 1198 373
rect 1132 323 1198 339
rect 1246 428 1408 444
rect 1246 394 1262 428
rect 1296 414 1408 428
rect 1296 394 1358 414
rect 1246 380 1358 394
rect 1392 380 1408 414
rect 1448 556 1498 649
rect 1482 522 1498 556
rect 1448 456 1498 522
rect 1482 422 1498 456
rect 1448 406 1498 422
rect 1533 580 1614 596
rect 1533 546 1549 580
rect 1583 546 1614 580
rect 1533 456 1614 546
rect 1533 422 1549 456
rect 1583 422 1614 456
rect 1533 406 1614 422
rect 1246 372 1408 380
rect 1246 360 1546 372
rect 1246 326 1262 360
rect 1296 338 1546 360
rect 1296 326 1312 338
rect 1246 310 1312 326
rect 1460 320 1546 338
rect 1360 288 1426 304
rect 1360 276 1376 288
rect 765 224 781 258
rect 815 237 924 258
rect 1064 254 1376 276
rect 1410 254 1426 288
rect 1064 242 1426 254
rect 815 224 980 237
rect 1064 224 1118 242
rect 1360 238 1426 242
rect 1460 286 1496 320
rect 1530 286 1546 320
rect 1460 270 1546 286
rect 765 218 980 224
rect 765 203 930 218
rect 914 184 930 203
rect 964 184 980 218
rect 1025 208 1118 224
rect 1025 174 1041 208
rect 1075 174 1118 208
rect 1025 158 1118 174
rect 1216 192 1282 208
rect 1460 204 1494 270
rect 1580 226 1614 406
rect 1216 158 1232 192
rect 1266 158 1282 192
rect 697 124 930 150
rect 697 116 1143 124
rect 697 85 731 116
rect 475 51 731 85
rect 896 108 1143 116
rect 796 48 812 82
rect 846 48 862 82
rect 896 74 1093 108
rect 1127 74 1143 108
rect 896 58 1143 74
rect 796 17 862 48
rect 1216 17 1282 158
rect 1328 170 1494 204
rect 1528 210 1614 226
rect 1528 176 1544 210
rect 1578 176 1614 210
rect 1328 146 1394 170
rect 1328 112 1344 146
rect 1378 112 1394 146
rect 1328 88 1394 112
rect 1428 120 1494 136
rect 1428 86 1444 120
rect 1478 86 1494 120
rect 1428 17 1494 86
rect 1528 120 1614 176
rect 1656 524 1691 540
rect 1656 490 1657 524
rect 1656 414 1691 490
rect 1656 380 1657 414
rect 1656 326 1691 380
rect 1731 524 1797 649
rect 1731 490 1747 524
rect 1781 490 1797 524
rect 1731 414 1797 490
rect 1731 380 1747 414
rect 1781 380 1797 414
rect 1731 364 1797 380
rect 1832 580 1903 596
rect 1832 546 1848 580
rect 1882 546 1903 580
rect 1832 497 1903 546
rect 1832 463 1848 497
rect 1882 463 1903 497
rect 1832 414 1903 463
rect 1832 380 1848 414
rect 1882 380 1903 414
rect 1832 364 1903 380
rect 1656 310 1835 326
rect 1656 276 1795 310
rect 1829 276 1835 310
rect 1656 260 1835 276
rect 1656 184 1706 260
rect 1869 226 1903 364
rect 1690 150 1706 184
rect 1656 125 1706 150
rect 1742 210 1792 226
rect 1742 176 1758 210
rect 1528 86 1544 120
rect 1578 86 1614 120
rect 1528 70 1614 86
rect 1742 120 1792 176
rect 1742 86 1758 120
rect 1742 17 1792 86
rect 1828 210 1903 226
rect 1828 176 1844 210
rect 1878 176 1903 210
rect 1828 120 1903 176
rect 1828 86 1844 120
rect 1878 86 1903 120
rect 1828 70 1903 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
<< metal1 >>
rect 0 683 1920 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 0 617 1920 649
rect 0 17 1920 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
rect 0 -49 1920 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dfxbp_1
flabel pwell s 0 0 1920 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nwell s 0 617 1920 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 0 617 1920 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 1920 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 415 242 449 276 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 1567 464 1601 498 0 FreeSans 340 0 0 0 Q
port 7 nsew
flabel corelocali s 1567 538 1601 572 0 FreeSans 340 0 0 0 Q
port 7 nsew
flabel corelocali s 1855 390 1889 424 0 FreeSans 340 0 0 0 Q_N
port 8 nsew
flabel corelocali s 1855 464 1889 498 0 FreeSans 340 0 0 0 Q_N
port 8 nsew
flabel corelocali s 1855 538 1889 572 0 FreeSans 340 0 0 0 Q_N
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 1920 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2696264
string GDS_START 2681298
<< end >>
