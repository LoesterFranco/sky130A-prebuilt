magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 1094 704
<< pwell >>
rect 0 0 1056 49
<< scnmos >>
rect 95 74 125 222
rect 240 74 270 222
rect 318 74 348 222
rect 459 74 489 222
rect 729 74 759 184
rect 842 74 872 222
rect 928 74 958 222
<< pmoshvt >>
rect 86 368 116 568
rect 176 368 206 568
rect 378 392 408 592
rect 488 392 518 592
rect 730 368 760 536
rect 839 368 869 592
rect 929 368 959 592
<< ndiff >>
rect 38 196 95 222
rect 38 162 50 196
rect 84 162 95 196
rect 38 120 95 162
rect 38 86 50 120
rect 84 86 95 120
rect 38 74 95 86
rect 125 186 240 222
rect 125 152 167 186
rect 201 152 240 186
rect 125 74 240 152
rect 270 74 318 222
rect 348 209 459 222
rect 348 175 359 209
rect 393 175 459 209
rect 348 74 459 175
rect 489 116 548 222
rect 792 184 842 222
rect 489 82 500 116
rect 534 82 548 116
rect 489 74 548 82
rect 672 146 729 184
rect 672 112 684 146
rect 718 112 729 146
rect 672 74 729 112
rect 759 120 842 184
rect 759 86 790 120
rect 824 86 842 120
rect 759 74 842 86
rect 872 207 928 222
rect 872 173 883 207
rect 917 173 928 207
rect 872 74 928 173
rect 958 210 1029 222
rect 958 176 983 210
rect 1017 176 1029 210
rect 958 120 1029 176
rect 958 86 983 120
rect 1017 86 1029 120
rect 958 74 1029 86
<< pdiff >>
rect 319 580 378 592
rect 27 556 86 568
rect 27 522 39 556
rect 73 522 86 556
rect 27 488 86 522
rect 27 454 39 488
rect 73 454 86 488
rect 27 415 86 454
rect 27 381 39 415
rect 73 381 86 415
rect 27 368 86 381
rect 116 529 176 568
rect 116 495 129 529
rect 163 495 176 529
rect 116 421 176 495
rect 116 387 129 421
rect 163 387 176 421
rect 116 368 176 387
rect 206 521 265 568
rect 206 487 219 521
rect 253 487 265 521
rect 206 368 265 487
rect 319 546 331 580
rect 365 546 378 580
rect 319 392 378 546
rect 408 580 488 592
rect 408 546 431 580
rect 465 546 488 580
rect 408 392 488 546
rect 518 580 577 592
rect 518 546 531 580
rect 565 546 577 580
rect 778 580 839 592
rect 518 512 577 546
rect 778 546 791 580
rect 825 546 839 580
rect 778 536 839 546
rect 518 478 531 512
rect 565 478 577 512
rect 518 392 577 478
rect 671 421 730 536
rect 671 387 683 421
rect 717 387 730 421
rect 671 368 730 387
rect 760 368 839 536
rect 869 421 929 592
rect 869 387 882 421
rect 916 387 929 421
rect 869 368 929 387
rect 959 580 1029 592
rect 959 546 977 580
rect 1011 546 1029 580
rect 959 368 1029 546
<< ndiffc >>
rect 50 162 84 196
rect 50 86 84 120
rect 167 152 201 186
rect 359 175 393 209
rect 500 82 534 116
rect 684 112 718 146
rect 790 86 824 120
rect 883 173 917 207
rect 983 176 1017 210
rect 983 86 1017 120
<< pdiffc >>
rect 39 522 73 556
rect 39 454 73 488
rect 39 381 73 415
rect 129 495 163 529
rect 129 387 163 421
rect 219 487 253 521
rect 331 546 365 580
rect 431 546 465 580
rect 531 546 565 580
rect 791 546 825 580
rect 531 478 565 512
rect 683 387 717 421
rect 882 387 916 421
rect 977 546 1011 580
<< poly >>
rect 86 568 116 594
rect 176 568 206 594
rect 378 592 408 618
rect 488 592 518 618
rect 839 592 869 618
rect 929 592 959 618
rect 730 536 760 562
rect 378 377 408 392
rect 488 377 518 392
rect 86 353 116 368
rect 176 353 206 368
rect 375 356 411 377
rect 83 310 119 353
rect 173 310 209 353
rect 318 340 411 356
rect 21 294 125 310
rect 21 260 37 294
rect 71 260 125 294
rect 21 244 125 260
rect 173 294 270 310
rect 173 260 189 294
rect 223 260 270 294
rect 173 244 270 260
rect 95 222 125 244
rect 240 222 270 244
rect 318 306 359 340
rect 393 306 411 340
rect 485 360 521 377
rect 485 344 577 360
rect 730 353 760 368
rect 839 353 869 368
rect 929 353 959 368
rect 485 324 527 344
rect 318 290 411 306
rect 459 310 527 324
rect 561 310 577 344
rect 459 294 577 310
rect 318 222 348 290
rect 459 222 489 294
rect 727 292 763 353
rect 625 276 763 292
rect 836 318 872 353
rect 926 326 962 353
rect 926 318 1033 326
rect 836 310 1033 318
rect 836 290 983 310
rect 625 242 641 276
rect 675 242 763 276
rect 625 226 763 242
rect 842 276 983 290
rect 1017 276 1033 310
rect 842 260 1033 276
rect 729 184 759 226
rect 842 222 872 260
rect 928 222 958 260
rect 95 48 125 74
rect 240 48 270 74
rect 318 48 348 74
rect 459 48 489 74
rect 729 48 759 74
rect 842 48 872 74
rect 928 48 958 74
<< polycont >>
rect 37 260 71 294
rect 189 260 223 294
rect 359 306 393 340
rect 527 310 561 344
rect 641 242 675 276
rect 983 276 1017 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 23 581 381 615
rect 23 556 89 581
rect 23 522 39 556
rect 73 522 89 556
rect 315 580 381 581
rect 23 488 89 522
rect 23 454 39 488
rect 73 454 89 488
rect 23 415 89 454
rect 23 381 39 415
rect 73 381 89 415
rect 23 365 89 381
rect 124 529 168 545
rect 124 495 129 529
rect 163 495 168 529
rect 124 428 168 495
rect 203 521 269 547
rect 315 546 331 580
rect 365 546 381 580
rect 315 530 381 546
rect 415 580 481 649
rect 415 546 431 580
rect 465 546 481 580
rect 415 530 481 546
rect 515 580 565 596
rect 515 546 531 580
rect 203 487 219 521
rect 253 496 269 521
rect 515 512 565 546
rect 774 580 842 649
rect 774 546 791 580
rect 825 546 842 580
rect 774 530 842 546
rect 956 580 1033 649
rect 956 546 977 580
rect 1011 546 1033 580
rect 956 530 1033 546
rect 515 496 531 512
rect 253 487 531 496
rect 203 478 531 487
rect 203 462 565 478
rect 599 462 1033 496
rect 599 428 633 462
rect 124 421 633 428
rect 124 387 129 421
rect 163 394 633 421
rect 667 421 759 428
rect 163 387 307 394
rect 124 364 307 387
rect 21 294 87 310
rect 21 260 37 294
rect 71 260 87 294
rect 21 236 87 260
rect 121 294 239 310
rect 121 260 189 294
rect 223 260 239 294
rect 121 236 239 260
rect 273 202 307 364
rect 667 387 683 421
rect 717 387 759 421
rect 667 360 759 387
rect 343 340 477 356
rect 343 306 359 340
rect 393 306 477 340
rect 343 290 477 306
rect 511 344 759 360
rect 511 310 527 344
rect 561 326 759 344
rect 561 310 577 326
rect 511 294 577 310
rect 443 260 477 290
rect 625 276 691 292
rect 625 260 641 276
rect 443 242 641 260
rect 675 242 691 276
rect 443 226 691 242
rect 34 196 100 202
rect 34 162 50 196
rect 84 162 100 196
rect 34 120 100 162
rect 134 186 307 202
rect 134 152 167 186
rect 201 152 307 186
rect 343 209 409 226
rect 343 175 359 209
rect 393 192 409 209
rect 393 175 634 192
rect 725 188 759 326
rect 343 158 634 175
rect 134 136 307 152
rect 34 86 50 120
rect 84 92 100 120
rect 484 116 550 124
rect 484 92 500 116
rect 84 86 500 92
rect 34 82 500 86
rect 534 82 550 116
rect 34 58 550 82
rect 600 17 634 158
rect 668 154 759 188
rect 793 421 933 428
rect 793 387 882 421
rect 916 387 933 421
rect 793 207 933 387
rect 967 310 1033 462
rect 967 276 983 310
rect 1017 276 1033 310
rect 967 260 1033 276
rect 793 173 883 207
rect 917 173 933 207
rect 793 154 933 173
rect 967 210 1033 226
rect 967 176 983 210
rect 1017 176 1033 210
rect 668 146 734 154
rect 668 112 684 146
rect 718 112 734 146
rect 967 120 1033 176
rect 668 70 734 112
rect 768 86 790 120
rect 824 86 846 120
rect 768 17 846 86
rect 967 86 983 120
rect 1017 86 1033 120
rect 967 17 1033 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 683 1056 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 0 617 1056 649
rect 0 17 1056 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -49 1056 -17
<< labels >>
rlabel comment s 0 0 0 0 4 mux2_2
flabel pwell s 0 0 1056 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 1056 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 1056 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 1056 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 S
port 3 nsew
flabel corelocali s 127 242 161 276 0 FreeSans 340 0 0 0 A1
port 2 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 A0
port 1 nsew
flabel corelocali s 799 168 833 202 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 799 242 833 276 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 X
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 1056 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2455354
string GDS_START 2447354
<< end >>
