magic
tech sky130A
magscale 1 2
timestamp 1601050082
<< locali >>
rect 183 275 263 356
rect 788 270 854 356
rect 1356 270 1422 356
rect 1656 368 1728 596
rect 1694 325 1728 368
rect 1836 325 1907 596
rect 1694 284 1907 325
rect 1694 234 1735 284
rect 1669 94 1735 234
rect 1841 88 1907 284
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 17 369 73 577
rect 113 458 179 649
rect 213 581 736 615
rect 213 424 279 581
rect 107 390 279 424
rect 313 513 545 547
rect 670 542 736 581
rect 878 546 944 649
rect 1097 581 1463 615
rect 1097 546 1163 581
rect 17 173 57 369
rect 107 293 141 390
rect 91 241 141 293
rect 313 275 353 513
rect 461 458 545 513
rect 1204 512 1254 547
rect 579 508 629 509
rect 888 508 1254 512
rect 579 478 1254 508
rect 579 474 922 478
rect 387 424 427 431
rect 387 335 449 424
rect 579 375 629 474
rect 720 390 854 440
rect 720 341 754 390
rect 387 301 551 335
rect 319 267 353 275
rect 91 207 285 241
rect 319 233 477 267
rect 17 73 99 173
rect 133 17 199 173
rect 235 85 285 207
rect 325 153 391 199
rect 427 187 477 233
rect 511 241 551 301
rect 599 275 754 341
rect 511 191 604 241
rect 720 225 754 275
rect 720 191 818 225
rect 888 206 922 474
rect 956 390 1056 444
rect 1204 394 1254 478
rect 1288 398 1392 500
rect 1426 424 1463 581
rect 1497 458 1622 649
rect 956 276 990 390
rect 1024 344 1090 356
rect 1288 344 1322 398
rect 1426 390 1498 424
rect 1024 310 1322 344
rect 956 242 1232 276
rect 1081 236 1232 242
rect 888 157 1032 206
rect 511 153 1032 157
rect 325 123 1032 153
rect 325 119 545 123
rect 640 85 706 89
rect 235 51 706 85
rect 854 17 920 89
rect 966 70 1032 123
rect 1066 85 1132 202
rect 1166 119 1232 236
rect 1278 234 1322 310
rect 1464 334 1498 390
rect 1537 368 1622 458
rect 1464 268 1660 334
rect 1762 364 1796 649
rect 1942 364 1992 649
rect 1464 236 1498 268
rect 1278 200 1344 234
rect 1378 202 1498 236
rect 1378 166 1412 202
rect 1583 168 1633 234
rect 1266 132 1412 166
rect 1266 85 1300 132
rect 1446 98 1633 168
rect 1066 51 1300 85
rect 1380 17 1633 98
rect 1771 17 1805 250
rect 1943 17 1993 250
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< obsm1 >>
rect 19 421 77 430
rect 307 421 365 430
rect 19 393 365 421
rect 19 384 77 393
rect 307 384 365 393
rect 403 421 461 430
rect 979 421 1037 430
rect 403 393 1037 421
rect 403 384 461 393
rect 979 384 1037 393
<< labels >>
rlabel locali s 183 275 263 356 6 A
port 1 nsew signal input
rlabel locali s 788 270 854 356 6 B
port 2 nsew signal input
rlabel locali s 1356 270 1422 356 6 C
port 3 nsew signal input
rlabel locali s 1841 88 1907 284 6 X
port 4 nsew signal output
rlabel locali s 1836 325 1907 596 6 X
port 4 nsew signal output
rlabel locali s 1694 325 1728 368 6 X
port 4 nsew signal output
rlabel locali s 1694 284 1907 325 6 X
port 4 nsew signal output
rlabel locali s 1694 234 1735 284 6 X
port 4 nsew signal output
rlabel locali s 1669 94 1735 234 6 X
port 4 nsew signal output
rlabel locali s 1656 368 1728 596 6 X
port 4 nsew signal output
rlabel metal1 s 0 -49 2016 49 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 617 2016 715 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2016 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 644484
string GDS_START 628746
<< end >>
