magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 217 294 331 360
rect 481 355 551 430
rect 653 270 737 356
rect 85 180 415 246
rect 313 162 415 180
rect 2118 394 2168 596
rect 2118 360 2190 394
rect 2156 226 2190 360
rect 2511 430 2567 596
rect 2511 364 2663 430
rect 2124 70 2190 226
rect 2615 230 2663 364
rect 2510 180 2663 230
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2688 683
rect 17 360 104 585
rect 145 462 211 649
rect 330 508 396 585
rect 534 542 618 649
rect 815 542 881 649
rect 1315 591 1381 649
rect 1017 533 1067 587
rect 915 508 1067 533
rect 330 499 1067 508
rect 330 474 949 499
rect 1101 495 1173 587
rect 1207 523 1547 557
rect 330 462 396 474
rect 149 394 439 428
rect 149 360 183 394
rect 17 294 183 360
rect 373 345 439 394
rect 585 304 619 474
rect 659 390 819 440
rect 17 146 51 294
rect 449 270 619 304
rect 771 270 819 390
rect 853 330 887 474
rect 1001 440 1067 465
rect 921 401 1067 440
rect 921 364 971 401
rect 853 296 980 330
rect 17 70 98 146
rect 132 17 198 146
rect 449 128 483 270
rect 771 236 805 270
rect 296 78 483 128
rect 539 17 589 226
rect 625 202 805 236
rect 625 70 691 202
rect 737 17 803 168
rect 839 85 889 226
rect 930 119 980 296
rect 1014 85 1048 401
rect 1101 349 1135 495
rect 1207 449 1241 523
rect 1169 383 1241 449
rect 1422 423 1479 489
rect 1346 349 1402 389
rect 1082 315 1402 349
rect 1082 175 1116 315
rect 1436 281 1470 423
rect 1513 386 1547 523
rect 1581 420 1647 596
rect 1772 530 1886 649
rect 1920 476 1990 596
rect 1513 320 1579 386
rect 1613 378 1647 420
rect 1742 412 1990 476
rect 1920 388 1990 412
rect 1613 344 1804 378
rect 1150 209 1216 275
rect 1250 222 1470 281
rect 1670 279 1736 310
rect 1182 188 1216 209
rect 1082 119 1148 175
rect 1182 154 1402 188
rect 1182 85 1216 154
rect 839 51 1216 85
rect 1268 17 1334 120
rect 1368 85 1402 154
rect 1436 119 1470 222
rect 1504 245 1736 279
rect 1770 245 1804 344
rect 1956 326 1990 388
rect 2028 364 2078 649
rect 2208 428 2274 649
rect 2224 364 2274 428
rect 1856 245 1922 310
rect 1504 206 1556 245
rect 1770 211 1922 245
rect 1956 260 2122 326
rect 1504 85 1538 206
rect 1604 177 1804 211
rect 1956 177 1990 260
rect 2316 330 2382 572
rect 2421 364 2471 649
rect 2601 464 2667 649
rect 2316 264 2547 330
rect 1604 162 1638 177
rect 1368 51 1538 85
rect 1572 70 1638 162
rect 1736 17 1878 143
rect 1912 70 1990 177
rect 2024 17 2090 226
rect 2226 17 2276 226
rect 2316 112 2388 264
rect 2424 146 2476 230
rect 2424 17 2490 146
rect 2599 17 2665 146
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2688 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
<< metal1 >>
rect 0 683 2688 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2688 683
rect 0 617 2688 649
rect 0 17 2688 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2688 17
rect 0 -49 2688 -17
<< labels >>
rlabel locali s 217 294 331 360 6 D
port 1 nsew signal input
rlabel locali s 2156 226 2190 360 6 Q
port 2 nsew signal output
rlabel locali s 2124 70 2190 226 6 Q
port 2 nsew signal output
rlabel locali s 2118 394 2168 596 6 Q
port 2 nsew signal output
rlabel locali s 2118 360 2190 394 6 Q
port 2 nsew signal output
rlabel locali s 2615 230 2663 364 6 Q_N
port 3 nsew signal output
rlabel locali s 2511 430 2567 596 6 Q_N
port 3 nsew signal output
rlabel locali s 2511 364 2663 430 6 Q_N
port 3 nsew signal output
rlabel locali s 2510 180 2663 230 6 Q_N
port 3 nsew signal output
rlabel locali s 481 355 551 430 6 SCD
port 4 nsew signal input
rlabel locali s 313 162 415 180 6 SCE
port 5 nsew signal input
rlabel locali s 85 180 415 246 6 SCE
port 5 nsew signal input
rlabel locali s 653 270 737 356 6 CLK
port 6 nsew clock input
rlabel metal1 s 0 -49 2688 49 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 617 2688 715 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2688 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 277842
string GDS_START 258190
<< end >>
