magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 1050 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 83 47 113 177
rect 187 47 217 177
rect 271 47 301 177
rect 375 47 405 177
rect 571 47 601 177
rect 675 47 705 177
rect 759 47 789 177
rect 863 47 893 177
<< pmoshvt >>
rect 85 297 121 497
rect 179 297 215 497
rect 273 297 309 497
rect 367 297 403 497
rect 573 297 609 497
rect 667 297 703 497
rect 761 297 797 497
rect 855 297 891 497
<< ndiff >>
rect 27 163 83 177
rect 27 129 39 163
rect 73 129 83 163
rect 27 95 83 129
rect 27 61 39 95
rect 73 61 83 95
rect 27 47 83 61
rect 113 163 187 177
rect 113 129 133 163
rect 167 129 187 163
rect 113 95 187 129
rect 113 61 133 95
rect 167 61 187 95
rect 113 47 187 61
rect 217 95 271 177
rect 217 61 227 95
rect 261 61 271 95
rect 217 47 271 61
rect 301 163 375 177
rect 301 129 321 163
rect 355 129 375 163
rect 301 95 375 129
rect 301 61 321 95
rect 355 61 375 95
rect 301 47 375 61
rect 405 95 461 177
rect 405 61 415 95
rect 449 61 461 95
rect 405 47 461 61
rect 515 95 571 177
rect 515 61 527 95
rect 561 61 571 95
rect 515 47 571 61
rect 601 163 675 177
rect 601 129 621 163
rect 655 129 675 163
rect 601 95 675 129
rect 601 61 621 95
rect 655 61 675 95
rect 601 47 675 61
rect 705 95 759 177
rect 705 61 715 95
rect 749 61 759 95
rect 705 47 759 61
rect 789 163 863 177
rect 789 129 809 163
rect 843 129 863 163
rect 789 95 863 129
rect 789 61 809 95
rect 843 61 863 95
rect 789 47 863 61
rect 893 95 945 177
rect 893 61 903 95
rect 937 61 945 95
rect 893 47 945 61
<< pdiff >>
rect 27 477 85 497
rect 27 443 39 477
rect 73 443 85 477
rect 27 409 85 443
rect 27 375 39 409
rect 73 375 85 409
rect 27 341 85 375
rect 27 307 39 341
rect 73 307 85 341
rect 27 297 85 307
rect 121 477 179 497
rect 121 443 133 477
rect 167 443 179 477
rect 121 409 179 443
rect 121 375 133 409
rect 167 375 179 409
rect 121 297 179 375
rect 215 477 273 497
rect 215 443 227 477
rect 261 443 273 477
rect 215 409 273 443
rect 215 375 227 409
rect 261 375 273 409
rect 215 341 273 375
rect 215 307 227 341
rect 261 307 273 341
rect 215 297 273 307
rect 309 477 367 497
rect 309 443 321 477
rect 355 443 367 477
rect 309 409 367 443
rect 309 375 321 409
rect 355 375 367 409
rect 309 297 367 375
rect 403 409 461 497
rect 403 375 415 409
rect 449 375 461 409
rect 403 341 461 375
rect 403 307 415 341
rect 449 307 461 341
rect 403 297 461 307
rect 515 409 573 497
rect 515 375 527 409
rect 561 375 573 409
rect 515 341 573 375
rect 515 307 527 341
rect 561 307 573 341
rect 515 297 573 307
rect 609 477 667 497
rect 609 443 621 477
rect 655 443 667 477
rect 609 409 667 443
rect 609 375 621 409
rect 655 375 667 409
rect 609 297 667 375
rect 703 477 761 497
rect 703 443 715 477
rect 749 443 761 477
rect 703 409 761 443
rect 703 375 715 409
rect 749 375 761 409
rect 703 341 761 375
rect 703 307 715 341
rect 749 307 761 341
rect 703 297 761 307
rect 797 409 855 497
rect 797 375 809 409
rect 843 375 855 409
rect 797 341 855 375
rect 797 307 809 341
rect 843 307 855 341
rect 797 297 855 307
rect 891 477 945 497
rect 891 443 903 477
rect 937 443 945 477
rect 891 409 945 443
rect 891 375 903 409
rect 937 375 945 409
rect 891 297 945 375
<< ndiffc >>
rect 39 129 73 163
rect 39 61 73 95
rect 133 129 167 163
rect 133 61 167 95
rect 227 61 261 95
rect 321 129 355 163
rect 321 61 355 95
rect 415 61 449 95
rect 527 61 561 95
rect 621 129 655 163
rect 621 61 655 95
rect 715 61 749 95
rect 809 129 843 163
rect 809 61 843 95
rect 903 61 937 95
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 133 443 167 477
rect 133 375 167 409
rect 227 443 261 477
rect 227 375 261 409
rect 227 307 261 341
rect 321 443 355 477
rect 321 375 355 409
rect 415 375 449 409
rect 415 307 449 341
rect 527 375 561 409
rect 527 307 561 341
rect 621 443 655 477
rect 621 375 655 409
rect 715 443 749 477
rect 715 375 749 409
rect 715 307 749 341
rect 809 375 843 409
rect 809 307 843 341
rect 903 443 937 477
rect 903 375 937 409
<< poly >>
rect 85 497 121 523
rect 179 497 215 523
rect 273 497 309 523
rect 367 497 403 523
rect 573 497 609 523
rect 667 497 703 523
rect 761 497 797 523
rect 855 497 891 523
rect 85 282 121 297
rect 179 282 215 297
rect 273 282 309 297
rect 367 282 403 297
rect 573 282 609 297
rect 667 282 703 297
rect 761 282 797 297
rect 855 282 891 297
rect 83 265 123 282
rect 177 265 217 282
rect 83 249 217 265
rect 83 215 112 249
rect 146 215 217 249
rect 83 199 217 215
rect 83 177 113 199
rect 187 177 217 199
rect 271 265 311 282
rect 365 265 405 282
rect 271 249 405 265
rect 271 215 318 249
rect 352 215 405 249
rect 271 199 405 215
rect 271 177 301 199
rect 375 177 405 199
rect 571 265 611 282
rect 665 265 705 282
rect 571 249 705 265
rect 571 215 621 249
rect 655 215 705 249
rect 571 199 705 215
rect 571 177 601 199
rect 675 177 705 199
rect 759 265 799 282
rect 853 265 893 282
rect 759 249 893 265
rect 759 215 805 249
rect 839 215 893 249
rect 759 199 893 215
rect 759 177 789 199
rect 863 177 893 199
rect 83 21 113 47
rect 187 21 217 47
rect 271 21 301 47
rect 375 21 405 47
rect 571 21 601 47
rect 675 21 705 47
rect 759 21 789 47
rect 863 21 893 47
<< polycont >>
rect 112 215 146 249
rect 318 215 352 249
rect 621 215 655 249
rect 805 215 839 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 30 477 81 493
rect 30 443 39 477
rect 73 443 81 477
rect 30 409 81 443
rect 30 375 39 409
rect 73 375 81 409
rect 30 341 81 375
rect 125 477 175 527
rect 125 443 133 477
rect 167 443 175 477
rect 125 409 175 443
rect 125 375 133 409
rect 167 375 175 409
rect 125 359 175 375
rect 219 477 269 493
rect 219 443 227 477
rect 261 443 269 477
rect 219 409 269 443
rect 219 375 227 409
rect 261 375 269 409
rect 30 307 39 341
rect 73 325 81 341
rect 219 341 269 375
rect 313 477 663 493
rect 313 443 321 477
rect 355 459 621 477
rect 355 443 363 459
rect 313 409 363 443
rect 613 443 621 459
rect 655 443 663 477
rect 313 375 321 409
rect 355 375 363 409
rect 313 359 363 375
rect 407 409 457 425
rect 407 375 415 409
rect 449 375 457 409
rect 219 325 227 341
rect 73 307 227 325
rect 261 325 269 341
rect 407 341 457 375
rect 407 325 415 341
rect 261 307 415 325
rect 449 307 457 341
rect 30 291 457 307
rect 519 409 569 425
rect 519 375 527 409
rect 561 375 569 409
rect 519 341 569 375
rect 613 409 663 443
rect 613 375 621 409
rect 655 375 663 409
rect 613 359 663 375
rect 707 477 945 493
rect 707 443 715 477
rect 749 459 903 477
rect 749 443 757 459
rect 707 409 757 443
rect 895 443 903 459
rect 937 443 945 477
rect 707 375 715 409
rect 749 375 757 409
rect 519 307 527 341
rect 561 325 569 341
rect 707 341 757 375
rect 707 325 715 341
rect 561 307 715 325
rect 749 307 757 341
rect 519 291 757 307
rect 808 409 858 425
rect 808 375 809 409
rect 843 375 858 409
rect 808 341 858 375
rect 895 409 945 443
rect 895 375 903 409
rect 937 375 945 409
rect 895 359 945 375
rect 808 307 809 341
rect 843 325 858 341
rect 843 307 990 325
rect 808 291 990 307
rect 40 249 203 257
rect 40 215 112 249
rect 146 215 203 249
rect 247 249 428 257
rect 247 215 318 249
rect 352 215 428 249
rect 482 249 671 257
rect 482 215 621 249
rect 655 215 671 249
rect 728 249 855 257
rect 728 215 805 249
rect 839 215 855 249
rect 923 181 990 291
rect 18 163 73 181
rect 18 129 39 163
rect 18 95 73 129
rect 18 61 39 95
rect 18 17 73 61
rect 114 163 990 181
rect 114 129 133 163
rect 167 145 321 163
rect 167 129 190 145
rect 114 95 190 129
rect 302 129 321 145
rect 355 145 621 163
rect 355 129 378 145
rect 114 61 133 95
rect 167 61 190 95
rect 114 51 190 61
rect 227 95 261 111
rect 227 17 261 61
rect 302 95 378 129
rect 602 129 621 145
rect 655 145 809 163
rect 655 129 678 145
rect 302 61 321 95
rect 355 61 378 95
rect 302 51 378 61
rect 415 95 561 111
rect 449 61 527 95
rect 415 17 561 61
rect 602 95 678 129
rect 790 129 809 145
rect 843 145 990 163
rect 843 129 866 145
rect 602 61 621 95
rect 655 61 678 95
rect 602 51 678 61
rect 715 95 749 111
rect 715 17 749 61
rect 790 95 866 129
rect 790 61 809 95
rect 843 61 866 95
rect 790 51 866 61
rect 903 95 961 111
rect 937 61 961 95
rect 903 17 961 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
flabel corelocali s 534 221 568 255 0 FreeSans 400 0 0 0 C
port 3 nsew
flabel corelocali s 738 221 772 255 0 FreeSans 400 0 0 0 D
port 4 nsew
flabel corelocali s 942 153 976 187 0 FreeSans 400 0 0 0 Y
port 9 nsew
flabel corelocali s 132 221 166 255 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 323 238 323 238 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
rlabel comment s 0 0 0 0 4 nor4_2
<< properties >>
string FIXED_BBOX 0 0 1012 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2487712
string GDS_START 2479646
<< end >>
