magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 736 561
rect 17 299 94 491
rect 137 367 195 527
rect 17 165 52 299
rect 297 265 362 425
rect 201 215 251 265
rect 201 199 235 215
rect 293 199 362 265
rect 396 199 451 332
rect 488 199 559 332
rect 661 299 719 527
rect 664 199 719 265
rect 17 51 119 165
rect 153 17 187 129
rect 329 17 395 97
rect 0 -17 736 17
<< obsli1 >>
rect 229 459 502 493
rect 229 333 263 459
rect 128 299 263 333
rect 128 265 162 299
rect 436 417 502 459
rect 436 367 627 417
rect 89 215 162 265
rect 89 199 127 215
rect 593 165 627 367
rect 228 131 508 165
rect 228 51 294 131
rect 442 93 508 131
rect 542 127 627 165
rect 661 93 719 147
rect 442 51 719 93
<< metal1 >>
rect 0 496 736 592
rect 0 -48 736 48
<< labels >>
rlabel locali s 201 215 251 265 6 A1
port 1 nsew signal input
rlabel locali s 201 199 235 215 6 A1
port 1 nsew signal input
rlabel locali s 297 265 362 425 6 A2
port 2 nsew signal input
rlabel locali s 293 199 362 265 6 A2
port 2 nsew signal input
rlabel locali s 396 199 451 332 6 A3
port 3 nsew signal input
rlabel locali s 664 199 719 265 6 B1
port 4 nsew signal input
rlabel locali s 488 199 559 332 6 B2
port 5 nsew signal input
rlabel locali s 17 299 94 491 6 X
port 6 nsew signal output
rlabel locali s 17 165 52 299 6 X
port 6 nsew signal output
rlabel locali s 17 51 119 165 6 X
port 6 nsew signal output
rlabel locali s 329 17 395 97 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 153 17 187 129 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 736 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 736 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 661 299 719 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 137 367 195 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 736 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 736 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 939794
string GDS_START 932750
<< end >>
