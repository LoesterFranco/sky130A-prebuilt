magic
tech sky130A
magscale 1 2
timestamp 1599588209
<< nwell >>
rect -38 332 3302 704
rect 1240 328 1461 332
<< pwell >>
rect 0 0 3264 49
<< scpmos >>
rect 99 464 129 592
rect 183 464 213 592
rect 409 463 439 591
rect 545 463 575 591
rect 623 463 653 591
rect 713 463 743 591
rect 913 455 943 583
rect 1049 455 1079 583
rect 1133 455 1163 583
rect 1336 364 1366 588
rect 1614 368 1644 592
rect 1816 508 1846 592
rect 1906 508 1936 592
rect 2016 508 2046 592
rect 2123 398 2153 566
rect 2327 392 2357 592
rect 2519 392 2549 592
rect 2627 508 2657 592
rect 2711 508 2741 592
rect 2853 464 2883 592
rect 3055 368 3085 592
rect 3148 368 3178 592
<< nmoslvt >>
rect 108 74 138 158
rect 186 74 216 158
rect 384 113 414 197
rect 470 113 500 197
rect 548 113 578 197
rect 663 113 693 197
rect 938 125 968 209
rect 1038 125 1068 209
rect 1110 125 1140 209
rect 1310 74 1340 222
rect 1508 74 1538 222
rect 1706 97 1736 181
rect 1842 97 1872 181
rect 1979 97 2009 181
rect 2134 74 2164 202
rect 2372 74 2402 202
rect 2444 74 2474 202
rect 2539 74 2569 158
rect 2617 74 2647 158
rect 2838 74 2868 158
rect 3050 74 3080 222
rect 3136 74 3166 222
<< ndiff >>
rect 327 172 384 197
rect 51 133 108 158
rect 51 99 63 133
rect 97 99 108 133
rect 51 74 108 99
rect 138 74 186 158
rect 216 133 273 158
rect 216 99 227 133
rect 261 99 273 133
rect 327 138 339 172
rect 373 138 384 172
rect 327 113 384 138
rect 414 172 470 197
rect 414 138 425 172
rect 459 138 470 172
rect 414 113 470 138
rect 500 113 548 197
rect 578 185 663 197
rect 578 151 603 185
rect 637 151 663 185
rect 578 113 663 151
rect 693 172 764 197
rect 693 138 718 172
rect 752 138 764 172
rect 693 113 764 138
rect 216 74 273 99
rect 881 178 938 209
rect 881 144 893 178
rect 927 144 938 178
rect 881 125 938 144
rect 968 178 1038 209
rect 968 144 993 178
rect 1027 144 1038 178
rect 968 125 1038 144
rect 1068 125 1110 209
rect 1140 184 1197 209
rect 1140 150 1151 184
rect 1185 150 1197 184
rect 1140 125 1197 150
rect 1251 120 1310 222
rect 1251 86 1264 120
rect 1298 86 1310 120
rect 1251 74 1310 86
rect 1340 202 1397 222
rect 1340 168 1351 202
rect 1385 168 1397 202
rect 1340 120 1397 168
rect 1340 86 1351 120
rect 1385 86 1397 120
rect 1340 74 1397 86
rect 1451 210 1508 222
rect 1451 176 1463 210
rect 1497 176 1508 210
rect 1451 120 1508 176
rect 1451 86 1463 120
rect 1497 86 1508 120
rect 1451 74 1508 86
rect 1538 210 1595 222
rect 1538 176 1549 210
rect 1583 176 1595 210
rect 2084 181 2134 202
rect 1538 120 1595 176
rect 1538 86 1549 120
rect 1583 86 1595 120
rect 1649 169 1706 181
rect 1649 135 1661 169
rect 1695 135 1706 169
rect 1649 97 1706 135
rect 1736 169 1842 181
rect 1736 135 1797 169
rect 1831 135 1842 169
rect 1736 97 1842 135
rect 1872 97 1979 181
rect 2009 120 2134 181
rect 2009 97 2037 120
rect 1538 74 1595 86
rect 2024 86 2037 97
rect 2071 86 2134 120
rect 2024 74 2134 86
rect 2164 179 2221 202
rect 2164 145 2175 179
rect 2209 145 2221 179
rect 2164 74 2221 145
rect 2315 120 2372 202
rect 2315 86 2327 120
rect 2361 86 2372 120
rect 2315 74 2372 86
rect 2402 74 2444 202
rect 2474 158 2524 202
rect 2979 190 3050 222
rect 2474 133 2539 158
rect 2474 99 2494 133
rect 2528 99 2539 133
rect 2474 74 2539 99
rect 2569 74 2617 158
rect 2647 120 2838 158
rect 2647 86 2658 120
rect 2692 86 2779 120
rect 2813 86 2838 120
rect 2647 74 2838 86
rect 2868 133 2925 158
rect 2868 99 2879 133
rect 2913 99 2925 133
rect 2868 74 2925 99
rect 2979 156 2991 190
rect 3025 156 3050 190
rect 2979 120 3050 156
rect 2979 86 2991 120
rect 3025 86 3050 120
rect 2979 74 3050 86
rect 3080 210 3136 222
rect 3080 176 3091 210
rect 3125 176 3136 210
rect 3080 120 3136 176
rect 3080 86 3091 120
rect 3125 86 3136 120
rect 3080 74 3136 86
rect 3166 210 3237 222
rect 3166 176 3191 210
rect 3225 176 3237 210
rect 3166 120 3237 176
rect 3166 86 3191 120
rect 3225 86 3237 120
rect 3166 74 3237 86
<< pdiff >>
rect 40 580 99 592
rect 40 546 52 580
rect 86 546 99 580
rect 40 510 99 546
rect 40 476 52 510
rect 86 476 99 510
rect 40 464 99 476
rect 129 464 183 592
rect 213 578 272 592
rect 213 544 226 578
rect 260 544 272 578
rect 213 464 272 544
rect 350 520 409 591
rect 350 486 362 520
rect 396 486 409 520
rect 350 463 409 486
rect 439 577 545 591
rect 439 543 498 577
rect 532 543 545 577
rect 439 463 545 543
rect 575 463 623 591
rect 653 579 713 591
rect 653 545 666 579
rect 700 545 713 579
rect 653 509 713 545
rect 653 475 666 509
rect 700 475 713 509
rect 653 463 713 475
rect 743 579 801 591
rect 743 545 756 579
rect 790 545 801 579
rect 743 509 801 545
rect 743 475 756 509
rect 790 475 801 509
rect 743 463 801 475
rect 855 516 913 583
rect 855 482 866 516
rect 900 482 913 516
rect 855 455 913 482
rect 943 570 1049 583
rect 943 536 1002 570
rect 1036 536 1049 570
rect 943 455 1049 536
rect 1079 455 1133 583
rect 1163 571 1222 583
rect 1163 537 1176 571
rect 1210 537 1222 571
rect 1163 501 1222 537
rect 1163 467 1176 501
rect 1210 467 1222 501
rect 1163 455 1222 467
rect 1276 576 1336 588
rect 1276 542 1288 576
rect 1322 542 1336 576
rect 1276 364 1336 542
rect 1366 417 1425 588
rect 1555 578 1614 592
rect 1555 544 1567 578
rect 1601 544 1614 578
rect 1366 383 1379 417
rect 1413 383 1425 417
rect 1366 364 1425 383
rect 1555 368 1614 544
rect 1644 419 1703 592
rect 1757 567 1816 592
rect 1757 533 1769 567
rect 1803 533 1816 567
rect 1757 508 1816 533
rect 1846 567 1906 592
rect 1846 533 1859 567
rect 1893 533 1906 567
rect 1846 508 1906 533
rect 1936 508 2016 592
rect 2046 580 2105 592
rect 2046 546 2059 580
rect 2093 566 2105 580
rect 2266 580 2327 592
rect 2093 546 2123 566
rect 2046 508 2123 546
rect 1644 385 1657 419
rect 1691 385 1703 419
rect 1644 368 1703 385
rect 2070 398 2123 508
rect 2153 444 2212 566
rect 2153 410 2166 444
rect 2200 410 2212 444
rect 2153 398 2212 410
rect 2266 546 2279 580
rect 2313 546 2327 580
rect 2266 392 2327 546
rect 2357 392 2519 592
rect 2549 567 2627 592
rect 2549 533 2580 567
rect 2614 533 2627 567
rect 2549 508 2627 533
rect 2657 508 2711 592
rect 2741 580 2853 592
rect 2741 546 2775 580
rect 2809 546 2853 580
rect 2741 508 2853 546
rect 2549 392 2602 508
rect 2800 464 2853 508
rect 2883 580 2942 592
rect 2883 546 2896 580
rect 2930 546 2942 580
rect 2883 510 2942 546
rect 2883 476 2896 510
rect 2930 476 2942 510
rect 2883 464 2942 476
rect 2996 580 3055 592
rect 2996 546 3008 580
rect 3042 546 3055 580
rect 2996 501 3055 546
rect 2996 467 3008 501
rect 3042 467 3055 501
rect 2996 424 3055 467
rect 2996 390 3008 424
rect 3042 390 3055 424
rect 2996 368 3055 390
rect 3085 580 3148 592
rect 3085 546 3099 580
rect 3133 546 3148 580
rect 3085 499 3148 546
rect 3085 465 3099 499
rect 3133 465 3148 499
rect 3085 414 3148 465
rect 3085 380 3099 414
rect 3133 380 3148 414
rect 3085 368 3148 380
rect 3178 580 3237 592
rect 3178 546 3191 580
rect 3225 546 3237 580
rect 3178 498 3237 546
rect 3178 464 3191 498
rect 3225 464 3237 498
rect 3178 368 3237 464
<< ndiffc >>
rect 63 99 97 133
rect 227 99 261 133
rect 339 138 373 172
rect 425 138 459 172
rect 603 151 637 185
rect 718 138 752 172
rect 893 144 927 178
rect 993 144 1027 178
rect 1151 150 1185 184
rect 1264 86 1298 120
rect 1351 168 1385 202
rect 1351 86 1385 120
rect 1463 176 1497 210
rect 1463 86 1497 120
rect 1549 176 1583 210
rect 1549 86 1583 120
rect 1661 135 1695 169
rect 1797 135 1831 169
rect 2037 86 2071 120
rect 2175 145 2209 179
rect 2327 86 2361 120
rect 2494 99 2528 133
rect 2658 86 2692 120
rect 2779 86 2813 120
rect 2879 99 2913 133
rect 2991 156 3025 190
rect 2991 86 3025 120
rect 3091 176 3125 210
rect 3091 86 3125 120
rect 3191 176 3225 210
rect 3191 86 3225 120
<< pdiffc >>
rect 52 546 86 580
rect 52 476 86 510
rect 226 544 260 578
rect 362 486 396 520
rect 498 543 532 577
rect 666 545 700 579
rect 666 475 700 509
rect 756 545 790 579
rect 756 475 790 509
rect 866 482 900 516
rect 1002 536 1036 570
rect 1176 537 1210 571
rect 1176 467 1210 501
rect 1288 542 1322 576
rect 1567 544 1601 578
rect 1379 383 1413 417
rect 1769 533 1803 567
rect 1859 533 1893 567
rect 2059 546 2093 580
rect 1657 385 1691 419
rect 2166 410 2200 444
rect 2279 546 2313 580
rect 2580 533 2614 567
rect 2775 546 2809 580
rect 2896 546 2930 580
rect 2896 476 2930 510
rect 3008 546 3042 580
rect 3008 467 3042 501
rect 3008 390 3042 424
rect 3099 546 3133 580
rect 3099 465 3133 499
rect 3099 380 3133 414
rect 3191 546 3225 580
rect 3191 464 3225 498
<< poly >>
rect 99 592 129 618
rect 183 592 213 618
rect 409 591 439 617
rect 545 591 575 617
rect 623 591 653 617
rect 710 606 946 636
rect 713 591 743 606
rect 910 598 946 606
rect 99 449 129 464
rect 183 449 213 464
rect 913 583 943 598
rect 1049 583 1079 609
rect 1133 583 1163 609
rect 1336 588 1366 614
rect 1614 592 1644 618
rect 1816 592 1846 618
rect 1906 592 1936 618
rect 2016 592 2046 618
rect 2327 592 2357 618
rect 2519 592 2549 618
rect 2627 592 2657 618
rect 2711 592 2741 618
rect 2853 592 2883 618
rect 3055 592 3085 618
rect 3148 592 3178 618
rect 96 398 132 449
rect 180 424 216 449
rect 409 448 439 463
rect 545 448 575 463
rect 623 448 653 463
rect 180 408 261 424
rect 72 382 138 398
rect 72 348 88 382
rect 122 348 138 382
rect 72 314 138 348
rect 72 280 88 314
rect 122 280 138 314
rect 180 374 211 408
rect 245 374 261 408
rect 180 340 261 374
rect 180 306 211 340
rect 245 306 261 340
rect 333 418 578 448
rect 333 330 363 418
rect 411 354 500 370
rect 620 369 656 448
rect 713 437 743 463
rect 913 440 943 455
rect 1049 440 1079 455
rect 1133 440 1163 455
rect 180 290 261 306
rect 303 314 369 330
rect 72 246 138 280
rect 72 212 88 246
rect 122 212 138 246
rect 303 280 319 314
rect 353 280 369 314
rect 411 320 427 354
rect 461 320 500 354
rect 411 304 500 320
rect 303 242 369 280
rect 72 196 138 212
rect 108 158 138 196
rect 186 212 414 242
rect 186 158 216 212
rect 384 197 414 212
rect 470 197 500 304
rect 548 353 656 369
rect 548 319 564 353
rect 598 319 656 353
rect 548 303 656 319
rect 793 373 859 389
rect 793 339 809 373
rect 843 339 859 373
rect 793 305 859 339
rect 548 197 578 303
rect 793 271 809 305
rect 843 271 859 305
rect 910 302 946 440
rect 1046 349 1082 440
rect 1130 417 1166 440
rect 1016 333 1082 349
rect 793 242 859 271
rect 663 237 859 242
rect 663 212 809 237
rect 663 197 693 212
rect 793 203 809 212
rect 843 203 859 237
rect 901 286 968 302
rect 901 252 917 286
rect 951 252 968 286
rect 1016 299 1032 333
rect 1066 299 1082 333
rect 1016 283 1082 299
rect 1124 401 1190 417
rect 1124 367 1140 401
rect 1174 367 1190 401
rect 1124 333 1190 367
rect 1457 424 1538 440
rect 1457 390 1473 424
rect 1507 390 1538 424
rect 1336 349 1366 364
rect 1457 356 1538 390
rect 2123 566 2153 592
rect 1816 493 1846 508
rect 1906 493 1936 508
rect 2016 493 2046 508
rect 1813 470 1849 493
rect 1903 470 1939 493
rect 1735 454 1849 470
rect 1735 420 1751 454
rect 1785 440 1849 454
rect 1901 454 1971 470
rect 1785 420 1801 440
rect 1735 404 1801 420
rect 1901 420 1921 454
rect 1955 420 1971 454
rect 1901 404 1971 420
rect 1124 299 1140 333
rect 1174 299 1190 333
rect 1333 310 1369 349
rect 1124 283 1190 299
rect 1279 294 1369 310
rect 1457 322 1473 356
rect 1507 353 1538 356
rect 1614 353 1644 368
rect 1901 353 1931 404
rect 1507 323 1931 353
rect 1507 322 1736 323
rect 1457 309 1736 322
rect 1457 306 1538 309
rect 901 236 968 252
rect 938 209 968 236
rect 1038 209 1068 283
rect 1279 260 1295 294
rect 1329 260 1369 294
rect 1279 244 1369 260
rect 1110 209 1140 235
rect 1310 222 1340 244
rect 1508 222 1538 306
rect 793 169 859 203
rect 793 135 809 169
rect 843 135 859 169
rect 384 87 414 113
rect 470 87 500 113
rect 548 87 578 113
rect 663 87 693 113
rect 793 101 859 135
rect 108 48 138 74
rect 186 48 216 74
rect 793 67 809 101
rect 843 67 859 101
rect 793 51 859 67
rect 938 51 968 125
rect 1038 99 1068 125
rect 1110 51 1140 125
rect 1706 181 1736 309
rect 2013 301 2049 493
rect 2123 383 2153 398
rect 2627 493 2657 508
rect 2711 493 2741 508
rect 2120 366 2156 383
rect 2327 377 2357 392
rect 2519 377 2549 392
rect 1979 285 2049 301
rect 2091 350 2164 366
rect 2091 316 2107 350
rect 2141 316 2164 350
rect 2091 300 2164 316
rect 2324 304 2360 377
rect 2516 360 2552 377
rect 1842 253 1931 269
rect 1842 219 1881 253
rect 1915 219 1931 253
rect 1842 203 1931 219
rect 1979 251 1999 285
rect 2033 251 2049 285
rect 1979 235 2049 251
rect 1842 181 1872 203
rect 1979 181 2009 235
rect 2134 202 2164 300
rect 2226 288 2360 304
rect 2408 344 2474 360
rect 2408 310 2424 344
rect 2458 310 2474 344
rect 2408 294 2474 310
rect 2516 344 2582 360
rect 2516 310 2532 344
rect 2566 310 2582 344
rect 2516 294 2582 310
rect 2624 317 2660 493
rect 2708 476 2744 493
rect 2702 460 2768 476
rect 2702 426 2718 460
rect 2752 426 2768 460
rect 2853 449 2883 464
rect 2850 426 2886 449
rect 2702 410 2768 426
rect 2624 301 2690 317
rect 2226 254 2242 288
rect 2276 254 2310 288
rect 2344 254 2360 288
rect 2226 252 2360 254
rect 2226 222 2402 252
rect 2372 202 2402 222
rect 2444 202 2474 294
rect 938 21 1140 51
rect 1310 48 1340 74
rect 1508 48 1538 74
rect 1706 71 1736 97
rect 1842 71 1872 97
rect 1979 71 2009 97
rect 2539 158 2569 294
rect 2624 267 2640 301
rect 2674 267 2690 301
rect 2624 251 2690 267
rect 2738 203 2768 410
rect 2816 410 2886 426
rect 2816 376 2832 410
rect 2866 376 2886 410
rect 2816 342 2886 376
rect 3055 353 3085 368
rect 3148 353 3178 368
rect 2816 308 2832 342
rect 2866 322 2886 342
rect 3052 322 3088 353
rect 3145 322 3181 353
rect 2866 308 3181 322
rect 2816 292 3181 308
rect 2617 173 2768 203
rect 2838 272 3166 292
rect 2617 158 2647 173
rect 2838 158 2868 272
rect 3050 222 3080 272
rect 3136 222 3166 272
rect 2134 48 2164 74
rect 2372 48 2402 74
rect 2444 48 2474 74
rect 2539 48 2569 74
rect 2617 48 2647 74
rect 2838 48 2868 74
rect 3050 48 3080 74
rect 3136 48 3166 74
<< polycont >>
rect 88 348 122 382
rect 88 280 122 314
rect 211 374 245 408
rect 211 306 245 340
rect 88 212 122 246
rect 319 280 353 314
rect 427 320 461 354
rect 564 319 598 353
rect 809 339 843 373
rect 809 271 843 305
rect 809 203 843 237
rect 917 252 951 286
rect 1032 299 1066 333
rect 1140 367 1174 401
rect 1473 390 1507 424
rect 1751 420 1785 454
rect 1921 420 1955 454
rect 1140 299 1174 333
rect 1473 322 1507 356
rect 1295 260 1329 294
rect 809 135 843 169
rect 809 67 843 101
rect 2107 316 2141 350
rect 1881 219 1915 253
rect 1999 251 2033 285
rect 2424 310 2458 344
rect 2532 310 2566 344
rect 2718 426 2752 460
rect 2242 254 2276 288
rect 2310 254 2344 288
rect 2640 267 2674 301
rect 2832 376 2866 410
rect 2832 308 2866 342
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3264 683
rect 17 580 102 596
rect 17 546 52 580
rect 86 546 102 580
rect 17 510 102 546
rect 210 578 260 649
rect 210 544 226 578
rect 210 526 260 544
rect 294 581 464 615
rect 17 476 52 510
rect 86 492 102 510
rect 294 492 328 581
rect 86 476 328 492
rect 17 458 328 476
rect 362 520 396 547
rect 17 162 51 458
rect 362 424 396 486
rect 430 492 464 581
rect 498 577 548 649
rect 532 543 548 577
rect 498 526 548 543
rect 650 579 700 595
rect 650 545 666 579
rect 650 509 700 545
rect 650 492 666 509
rect 430 475 666 492
rect 430 458 700 475
rect 195 408 477 424
rect 85 382 161 398
rect 85 348 88 382
rect 122 348 161 382
rect 85 314 161 348
rect 85 280 88 314
rect 122 280 161 314
rect 85 246 161 280
rect 85 212 88 246
rect 122 212 161 246
rect 85 196 161 212
rect 195 374 211 408
rect 245 390 477 408
rect 245 374 261 390
rect 195 340 261 374
rect 195 306 211 340
rect 245 306 261 340
rect 195 230 261 306
rect 303 314 369 356
rect 303 280 319 314
rect 353 280 369 314
rect 411 354 477 390
rect 411 320 427 354
rect 461 320 477 354
rect 411 304 477 320
rect 511 353 614 369
rect 511 350 564 353
rect 545 319 564 350
rect 598 319 614 353
rect 545 316 614 319
rect 511 303 614 316
rect 303 264 369 280
rect 666 269 700 458
rect 634 235 700 269
rect 734 581 968 615
rect 734 579 790 581
rect 734 545 756 579
rect 734 509 790 545
rect 734 475 756 509
rect 734 459 790 475
rect 825 516 900 547
rect 825 482 866 516
rect 195 196 373 230
rect 634 201 668 235
rect 734 201 768 459
rect 825 451 900 482
rect 934 485 968 581
rect 1002 570 1052 649
rect 1036 536 1052 570
rect 1002 519 1052 536
rect 1160 571 1226 587
rect 1160 537 1176 571
rect 1210 537 1226 571
rect 1272 576 1339 649
rect 1272 542 1288 576
rect 1322 542 1339 576
rect 1551 578 1617 649
rect 1551 544 1567 578
rect 1601 544 1617 578
rect 1551 542 1617 544
rect 1753 567 1803 596
rect 1753 538 1769 567
rect 1160 508 1226 537
rect 1651 533 1769 538
rect 1651 508 1803 533
rect 1160 504 1803 508
rect 1837 567 1909 596
rect 1837 533 1859 567
rect 1893 533 1909 567
rect 2043 580 2109 649
rect 2043 546 2059 580
rect 2093 546 2109 580
rect 2262 580 2330 649
rect 2262 546 2279 580
rect 2313 546 2330 580
rect 2580 567 2650 596
rect 1837 504 1909 533
rect 2614 533 2650 567
rect 1160 501 1685 504
rect 1160 485 1176 501
rect 934 467 1176 485
rect 1210 474 1685 501
rect 1210 467 1245 474
rect 934 451 1245 467
rect 825 417 859 451
rect 323 172 373 196
rect 17 133 113 162
rect 17 99 63 133
rect 97 99 113 133
rect 17 70 113 99
rect 211 133 277 162
rect 211 99 227 133
rect 261 99 277 133
rect 323 138 339 172
rect 323 109 373 138
rect 409 172 475 201
rect 409 138 425 172
rect 459 138 475 172
rect 211 17 277 99
rect 409 17 475 138
rect 573 185 668 201
rect 573 151 603 185
rect 637 151 668 185
rect 573 135 668 151
rect 702 172 768 201
rect 702 138 718 172
rect 752 138 768 172
rect 702 109 768 138
rect 802 401 1177 417
rect 802 383 1140 401
rect 802 373 859 383
rect 802 339 809 373
rect 843 339 859 373
rect 1124 367 1140 383
rect 1174 367 1177 401
rect 802 305 859 339
rect 802 271 809 305
rect 843 271 859 305
rect 991 333 1082 349
rect 802 237 859 271
rect 802 203 809 237
rect 843 203 859 237
rect 893 286 957 302
rect 893 252 917 286
rect 951 252 957 286
rect 893 236 957 252
rect 991 299 1032 333
rect 1066 299 1082 333
rect 991 236 1082 299
rect 1124 333 1177 367
rect 1124 299 1140 333
rect 1174 299 1177 333
rect 1124 283 1177 299
rect 1211 213 1245 451
rect 1379 424 1523 440
rect 1379 417 1473 424
rect 1413 390 1473 417
rect 1507 390 1523 424
rect 1413 383 1523 390
rect 1379 356 1523 383
rect 1379 322 1473 356
rect 1507 322 1523 356
rect 1279 294 1345 310
rect 1279 260 1295 294
rect 1329 260 1345 294
rect 1279 236 1345 260
rect 1379 306 1523 322
rect 1573 330 1607 474
rect 1729 454 1801 470
rect 1729 440 1751 454
rect 1641 420 1751 440
rect 1785 420 1801 454
rect 1641 419 1801 420
rect 1641 385 1657 419
rect 1691 404 1801 419
rect 1691 385 1763 404
rect 1641 364 1763 385
rect 1837 366 1871 504
rect 1943 478 2546 512
rect 1943 470 1977 478
rect 1905 454 1977 470
rect 1905 420 1921 454
rect 1955 420 1977 454
rect 1905 404 1977 420
rect 2150 410 2166 444
rect 2200 410 2225 444
rect 802 202 859 203
rect 802 178 943 202
rect 802 169 893 178
rect 802 135 809 169
rect 843 144 893 169
rect 927 144 943 178
rect 843 135 943 144
rect 802 121 943 135
rect 977 178 1043 202
rect 977 144 993 178
rect 1027 144 1043 178
rect 802 101 859 121
rect 802 67 809 101
rect 843 67 859 101
rect 802 51 859 67
rect 977 17 1043 144
rect 1135 184 1245 213
rect 1379 202 1413 306
rect 1573 296 1695 330
rect 1135 150 1151 184
rect 1185 179 1245 184
rect 1185 150 1201 179
rect 1135 121 1201 150
rect 1335 168 1351 202
rect 1385 168 1413 202
rect 1247 120 1299 136
rect 1247 86 1264 120
rect 1298 86 1299 120
rect 1247 17 1299 86
rect 1335 120 1413 168
rect 1335 86 1351 120
rect 1385 86 1413 120
rect 1335 70 1413 86
rect 1447 210 1497 226
rect 1447 176 1463 210
rect 1447 120 1497 176
rect 1447 86 1463 120
rect 1447 17 1497 86
rect 1533 210 1599 226
rect 1533 176 1549 210
rect 1583 176 1599 210
rect 1533 120 1599 176
rect 1533 86 1549 120
rect 1583 86 1599 120
rect 1645 169 1695 296
rect 1645 135 1661 169
rect 1645 119 1695 135
rect 1533 85 1599 86
rect 1729 85 1763 364
rect 1797 350 2157 366
rect 1797 332 2107 350
rect 1797 169 1831 332
rect 2091 316 2107 332
rect 2141 316 2157 350
rect 2091 306 2157 316
rect 2191 304 2225 410
rect 2408 344 2474 360
rect 2408 310 2424 344
rect 2458 310 2474 344
rect 1983 285 2049 298
rect 1797 119 1831 135
rect 1865 253 1931 269
rect 1865 219 1881 253
rect 1915 219 1931 253
rect 1983 251 1999 285
rect 2033 272 2049 285
rect 2191 288 2360 304
rect 2191 272 2242 288
rect 2033 254 2242 272
rect 2276 254 2310 288
rect 2344 254 2360 288
rect 2033 251 2360 254
rect 1983 238 2360 251
rect 2408 272 2474 310
rect 2512 351 2546 478
rect 2580 385 2650 533
rect 2738 580 2846 649
rect 2738 546 2775 580
rect 2809 546 2846 580
rect 2738 530 2846 546
rect 2880 580 2950 596
rect 2880 546 2896 580
rect 2930 546 2950 580
rect 2880 510 2950 546
rect 2880 494 2896 510
rect 2702 476 2896 494
rect 2930 476 2950 510
rect 2702 460 2950 476
rect 2702 426 2718 460
rect 2752 426 2768 460
rect 2702 419 2768 426
rect 2816 410 2882 426
rect 2816 385 2832 410
rect 2616 376 2832 385
rect 2866 376 2882 410
rect 2616 351 2882 376
rect 2512 344 2582 351
rect 2512 310 2532 344
rect 2566 310 2582 344
rect 2512 306 2582 310
rect 2624 301 2690 317
rect 2624 272 2640 301
rect 2408 267 2640 272
rect 2674 267 2690 301
rect 2408 238 2690 267
rect 1865 204 1931 219
rect 1865 170 2141 204
rect 1865 85 1899 170
rect 1533 51 1899 85
rect 2020 120 2073 136
rect 2020 86 2037 120
rect 2071 86 2073 120
rect 2020 17 2073 86
rect 2107 85 2141 170
rect 2175 179 2225 238
rect 2408 204 2442 238
rect 2724 204 2758 351
rect 2816 342 2882 351
rect 2816 308 2832 342
rect 2866 308 2882 342
rect 2816 292 2882 308
rect 2916 356 2950 460
rect 2992 580 3058 649
rect 2992 546 3008 580
rect 3042 546 3058 580
rect 2992 501 3058 546
rect 2992 467 3008 501
rect 3042 467 3058 501
rect 2992 424 3058 467
rect 2992 390 3008 424
rect 3042 390 3058 424
rect 3092 580 3141 596
rect 3092 546 3099 580
rect 3133 546 3141 580
rect 3092 499 3141 546
rect 3092 465 3099 499
rect 3133 465 3141 499
rect 3092 430 3141 465
rect 3175 580 3241 649
rect 3175 546 3191 580
rect 3225 546 3241 580
rect 3175 498 3241 546
rect 3175 464 3191 498
rect 3225 464 3241 498
rect 3092 414 3239 430
rect 3092 380 3099 414
rect 3133 380 3239 414
rect 2916 350 3047 356
rect 2916 316 3007 350
rect 3041 316 3047 350
rect 2916 310 3047 316
rect 3092 310 3239 380
rect 2916 258 2950 310
rect 2209 145 2225 179
rect 2175 119 2225 145
rect 2259 170 2442 204
rect 2478 170 2758 204
rect 2863 224 2950 258
rect 3092 226 3141 310
rect 2259 85 2293 170
rect 2107 51 2293 85
rect 2327 120 2377 136
rect 2361 86 2377 120
rect 2327 17 2377 86
rect 2478 133 2544 170
rect 2478 99 2494 133
rect 2528 99 2544 133
rect 2478 70 2544 99
rect 2642 120 2829 136
rect 2642 86 2658 120
rect 2692 86 2779 120
rect 2813 86 2829 120
rect 2642 17 2829 86
rect 2863 133 2929 224
rect 3075 210 3141 226
rect 2863 99 2879 133
rect 2913 99 2929 133
rect 2863 70 2929 99
rect 2975 156 2991 190
rect 3025 156 3041 190
rect 2975 120 3041 156
rect 2975 86 2991 120
rect 3025 86 3041 120
rect 2975 17 3041 86
rect 3075 176 3091 210
rect 3125 176 3141 210
rect 3075 120 3141 176
rect 3075 86 3091 120
rect 3125 86 3141 120
rect 3075 70 3141 86
rect 3175 210 3241 226
rect 3175 176 3191 210
rect 3225 176 3241 210
rect 3175 120 3241 176
rect 3175 86 3191 120
rect 3225 86 3241 120
rect 3175 17 3241 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3264 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 3199 649 3233 683
rect 511 316 545 350
rect 3007 316 3041 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
<< metal1 >>
rect 0 683 3264 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3264 683
rect 0 617 3264 649
rect 499 350 557 356
rect 499 316 511 350
rect 545 347 557 350
rect 2995 350 3053 356
rect 2995 347 3007 350
rect 545 319 3007 347
rect 545 316 557 319
rect 499 310 557 316
rect 2995 316 3007 319
rect 3041 316 3053 350
rect 2995 310 3053 316
rect 0 17 3264 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3264 17
rect 0 -49 3264 -17
<< labels >>
rlabel comment s 0 0 0 0 4 sedfxtp_2
flabel comment s 1711 344 1711 344 0 FreeSans 200 0 0 0 no_jumper_check
flabel pwell s 0 0 3264 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nwell s 0 617 3264 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 0 617 3264 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 3264 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 895 242 929 276 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 1279 242 1313 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 127 242 161 276 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 DE
port 3 nsew
flabel corelocali s 991 242 1025 276 0 FreeSans 340 0 0 0 SCD
port 4 nsew
flabel corelocali s 3103 316 3137 350 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 3199 316 3233 350 0 FreeSans 340 0 0 0 Q
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 3264 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 436894
string GDS_START 414684
<< end >>
