magic
tech sky130A
magscale 1 2
timestamp 1601050047
<< nwell >>
rect -38 332 1190 704
<< pwell >>
rect 0 0 1152 49
<< scpmos >>
rect 97 368 127 592
rect 187 368 217 592
rect 277 368 307 592
rect 367 368 397 592
rect 463 368 493 592
rect 553 368 583 592
rect 747 368 777 592
rect 837 368 867 592
rect 927 368 957 592
rect 1017 368 1047 592
<< nmoslvt >>
rect 98 74 128 222
rect 184 74 214 222
rect 270 74 300 222
rect 356 74 386 222
rect 572 74 602 222
rect 658 74 688 222
rect 744 74 774 222
rect 912 74 942 222
<< ndiff >>
rect 45 194 98 222
rect 45 160 53 194
rect 87 160 98 194
rect 45 120 98 160
rect 45 86 53 120
rect 87 86 98 120
rect 45 74 98 86
rect 128 127 184 222
rect 128 93 139 127
rect 173 93 184 127
rect 128 74 184 93
rect 214 186 270 222
rect 214 152 225 186
rect 259 152 270 186
rect 214 116 270 152
rect 214 82 225 116
rect 259 82 270 116
rect 214 74 270 82
rect 300 120 356 222
rect 300 86 311 120
rect 345 86 356 120
rect 300 74 356 86
rect 386 191 439 222
rect 386 157 397 191
rect 431 157 439 191
rect 386 74 439 157
rect 519 207 572 222
rect 519 173 527 207
rect 561 173 572 207
rect 519 74 572 173
rect 602 120 658 222
rect 602 86 613 120
rect 647 86 658 120
rect 602 74 658 86
rect 688 210 744 222
rect 688 176 699 210
rect 733 176 744 210
rect 688 120 744 176
rect 688 86 699 120
rect 733 86 744 120
rect 688 74 744 86
rect 774 152 912 222
rect 774 118 785 152
rect 819 118 867 152
rect 901 118 912 152
rect 774 74 912 118
rect 942 210 995 222
rect 942 176 953 210
rect 987 176 995 210
rect 942 120 995 176
rect 942 86 953 120
rect 987 86 995 120
rect 942 74 995 86
<< pdiff >>
rect 42 580 97 592
rect 42 546 50 580
rect 84 546 97 580
rect 42 497 97 546
rect 42 463 50 497
rect 84 463 97 497
rect 42 414 97 463
rect 42 380 50 414
rect 84 380 97 414
rect 42 368 97 380
rect 127 580 187 592
rect 127 546 140 580
rect 174 546 187 580
rect 127 497 187 546
rect 127 463 140 497
rect 174 463 187 497
rect 127 414 187 463
rect 127 380 140 414
rect 174 380 187 414
rect 127 368 187 380
rect 217 580 277 592
rect 217 546 230 580
rect 264 546 277 580
rect 217 462 277 546
rect 217 428 230 462
rect 264 428 277 462
rect 217 368 277 428
rect 307 580 367 592
rect 307 546 320 580
rect 354 546 367 580
rect 307 497 367 546
rect 307 463 320 497
rect 354 463 367 497
rect 307 414 367 463
rect 307 380 320 414
rect 354 380 367 414
rect 307 368 367 380
rect 397 580 463 592
rect 397 546 413 580
rect 447 546 463 580
rect 397 462 463 546
rect 397 428 413 462
rect 447 428 463 462
rect 397 368 463 428
rect 493 580 553 592
rect 493 546 506 580
rect 540 546 553 580
rect 493 497 553 546
rect 493 463 506 497
rect 540 463 553 497
rect 493 414 553 463
rect 493 380 506 414
rect 540 380 553 414
rect 493 368 553 380
rect 583 580 638 592
rect 583 546 596 580
rect 630 546 638 580
rect 583 498 638 546
rect 583 464 596 498
rect 630 464 638 498
rect 583 368 638 464
rect 692 576 747 592
rect 692 542 700 576
rect 734 542 747 576
rect 692 497 747 542
rect 692 463 700 497
rect 734 463 747 497
rect 692 368 747 463
rect 777 531 837 592
rect 777 497 790 531
rect 824 497 837 531
rect 777 440 837 497
rect 777 406 790 440
rect 824 406 837 440
rect 777 368 837 406
rect 867 580 927 592
rect 867 546 880 580
rect 914 546 927 580
rect 867 507 927 546
rect 867 473 880 507
rect 914 473 927 507
rect 867 431 927 473
rect 867 397 880 431
rect 914 397 927 431
rect 867 368 927 397
rect 957 531 1017 592
rect 957 497 970 531
rect 1004 497 1017 531
rect 957 440 1017 497
rect 957 406 970 440
rect 1004 406 1017 440
rect 957 368 1017 406
rect 1047 580 1102 592
rect 1047 546 1060 580
rect 1094 546 1102 580
rect 1047 502 1102 546
rect 1047 468 1060 502
rect 1094 468 1102 502
rect 1047 368 1102 468
<< ndiffc >>
rect 53 160 87 194
rect 53 86 87 120
rect 139 93 173 127
rect 225 152 259 186
rect 225 82 259 116
rect 311 86 345 120
rect 397 157 431 191
rect 527 173 561 207
rect 613 86 647 120
rect 699 176 733 210
rect 699 86 733 120
rect 785 118 819 152
rect 867 118 901 152
rect 953 176 987 210
rect 953 86 987 120
<< pdiffc >>
rect 50 546 84 580
rect 50 463 84 497
rect 50 380 84 414
rect 140 546 174 580
rect 140 463 174 497
rect 140 380 174 414
rect 230 546 264 580
rect 230 428 264 462
rect 320 546 354 580
rect 320 463 354 497
rect 320 380 354 414
rect 413 546 447 580
rect 413 428 447 462
rect 506 546 540 580
rect 506 463 540 497
rect 506 380 540 414
rect 596 546 630 580
rect 596 464 630 498
rect 700 542 734 576
rect 700 463 734 497
rect 790 497 824 531
rect 790 406 824 440
rect 880 546 914 580
rect 880 473 914 507
rect 880 397 914 431
rect 970 497 1004 531
rect 970 406 1004 440
rect 1060 546 1094 580
rect 1060 468 1094 502
<< poly >>
rect 97 592 127 618
rect 187 592 217 618
rect 277 592 307 618
rect 367 592 397 618
rect 463 592 493 618
rect 553 592 583 618
rect 747 592 777 618
rect 837 592 867 618
rect 927 592 957 618
rect 1017 592 1047 618
rect 97 353 127 368
rect 187 353 217 368
rect 277 353 307 368
rect 367 353 397 368
rect 463 353 493 368
rect 553 353 583 368
rect 747 353 777 368
rect 837 353 867 368
rect 927 353 957 368
rect 1017 353 1047 368
rect 94 310 130 353
rect 184 310 220 353
rect 274 310 310 353
rect 364 310 400 353
rect 460 336 496 353
rect 550 336 586 353
rect 744 336 780 353
rect 834 336 870 353
rect 924 336 960 353
rect 1014 336 1050 353
rect 460 320 640 336
rect 460 310 590 320
rect 94 294 214 310
rect 94 260 110 294
rect 144 260 214 294
rect 274 294 418 310
rect 274 274 290 294
rect 94 244 214 260
rect 98 222 128 244
rect 184 222 214 244
rect 270 260 290 274
rect 324 260 368 294
rect 402 260 418 294
rect 460 276 476 310
rect 510 286 590 310
rect 624 300 640 320
rect 736 320 870 336
rect 624 286 688 300
rect 510 276 688 286
rect 460 270 688 276
rect 736 286 752 320
rect 786 286 820 320
rect 854 286 870 320
rect 736 270 870 286
rect 912 320 1050 336
rect 912 286 985 320
rect 1019 286 1050 320
rect 912 270 1050 286
rect 460 260 602 270
rect 270 244 418 260
rect 270 222 300 244
rect 356 222 386 244
rect 572 222 602 260
rect 658 222 688 270
rect 744 222 774 270
rect 912 222 942 270
rect 98 48 128 74
rect 184 48 214 74
rect 270 48 300 74
rect 356 48 386 74
rect 572 48 602 74
rect 658 48 688 74
rect 744 48 774 74
rect 912 48 942 74
<< polycont >>
rect 110 260 144 294
rect 290 260 324 294
rect 368 260 402 294
rect 476 276 510 310
rect 590 286 624 320
rect 752 286 786 320
rect 820 286 854 320
rect 985 286 1019 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 34 580 84 649
rect 34 546 50 580
rect 34 497 84 546
rect 34 463 50 497
rect 34 414 84 463
rect 34 380 50 414
rect 34 364 84 380
rect 124 580 190 596
rect 124 546 140 580
rect 174 546 190 580
rect 124 497 190 546
rect 124 463 140 497
rect 174 463 190 497
rect 124 414 190 463
rect 124 380 140 414
rect 174 380 190 414
rect 230 580 264 649
rect 230 462 264 546
rect 230 412 264 428
rect 304 580 370 596
rect 304 546 320 580
rect 354 546 370 580
rect 304 497 370 546
rect 304 463 320 497
rect 354 463 370 497
rect 304 414 370 463
rect 124 378 190 380
rect 304 380 320 414
rect 354 380 370 414
rect 410 580 466 649
rect 410 546 413 580
rect 447 546 466 580
rect 410 462 466 546
rect 410 428 413 462
rect 447 428 466 462
rect 410 412 466 428
rect 506 580 540 596
rect 506 497 540 546
rect 506 424 540 463
rect 580 580 646 649
rect 580 546 596 580
rect 630 546 646 580
rect 580 498 646 546
rect 580 464 596 498
rect 630 464 646 498
rect 580 458 646 464
rect 684 581 1110 615
rect 684 576 751 581
rect 684 542 700 576
rect 734 542 751 576
rect 864 580 930 581
rect 684 497 751 542
rect 684 463 700 497
rect 734 463 751 497
rect 684 458 751 463
rect 785 531 824 547
rect 785 497 790 531
rect 785 440 824 497
rect 785 424 790 440
rect 506 414 790 424
rect 304 378 370 380
rect 540 406 790 414
rect 540 390 824 406
rect 864 546 880 580
rect 914 546 930 580
rect 1044 580 1110 581
rect 864 507 930 546
rect 864 473 880 507
rect 914 473 930 507
rect 864 431 930 473
rect 864 397 880 431
rect 914 397 930 431
rect 864 390 930 397
rect 970 531 1004 547
rect 970 440 1004 497
rect 1044 546 1060 580
rect 1094 546 1110 580
rect 1044 502 1110 546
rect 1044 468 1060 502
rect 1094 468 1110 502
rect 1044 458 1110 468
rect 1004 406 1127 424
rect 970 390 1127 406
rect 506 378 540 380
rect 124 344 540 378
rect 574 320 647 356
rect 574 310 590 320
rect 94 294 167 310
rect 94 260 110 294
rect 144 260 167 294
rect 94 244 167 260
rect 121 236 167 244
rect 217 294 418 310
rect 217 260 290 294
rect 324 260 368 294
rect 402 260 418 294
rect 460 276 476 310
rect 510 286 590 310
rect 624 286 647 320
rect 510 276 647 286
rect 460 270 647 276
rect 697 320 935 356
rect 697 286 752 320
rect 786 286 820 320
rect 854 286 935 320
rect 697 270 935 286
rect 969 320 1035 356
rect 969 286 985 320
rect 1019 286 1035 320
rect 969 270 1035 286
rect 217 244 418 260
rect 217 236 263 244
rect 1081 236 1127 390
rect 511 210 1127 236
rect 37 202 87 210
rect 381 202 447 210
rect 37 194 447 202
rect 37 160 53 194
rect 87 191 447 194
rect 87 186 397 191
rect 87 168 225 186
rect 37 120 87 160
rect 259 157 397 186
rect 431 157 447 191
rect 511 207 699 210
rect 511 173 527 207
rect 561 176 699 207
rect 733 202 953 210
rect 733 176 749 202
rect 561 173 749 176
rect 511 170 749 173
rect 259 154 447 157
rect 37 86 53 120
rect 37 70 87 86
rect 123 127 189 134
rect 123 93 139 127
rect 173 93 189 127
rect 123 17 189 93
rect 225 116 259 152
rect 597 120 663 136
rect 225 66 259 82
rect 295 86 311 120
rect 345 86 613 120
rect 647 86 663 120
rect 295 70 663 86
rect 699 120 749 170
rect 937 176 953 202
rect 987 176 1127 210
rect 733 86 749 120
rect 699 70 749 86
rect 783 152 903 168
rect 783 118 785 152
rect 819 118 867 152
rect 901 118 903 152
rect 783 17 903 118
rect 937 120 1127 176
rect 937 86 953 120
rect 987 86 1127 120
rect 937 70 1127 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a311oi_2
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 1087 94 1121 128 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 1087 168 1121 202 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 1087 242 1121 276 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 1087 316 1121 350 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 C1
port 5 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 B1
port 4 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 B1
port 4 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 B1
port 4 nsew
flabel corelocali s 127 242 161 276 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 223 242 257 276 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 1152 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3699648
string GDS_START 3689400
<< end >>
