magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 19 195 89 325
rect 359 153 431 344
rect 465 237 505 274
rect 465 153 553 237
rect 1121 221 1177 323
rect 1289 221 1390 333
rect 2592 51 2663 493
rect 2931 51 3014 484
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3036 561
rect 35 393 69 493
rect 103 427 179 527
rect 35 359 179 393
rect 133 161 179 359
rect 35 127 179 161
rect 35 69 69 127
rect 103 17 179 93
rect 223 69 257 493
rect 291 378 377 493
rect 477 378 553 527
rect 291 103 325 378
rect 591 344 657 485
rect 703 365 742 527
rect 885 404 961 493
rect 1007 442 1073 493
rect 885 364 973 404
rect 539 271 657 344
rect 596 235 657 271
rect 821 264 905 330
rect 596 169 777 235
rect 291 51 377 103
rect 477 17 553 103
rect 596 51 641 169
rect 821 137 855 264
rect 939 230 973 364
rect 889 196 973 230
rect 1017 357 1073 442
rect 1158 401 1226 493
rect 1270 435 1339 527
rect 1492 430 1558 493
rect 1600 435 1838 475
rect 1158 367 1474 401
rect 677 17 753 122
rect 889 51 953 196
rect 1017 165 1051 357
rect 1211 187 1245 367
rect 1424 271 1474 367
rect 1508 373 1558 430
rect 1508 237 1542 373
rect 999 129 1051 165
rect 999 51 1039 129
rect 1179 103 1245 187
rect 1073 51 1245 103
rect 1289 17 1339 181
rect 1460 113 1542 237
rect 1576 225 1623 344
rect 1657 331 1760 401
rect 1657 191 1691 331
rect 1794 315 1838 435
rect 1872 367 1919 527
rect 1794 297 1919 315
rect 1580 147 1691 191
rect 1739 263 1919 297
rect 1739 113 1773 263
rect 1885 249 1919 263
rect 1953 275 2029 493
rect 2071 421 2129 527
rect 2252 433 2475 471
rect 1811 213 1861 219
rect 1953 213 2146 275
rect 2225 249 2273 393
rect 1811 209 2146 213
rect 1811 153 2044 209
rect 2307 207 2381 399
rect 1460 51 1584 113
rect 1628 51 1773 113
rect 1836 17 1915 112
rect 1953 51 2044 153
rect 2275 141 2381 207
rect 2090 17 2145 123
rect 2425 107 2475 433
rect 2519 299 2553 527
rect 2282 66 2475 107
rect 2509 17 2558 180
rect 2721 244 2789 493
rect 2833 293 2880 527
rect 2697 178 2789 244
rect 2823 214 2889 259
rect 2721 51 2789 178
rect 2833 17 2880 180
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3036 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 2881 527 2915 561
rect 2973 527 3007 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
rect 2881 -17 2915 17
rect 2973 -17 3007 17
<< metal1 >>
rect 0 561 3036 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3036 561
rect 0 496 3036 527
rect 0 17 3036 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3036 17
rect 0 -48 3036 -17
<< obsm1 >>
rect 125 388 183 397
rect 1657 388 1725 397
rect 2215 388 2283 397
rect 125 360 2283 388
rect 125 351 183 360
rect 1657 351 1725 360
rect 2215 351 2283 360
rect 201 320 269 329
rect 1565 320 1633 329
rect 2309 320 2377 329
rect 201 292 2377 320
rect 201 283 269 292
rect 1565 283 1633 292
rect 2309 283 2377 292
rect 2421 252 2479 261
rect 2827 252 2885 261
rect 2421 224 2885 252
rect 2421 215 2479 224
rect 2827 215 2885 224
rect 809 184 867 193
rect 2728 184 2786 193
rect 809 156 2786 184
rect 809 147 867 156
rect 2728 147 2786 156
rect 279 116 337 125
rect 885 116 953 125
rect 279 79 953 116
rect 981 116 1049 125
rect 1441 116 1509 125
rect 981 79 1509 116
<< labels >>
rlabel locali s 19 195 89 325 6 CLK
port 1 nsew signal input
rlabel locali s 359 153 431 344 6 D
port 2 nsew signal input
rlabel locali s 465 237 505 274 6 DE
port 3 nsew signal input
rlabel locali s 465 153 553 237 6 DE
port 3 nsew signal input
rlabel locali s 2931 51 3014 484 6 Q
port 4 nsew signal output
rlabel locali s 2592 51 2663 493 6 Q_N
port 5 nsew signal output
rlabel locali s 1289 221 1390 333 6 SCD
port 6 nsew signal input
rlabel locali s 1121 221 1177 323 6 SCE
port 7 nsew signal input
rlabel metal1 s 0 -48 3036 48 8 VGND
port 8 nsew ground bidirectional
rlabel metal1 s 0 496 3036 592 6 VPWR
port 9 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 3036 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 429640
string GDS_START 407262
<< end >>
