magic
tech sky130A
magscale 1 2
timestamp 1604502693
<< nwell >>
rect -38 261 1694 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 251 47 281 177
rect 335 47 365 177
rect 419 47 449 177
rect 503 47 533 177
rect 587 47 617 177
rect 671 47 701 177
rect 755 47 785 177
rect 950 47 980 177
rect 1034 47 1064 177
rect 1118 47 1148 177
rect 1202 47 1232 177
rect 1286 47 1316 177
rect 1370 47 1400 177
rect 1454 47 1484 177
rect 1538 47 1568 177
<< pmoshvt >>
rect 79 297 109 497
rect 267 309 297 497
rect 351 309 381 497
rect 435 309 465 497
rect 519 309 549 497
rect 603 309 633 497
rect 687 309 717 497
rect 771 309 801 497
rect 855 309 885 497
rect 950 297 980 497
rect 1034 297 1064 497
rect 1118 297 1148 497
rect 1202 297 1232 497
rect 1286 297 1316 497
rect 1370 297 1400 497
rect 1454 297 1484 497
rect 1538 297 1568 497
<< ndiff >>
rect 27 106 79 177
rect 27 72 35 106
rect 69 72 79 106
rect 27 47 79 72
rect 109 89 163 177
rect 109 55 119 89
rect 153 55 163 89
rect 109 47 163 55
rect 193 124 251 177
rect 193 90 207 124
rect 241 90 251 124
rect 193 47 251 90
rect 281 89 335 177
rect 281 55 291 89
rect 325 55 335 89
rect 281 47 335 55
rect 365 124 419 177
rect 365 90 375 124
rect 409 90 419 124
rect 365 47 419 90
rect 449 89 503 177
rect 449 55 459 89
rect 493 55 503 89
rect 449 47 503 55
rect 533 124 587 177
rect 533 90 543 124
rect 577 90 587 124
rect 533 47 587 90
rect 617 89 671 177
rect 617 55 627 89
rect 661 55 671 89
rect 617 47 671 55
rect 701 124 755 177
rect 701 90 711 124
rect 745 90 755 124
rect 701 47 755 90
rect 785 89 841 177
rect 785 55 795 89
rect 829 55 841 89
rect 785 47 841 55
rect 898 124 950 177
rect 898 90 906 124
rect 940 90 950 124
rect 898 47 950 90
rect 980 169 1034 177
rect 980 135 990 169
rect 1024 135 1034 169
rect 980 47 1034 135
rect 1064 89 1118 177
rect 1064 55 1074 89
rect 1108 55 1118 89
rect 1064 47 1118 55
rect 1148 169 1202 177
rect 1148 135 1158 169
rect 1192 135 1202 169
rect 1148 47 1202 135
rect 1232 89 1286 177
rect 1232 55 1242 89
rect 1276 55 1286 89
rect 1232 47 1286 55
rect 1316 169 1370 177
rect 1316 135 1326 169
rect 1360 135 1370 169
rect 1316 47 1370 135
rect 1400 89 1454 177
rect 1400 55 1410 89
rect 1444 55 1454 89
rect 1400 47 1454 55
rect 1484 169 1538 177
rect 1484 135 1494 169
rect 1528 135 1538 169
rect 1484 47 1538 135
rect 1568 89 1624 177
rect 1568 55 1578 89
rect 1612 55 1624 89
rect 1568 47 1624 55
<< pdiff >>
rect 27 450 79 497
rect 27 416 35 450
rect 69 416 79 450
rect 27 297 79 416
rect 109 485 161 497
rect 109 451 119 485
rect 153 451 161 485
rect 109 297 161 451
rect 215 465 267 497
rect 215 431 223 465
rect 257 431 267 465
rect 215 309 267 431
rect 297 489 351 497
rect 297 455 307 489
rect 341 455 351 489
rect 297 421 351 455
rect 297 387 307 421
rect 341 387 351 421
rect 297 309 351 387
rect 381 477 435 497
rect 381 443 391 477
rect 425 443 435 477
rect 381 409 435 443
rect 381 375 391 409
rect 425 375 435 409
rect 381 309 435 375
rect 465 489 519 497
rect 465 455 475 489
rect 509 455 519 489
rect 465 421 519 455
rect 465 387 475 421
rect 509 387 519 421
rect 465 309 519 387
rect 549 477 603 497
rect 549 443 559 477
rect 593 443 603 477
rect 549 409 603 443
rect 549 375 559 409
rect 593 375 603 409
rect 549 309 603 375
rect 633 489 687 497
rect 633 455 643 489
rect 677 455 687 489
rect 633 421 687 455
rect 633 387 643 421
rect 677 387 687 421
rect 633 309 687 387
rect 717 477 771 497
rect 717 443 727 477
rect 761 443 771 477
rect 717 409 771 443
rect 717 375 727 409
rect 761 375 771 409
rect 717 309 771 375
rect 801 489 855 497
rect 801 455 811 489
rect 845 455 855 489
rect 801 421 855 455
rect 801 387 811 421
rect 845 387 855 421
rect 801 309 855 387
rect 885 477 950 497
rect 885 443 901 477
rect 935 443 950 477
rect 885 409 950 443
rect 885 375 901 409
rect 935 375 950 409
rect 885 309 950 375
rect 900 297 950 309
rect 980 407 1034 497
rect 980 373 990 407
rect 1024 373 1034 407
rect 980 339 1034 373
rect 980 305 990 339
rect 1024 305 1034 339
rect 980 297 1034 305
rect 1064 477 1118 497
rect 1064 443 1074 477
rect 1108 443 1118 477
rect 1064 409 1118 443
rect 1064 375 1074 409
rect 1108 375 1118 409
rect 1064 297 1118 375
rect 1148 407 1202 497
rect 1148 373 1158 407
rect 1192 373 1202 407
rect 1148 339 1202 373
rect 1148 305 1158 339
rect 1192 305 1202 339
rect 1148 297 1202 305
rect 1232 477 1286 497
rect 1232 443 1242 477
rect 1276 443 1286 477
rect 1232 409 1286 443
rect 1232 375 1242 409
rect 1276 375 1286 409
rect 1232 297 1286 375
rect 1316 407 1370 497
rect 1316 373 1326 407
rect 1360 373 1370 407
rect 1316 339 1370 373
rect 1316 305 1326 339
rect 1360 305 1370 339
rect 1316 297 1370 305
rect 1400 477 1454 497
rect 1400 443 1410 477
rect 1444 443 1454 477
rect 1400 409 1454 443
rect 1400 375 1410 409
rect 1444 375 1454 409
rect 1400 297 1454 375
rect 1484 407 1538 497
rect 1484 373 1494 407
rect 1528 373 1538 407
rect 1484 339 1538 373
rect 1484 305 1494 339
rect 1528 305 1538 339
rect 1484 297 1538 305
rect 1568 477 1620 497
rect 1568 443 1578 477
rect 1612 443 1620 477
rect 1568 409 1620 443
rect 1568 375 1578 409
rect 1612 375 1620 409
rect 1568 297 1620 375
<< ndiffc >>
rect 35 72 69 106
rect 119 55 153 89
rect 207 90 241 124
rect 291 55 325 89
rect 375 90 409 124
rect 459 55 493 89
rect 543 90 577 124
rect 627 55 661 89
rect 711 90 745 124
rect 795 55 829 89
rect 906 90 940 124
rect 990 135 1024 169
rect 1074 55 1108 89
rect 1158 135 1192 169
rect 1242 55 1276 89
rect 1326 135 1360 169
rect 1410 55 1444 89
rect 1494 135 1528 169
rect 1578 55 1612 89
<< pdiffc >>
rect 35 416 69 450
rect 119 451 153 485
rect 223 431 257 465
rect 307 455 341 489
rect 307 387 341 421
rect 391 443 425 477
rect 391 375 425 409
rect 475 455 509 489
rect 475 387 509 421
rect 559 443 593 477
rect 559 375 593 409
rect 643 455 677 489
rect 643 387 677 421
rect 727 443 761 477
rect 727 375 761 409
rect 811 455 845 489
rect 811 387 845 421
rect 901 443 935 477
rect 901 375 935 409
rect 990 373 1024 407
rect 990 305 1024 339
rect 1074 443 1108 477
rect 1074 375 1108 409
rect 1158 373 1192 407
rect 1158 305 1192 339
rect 1242 443 1276 477
rect 1242 375 1276 409
rect 1326 373 1360 407
rect 1326 305 1360 339
rect 1410 443 1444 477
rect 1410 375 1444 409
rect 1494 373 1528 407
rect 1494 305 1528 339
rect 1578 443 1612 477
rect 1578 375 1612 409
<< poly >>
rect 79 497 109 523
rect 267 497 297 523
rect 351 497 381 523
rect 435 497 465 523
rect 519 497 549 523
rect 603 497 633 523
rect 687 497 717 523
rect 771 497 801 523
rect 855 497 885 523
rect 950 497 980 523
rect 1034 497 1064 523
rect 1118 497 1148 523
rect 1202 497 1232 523
rect 1286 497 1316 523
rect 1370 497 1400 523
rect 1454 497 1484 523
rect 1538 497 1568 523
rect 79 265 109 297
rect 22 249 109 265
rect 267 294 297 309
rect 351 294 381 309
rect 435 294 465 309
rect 519 294 549 309
rect 603 294 633 309
rect 687 294 717 309
rect 771 294 801 309
rect 855 294 885 309
rect 267 264 885 294
rect 22 215 32 249
rect 66 222 109 249
rect 831 249 885 264
rect 66 215 785 222
rect 22 199 785 215
rect 831 215 841 249
rect 875 215 885 249
rect 831 199 885 215
rect 950 265 980 297
rect 1034 265 1064 297
rect 950 259 1064 265
rect 1118 259 1148 297
rect 1202 259 1232 297
rect 1286 265 1316 297
rect 1370 265 1400 297
rect 1286 259 1400 265
rect 1454 259 1484 297
rect 1538 261 1568 297
rect 1538 259 1626 261
rect 950 249 1626 259
rect 950 215 1100 249
rect 1134 215 1168 249
rect 1202 215 1236 249
rect 1270 215 1304 249
rect 1338 215 1372 249
rect 1406 215 1440 249
rect 1474 215 1508 249
rect 1542 215 1576 249
rect 1610 215 1626 249
rect 950 205 1626 215
rect 950 199 1064 205
rect 79 192 785 199
rect 79 177 109 192
rect 163 177 193 192
rect 251 177 281 192
rect 335 177 365 192
rect 419 177 449 192
rect 503 177 533 192
rect 587 177 617 192
rect 671 177 701 192
rect 755 177 785 192
rect 950 177 980 199
rect 1034 177 1064 199
rect 1118 177 1148 205
rect 1202 177 1232 205
rect 1286 199 1400 205
rect 1286 177 1316 199
rect 1370 177 1400 199
rect 1454 177 1484 205
rect 1538 203 1626 205
rect 1538 177 1568 203
rect 79 21 109 47
rect 163 21 193 47
rect 251 21 281 47
rect 335 21 365 47
rect 419 21 449 47
rect 503 21 533 47
rect 587 21 617 47
rect 671 21 701 47
rect 755 21 785 47
rect 950 21 980 47
rect 1034 21 1064 47
rect 1118 21 1148 47
rect 1202 21 1232 47
rect 1286 21 1316 47
rect 1370 21 1400 47
rect 1454 21 1484 47
rect 1538 21 1568 47
<< polycont >>
rect 32 215 66 249
rect 841 215 875 249
rect 1100 215 1134 249
rect 1168 215 1202 249
rect 1236 215 1270 249
rect 1304 215 1338 249
rect 1372 215 1406 249
rect 1440 215 1474 249
rect 1508 215 1542 249
rect 1576 215 1610 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 17 450 69 493
rect 17 416 35 450
rect 103 485 175 527
rect 103 451 119 485
rect 153 451 175 485
rect 103 425 175 451
rect 215 465 257 493
rect 215 431 223 465
rect 17 391 69 416
rect 17 357 175 391
rect 17 249 66 323
rect 17 215 32 249
rect 17 199 66 215
rect 100 265 175 357
rect 215 345 257 431
rect 291 489 357 527
rect 291 455 307 489
rect 341 455 357 489
rect 291 421 357 455
rect 291 387 307 421
rect 341 387 357 421
rect 291 379 357 387
rect 391 477 425 493
rect 391 409 425 443
rect 459 489 525 527
rect 459 455 475 489
rect 509 455 525 489
rect 459 421 525 455
rect 459 387 475 421
rect 509 387 525 421
rect 459 379 525 387
rect 559 477 593 493
rect 559 409 593 443
rect 391 345 425 375
rect 627 489 693 527
rect 627 455 643 489
rect 677 455 693 489
rect 627 421 693 455
rect 627 387 643 421
rect 677 387 693 421
rect 627 379 693 387
rect 727 477 761 493
rect 727 409 761 443
rect 559 345 593 375
rect 795 489 861 527
rect 795 455 811 489
rect 845 455 861 489
rect 795 421 861 455
rect 795 387 811 421
rect 845 387 861 421
rect 795 379 861 387
rect 895 477 1639 493
rect 895 443 901 477
rect 935 459 1074 477
rect 935 443 940 459
rect 895 409 940 443
rect 1108 459 1242 477
rect 727 345 761 375
rect 895 375 901 409
rect 935 375 940 409
rect 895 345 940 375
rect 215 311 940 345
rect 974 407 1040 425
rect 974 373 990 407
rect 1024 373 1040 407
rect 974 339 1040 373
rect 1074 409 1108 443
rect 1276 459 1410 477
rect 1074 357 1108 375
rect 1142 407 1208 425
rect 1142 373 1158 407
rect 1192 373 1208 407
rect 974 305 990 339
rect 1024 323 1040 339
rect 1142 339 1208 373
rect 1242 409 1276 443
rect 1444 459 1578 477
rect 1242 357 1276 375
rect 1310 407 1376 425
rect 1310 373 1326 407
rect 1360 373 1376 407
rect 1142 323 1158 339
rect 1024 305 1158 323
rect 1192 323 1208 339
rect 1310 339 1376 373
rect 1410 409 1444 443
rect 1612 443 1639 477
rect 1410 357 1444 375
rect 1478 407 1544 425
rect 1478 373 1494 407
rect 1528 373 1544 407
rect 1310 323 1326 339
rect 1192 305 1326 323
rect 1360 323 1376 339
rect 1478 339 1544 373
rect 1478 323 1494 339
rect 1360 305 1494 323
rect 1528 305 1544 339
rect 974 289 1544 305
rect 1578 409 1639 443
rect 1612 375 1639 409
rect 1578 289 1639 375
rect 100 249 940 265
rect 100 215 841 249
rect 875 215 940 249
rect 100 199 940 215
rect 100 165 139 199
rect 974 170 1050 289
rect 1084 249 1639 255
rect 1084 215 1100 249
rect 1134 215 1168 249
rect 1202 215 1236 249
rect 1270 215 1304 249
rect 1338 215 1372 249
rect 1406 215 1440 249
rect 1474 215 1508 249
rect 1542 215 1576 249
rect 1610 215 1639 249
rect 1084 204 1639 215
rect 974 169 1639 170
rect 17 131 139 165
rect 207 131 940 165
rect 17 106 69 131
rect 17 72 35 106
rect 207 124 241 131
rect 17 51 69 72
rect 103 89 169 97
rect 103 55 119 89
rect 153 55 169 89
rect 103 17 169 55
rect 375 124 409 131
rect 207 51 241 90
rect 275 89 341 97
rect 275 55 291 89
rect 325 55 341 89
rect 275 17 341 55
rect 543 124 577 131
rect 375 51 409 90
rect 443 89 509 97
rect 443 55 459 89
rect 493 55 509 89
rect 443 17 509 55
rect 711 124 745 131
rect 543 51 577 90
rect 611 89 677 97
rect 611 55 627 89
rect 661 55 677 89
rect 611 17 677 55
rect 881 124 940 131
rect 974 135 990 169
rect 1024 135 1158 169
rect 1192 135 1326 169
rect 1360 135 1494 169
rect 1528 135 1639 169
rect 974 127 1639 135
rect 711 51 745 90
rect 779 89 847 97
rect 779 55 795 89
rect 829 55 847 89
rect 779 17 847 55
rect 881 90 906 124
rect 940 90 1639 93
rect 881 89 1639 90
rect 881 55 1074 89
rect 1108 55 1242 89
rect 1276 55 1410 89
rect 1444 55 1578 89
rect 1612 55 1639 89
rect 881 51 1639 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
<< metal1 >>
rect 0 561 1656 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 0 496 1656 527
rect 0 17 1656 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
rect 0 -48 1656 -17
<< labels >>
flabel corelocali s 1322 221 1356 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 1230 221 1264 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 1138 221 1172 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 1598 221 1632 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 1506 221 1540 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 1414 221 1448 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 1322 357 1356 391 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 1506 357 1540 391 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 1506 289 1540 323 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 1414 289 1448 323 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 200 0 0 0 TE
port 2 nsew
flabel corelocali s 30 289 64 323 0 FreeSans 200 0 0 0 TE
port 2 nsew
flabel corelocali s 1138 289 1172 323 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 1046 289 1080 323 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 1322 289 1356 323 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 1230 289 1264 323 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew
rlabel comment s 0 0 0 0 4 einvp_8
<< properties >>
string FIXED_BBOX 0 0 1656 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2006066
string GDS_START 1993444
string path 0.000 13.600 41.400 13.600 
<< end >>
