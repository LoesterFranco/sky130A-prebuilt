magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 2024 561
rect 114 435 164 527
rect 282 435 332 527
rect 890 435 940 527
rect 1058 435 1108 527
rect 1226 435 1276 527
rect 1394 435 1444 527
rect 526 289 1233 323
rect 1576 333 1634 425
rect 1752 333 1802 425
rect 1576 325 1802 333
rect 1920 325 2007 493
rect 1576 289 2007 325
rect 526 255 560 289
rect 1199 255 1233 289
rect 85 215 560 255
rect 594 221 1148 255
rect 594 215 1000 221
rect 1199 215 1474 255
rect 1030 181 1116 187
rect 1570 181 1661 187
rect 1947 181 2007 289
rect 17 17 72 113
rect 206 17 240 111
rect 374 17 408 111
rect 542 17 576 111
rect 710 17 764 179
rect 833 129 1116 181
rect 1570 147 2007 181
rect 1570 145 1726 147
rect 1234 17 1268 111
rect 1402 17 1436 111
rect 1592 17 1626 111
rect 1660 51 1726 145
rect 1760 17 1794 111
rect 1828 51 1894 147
rect 1928 17 1962 111
rect 0 -17 2024 17
<< obsli1 >>
rect 17 401 80 493
rect 198 401 248 493
rect 366 459 752 493
rect 366 401 416 459
rect 534 425 584 459
rect 17 357 416 401
rect 450 391 500 425
rect 618 391 668 425
rect 450 357 668 391
rect 702 359 752 459
rect 806 401 856 493
rect 974 401 1024 493
rect 1142 401 1192 493
rect 1310 401 1360 493
rect 1478 459 1886 493
rect 1478 401 1528 459
rect 806 357 1528 401
rect 450 323 484 357
rect 17 289 397 323
rect 431 289 484 323
rect 1310 291 1360 357
rect 1668 367 1718 459
rect 1836 359 1886 459
rect 1452 289 1501 323
rect 1535 289 1542 323
rect 17 181 51 289
rect 1508 255 1542 289
rect 1508 221 1913 255
rect 1708 215 1913 221
rect 17 147 676 181
rect 106 145 676 147
rect 106 51 172 145
rect 274 51 340 145
rect 442 51 508 145
rect 610 51 676 145
rect 1150 145 1536 181
rect 1150 95 1200 145
rect 798 51 1200 95
rect 1302 51 1368 145
rect 1470 51 1536 145
<< obsli1c >>
rect 397 289 431 323
rect 1501 289 1535 323
<< metal1 >>
rect 0 496 2024 592
rect 1029 184 1087 193
rect 1581 184 1639 193
rect 1029 156 1639 184
rect 1029 147 1087 156
rect 1581 147 1639 156
rect 0 -48 2024 48
<< obsm1 >>
rect 385 323 443 329
rect 385 289 397 323
rect 431 320 443 323
rect 1489 323 1547 329
rect 1489 320 1501 323
rect 431 292 1501 320
rect 431 289 443 292
rect 385 283 443 289
rect 1489 289 1501 292
rect 1535 289 1547 323
rect 1489 283 1547 289
<< labels >>
rlabel locali s 1199 255 1233 289 6 A
port 1 nsew signal input
rlabel locali s 1199 215 1474 255 6 A
port 1 nsew signal input
rlabel locali s 526 289 1233 323 6 A
port 1 nsew signal input
rlabel locali s 526 255 560 289 6 A
port 1 nsew signal input
rlabel locali s 85 215 560 255 6 A
port 1 nsew signal input
rlabel locali s 594 221 1148 255 6 B
port 2 nsew signal input
rlabel locali s 594 215 1000 221 6 B
port 2 nsew signal input
rlabel locali s 1030 181 1116 187 6 X
port 3 nsew signal output
rlabel locali s 833 129 1116 181 6 X
port 3 nsew signal output
rlabel locali s 1947 181 2007 289 6 X
port 3 nsew signal output
rlabel locali s 1920 325 2007 493 6 X
port 3 nsew signal output
rlabel locali s 1828 51 1894 147 6 X
port 3 nsew signal output
rlabel locali s 1752 333 1802 425 6 X
port 3 nsew signal output
rlabel locali s 1660 51 1726 145 6 X
port 3 nsew signal output
rlabel locali s 1576 333 1634 425 6 X
port 3 nsew signal output
rlabel locali s 1576 325 1802 333 6 X
port 3 nsew signal output
rlabel locali s 1576 289 2007 325 6 X
port 3 nsew signal output
rlabel locali s 1570 181 1661 187 6 X
port 3 nsew signal output
rlabel locali s 1570 147 2007 181 6 X
port 3 nsew signal output
rlabel locali s 1570 145 1726 147 6 X
port 3 nsew signal output
rlabel metal1 s 1581 184 1639 193 6 X
port 3 nsew signal output
rlabel metal1 s 1581 147 1639 156 6 X
port 3 nsew signal output
rlabel metal1 s 1029 184 1087 193 6 X
port 3 nsew signal output
rlabel metal1 s 1029 156 1639 184 6 X
port 3 nsew signal output
rlabel metal1 s 1029 147 1087 156 6 X
port 3 nsew signal output
rlabel locali s 1928 17 1962 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 1760 17 1794 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 1592 17 1626 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 1402 17 1436 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 1234 17 1268 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 710 17 764 179 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 542 17 576 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 374 17 408 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 206 17 240 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 17 17 72 113 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 2024 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 2024 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 1394 435 1444 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 1226 435 1276 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 1058 435 1108 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 890 435 940 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 282 435 332 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 114 435 164 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 2024 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 2024 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2024 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 661364
string GDS_START 646958
<< end >>
