magic
tech sky130A
magscale 1 2
timestamp 1599588218
<< nwell >>
rect -38 332 1190 704
<< pwell >>
rect 0 0 1152 49
<< scpmos >>
rect 100 387 136 555
rect 190 387 226 555
rect 314 387 350 555
rect 423 368 459 536
rect 562 368 598 592
rect 655 368 691 592
rect 763 368 799 592
rect 853 368 889 592
rect 943 368 979 592
rect 1033 368 1069 592
<< nmoslvt >>
rect 104 74 134 202
rect 190 74 220 202
rect 291 74 321 202
rect 377 74 407 202
rect 575 74 605 222
rect 661 74 691 222
rect 753 74 783 222
rect 853 74 883 222
rect 949 74 979 222
rect 1038 74 1068 222
<< ndiff >>
rect 33 190 104 202
rect 33 156 45 190
rect 79 156 104 190
rect 33 120 104 156
rect 33 86 45 120
rect 79 86 104 120
rect 33 74 104 86
rect 134 187 190 202
rect 134 153 145 187
rect 179 153 190 187
rect 134 116 190 153
rect 134 82 145 116
rect 179 82 190 116
rect 134 74 190 82
rect 220 173 291 202
rect 220 139 231 173
rect 265 139 291 173
rect 220 74 291 139
rect 321 149 377 202
rect 321 115 332 149
rect 366 115 377 149
rect 321 74 377 115
rect 407 149 464 202
rect 407 115 418 149
rect 452 115 464 149
rect 407 74 464 115
rect 518 149 575 222
rect 518 115 530 149
rect 564 115 575 149
rect 518 74 575 115
rect 605 189 661 222
rect 605 155 616 189
rect 650 155 661 189
rect 605 74 661 155
rect 691 210 753 222
rect 691 176 708 210
rect 742 176 753 210
rect 691 120 753 176
rect 691 86 708 120
rect 742 86 753 120
rect 691 74 753 86
rect 783 127 853 222
rect 783 93 808 127
rect 842 93 853 127
rect 783 74 853 93
rect 883 202 949 222
rect 883 168 899 202
rect 933 168 949 202
rect 883 120 949 168
rect 883 86 899 120
rect 933 86 949 120
rect 883 74 949 86
rect 979 120 1038 222
rect 979 86 991 120
rect 1025 86 1038 120
rect 979 74 1038 86
rect 1068 207 1125 222
rect 1068 173 1079 207
rect 1113 173 1125 207
rect 1068 120 1125 173
rect 1068 86 1079 120
rect 1113 86 1125 120
rect 1068 74 1125 86
<< pdiff >>
rect 27 585 85 597
rect 27 551 39 585
rect 73 555 85 585
rect 241 592 299 604
rect 241 558 253 592
rect 287 558 299 592
rect 241 555 299 558
rect 505 580 562 592
rect 73 551 100 555
rect 27 387 100 551
rect 136 433 190 555
rect 136 399 146 433
rect 180 399 190 433
rect 136 387 190 399
rect 226 387 314 555
rect 350 536 400 555
rect 505 546 517 580
rect 551 546 562 580
rect 505 536 562 546
rect 350 440 423 536
rect 350 406 362 440
rect 396 406 423 440
rect 350 387 423 406
rect 373 368 423 387
rect 459 497 562 536
rect 459 463 517 497
rect 551 463 562 497
rect 459 414 562 463
rect 459 380 517 414
rect 551 380 562 414
rect 459 368 562 380
rect 598 580 655 592
rect 598 546 608 580
rect 642 546 655 580
rect 598 497 655 546
rect 598 463 608 497
rect 642 463 655 497
rect 598 414 655 463
rect 598 380 608 414
rect 642 380 655 414
rect 598 368 655 380
rect 691 582 763 592
rect 691 548 708 582
rect 742 548 763 582
rect 691 514 763 548
rect 691 480 708 514
rect 742 480 763 514
rect 691 368 763 480
rect 799 582 853 592
rect 799 548 809 582
rect 843 548 853 582
rect 799 514 853 548
rect 799 480 809 514
rect 843 480 853 514
rect 799 368 853 480
rect 889 531 943 592
rect 889 497 899 531
rect 933 497 943 531
rect 889 462 943 497
rect 889 428 899 462
rect 933 428 943 462
rect 889 368 943 428
rect 979 582 1033 592
rect 979 548 989 582
rect 1023 548 1033 582
rect 979 514 1033 548
rect 979 480 989 514
rect 1023 480 1033 514
rect 979 446 1033 480
rect 979 412 989 446
rect 1023 412 1033 446
rect 979 368 1033 412
rect 1069 580 1125 592
rect 1069 546 1079 580
rect 1113 546 1125 580
rect 1069 510 1125 546
rect 1069 476 1079 510
rect 1113 476 1125 510
rect 1069 440 1125 476
rect 1069 406 1079 440
rect 1113 406 1125 440
rect 1069 368 1125 406
<< ndiffc >>
rect 45 156 79 190
rect 45 86 79 120
rect 145 153 179 187
rect 145 82 179 116
rect 231 139 265 173
rect 332 115 366 149
rect 418 115 452 149
rect 530 115 564 149
rect 616 155 650 189
rect 708 176 742 210
rect 708 86 742 120
rect 808 93 842 127
rect 899 168 933 202
rect 899 86 933 120
rect 991 86 1025 120
rect 1079 173 1113 207
rect 1079 86 1113 120
<< pdiffc >>
rect 39 551 73 585
rect 253 558 287 592
rect 146 399 180 433
rect 517 546 551 580
rect 362 406 396 440
rect 517 463 551 497
rect 517 380 551 414
rect 608 546 642 580
rect 608 463 642 497
rect 608 380 642 414
rect 708 548 742 582
rect 708 480 742 514
rect 809 548 843 582
rect 809 480 843 514
rect 899 497 933 531
rect 899 428 933 462
rect 989 548 1023 582
rect 989 480 1023 514
rect 989 412 1023 446
rect 1079 546 1113 580
rect 1079 476 1113 510
rect 1079 406 1113 440
<< poly >>
rect 562 592 598 618
rect 655 592 691 618
rect 763 592 799 618
rect 853 592 889 618
rect 943 592 979 618
rect 1033 592 1069 618
rect 100 555 136 581
rect 190 555 226 581
rect 314 555 350 581
rect 423 536 459 562
rect 100 326 136 387
rect 190 355 226 387
rect 314 355 350 387
rect 190 339 350 355
rect 30 310 134 326
rect 30 276 46 310
rect 80 276 134 310
rect 30 260 134 276
rect 104 202 134 260
rect 190 305 291 339
rect 325 305 350 339
rect 423 336 459 368
rect 190 289 350 305
rect 393 320 459 336
rect 562 326 598 368
rect 190 202 220 289
rect 291 202 321 289
rect 393 286 409 320
rect 443 286 459 320
rect 393 270 459 286
rect 501 321 598 326
rect 655 321 691 368
rect 763 336 799 368
rect 501 310 691 321
rect 501 276 517 310
rect 551 276 691 310
rect 393 247 423 270
rect 501 260 691 276
rect 739 320 805 336
rect 739 286 755 320
rect 789 286 805 320
rect 739 270 805 286
rect 853 310 889 368
rect 943 310 979 368
rect 853 294 979 310
rect 377 217 423 247
rect 575 222 605 260
rect 661 222 691 260
rect 753 222 783 270
rect 853 260 885 294
rect 919 260 979 294
rect 1033 336 1069 368
rect 1033 320 1099 336
rect 1033 286 1049 320
rect 1083 286 1099 320
rect 1033 270 1099 286
rect 853 244 979 260
rect 853 222 883 244
rect 949 222 979 244
rect 1038 222 1068 270
rect 377 202 407 217
rect 104 48 134 74
rect 190 48 220 74
rect 291 48 321 74
rect 377 48 407 74
rect 575 48 605 74
rect 661 48 691 74
rect 753 48 783 74
rect 853 48 883 74
rect 949 48 979 74
rect 1038 48 1068 74
<< polycont >>
rect 46 276 80 310
rect 291 305 325 339
rect 409 286 443 320
rect 517 276 551 310
rect 755 286 789 320
rect 885 260 919 294
rect 1049 286 1083 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 23 585 89 649
rect 23 551 39 585
rect 73 551 89 585
rect 237 592 303 649
rect 237 558 253 592
rect 287 558 303 592
rect 501 580 567 649
rect 501 546 517 580
rect 551 546 567 580
rect 130 517 467 524
rect 25 490 467 517
rect 25 483 164 490
rect 25 326 71 483
rect 344 449 399 456
rect 130 440 399 449
rect 130 433 362 440
rect 130 399 146 433
rect 180 406 362 433
rect 396 406 399 440
rect 180 399 399 406
rect 130 390 399 399
rect 25 310 96 326
rect 25 276 46 310
rect 80 276 96 310
rect 25 260 96 276
rect 130 255 196 390
rect 275 339 359 356
rect 275 305 291 339
rect 325 305 359 339
rect 433 336 467 490
rect 501 497 567 546
rect 501 463 517 497
rect 551 463 567 497
rect 501 414 567 463
rect 501 380 517 414
rect 551 380 567 414
rect 501 364 567 380
rect 601 580 658 596
rect 601 546 608 580
rect 642 546 658 580
rect 601 497 658 546
rect 601 463 608 497
rect 642 463 658 497
rect 692 582 758 649
rect 692 548 708 582
rect 742 548 758 582
rect 692 514 758 548
rect 692 480 708 514
rect 742 480 758 514
rect 793 582 1039 615
rect 793 548 809 582
rect 843 581 989 582
rect 843 548 859 581
rect 793 514 859 548
rect 973 548 989 581
rect 1023 548 1039 582
rect 793 480 809 514
rect 843 480 859 514
rect 893 531 939 547
rect 893 497 899 531
rect 933 497 939 531
rect 601 446 658 463
rect 893 462 939 497
rect 893 446 899 462
rect 601 428 899 446
rect 933 428 939 462
rect 601 414 939 428
rect 601 380 608 414
rect 642 412 939 414
rect 973 514 1039 548
rect 973 480 989 514
rect 1023 480 1039 514
rect 973 446 1039 480
rect 973 412 989 446
rect 1023 412 1039 446
rect 1079 580 1129 649
rect 1113 546 1129 580
rect 1079 510 1129 546
rect 1113 476 1129 510
rect 1079 440 1129 476
rect 642 380 658 412
rect 1113 406 1129 440
rect 1079 390 1129 406
rect 275 289 359 305
rect 393 320 467 336
rect 393 286 409 320
rect 443 286 467 320
rect 393 270 467 286
rect 501 310 567 326
rect 501 276 517 310
rect 551 276 567 310
rect 501 260 567 276
rect 130 236 281 255
rect 501 236 535 260
rect 130 221 535 236
rect 601 226 658 380
rect 739 356 1019 378
rect 739 344 1099 356
rect 739 320 805 344
rect 739 286 755 320
rect 789 286 805 320
rect 985 320 1099 344
rect 739 270 805 286
rect 869 294 935 310
rect 869 260 885 294
rect 919 260 935 294
rect 985 286 1049 320
rect 1083 286 1099 320
rect 985 270 1099 286
rect 869 236 935 260
rect 29 190 95 206
rect 29 156 45 190
rect 79 156 95 190
rect 231 202 535 221
rect 29 120 95 156
rect 29 86 45 120
rect 79 86 95 120
rect 29 17 95 86
rect 129 153 145 187
rect 179 153 195 187
rect 129 116 195 153
rect 231 173 281 202
rect 265 139 281 173
rect 600 189 658 226
rect 231 121 281 139
rect 316 149 382 165
rect 129 82 145 116
rect 179 85 195 116
rect 316 115 332 149
rect 366 115 382 149
rect 316 85 382 115
rect 179 82 382 85
rect 129 51 382 82
rect 416 149 468 165
rect 416 115 418 149
rect 452 115 468 149
rect 416 17 468 115
rect 514 149 564 165
rect 514 115 530 149
rect 600 155 616 189
rect 650 155 658 189
rect 600 119 658 155
rect 692 210 758 226
rect 692 176 708 210
rect 742 202 758 210
rect 1063 207 1129 226
rect 1063 202 1079 207
rect 742 176 899 202
rect 692 168 899 176
rect 933 173 1079 202
rect 1113 173 1129 207
rect 933 168 1129 173
rect 692 120 758 168
rect 894 154 1129 168
rect 514 85 564 115
rect 692 86 708 120
rect 742 86 758 120
rect 692 85 758 86
rect 514 51 758 85
rect 792 127 858 134
rect 792 93 808 127
rect 842 93 858 127
rect 792 17 858 93
rect 894 120 938 154
rect 1079 120 1129 154
rect 894 86 899 120
rect 933 86 938 120
rect 894 70 938 86
rect 974 86 991 120
rect 1025 86 1043 120
rect 974 17 1043 86
rect 1113 86 1129 120
rect 1079 70 1129 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
rlabel comment s 0 0 0 0 4 o2bb2ai_2
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 895 242 929 276 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A2_N
port 2 nsew
flabel corelocali s 607 168 641 202 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 607 242 641 276 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 607 390 641 424 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 A1_N
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 1152 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1251040
string GDS_START 1241500
<< end >>
