magic
tech sky130A
magscale 1 2
timestamp 1599588232
<< locali >>
rect 1555 270 2087 356
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 23 364 73 649
rect 112 424 163 596
rect 112 390 127 424
rect 161 390 163 424
rect 219 393 253 649
rect 293 424 344 596
rect 26 17 76 226
rect 112 70 163 390
rect 293 390 303 424
rect 337 390 344 424
rect 393 393 443 649
rect 483 424 535 596
rect 197 350 259 356
rect 197 316 211 350
rect 245 316 259 350
rect 197 260 259 316
rect 198 17 257 226
rect 293 70 344 390
rect 483 390 494 424
rect 528 390 535 424
rect 589 393 623 649
rect 662 424 713 596
rect 378 350 435 356
rect 378 316 390 350
rect 424 316 435 350
rect 378 260 435 316
rect 483 271 535 390
rect 662 390 672 424
rect 706 390 713 424
rect 769 393 803 649
rect 843 424 909 596
rect 662 364 713 390
rect 843 390 860 424
rect 894 390 909 424
rect 949 393 983 649
rect 1023 424 1082 596
rect 843 380 909 390
rect 1023 390 1039 424
rect 1073 390 1082 424
rect 1129 393 1163 649
rect 1212 424 1266 596
rect 469 237 535 271
rect 569 350 628 356
rect 569 316 582 350
rect 616 316 628 350
rect 569 260 628 316
rect 379 17 420 226
rect 469 70 522 237
rect 662 226 696 364
rect 747 350 809 356
rect 747 331 760 350
rect 731 316 760 331
rect 794 316 809 350
rect 731 260 809 316
rect 843 226 877 380
rect 935 350 973 356
rect 935 346 936 350
rect 911 316 936 346
rect 970 316 973 350
rect 911 260 973 316
rect 1023 275 1082 390
rect 1212 390 1219 424
rect 1253 390 1266 424
rect 1309 393 1343 649
rect 1396 424 1449 596
rect 1489 458 1539 649
rect 1573 424 1639 596
rect 1679 458 1713 649
rect 1753 424 1819 596
rect 1859 458 1893 649
rect 1933 424 1999 596
rect 1007 241 1082 275
rect 1116 350 1178 356
rect 1116 316 1130 350
rect 1164 316 1178 350
rect 1116 260 1178 316
rect 558 17 592 203
rect 644 70 696 226
rect 730 17 764 226
rect 800 70 877 226
rect 911 17 966 226
rect 1007 70 1066 241
rect 1212 226 1266 390
rect 1396 390 1405 424
rect 1439 390 1449 424
rect 1300 350 1362 356
rect 1300 316 1313 350
rect 1347 316 1362 350
rect 1300 260 1362 316
rect 1396 250 1449 390
rect 1484 390 1999 424
rect 2039 390 2089 649
rect 1484 350 1518 390
rect 1100 17 1166 207
rect 1200 70 1266 226
rect 1300 17 1366 226
rect 1400 70 1450 250
rect 1484 236 1518 316
rect 1484 202 1989 236
rect 1486 17 1552 168
rect 1588 70 1622 202
rect 1658 17 1724 168
rect 1760 70 1794 202
rect 1830 17 1896 168
rect 1939 70 1989 202
rect 2023 17 2089 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 127 390 161 424
rect 303 390 337 424
rect 211 316 245 350
rect 494 390 528 424
rect 390 316 424 350
rect 672 390 706 424
rect 860 390 894 424
rect 1039 390 1073 424
rect 582 316 616 350
rect 760 316 794 350
rect 936 316 970 350
rect 1219 390 1253 424
rect 1130 316 1164 350
rect 1405 390 1439 424
rect 1313 316 1347 350
rect 1484 316 1518 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
<< metal1 >>
rect 0 683 2112 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 0 617 2112 649
rect 0 616 50 617
rect 115 424 1451 430
rect 115 390 127 424
rect 161 390 303 424
rect 337 390 494 424
rect 528 390 672 424
rect 706 390 860 424
rect 894 390 1039 424
rect 1073 390 1219 424
rect 1253 390 1405 424
rect 1439 390 1451 424
rect 115 384 1451 390
rect 0 49 50 50
rect 0 17 2112 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
rect 0 -49 2112 -17
<< obsm1 >>
rect 197 350 1530 356
rect 197 316 211 350
rect 245 316 390 350
rect 424 316 582 350
rect 616 316 760 350
rect 794 316 936 350
rect 970 316 1130 350
rect 1164 316 1313 350
rect 1347 316 1484 350
rect 1518 316 1530 350
rect 197 310 1530 316
<< labels >>
rlabel locali s 1555 270 2087 356 6 A
port 1 nsew signal input
rlabel metal1 s 115 384 1451 430 6 X
port 2 nsew signal output
rlabel metal1 s 0 -49 2112 49 8 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 4 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 617 2112 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2112 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3299012
string GDS_START 3280532
<< end >>
