magic
tech sky130A
magscale 1 2
timestamp 1604502710
<< nwell >>
rect -38 332 1190 704
<< pwell >>
rect 0 0 1152 49
<< scpmos >>
rect 83 368 119 592
rect 173 368 209 592
rect 263 368 299 592
rect 353 368 389 592
rect 443 368 479 592
rect 533 368 569 592
rect 752 368 788 592
rect 852 368 888 592
rect 942 368 978 592
rect 1032 368 1068 592
<< nmoslvt >>
rect 84 74 114 222
rect 170 74 200 222
rect 256 74 286 222
rect 345 74 375 222
rect 431 74 461 222
rect 517 74 547 222
rect 603 74 633 222
rect 689 74 719 222
rect 780 74 810 222
rect 866 74 896 222
rect 952 74 982 222
rect 1038 74 1068 222
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 141 170 222
rect 114 107 125 141
rect 159 107 170 141
rect 114 74 170 107
rect 200 210 256 222
rect 200 176 211 210
rect 245 176 256 210
rect 200 120 256 176
rect 200 86 211 120
rect 245 86 256 120
rect 200 74 256 86
rect 286 127 345 222
rect 286 93 297 127
rect 331 93 345 127
rect 286 74 345 93
rect 375 186 431 222
rect 375 152 386 186
rect 420 152 431 186
rect 375 116 431 152
rect 375 82 386 116
rect 420 82 431 116
rect 375 74 431 82
rect 461 177 517 222
rect 461 143 472 177
rect 506 143 517 177
rect 461 74 517 143
rect 547 127 603 222
rect 547 93 558 127
rect 592 93 603 127
rect 547 74 603 93
rect 633 177 689 222
rect 633 143 644 177
rect 678 143 689 177
rect 633 74 689 143
rect 719 210 780 222
rect 719 176 735 210
rect 769 176 780 210
rect 719 120 780 176
rect 719 86 735 120
rect 769 86 780 120
rect 719 74 780 86
rect 810 136 866 222
rect 810 102 821 136
rect 855 102 866 136
rect 810 74 866 102
rect 896 210 952 222
rect 896 176 907 210
rect 941 176 952 210
rect 896 120 952 176
rect 896 86 907 120
rect 941 86 952 120
rect 896 74 952 86
rect 982 136 1038 222
rect 982 102 993 136
rect 1027 102 1038 136
rect 982 74 1038 102
rect 1068 210 1125 222
rect 1068 176 1079 210
rect 1113 176 1125 210
rect 1068 120 1125 176
rect 1068 86 1079 120
rect 1113 86 1125 120
rect 1068 74 1125 86
<< pdiff >>
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 497 83 546
rect 27 463 39 497
rect 73 463 83 497
rect 27 414 83 463
rect 27 380 39 414
rect 73 380 83 414
rect 27 368 83 380
rect 119 580 173 592
rect 119 546 129 580
rect 163 546 173 580
rect 119 497 173 546
rect 119 463 129 497
rect 163 463 173 497
rect 119 414 173 463
rect 119 380 129 414
rect 163 380 173 414
rect 119 368 173 380
rect 209 580 263 592
rect 209 546 219 580
rect 253 546 263 580
rect 209 508 263 546
rect 209 474 219 508
rect 253 474 263 508
rect 209 368 263 474
rect 299 580 353 592
rect 299 546 309 580
rect 343 546 353 580
rect 299 510 353 546
rect 299 476 309 510
rect 343 476 353 510
rect 299 440 353 476
rect 299 406 309 440
rect 343 406 353 440
rect 299 368 353 406
rect 389 578 443 592
rect 389 544 399 578
rect 433 544 443 578
rect 389 368 443 544
rect 479 419 533 592
rect 479 385 489 419
rect 523 385 533 419
rect 479 368 533 385
rect 569 578 642 592
rect 569 544 596 578
rect 630 544 642 578
rect 569 368 642 544
rect 696 580 752 592
rect 696 546 708 580
rect 742 546 752 580
rect 696 508 752 546
rect 696 474 708 508
rect 742 474 752 508
rect 696 368 752 474
rect 788 531 852 592
rect 788 497 808 531
rect 842 497 852 531
rect 788 440 852 497
rect 788 406 808 440
rect 842 406 852 440
rect 788 368 852 406
rect 888 580 942 592
rect 888 546 898 580
rect 932 546 942 580
rect 888 508 942 546
rect 888 474 898 508
rect 932 474 942 508
rect 888 368 942 474
rect 978 531 1032 592
rect 978 497 988 531
rect 1022 497 1032 531
rect 978 440 1032 497
rect 978 406 988 440
rect 1022 406 1032 440
rect 978 368 1032 406
rect 1068 580 1124 592
rect 1068 546 1078 580
rect 1112 546 1124 580
rect 1068 510 1124 546
rect 1068 476 1078 510
rect 1112 476 1124 510
rect 1068 440 1124 476
rect 1068 406 1078 440
rect 1112 406 1124 440
rect 1068 368 1124 406
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 125 107 159 141
rect 211 176 245 210
rect 211 86 245 120
rect 297 93 331 127
rect 386 152 420 186
rect 386 82 420 116
rect 472 143 506 177
rect 558 93 592 127
rect 644 143 678 177
rect 735 176 769 210
rect 735 86 769 120
rect 821 102 855 136
rect 907 176 941 210
rect 907 86 941 120
rect 993 102 1027 136
rect 1079 176 1113 210
rect 1079 86 1113 120
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 129 546 163 580
rect 129 463 163 497
rect 129 380 163 414
rect 219 546 253 580
rect 219 474 253 508
rect 309 546 343 580
rect 309 476 343 510
rect 309 406 343 440
rect 399 544 433 578
rect 489 385 523 419
rect 596 544 630 578
rect 708 546 742 580
rect 708 474 742 508
rect 808 497 842 531
rect 808 406 842 440
rect 898 546 932 580
rect 898 474 932 508
rect 988 497 1022 531
rect 988 406 1022 440
rect 1078 546 1112 580
rect 1078 476 1112 510
rect 1078 406 1112 440
<< poly >>
rect 83 592 119 618
rect 173 592 209 618
rect 263 592 299 618
rect 353 592 389 618
rect 443 592 479 618
rect 533 592 569 618
rect 752 592 788 618
rect 852 592 888 618
rect 942 592 978 618
rect 1032 592 1068 618
rect 83 330 119 368
rect 173 330 209 368
rect 263 330 299 368
rect 353 330 389 368
rect 83 314 389 330
rect 83 280 105 314
rect 139 280 173 314
rect 207 280 241 314
rect 275 280 309 314
rect 343 280 389 314
rect 443 310 479 368
rect 533 310 569 368
rect 752 345 788 368
rect 852 345 888 368
rect 942 345 978 368
rect 1032 345 1068 368
rect 752 320 1068 345
rect 752 315 809 320
rect 83 264 389 280
rect 431 294 633 310
rect 84 222 114 264
rect 170 222 200 264
rect 256 222 286 264
rect 345 222 375 264
rect 431 260 447 294
rect 481 260 515 294
rect 549 260 583 294
rect 617 267 633 294
rect 780 286 809 315
rect 843 286 877 320
rect 911 286 945 320
rect 979 286 1013 320
rect 1047 286 1068 320
rect 780 270 1068 286
rect 617 260 719 267
rect 431 237 719 260
rect 431 222 461 237
rect 517 222 547 237
rect 603 222 633 237
rect 689 222 719 237
rect 780 222 810 270
rect 866 222 896 270
rect 952 222 982 270
rect 1038 222 1068 270
rect 84 48 114 74
rect 170 48 200 74
rect 256 48 286 74
rect 345 48 375 74
rect 431 48 461 74
rect 517 48 547 74
rect 603 48 633 74
rect 689 48 719 74
rect 780 48 810 74
rect 866 48 896 74
rect 952 48 982 74
rect 1038 48 1068 74
<< polycont >>
rect 105 280 139 314
rect 173 280 207 314
rect 241 280 275 314
rect 309 280 343 314
rect 447 260 481 294
rect 515 260 549 294
rect 583 260 617 294
rect 809 286 843 320
rect 877 286 911 320
rect 945 286 979 320
rect 1013 286 1047 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 23 580 73 649
rect 23 546 39 580
rect 23 497 73 546
rect 23 463 39 497
rect 23 414 73 463
rect 23 380 39 414
rect 23 364 73 380
rect 113 580 179 596
rect 113 546 129 580
rect 163 546 179 580
rect 113 497 179 546
rect 113 463 129 497
rect 163 463 179 497
rect 113 424 179 463
rect 219 580 253 649
rect 219 508 253 546
rect 219 458 253 474
rect 293 580 359 596
rect 293 546 309 580
rect 343 546 359 580
rect 293 510 359 546
rect 399 578 449 649
rect 433 544 449 578
rect 399 526 449 544
rect 580 578 646 649
rect 580 544 596 578
rect 630 544 646 578
rect 580 526 646 544
rect 692 581 1128 615
rect 692 580 758 581
rect 692 546 708 580
rect 742 546 758 580
rect 898 580 932 581
rect 293 476 309 510
rect 343 492 359 510
rect 692 508 758 546
rect 692 492 708 508
rect 343 476 708 492
rect 293 474 708 476
rect 742 474 758 508
rect 293 458 758 474
rect 792 531 858 547
rect 792 497 808 531
rect 842 497 858 531
rect 293 440 359 458
rect 293 424 309 440
rect 113 414 309 424
rect 113 380 129 414
rect 163 406 309 414
rect 343 406 359 440
rect 792 440 858 497
rect 1078 580 1128 581
rect 898 508 932 546
rect 898 458 932 474
rect 972 531 1038 547
rect 972 497 988 531
rect 1022 497 1038 531
rect 792 424 808 440
rect 163 390 359 406
rect 473 419 808 424
rect 163 380 179 390
rect 113 364 179 380
rect 473 385 489 419
rect 523 406 808 419
rect 842 424 858 440
rect 972 440 1038 497
rect 972 424 988 440
rect 842 406 988 424
rect 1022 406 1038 440
rect 523 390 1038 406
rect 1112 546 1128 580
rect 1078 510 1128 546
rect 1112 476 1128 510
rect 1078 440 1128 476
rect 1112 406 1128 440
rect 1078 390 1128 406
rect 523 385 743 390
rect 473 364 743 385
rect 217 330 359 356
rect 89 314 359 330
rect 89 280 105 314
rect 139 280 173 314
rect 207 280 241 314
rect 275 280 309 314
rect 343 280 359 314
rect 667 310 743 364
rect 793 320 1127 356
rect 89 264 359 280
rect 409 294 633 310
rect 409 260 447 294
rect 481 260 515 294
rect 549 260 583 294
rect 617 260 633 294
rect 409 236 633 260
rect 23 210 245 230
rect 23 176 39 210
rect 73 196 211 210
rect 23 120 73 176
rect 667 202 701 310
rect 793 286 809 320
rect 843 286 877 320
rect 911 286 945 320
rect 979 286 1013 320
rect 1047 286 1127 320
rect 793 270 1127 286
rect 245 186 420 202
rect 245 176 386 186
rect 211 168 386 176
rect 23 86 39 120
rect 23 70 73 86
rect 109 141 175 162
rect 109 107 125 141
rect 159 107 175 141
rect 109 17 175 107
rect 211 120 245 168
rect 211 70 245 86
rect 281 127 347 134
rect 281 93 297 127
rect 331 93 347 127
rect 281 17 347 93
rect 386 116 420 152
rect 456 177 701 202
rect 456 143 472 177
rect 506 168 644 177
rect 456 119 506 143
rect 678 143 701 177
rect 542 127 608 134
rect 542 93 558 127
rect 592 93 608 127
rect 644 119 701 143
rect 735 210 1129 236
rect 769 202 907 210
rect 735 120 769 176
rect 941 202 1079 210
rect 542 85 608 93
rect 735 85 769 86
rect 420 82 769 85
rect 386 51 769 82
rect 805 136 871 168
rect 805 102 821 136
rect 855 102 871 136
rect 805 17 871 102
rect 907 120 941 176
rect 1113 176 1129 210
rect 907 70 941 86
rect 977 136 1043 168
rect 977 102 993 136
rect 1027 102 1043 136
rect 977 17 1043 102
rect 1079 120 1129 176
rect 1113 86 1129 120
rect 1079 70 1129 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
rlabel comment s 0 0 0 0 4 o21ai_4
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 415 242 449 276 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 511 242 545 276 0 FreeSans 340 0 0 0 B1
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 1152 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1080240
string GDS_START 1070500
<< end >>
