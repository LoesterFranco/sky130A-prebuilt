magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1564 561
rect 103 427 169 527
rect 18 197 66 325
rect 290 439 363 527
rect 667 435 739 527
rect 103 17 169 93
rect 859 402 916 527
rect 1115 367 1168 527
rect 1208 401 1274 491
rect 1308 435 1360 527
rect 1394 401 1460 493
rect 1208 367 1460 401
rect 1317 357 1460 367
rect 306 153 390 203
rect 1046 211 1148 265
rect 1350 177 1460 357
rect 1494 297 1547 527
rect 290 17 357 93
rect 663 17 730 106
rect 1258 143 1460 177
rect 859 17 916 143
rect 1258 109 1292 143
rect 1118 17 1174 109
rect 1208 51 1292 109
rect 1326 17 1360 109
rect 1394 51 1460 143
rect 1494 17 1547 177
rect 0 -17 1564 17
<< obsli1 >>
rect 17 393 69 493
rect 17 391 156 393
rect 17 359 122 391
rect 122 280 156 357
rect 203 317 248 493
rect 495 439 633 485
rect 583 421 633 439
rect 583 418 636 421
rect 583 412 637 418
rect 305 391 547 405
rect 596 403 637 412
rect 339 381 547 391
rect 339 371 569 381
rect 409 317 467 337
rect 122 214 168 280
rect 203 271 467 317
rect 501 315 569 371
rect 122 161 156 214
rect 17 127 156 161
rect 17 69 69 127
rect 203 69 256 271
rect 513 207 547 315
rect 603 265 637 403
rect 779 373 823 487
rect 671 307 823 373
rect 789 265 823 307
rect 950 333 1007 493
rect 950 299 1228 333
rect 603 233 755 265
rect 458 141 547 207
rect 581 199 755 233
rect 789 199 944 265
rect 581 107 615 199
rect 789 149 823 199
rect 978 177 1012 299
rect 1182 258 1228 299
rect 1182 211 1316 258
rect 1182 177 1224 211
rect 978 165 1224 177
rect 483 73 615 107
rect 779 83 823 149
rect 950 143 1224 165
rect 950 58 1012 143
<< obsli1c >>
rect 122 357 156 391
rect 305 357 339 391
<< metal1 >>
rect 0 496 1564 592
rect 18 252 76 261
rect 1034 252 1092 261
rect 18 224 1092 252
rect 18 215 76 224
rect 1034 215 1092 224
rect 0 -48 1564 48
<< obsm1 >>
rect 110 391 168 397
rect 110 357 122 391
rect 156 388 168 391
rect 293 391 351 397
rect 293 388 305 391
rect 156 360 305 388
rect 156 357 168 360
rect 110 351 168 357
rect 293 357 305 360
rect 339 357 351 391
rect 293 351 351 357
<< labels >>
rlabel locali s 306 153 390 203 6 GATE
port 1 nsew signal input
rlabel locali s 1394 401 1460 493 6 GCLK
port 2 nsew signal output
rlabel locali s 1394 51 1460 143 6 GCLK
port 2 nsew signal output
rlabel locali s 1350 177 1460 357 6 GCLK
port 2 nsew signal output
rlabel locali s 1317 357 1460 367 6 GCLK
port 2 nsew signal output
rlabel locali s 1258 143 1460 177 6 GCLK
port 2 nsew signal output
rlabel locali s 1258 109 1292 143 6 GCLK
port 2 nsew signal output
rlabel locali s 1208 401 1274 491 6 GCLK
port 2 nsew signal output
rlabel locali s 1208 367 1460 401 6 GCLK
port 2 nsew signal output
rlabel locali s 1208 51 1292 109 6 GCLK
port 2 nsew signal output
rlabel locali s 18 197 66 325 6 CLK
port 3 nsew clock input
rlabel locali s 1046 211 1148 265 6 CLK
port 3 nsew clock input
rlabel metal1 s 1034 252 1092 261 6 CLK
port 3 nsew clock input
rlabel metal1 s 1034 215 1092 224 6 CLK
port 3 nsew clock input
rlabel metal1 s 18 252 76 261 6 CLK
port 3 nsew clock input
rlabel metal1 s 18 224 1092 252 6 CLK
port 3 nsew clock input
rlabel metal1 s 18 215 76 224 6 CLK
port 3 nsew clock input
rlabel locali s 1494 17 1547 177 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 1326 17 1360 109 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 1118 17 1174 109 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 859 17 916 143 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 663 17 730 106 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 290 17 357 93 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 103 17 169 93 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 1564 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1564 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 1494 297 1547 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 1308 435 1360 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 1115 367 1168 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 859 402 916 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 667 435 739 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 290 439 363 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 103 427 169 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 1564 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 1564 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1564 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2598802
string GDS_START 2586004
<< end >>
