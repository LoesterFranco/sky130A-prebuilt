magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 28 195 98 325
rect 317 267 444 349
rect 317 214 398 267
rect 624 271 731 493
rect 922 142 991 340
rect 2484 53 2557 465
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2576 561
rect 18 393 69 493
rect 106 427 182 527
rect 18 391 183 393
rect 18 359 145 391
rect 142 357 145 359
rect 179 357 183 391
rect 142 265 183 357
rect 227 346 273 493
rect 422 417 476 480
rect 520 451 586 527
rect 422 383 546 417
rect 142 199 205 265
rect 239 255 273 346
rect 142 161 177 199
rect 19 127 177 161
rect 239 135 273 221
rect 495 237 546 383
rect 774 421 808 493
rect 971 455 1041 527
rect 1096 437 1170 487
rect 1096 421 1130 437
rect 1219 427 1292 493
rect 774 387 1130 421
rect 495 233 689 237
rect 453 199 689 233
rect 774 215 809 387
rect 453 180 487 199
rect 19 69 69 127
rect 103 17 179 93
rect 223 69 273 135
rect 339 146 487 180
rect 339 79 373 146
rect 407 17 483 112
rect 531 17 607 165
rect 655 85 689 199
rect 733 135 809 215
rect 853 85 887 337
rect 1028 179 1062 387
rect 1164 357 1190 391
rect 1164 315 1224 357
rect 1096 255 1130 279
rect 1096 213 1130 221
rect 1180 207 1224 315
rect 1258 277 1292 427
rect 1336 421 1370 475
rect 1427 471 1493 527
rect 1554 421 1588 475
rect 1630 435 1714 527
rect 1336 387 1588 421
rect 1763 401 1797 493
rect 1839 425 2043 493
rect 2083 439 2133 527
rect 1646 367 1797 401
rect 1646 353 1708 367
rect 1392 319 1708 353
rect 1837 357 1913 391
rect 1947 357 1969 391
rect 1837 333 1969 357
rect 1258 243 1630 277
rect 1028 143 1144 179
rect 655 51 887 85
rect 1001 17 1070 108
rect 1110 101 1144 143
rect 1180 141 1330 207
rect 1110 67 1178 101
rect 1368 95 1402 243
rect 1446 187 1562 209
rect 1596 201 1630 243
rect 1446 153 1451 187
rect 1485 153 1523 187
rect 1557 153 1562 187
rect 1674 167 1708 319
rect 1222 61 1402 95
rect 1538 17 1604 109
rect 1646 89 1708 167
rect 1742 332 1969 333
rect 2008 349 2043 425
rect 2182 417 2216 475
rect 2251 451 2327 527
rect 2182 383 2346 417
rect 1742 299 1889 332
rect 2008 315 2274 349
rect 1742 141 1794 299
rect 2008 297 2057 315
rect 1847 255 1881 265
rect 1847 184 1881 221
rect 1934 263 2057 297
rect 2312 265 2346 383
rect 2381 299 2438 527
rect 1934 107 1978 263
rect 2030 173 2074 229
rect 2120 213 2274 255
rect 2213 187 2274 213
rect 2030 139 2146 173
rect 1646 55 1722 89
rect 1756 51 1978 107
rect 2022 17 2066 105
rect 2112 93 2146 139
rect 2213 153 2235 187
rect 2269 153 2274 187
rect 2213 127 2274 153
rect 2312 199 2441 265
rect 2312 93 2347 199
rect 2112 59 2347 93
rect 2381 17 2438 142
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2576 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 145 357 179 391
rect 239 221 273 255
rect 1190 357 1224 391
rect 1096 221 1130 255
rect 1913 357 1947 391
rect 1451 153 1485 187
rect 1523 153 1557 187
rect 1847 221 1881 255
rect 2235 153 2269 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
<< metal1 >>
rect 0 561 2576 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2576 561
rect 0 496 2576 527
rect 1429 187 1580 193
rect 1429 153 1451 187
rect 1485 153 1523 187
rect 1557 184 1580 187
rect 2223 187 2281 193
rect 2223 184 2235 187
rect 1557 156 2235 184
rect 1557 153 1580 156
rect 1429 147 1580 153
rect 2223 153 2235 156
rect 2269 153 2281 187
rect 2223 147 2281 153
rect 0 17 2576 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2576 17
rect 0 -48 2576 -17
<< obsm1 >>
rect 132 391 192 397
rect 132 357 145 391
rect 179 388 192 391
rect 1178 391 1236 397
rect 1178 388 1190 391
rect 179 360 1190 388
rect 179 357 192 360
rect 132 351 192 357
rect 1178 357 1190 360
rect 1224 388 1236 391
rect 1900 391 1959 397
rect 1900 388 1913 391
rect 1224 360 1913 388
rect 1224 357 1236 360
rect 1178 351 1236 357
rect 1900 357 1913 360
rect 1947 357 1959 391
rect 1900 351 1959 357
rect 227 255 285 261
rect 227 221 239 255
rect 273 252 285 255
rect 1084 255 1142 261
rect 1084 252 1096 255
rect 273 224 1096 252
rect 273 221 285 224
rect 227 215 285 221
rect 1084 221 1096 224
rect 1130 252 1142 255
rect 1831 255 1893 261
rect 1831 252 1847 255
rect 1130 224 1847 252
rect 1130 221 1142 224
rect 1084 215 1142 221
rect 1831 221 1847 224
rect 1881 221 1893 255
rect 1831 215 1893 221
<< labels >>
rlabel locali s 28 195 98 325 6 CLK_N
port 1 nsew signal input
rlabel locali s 624 271 731 493 6 D
port 2 nsew signal input
rlabel locali s 2484 53 2557 465 6 Q
port 3 nsew signal output
rlabel metal1 s 2223 184 2281 193 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 2223 147 2281 156 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 1429 184 1580 193 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 1429 156 2281 184 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 1429 147 1580 156 6 RESET_B
port 4 nsew signal input
rlabel locali s 922 142 991 340 6 SCD
port 5 nsew signal input
rlabel locali s 317 267 444 349 6 SCE
port 6 nsew signal input
rlabel locali s 317 214 398 267 6 SCE
port 6 nsew signal input
rlabel metal1 s 0 -48 2576 48 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 496 2576 592 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2576 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 82818
string GDS_START 64726
<< end >>
