magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 29 299 426 335
rect 29 207 139 299
rect 179 199 315 265
rect 351 215 426 299
rect 503 266 573 423
rect 482 157 573 266
rect 607 199 707 325
rect 201 123 573 157
rect 201 51 280 123
rect 509 51 573 123
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 22 421 74 493
rect 108 455 184 527
rect 230 421 264 493
rect 325 439 359 527
rect 403 457 678 493
rect 22 405 264 421
rect 403 405 469 457
rect 22 371 469 405
rect 617 359 678 457
rect 20 17 79 173
rect 382 17 458 89
rect 619 17 685 165
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel locali s 179 199 315 265 6 A1
port 1 nsew signal input
rlabel locali s 351 215 426 299 6 A2
port 2 nsew signal input
rlabel locali s 29 299 426 335 6 A2
port 2 nsew signal input
rlabel locali s 29 207 139 299 6 A2
port 2 nsew signal input
rlabel locali s 607 199 707 325 6 B1
port 3 nsew signal input
rlabel locali s 509 51 573 123 6 Y
port 4 nsew signal output
rlabel locali s 503 266 573 423 6 Y
port 4 nsew signal output
rlabel locali s 482 157 573 266 6 Y
port 4 nsew signal output
rlabel locali s 201 123 573 157 6 Y
port 4 nsew signal output
rlabel locali s 201 51 280 123 6 Y
port 4 nsew signal output
rlabel metal1 s 0 -48 736 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 736 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1205780
string GDS_START 1199644
<< end >>
