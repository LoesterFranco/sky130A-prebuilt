magic
tech sky130A
magscale 1 2
timestamp 1604502697
<< nwell >>
rect -38 261 1510 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 89 47 119 131
rect 174 47 204 131
rect 269 47 299 119
rect 385 47 415 119
rect 516 47 546 131
rect 635 47 665 177
rect 823 47 853 131
rect 943 47 973 131
rect 1151 47 1181 131
rect 1247 47 1277 131
rect 1352 47 1382 177
<< pmoshvt >>
rect 81 369 117 497
rect 163 369 199 497
rect 268 413 304 497
rect 374 413 410 497
rect 486 413 522 497
rect 627 297 663 497
rect 825 303 861 431
rect 945 303 981 431
rect 1143 369 1179 497
rect 1239 369 1275 497
rect 1344 297 1380 497
<< ndiff >>
rect 27 103 89 131
rect 27 69 35 103
rect 69 69 89 103
rect 27 47 89 69
rect 119 89 174 131
rect 119 55 129 89
rect 163 55 174 89
rect 119 47 174 55
rect 204 119 254 131
rect 570 131 635 177
rect 466 119 516 131
rect 204 101 269 119
rect 204 67 223 101
rect 257 67 269 101
rect 204 47 269 67
rect 299 89 385 119
rect 299 55 329 89
rect 363 55 385 89
rect 299 47 385 55
rect 415 47 516 119
rect 546 119 635 131
rect 546 85 582 119
rect 616 85 635 119
rect 546 47 635 85
rect 665 101 717 177
rect 1292 131 1352 177
rect 665 67 675 101
rect 709 67 717 101
rect 665 47 717 67
rect 771 110 823 131
rect 771 76 779 110
rect 813 76 823 110
rect 771 47 823 76
rect 853 89 943 131
rect 853 55 873 89
rect 907 55 943 89
rect 853 47 943 55
rect 973 110 1035 131
rect 973 76 993 110
rect 1027 76 1035 110
rect 973 47 1035 76
rect 1089 109 1151 131
rect 1089 75 1107 109
rect 1141 75 1151 109
rect 1089 47 1151 75
rect 1181 47 1247 131
rect 1277 89 1352 131
rect 1277 55 1287 89
rect 1321 55 1352 89
rect 1277 47 1352 55
rect 1382 145 1439 177
rect 1382 111 1397 145
rect 1431 111 1439 145
rect 1382 47 1439 111
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 369 81 383
rect 117 369 163 497
rect 199 475 268 497
rect 199 441 222 475
rect 256 441 268 475
rect 199 413 268 441
rect 304 475 374 497
rect 304 441 322 475
rect 356 441 374 475
rect 304 413 374 441
rect 410 413 486 497
rect 522 489 627 497
rect 522 455 560 489
rect 594 455 627 489
rect 522 413 627 455
rect 199 369 251 413
rect 575 297 627 413
rect 663 458 717 497
rect 663 424 675 458
rect 709 424 717 458
rect 878 485 928 497
rect 878 451 886 485
rect 920 451 928 485
rect 1089 485 1143 497
rect 878 431 928 451
rect 1089 451 1097 485
rect 1131 451 1143 485
rect 663 297 717 424
rect 771 349 825 431
rect 771 315 779 349
rect 813 315 825 349
rect 771 303 825 315
rect 861 303 945 431
rect 981 349 1035 431
rect 1089 369 1143 451
rect 1179 442 1239 497
rect 1179 408 1191 442
rect 1225 408 1239 442
rect 1179 369 1239 408
rect 1275 489 1344 497
rect 1275 455 1293 489
rect 1327 455 1344 489
rect 1275 369 1344 455
rect 981 315 993 349
rect 1027 315 1035 349
rect 981 303 1035 315
rect 1292 297 1344 369
rect 1380 448 1439 497
rect 1380 414 1397 448
rect 1431 414 1439 448
rect 1380 380 1439 414
rect 1380 346 1397 380
rect 1431 346 1439 380
rect 1380 297 1439 346
<< ndiffc >>
rect 35 69 69 103
rect 129 55 163 89
rect 223 67 257 101
rect 329 55 363 89
rect 582 85 616 119
rect 675 67 709 101
rect 779 76 813 110
rect 873 55 907 89
rect 993 76 1027 110
rect 1107 75 1141 109
rect 1287 55 1321 89
rect 1397 111 1431 145
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 222 441 256 475
rect 322 441 356 475
rect 560 455 594 489
rect 675 424 709 458
rect 886 451 920 485
rect 1097 451 1131 485
rect 779 315 813 349
rect 1191 408 1225 442
rect 1293 455 1327 489
rect 993 315 1027 349
rect 1397 414 1431 448
rect 1397 346 1431 380
<< poly >>
rect 81 497 117 523
rect 163 497 199 523
rect 268 497 304 523
rect 374 497 410 523
rect 486 497 522 523
rect 627 497 663 523
rect 268 398 304 413
rect 374 398 410 413
rect 486 398 522 413
rect 81 354 117 369
rect 163 354 199 369
rect 79 265 119 354
rect 22 249 119 265
rect 22 215 32 249
rect 66 215 119 249
rect 22 199 119 215
rect 161 265 201 354
rect 266 273 306 398
rect 372 381 412 398
rect 348 365 412 381
rect 348 331 358 365
rect 392 331 412 365
rect 348 315 412 331
rect 484 381 524 398
rect 484 365 546 381
rect 484 331 494 365
rect 528 331 546 365
rect 484 315 546 331
rect 161 249 222 265
rect 161 215 171 249
rect 205 215 222 249
rect 266 243 424 273
rect 161 199 222 215
rect 385 207 424 243
rect 89 131 119 199
rect 174 131 204 199
rect 269 191 343 201
rect 269 157 293 191
rect 327 157 343 191
rect 269 147 343 157
rect 385 191 439 207
rect 385 157 395 191
rect 429 157 439 191
rect 269 119 299 147
rect 385 141 439 157
rect 385 119 415 141
rect 516 131 546 315
rect 823 457 863 523
rect 825 431 861 457
rect 943 457 983 523
rect 1143 497 1179 523
rect 1239 497 1275 523
rect 1344 497 1380 523
rect 945 431 981 457
rect 1143 354 1179 369
rect 1239 354 1275 369
rect 627 282 663 297
rect 825 288 861 303
rect 945 288 981 303
rect 625 265 665 282
rect 597 249 665 265
rect 597 215 607 249
rect 641 215 665 249
rect 597 199 665 215
rect 635 177 665 199
rect 823 265 863 288
rect 943 265 983 288
rect 1141 265 1181 354
rect 1237 265 1277 354
rect 1344 282 1380 297
rect 1342 265 1382 282
rect 823 255 889 265
rect 823 221 839 255
rect 873 221 889 255
rect 823 199 889 221
rect 943 249 1012 265
rect 943 215 968 249
rect 1002 215 1012 249
rect 943 199 1012 215
rect 1095 249 1181 265
rect 1095 215 1105 249
rect 1139 215 1181 249
rect 1095 199 1181 215
rect 1223 249 1277 265
rect 1223 215 1233 249
rect 1267 215 1277 249
rect 1223 199 1277 215
rect 1319 249 1382 265
rect 1319 215 1329 249
rect 1363 215 1382 249
rect 1319 199 1382 215
rect 823 131 853 199
rect 943 131 973 199
rect 1151 131 1181 199
rect 1247 131 1277 199
rect 1352 177 1382 199
rect 89 21 119 47
rect 174 21 204 47
rect 269 21 299 47
rect 385 21 415 47
rect 516 21 546 47
rect 635 21 665 47
rect 823 21 853 47
rect 943 21 973 47
rect 1151 21 1181 47
rect 1247 21 1277 47
rect 1352 21 1382 47
<< polycont >>
rect 32 215 66 249
rect 358 331 392 365
rect 494 331 528 365
rect 171 215 205 249
rect 293 157 327 191
rect 395 157 429 191
rect 607 215 641 249
rect 839 221 873 255
rect 968 215 1002 249
rect 1105 215 1139 249
rect 1233 215 1267 249
rect 1329 215 1363 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 17 485 69 527
rect 17 451 35 485
rect 17 417 69 451
rect 17 383 35 417
rect 17 367 69 383
rect 103 475 256 493
rect 103 441 222 475
rect 103 425 256 441
rect 322 475 460 493
rect 356 441 460 475
rect 322 425 460 441
rect 17 249 66 333
rect 17 215 32 249
rect 17 191 66 215
rect 103 157 137 425
rect 171 249 247 391
rect 205 215 247 249
rect 171 191 247 215
rect 293 365 392 391
rect 293 331 358 365
rect 293 323 392 331
rect 293 289 325 323
rect 359 289 392 323
rect 293 241 392 289
rect 426 275 460 425
rect 504 489 621 527
rect 504 455 560 489
rect 594 455 621 489
rect 504 415 621 455
rect 665 458 709 493
rect 665 424 675 458
rect 777 485 1147 527
rect 777 451 886 485
rect 920 451 1097 485
rect 1131 451 1147 485
rect 665 417 709 424
rect 1191 442 1225 493
rect 1277 489 1343 527
rect 1277 455 1293 489
rect 1327 455 1343 489
rect 1277 451 1343 455
rect 665 383 1147 417
rect 665 381 709 383
rect 494 365 709 381
rect 528 331 709 365
rect 494 327 709 331
rect 494 315 533 327
rect 426 249 641 275
rect 426 241 607 249
rect 293 191 360 241
rect 495 215 607 241
rect 327 157 360 191
rect 17 123 259 157
rect 293 141 360 157
rect 394 191 461 207
rect 394 157 395 191
rect 429 187 461 191
rect 394 153 427 157
rect 394 141 461 153
rect 495 199 641 215
rect 17 103 69 123
rect 17 69 35 103
rect 223 101 259 123
rect 495 107 529 199
rect 17 51 69 69
rect 103 55 129 89
rect 163 55 179 89
rect 103 17 179 55
rect 257 67 259 101
rect 223 51 259 67
rect 293 89 529 107
rect 293 55 329 89
rect 363 55 529 89
rect 293 51 529 55
rect 582 119 616 165
rect 582 17 616 85
rect 675 101 709 327
rect 675 51 709 67
rect 747 315 779 349
rect 813 315 829 349
rect 873 323 993 349
rect 747 187 781 315
rect 907 315 993 323
rect 1027 315 1043 349
rect 907 299 1043 315
rect 907 289 910 299
rect 815 221 839 255
rect 873 221 910 289
rect 747 153 760 187
rect 794 153 813 187
rect 747 110 813 153
rect 876 157 910 221
rect 949 255 1012 265
rect 949 221 961 255
rect 995 249 1012 255
rect 949 215 968 221
rect 1002 215 1012 249
rect 949 199 1012 215
rect 1077 249 1147 383
rect 1397 448 1447 493
rect 1225 408 1363 417
rect 1191 299 1363 408
rect 1077 215 1105 249
rect 1139 215 1147 249
rect 1077 199 1147 215
rect 1191 255 1279 265
rect 1191 221 1200 255
rect 1234 249 1279 255
rect 1191 215 1233 221
rect 1267 215 1279 249
rect 1191 199 1279 215
rect 1329 249 1363 299
rect 1329 157 1363 215
rect 876 123 1043 157
rect 747 76 779 110
rect 993 110 1043 123
rect 747 51 813 76
rect 857 55 873 89
rect 907 55 923 89
rect 857 17 923 55
rect 1027 76 1043 110
rect 993 51 1043 76
rect 1107 123 1363 157
rect 1431 414 1447 448
rect 1397 380 1447 414
rect 1431 346 1447 380
rect 1397 145 1447 346
rect 1107 109 1141 123
rect 1431 111 1447 145
rect 1107 51 1141 75
rect 1265 55 1287 89
rect 1321 55 1337 89
rect 1265 17 1337 55
rect 1397 51 1447 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 325 289 359 323
rect 427 157 429 187
rect 429 157 461 187
rect 427 153 461 157
rect 873 289 907 323
rect 760 153 794 187
rect 961 249 995 255
rect 961 221 968 249
rect 968 221 995 249
rect 1200 249 1234 255
rect 1200 221 1233 249
rect 1233 221 1234 249
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 313 323 371 329
rect 313 289 325 323
rect 359 320 371 323
rect 861 323 919 329
rect 861 320 873 323
rect 359 292 873 320
rect 359 289 371 292
rect 313 283 371 289
rect 861 289 873 292
rect 907 289 919 323
rect 861 283 919 289
rect 949 255 1007 261
rect 949 221 961 255
rect 995 252 1007 255
rect 1188 255 1246 261
rect 1188 252 1200 255
rect 995 224 1200 252
rect 995 221 1007 224
rect 949 215 1007 221
rect 1188 221 1200 224
rect 1234 221 1246 255
rect 1188 215 1246 221
rect 415 187 473 193
rect 415 153 427 187
rect 461 184 473 187
rect 748 187 806 193
rect 748 184 760 187
rect 461 156 760 184
rect 461 153 473 156
rect 415 147 473 153
rect 748 153 760 156
rect 794 153 806 187
rect 748 147 806 153
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< labels >>
rlabel comment s 0 0 0 0 4 sdlclkp_2
flabel metal1 s 949 221 983 255 0 FreeSans 200 0 0 0 CLK
port 1 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
flabel corelocali s 30 289 64 323 0 FreeSans 200 0 0 0 SCE
port 3 nsew
flabel corelocali s 1409 425 1443 459 0 FreeSans 200 0 0 0 GCLK
port 8 nsew
flabel corelocali s 1409 357 1443 391 0 FreeSans 200 0 0 0 GCLK
port 8 nsew
flabel corelocali s 213 357 247 391 0 FreeSans 200 0 0 0 GATE
port 2 nsew
flabel corelocali s 1409 85 1443 119 0 FreeSans 200 0 0 0 GCLK
port 8 nsew
flabel corelocali s 213 289 247 323 0 FreeSans 200 0 0 0 GATE
port 2 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 200 0 0 0 SCE
port 3 nsew
flabel corelocali s 1409 221 1443 255 0 FreeSans 200 0 0 0 GCLK
port 8 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 1472 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 381274
string GDS_START 369770
<< end >>
