magic
tech sky130A
magscale 1 2
timestamp 1601050088
<< locali >>
rect 17 364 71 596
rect 17 226 51 364
rect 17 70 73 226
rect 177 244 243 308
rect 209 218 243 244
rect 660 218 726 291
rect 876 221 942 291
rect 1162 264 1242 315
rect 1162 221 1196 264
rect 1360 264 1494 356
rect 876 218 1196 221
rect 209 187 1196 218
rect 1657 226 1708 596
rect 209 184 942 187
rect 1642 70 1708 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 111 410 177 649
rect 416 424 482 551
rect 211 390 482 424
rect 522 492 572 551
rect 616 526 682 649
rect 720 492 786 551
rect 522 458 786 492
rect 821 461 887 649
rect 522 393 572 458
rect 1014 424 1099 551
rect 211 376 245 390
rect 107 342 245 376
rect 313 350 359 356
rect 107 326 141 342
rect 85 260 141 326
rect 313 316 319 350
rect 353 316 359 350
rect 416 349 482 390
rect 606 390 1099 424
rect 1133 451 1190 551
rect 1224 500 1365 649
rect 1400 451 1464 566
rect 1133 417 1464 451
rect 1398 390 1464 417
rect 606 359 640 390
rect 313 315 359 316
rect 516 325 640 359
rect 1065 383 1099 390
rect 768 350 839 356
rect 516 315 550 325
rect 107 150 141 260
rect 313 252 423 315
rect 465 252 550 315
rect 768 316 799 350
rect 833 316 839 350
rect 768 252 839 316
rect 985 350 1031 356
rect 985 316 991 350
rect 1025 316 1031 350
rect 1065 349 1310 383
rect 1551 364 1617 649
rect 985 315 1031 316
rect 985 255 1128 315
rect 1276 230 1310 349
rect 1542 230 1608 310
rect 1230 196 1608 230
rect 1230 153 1264 196
rect 107 116 454 150
rect 125 17 196 82
rect 388 71 454 116
rect 496 116 782 150
rect 496 84 578 116
rect 716 84 782 116
rect 614 17 680 82
rect 816 17 911 142
rect 1009 119 1264 153
rect 1298 128 1518 162
rect 1009 87 1075 119
rect 1298 85 1332 128
rect 1452 96 1518 128
rect 1111 51 1332 85
rect 1366 17 1416 94
rect 1556 17 1606 154
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 319 316 353 350
rect 799 316 833 350
rect 991 316 1025 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
<< metal1 >>
rect 0 683 1728 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 0 617 1728 649
rect 307 350 365 356
rect 307 316 319 350
rect 353 347 365 350
rect 787 350 845 356
rect 787 347 799 350
rect 353 319 799 347
rect 353 316 365 319
rect 307 310 365 316
rect 787 316 799 319
rect 833 347 845 350
rect 979 350 1037 356
rect 979 347 991 350
rect 833 319 991 347
rect 833 316 845 319
rect 787 310 845 316
rect 979 316 991 319
rect 1025 316 1037 350
rect 979 310 1037 316
rect 0 17 1728 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
rect 0 -49 1728 -17
<< labels >>
rlabel locali s 1162 264 1242 315 6 A
port 1 nsew signal input
rlabel locali s 1162 221 1196 264 6 A
port 1 nsew signal input
rlabel locali s 876 221 942 291 6 A
port 1 nsew signal input
rlabel locali s 876 218 1196 221 6 A
port 1 nsew signal input
rlabel locali s 660 218 726 291 6 A
port 1 nsew signal input
rlabel locali s 209 218 243 244 6 A
port 1 nsew signal input
rlabel locali s 209 187 1196 218 6 A
port 1 nsew signal input
rlabel locali s 209 184 942 187 6 A
port 1 nsew signal input
rlabel locali s 177 244 243 308 6 A
port 1 nsew signal input
rlabel locali s 1360 264 1494 356 6 B
port 2 nsew signal input
rlabel metal1 s 979 347 1037 356 6 CIN
port 3 nsew signal input
rlabel metal1 s 979 310 1037 319 6 CIN
port 3 nsew signal input
rlabel metal1 s 787 347 845 356 6 CIN
port 3 nsew signal input
rlabel metal1 s 787 310 845 319 6 CIN
port 3 nsew signal input
rlabel metal1 s 307 347 365 356 6 CIN
port 3 nsew signal input
rlabel metal1 s 307 319 1037 347 6 CIN
port 3 nsew signal input
rlabel metal1 s 307 310 365 319 6 CIN
port 3 nsew signal input
rlabel locali s 1657 226 1708 596 6 COUT
port 4 nsew signal output
rlabel locali s 1642 70 1708 226 6 COUT
port 4 nsew signal output
rlabel locali s 17 364 71 596 6 SUM
port 5 nsew signal output
rlabel locali s 17 226 51 364 6 SUM
port 5 nsew signal output
rlabel locali s 17 70 73 226 6 SUM
port 5 nsew signal output
rlabel metal1 s 0 -49 1728 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 1728 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1728 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 2402036
string GDS_START 2388574
<< end >>
