magic
tech sky130A
magscale 1 2
timestamp 1599588244
<< locali >>
rect 167 394 233 596
rect 347 394 413 596
rect 25 360 413 394
rect 25 226 130 360
rect 25 192 489 226
rect 677 252 743 356
rect 793 290 1031 356
rect 1081 290 1223 356
rect 1257 290 1415 356
rect 1449 252 1607 356
rect 283 70 333 192
rect 439 70 489 192
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 77 428 127 649
rect 273 428 307 649
rect 453 364 503 649
rect 541 581 967 615
rect 541 458 607 581
rect 647 424 681 547
rect 609 390 681 424
rect 721 390 787 581
rect 827 424 861 547
rect 901 458 967 581
rect 1005 581 1235 615
rect 1005 458 1061 581
rect 1095 424 1161 547
rect 827 390 1161 424
rect 1201 424 1235 581
rect 1275 458 1341 649
rect 1381 424 1415 596
rect 1455 458 1505 649
rect 1545 424 1611 596
rect 1201 390 1611 424
rect 609 326 643 390
rect 174 260 643 326
rect 609 218 643 260
rect 810 222 1354 256
rect 810 218 844 222
rect 181 17 247 158
rect 369 17 403 158
rect 525 17 575 206
rect 609 184 844 218
rect 609 70 670 184
rect 706 17 774 150
rect 810 70 844 184
rect 880 17 948 188
rect 984 70 1018 222
rect 1054 17 1120 188
rect 1202 91 1268 188
rect 1302 125 1354 222
rect 1390 184 1612 218
rect 1390 91 1424 184
rect 1202 57 1424 91
rect 1460 17 1526 150
rect 1562 70 1612 184
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
rlabel locali s 1257 290 1415 356 6 A1
port 1 nsew signal input
rlabel locali s 1449 252 1607 356 6 A2
port 2 nsew signal input
rlabel locali s 1081 290 1223 356 6 B1
port 3 nsew signal input
rlabel locali s 793 290 1031 356 6 C1
port 4 nsew signal input
rlabel locali s 677 252 743 356 6 D1
port 5 nsew signal input
rlabel locali s 439 70 489 192 6 X
port 6 nsew signal output
rlabel locali s 347 394 413 596 6 X
port 6 nsew signal output
rlabel locali s 283 70 333 192 6 X
port 6 nsew signal output
rlabel locali s 167 394 233 596 6 X
port 6 nsew signal output
rlabel locali s 25 360 413 394 6 X
port 6 nsew signal output
rlabel locali s 25 226 130 360 6 X
port 6 nsew signal output
rlabel locali s 25 192 489 226 6 X
port 6 nsew signal output
rlabel metal1 s 0 -49 1632 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 8 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 9 nsew power bidirectional
rlabel metal1 s 0 617 1632 715 6 VPWR
port 10 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3845918
string GDS_START 3832520
<< end >>
