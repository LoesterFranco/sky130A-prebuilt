magic
tech sky130A
magscale 1 2
timestamp 1604502741
<< locali >>
rect 217 291 331 357
rect 481 294 548 428
rect 85 191 450 257
rect 217 180 450 191
rect 650 236 737 310
rect 217 162 263 180
rect 2120 74 2187 596
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 17 425 111 596
rect 145 460 211 649
rect 319 496 385 596
rect 534 530 635 649
rect 771 546 873 649
rect 907 542 1075 596
rect 907 512 941 542
rect 669 496 941 512
rect 1109 508 1175 596
rect 1296 572 1362 649
rect 319 478 941 496
rect 319 462 879 478
rect 373 425 439 428
rect 17 391 439 425
rect 17 305 165 391
rect 17 157 51 305
rect 373 294 439 391
rect 582 260 616 462
rect 659 364 811 428
rect 484 226 616 260
rect 771 260 811 364
rect 845 330 879 462
rect 991 444 1045 476
rect 913 410 1045 444
rect 913 364 963 410
rect 845 296 957 330
rect 17 70 81 157
rect 117 17 183 157
rect 484 146 518 226
rect 771 192 805 260
rect 625 158 805 192
rect 297 80 518 146
rect 555 17 589 158
rect 625 70 691 158
rect 737 17 803 124
rect 839 85 889 226
rect 923 188 957 296
rect 923 119 977 188
rect 1011 85 1045 410
rect 1079 474 1175 508
rect 1209 504 1543 538
rect 1079 340 1113 474
rect 1209 440 1243 504
rect 1147 374 1243 440
rect 1403 420 1475 470
rect 1329 340 1395 386
rect 1079 306 1395 340
rect 1079 119 1113 306
rect 1429 272 1463 420
rect 1509 386 1543 504
rect 1577 483 1627 596
rect 1769 530 1884 649
rect 1577 449 1779 483
rect 1577 420 1627 449
rect 1509 320 1580 386
rect 1661 298 1711 415
rect 1614 272 1711 298
rect 1147 172 1197 272
rect 1239 206 1463 272
rect 1497 264 1711 272
rect 1745 386 1779 449
rect 1918 420 1987 596
rect 1745 320 1919 386
rect 1953 330 1987 420
rect 2030 364 2080 649
rect 1497 238 1648 264
rect 1497 206 1563 238
rect 1745 230 1779 320
rect 1953 272 2049 330
rect 1429 172 1463 206
rect 1147 138 1395 172
rect 1147 85 1181 138
rect 839 51 1181 85
rect 1277 17 1327 104
rect 1361 85 1395 138
rect 1429 119 1495 172
rect 1529 85 1563 206
rect 1682 196 1779 230
rect 1813 264 2049 272
rect 1813 206 1996 264
rect 1682 188 1716 196
rect 1597 154 1716 188
rect 1597 96 1663 154
rect 1361 51 1563 85
rect 1761 17 1896 162
rect 1930 70 1996 206
rect 2035 17 2085 230
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
<< metal1 >>
rect 0 683 2208 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 0 617 2208 649
rect 0 17 2208 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
rect 0 -49 2208 -17
<< labels >>
rlabel locali s 217 291 331 357 6 D
port 1 nsew signal input
rlabel locali s 2120 74 2187 596 6 Q
port 2 nsew signal output
rlabel locali s 481 294 548 428 6 SCD
port 3 nsew signal input
rlabel locali s 217 180 450 191 6 SCE
port 4 nsew signal input
rlabel locali s 217 162 263 180 6 SCE
port 4 nsew signal input
rlabel locali s 85 191 450 257 6 SCE
port 4 nsew signal input
rlabel locali s 650 236 737 310 6 CLK
port 5 nsew clock input
rlabel metal1 s 0 -49 2208 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 2208 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2208 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 292482
string GDS_START 276280
<< end >>
