magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 123 326 171 487
rect 311 326 359 487
rect 499 326 549 487
rect 686 326 735 487
rect 884 326 945 487
rect 1093 326 1141 487
rect 23 292 1266 326
rect 23 173 57 292
rect 91 207 1113 258
rect 1212 173 1266 292
rect 23 139 1266 173
rect 337 56 375 139
rect 529 56 567 139
rect 721 56 759 139
rect 933 56 971 139
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 27 360 79 527
rect 215 360 267 527
rect 403 360 455 527
rect 593 360 642 527
rect 779 360 840 527
rect 989 360 1049 527
rect 1185 360 1236 527
rect 227 17 293 105
rect 419 17 485 105
rect 611 17 687 105
rect 803 17 889 105
rect 1015 17 1101 105
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
rlabel locali s 91 207 1113 258 6 A
port 1 nsew signal input
rlabel locali s 1212 173 1266 292 6 Y
port 2 nsew signal output
rlabel locali s 1093 326 1141 487 6 Y
port 2 nsew signal output
rlabel locali s 933 56 971 139 6 Y
port 2 nsew signal output
rlabel locali s 884 326 945 487 6 Y
port 2 nsew signal output
rlabel locali s 721 56 759 139 6 Y
port 2 nsew signal output
rlabel locali s 686 326 735 487 6 Y
port 2 nsew signal output
rlabel locali s 529 56 567 139 6 Y
port 2 nsew signal output
rlabel locali s 499 326 549 487 6 Y
port 2 nsew signal output
rlabel locali s 337 56 375 139 6 Y
port 2 nsew signal output
rlabel locali s 311 326 359 487 6 Y
port 2 nsew signal output
rlabel locali s 123 326 171 487 6 Y
port 2 nsew signal output
rlabel locali s 23 292 1266 326 6 Y
port 2 nsew signal output
rlabel locali s 23 173 57 292 6 Y
port 2 nsew signal output
rlabel locali s 23 139 1266 173 6 Y
port 2 nsew signal output
rlabel metal1 s 0 -48 1288 48 8 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 496 1288 592 6 VPWR
port 4 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1288 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1817926
string GDS_START 1808192
<< end >>
