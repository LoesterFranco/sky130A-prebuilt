magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 103 319 175 493
rect 103 51 160 319
rect 427 282 615 325
rect 425 265 615 282
rect 384 256 615 265
rect 384 153 459 256
rect 506 155 615 221
rect 574 84 615 155
rect 671 151 709 325
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 18 299 69 527
rect 223 435 257 527
rect 291 451 572 485
rect 291 401 325 451
rect 692 435 736 527
rect 770 401 847 493
rect 219 367 325 401
rect 359 367 847 401
rect 18 17 69 177
rect 219 265 253 367
rect 359 333 393 367
rect 194 199 253 265
rect 287 299 393 333
rect 287 199 331 299
rect 219 161 253 199
rect 219 127 341 161
rect 307 119 341 127
rect 197 17 273 93
rect 307 53 450 119
rect 697 17 737 117
rect 797 51 847 367
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
rlabel locali s 427 282 615 325 6 A0
port 1 nsew signal input
rlabel locali s 425 265 615 282 6 A0
port 1 nsew signal input
rlabel locali s 384 256 615 265 6 A0
port 1 nsew signal input
rlabel locali s 384 153 459 256 6 A0
port 1 nsew signal input
rlabel locali s 574 84 615 155 6 A1
port 2 nsew signal input
rlabel locali s 506 155 615 221 6 A1
port 2 nsew signal input
rlabel locali s 671 151 709 325 6 S
port 3 nsew signal input
rlabel locali s 103 319 175 493 6 X
port 4 nsew signal output
rlabel locali s 103 51 160 319 6 X
port 4 nsew signal output
rlabel metal1 s 0 -48 920 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 920 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 920 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2136170
string GDS_START 2128756
<< end >>
