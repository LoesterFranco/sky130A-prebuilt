magic
tech sky130A
magscale 1 2
timestamp 1599588218
<< nwell >>
rect -38 332 998 704
<< pwell >>
rect 0 0 960 49
<< scpmos >>
rect 83 368 119 568
rect 299 368 335 568
rect 383 368 419 568
rect 497 368 533 568
rect 611 368 647 568
rect 751 368 787 592
rect 841 368 877 592
<< nmoslvt >>
rect 135 74 165 222
rect 234 74 264 222
rect 335 74 365 222
rect 533 74 563 222
rect 619 74 649 222
rect 733 74 763 222
rect 819 74 849 222
<< ndiff >>
rect 78 202 135 222
rect 78 168 90 202
rect 124 168 135 202
rect 78 120 135 168
rect 78 86 90 120
rect 124 86 135 120
rect 78 74 135 86
rect 165 210 234 222
rect 165 176 189 210
rect 223 176 234 210
rect 165 120 234 176
rect 165 86 189 120
rect 223 86 234 120
rect 165 74 234 86
rect 264 210 335 222
rect 264 176 282 210
rect 316 176 335 210
rect 264 74 335 176
rect 365 150 422 222
rect 365 116 376 150
rect 410 116 422 150
rect 365 74 422 116
rect 476 150 533 222
rect 476 116 488 150
rect 522 116 533 150
rect 476 74 533 116
rect 563 210 619 222
rect 563 176 574 210
rect 608 176 619 210
rect 563 120 619 176
rect 563 86 574 120
rect 608 86 619 120
rect 563 74 619 86
rect 649 210 733 222
rect 649 176 674 210
rect 708 176 733 210
rect 649 120 733 176
rect 649 86 674 120
rect 708 86 733 120
rect 649 74 733 86
rect 763 210 819 222
rect 763 176 774 210
rect 808 176 819 210
rect 763 120 819 176
rect 763 86 774 120
rect 808 86 819 120
rect 763 74 819 86
rect 849 210 933 222
rect 849 176 887 210
rect 921 176 933 210
rect 849 120 933 176
rect 849 86 887 120
rect 921 86 933 120
rect 849 74 933 86
<< pdiff >>
rect 685 580 751 592
rect 685 568 697 580
rect 27 556 83 568
rect 27 522 39 556
rect 73 522 83 556
rect 27 485 83 522
rect 27 451 39 485
rect 73 451 83 485
rect 27 414 83 451
rect 27 380 39 414
rect 73 380 83 414
rect 27 368 83 380
rect 119 560 299 568
rect 119 526 139 560
rect 173 526 255 560
rect 289 526 299 560
rect 119 492 299 526
rect 119 458 139 492
rect 173 458 255 492
rect 289 458 299 492
rect 119 368 299 458
rect 335 368 383 568
rect 419 560 497 568
rect 419 526 429 560
rect 463 526 497 560
rect 419 492 497 526
rect 419 458 429 492
rect 463 458 497 492
rect 419 424 497 458
rect 419 390 429 424
rect 463 390 497 424
rect 419 368 497 390
rect 533 368 611 568
rect 647 546 697 568
rect 731 546 751 580
rect 647 508 751 546
rect 647 474 697 508
rect 731 474 751 508
rect 647 368 751 474
rect 787 580 841 592
rect 787 546 797 580
rect 831 546 841 580
rect 787 497 841 546
rect 787 463 797 497
rect 831 463 841 497
rect 787 414 841 463
rect 787 380 797 414
rect 831 380 841 414
rect 787 368 841 380
rect 877 580 933 592
rect 877 546 887 580
rect 921 546 933 580
rect 877 497 933 546
rect 877 463 887 497
rect 921 463 933 497
rect 877 414 933 463
rect 877 380 887 414
rect 921 380 933 414
rect 877 368 933 380
<< ndiffc >>
rect 90 168 124 202
rect 90 86 124 120
rect 189 176 223 210
rect 189 86 223 120
rect 282 176 316 210
rect 376 116 410 150
rect 488 116 522 150
rect 574 176 608 210
rect 574 86 608 120
rect 674 176 708 210
rect 674 86 708 120
rect 774 176 808 210
rect 774 86 808 120
rect 887 176 921 210
rect 887 86 921 120
<< pdiffc >>
rect 39 522 73 556
rect 39 451 73 485
rect 39 380 73 414
rect 139 526 173 560
rect 255 526 289 560
rect 139 458 173 492
rect 255 458 289 492
rect 429 526 463 560
rect 429 458 463 492
rect 429 390 463 424
rect 697 546 731 580
rect 697 474 731 508
rect 797 546 831 580
rect 797 463 831 497
rect 797 380 831 414
rect 887 546 921 580
rect 887 463 921 497
rect 887 380 921 414
<< poly >>
rect 83 568 119 594
rect 299 568 335 594
rect 383 568 419 594
rect 497 568 533 594
rect 611 568 647 594
rect 751 592 787 618
rect 841 592 877 618
rect 83 310 119 368
rect 299 345 335 368
rect 213 320 335 345
rect 21 294 165 310
rect 21 260 37 294
rect 71 260 165 294
rect 213 286 229 320
rect 263 315 335 320
rect 383 336 419 368
rect 497 336 533 368
rect 611 336 647 368
rect 383 320 449 336
rect 263 286 279 315
rect 213 270 279 286
rect 383 286 399 320
rect 433 286 449 320
rect 21 244 165 260
rect 135 222 165 244
rect 234 222 264 270
rect 383 267 449 286
rect 497 320 563 336
rect 497 286 513 320
rect 547 286 563 320
rect 497 270 563 286
rect 611 320 677 336
rect 751 330 787 368
rect 611 286 627 320
rect 661 286 677 320
rect 611 270 677 286
rect 719 314 787 330
rect 719 280 735 314
rect 769 294 787 314
rect 841 294 877 368
rect 769 280 877 294
rect 335 237 449 267
rect 335 222 365 237
rect 533 222 563 270
rect 619 222 649 270
rect 719 264 877 280
rect 733 222 763 264
rect 819 222 849 264
rect 135 48 165 74
rect 234 48 264 74
rect 335 48 365 74
rect 533 48 563 74
rect 619 48 649 74
rect 733 48 763 74
rect 819 48 849 74
<< polycont >>
rect 37 260 71 294
rect 229 286 263 320
rect 399 286 433 320
rect 513 286 547 320
rect 627 286 661 320
rect 735 280 769 314
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 23 556 89 572
rect 23 522 39 556
rect 73 522 89 556
rect 23 485 89 522
rect 23 451 39 485
rect 73 451 89 485
rect 123 560 305 649
rect 681 580 747 649
rect 123 526 139 560
rect 173 526 255 560
rect 289 526 305 560
rect 123 492 305 526
rect 123 458 139 492
rect 173 458 255 492
rect 289 458 305 492
rect 413 560 479 572
rect 413 526 429 560
rect 463 526 479 560
rect 413 492 479 526
rect 413 458 429 492
rect 463 458 479 492
rect 681 546 697 580
rect 731 546 747 580
rect 681 508 747 546
rect 681 474 697 508
rect 731 474 747 508
rect 681 458 747 474
rect 781 580 853 596
rect 781 546 797 580
rect 831 546 853 580
rect 781 497 853 546
rect 781 463 797 497
rect 831 463 853 497
rect 23 424 89 451
rect 413 424 479 458
rect 23 414 429 424
rect 23 380 39 414
rect 73 390 429 414
rect 463 390 747 424
rect 73 380 155 390
rect 23 364 155 380
rect 21 294 87 310
rect 21 260 37 294
rect 71 260 87 294
rect 21 236 87 260
rect 121 202 155 364
rect 213 320 279 356
rect 213 286 229 320
rect 263 286 279 320
rect 213 270 279 286
rect 313 320 455 356
rect 313 286 399 320
rect 433 286 455 320
rect 313 270 455 286
rect 497 320 563 356
rect 497 286 513 320
rect 547 286 563 320
rect 497 270 563 286
rect 601 320 677 356
rect 601 286 627 320
rect 661 286 677 320
rect 601 270 677 286
rect 713 330 747 390
rect 781 414 853 463
rect 781 380 797 414
rect 831 380 853 414
rect 781 364 853 380
rect 887 580 937 649
rect 921 546 937 580
rect 887 497 937 546
rect 921 463 937 497
rect 887 414 937 463
rect 921 380 937 414
rect 887 364 937 380
rect 713 314 785 330
rect 713 280 735 314
rect 769 280 785 314
rect 713 264 785 280
rect 74 168 90 202
rect 124 168 155 202
rect 74 120 155 168
rect 74 86 90 120
rect 124 86 155 120
rect 74 70 155 86
rect 189 210 223 226
rect 189 120 223 176
rect 259 210 624 236
rect 819 226 853 364
rect 259 176 282 210
rect 316 202 574 210
rect 316 176 324 202
rect 259 160 324 176
rect 608 176 624 210
rect 360 150 426 166
rect 360 116 376 150
rect 410 116 426 150
rect 360 104 426 116
rect 223 86 426 104
rect 189 70 426 86
rect 472 150 538 166
rect 472 116 488 150
rect 522 116 538 150
rect 472 17 538 116
rect 574 120 624 176
rect 608 86 624 120
rect 574 70 624 86
rect 658 210 724 226
rect 658 176 674 210
rect 708 176 724 210
rect 658 120 724 176
rect 658 86 674 120
rect 708 86 724 120
rect 658 17 724 86
rect 758 210 853 226
rect 758 176 774 210
rect 808 176 853 210
rect 758 120 853 176
rect 758 86 774 120
rect 808 86 853 120
rect 758 70 853 86
rect 887 210 937 226
rect 921 176 937 210
rect 887 120 937 176
rect 921 86 937 120
rect 887 17 937 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
rlabel comment s 0 0 0 0 4 o221a_2
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 C1
port 5 nsew
flabel corelocali s 799 94 833 128 0 FreeSans 340 0 0 0 X
port 10 nsew
flabel corelocali s 799 168 833 202 0 FreeSans 340 0 0 0 X
port 10 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 960 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1142998
string GDS_START 1134888
<< end >>
