magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 552 561
rect 18 299 69 527
rect 108 417 347 483
rect 383 367 439 527
rect 481 299 535 493
rect 18 215 85 265
rect 501 152 535 299
rect 118 17 265 113
rect 367 17 443 97
rect 481 83 535 152
rect 0 -17 552 17
<< obsli1 >>
rect 119 265 153 377
rect 198 333 282 383
rect 198 299 447 333
rect 413 265 447 299
rect 119 199 267 265
rect 413 199 459 265
rect 119 181 169 199
rect 22 147 169 181
rect 413 165 447 199
rect 22 53 84 147
rect 299 131 447 165
rect 299 61 333 131
<< metal1 >>
rect 0 496 552 592
rect 0 -48 552 48
<< labels >>
rlabel locali s 108 417 347 483 6 A
port 1 nsew signal input
rlabel locali s 18 215 85 265 6 B_N
port 2 nsew signal input
rlabel locali s 501 152 535 299 6 X
port 3 nsew signal output
rlabel locali s 481 299 535 493 6 X
port 3 nsew signal output
rlabel locali s 481 83 535 152 6 X
port 3 nsew signal output
rlabel locali s 367 17 443 97 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 118 17 265 113 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 552 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 552 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 383 367 439 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 18 299 69 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 552 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 552 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 552 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1014130
string GDS_START 1009242
<< end >>
