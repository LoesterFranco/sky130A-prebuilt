magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 314 347 366 492
rect 506 347 558 492
rect 698 347 750 492
rect 890 347 942 492
rect 314 299 1046 347
rect 17 143 80 265
rect 832 181 1046 299
rect 314 147 1046 181
rect 314 56 366 147
rect 506 56 558 147
rect 698 56 750 147
rect 890 56 942 147
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 19 305 78 527
rect 124 265 174 492
rect 218 305 270 527
rect 410 381 462 527
rect 602 381 654 527
rect 794 381 846 527
rect 986 381 1045 527
rect 124 215 798 265
rect 29 17 78 109
rect 124 53 174 215
rect 218 17 270 122
rect 410 17 462 113
rect 602 17 654 113
rect 794 17 846 113
rect 986 17 1046 113
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
rlabel locali s 17 143 80 265 6 A
port 1 nsew signal input
rlabel locali s 890 347 942 492 6 X
port 2 nsew signal output
rlabel locali s 890 56 942 147 6 X
port 2 nsew signal output
rlabel locali s 832 181 1046 299 6 X
port 2 nsew signal output
rlabel locali s 698 347 750 492 6 X
port 2 nsew signal output
rlabel locali s 698 56 750 147 6 X
port 2 nsew signal output
rlabel locali s 506 347 558 492 6 X
port 2 nsew signal output
rlabel locali s 506 56 558 147 6 X
port 2 nsew signal output
rlabel locali s 314 347 366 492 6 X
port 2 nsew signal output
rlabel locali s 314 299 1046 347 6 X
port 2 nsew signal output
rlabel locali s 314 147 1046 181 6 X
port 2 nsew signal output
rlabel locali s 314 56 366 147 6 X
port 2 nsew signal output
rlabel metal1 s 0 -48 1104 48 8 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 496 1104 592 6 VPWR
port 4 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1104 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1779194
string GDS_START 1770988
<< end >>
