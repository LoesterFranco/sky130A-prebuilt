magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 276 561
rect 17 299 73 527
rect 107 297 173 493
rect 207 299 259 527
rect 19 211 86 265
rect 120 177 154 297
rect 188 215 255 265
rect 17 17 79 177
rect 120 51 259 177
rect 0 -17 276 17
<< metal1 >>
rect 0 496 276 592
rect 0 -48 276 48
<< labels >>
rlabel locali s 188 215 255 265 6 A
port 1 nsew signal input
rlabel locali s 19 211 86 265 6 B
port 2 nsew signal input
rlabel locali s 120 177 154 297 6 Y
port 3 nsew signal output
rlabel locali s 120 51 259 177 6 Y
port 3 nsew signal output
rlabel locali s 107 297 173 493 6 Y
port 3 nsew signal output
rlabel locali s 17 17 79 177 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 276 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 276 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 207 299 259 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 17 299 73 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 276 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 276 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 276 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1690806
string GDS_START 1686914
<< end >>
