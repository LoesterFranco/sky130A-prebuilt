magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 89 53 119 137
rect 279 53 309 137
rect 373 53 403 137
rect 481 47 511 177
<< pmoshvt >>
rect 81 297 117 381
rect 283 297 319 381
rect 365 297 401 381
rect 473 297 509 497
<< ndiff >>
rect 418 137 481 177
rect 27 106 89 137
rect 27 72 35 106
rect 69 72 89 106
rect 27 53 89 72
rect 119 97 279 137
rect 119 63 129 97
rect 163 63 225 97
rect 259 63 279 97
rect 119 53 279 63
rect 309 111 373 137
rect 309 77 319 111
rect 353 77 373 111
rect 309 53 373 77
rect 403 97 481 137
rect 403 63 423 97
rect 457 63 481 97
rect 403 53 481 63
rect 418 47 481 53
rect 511 135 565 177
rect 511 101 521 135
rect 555 101 565 135
rect 511 47 565 101
<< pdiff >>
rect 418 485 473 497
rect 418 451 426 485
rect 460 451 473 485
rect 418 417 473 451
rect 418 383 426 417
rect 460 383 473 417
rect 418 381 473 383
rect 27 349 81 381
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 341 175 381
rect 117 307 129 341
rect 163 307 175 341
rect 117 297 175 307
rect 229 354 283 381
rect 229 320 237 354
rect 271 320 283 354
rect 229 297 283 320
rect 319 297 365 381
rect 401 297 473 381
rect 509 454 565 497
rect 509 420 521 454
rect 555 420 565 454
rect 509 386 565 420
rect 509 352 521 386
rect 555 352 565 386
rect 509 297 565 352
<< ndiffc >>
rect 35 72 69 106
rect 129 63 163 97
rect 225 63 259 97
rect 319 77 353 111
rect 423 63 457 97
rect 521 101 555 135
<< pdiffc >>
rect 426 451 460 485
rect 426 383 460 417
rect 35 315 69 349
rect 129 307 163 341
rect 237 320 271 354
rect 521 420 555 454
rect 521 352 555 386
<< poly >>
rect 473 497 509 523
rect 179 473 403 483
rect 179 439 195 473
rect 229 453 403 473
rect 229 439 245 453
rect 179 429 245 439
rect 363 407 403 453
rect 81 381 117 407
rect 283 381 319 407
rect 365 381 401 407
rect 81 282 117 297
rect 283 282 319 297
rect 365 282 401 297
rect 473 282 509 297
rect 79 265 119 282
rect 281 265 321 282
rect 22 249 119 265
rect 22 215 35 249
rect 69 215 119 249
rect 22 199 119 215
rect 227 249 321 265
rect 227 215 237 249
rect 271 215 321 249
rect 363 227 403 282
rect 471 265 511 282
rect 227 199 321 215
rect 89 137 119 199
rect 279 137 309 199
rect 373 137 403 227
rect 445 249 511 265
rect 445 215 455 249
rect 489 215 511 249
rect 445 199 511 215
rect 481 177 511 199
rect 89 27 119 53
rect 279 27 309 53
rect 373 27 403 53
rect 481 21 511 47
<< polycont >>
rect 195 439 229 473
rect 35 215 69 249
rect 237 215 271 249
rect 455 215 489 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 644 561
rect 18 349 69 527
rect 413 485 469 527
rect 108 473 367 483
rect 108 439 195 473
rect 229 439 367 473
rect 108 417 367 439
rect 413 451 426 485
rect 460 451 469 485
rect 413 417 469 451
rect 413 383 426 417
rect 460 383 469 417
rect 18 315 35 349
rect 18 299 69 315
rect 129 341 163 377
rect 129 265 163 307
rect 208 354 292 383
rect 413 367 469 383
rect 521 454 618 493
rect 555 420 618 454
rect 521 386 618 420
rect 208 320 237 354
rect 271 333 292 354
rect 555 352 618 386
rect 271 320 477 333
rect 208 299 477 320
rect 521 299 618 352
rect 443 265 477 299
rect 18 249 85 265
rect 18 215 35 249
rect 69 215 85 249
rect 129 249 277 265
rect 129 215 237 249
rect 271 215 277 249
rect 129 199 277 215
rect 443 249 489 265
rect 443 215 455 249
rect 443 199 489 215
rect 129 181 179 199
rect 22 147 179 181
rect 443 165 477 199
rect 22 106 84 147
rect 319 131 477 165
rect 541 152 618 299
rect 521 135 618 152
rect 22 72 35 106
rect 69 72 84 106
rect 22 53 84 72
rect 128 97 275 113
rect 128 63 129 97
rect 163 63 225 97
rect 259 63 275 97
rect 128 17 275 63
rect 319 111 353 131
rect 555 101 618 135
rect 319 61 353 77
rect 387 63 423 97
rect 457 63 473 97
rect 521 83 618 101
rect 387 17 473 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel corelocali s 224 425 258 459 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 400 0 0 0 B_N
port 2 nsew
flabel corelocali s 578 357 612 391 0 FreeSans 400 0 0 0 X
port 7 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew
rlabel comment s 0 0 0 0 4 or2b_1
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 648822
string GDS_START 643726
<< end >>
