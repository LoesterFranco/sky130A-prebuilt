magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 2522 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 93 47 123 177
rect 177 47 207 177
rect 281 47 311 177
rect 365 47 395 177
rect 469 47 499 177
rect 553 47 583 177
rect 657 47 687 177
rect 741 47 771 177
rect 845 47 875 177
rect 929 47 959 177
rect 1033 47 1063 177
rect 1117 47 1147 177
rect 1325 47 1355 177
rect 1409 47 1439 177
rect 1513 47 1543 177
rect 1597 47 1627 177
rect 1701 47 1731 177
rect 1785 47 1815 177
rect 1889 47 1919 177
rect 1973 47 2003 177
rect 2077 47 2107 177
rect 2161 47 2191 177
rect 2265 47 2295 177
rect 2349 47 2379 177
<< pmoshvt >>
rect 85 297 121 497
rect 179 297 215 497
rect 273 297 309 497
rect 367 297 403 497
rect 461 297 497 497
rect 555 297 591 497
rect 649 297 685 497
rect 743 297 779 497
rect 837 297 873 497
rect 931 297 967 497
rect 1025 297 1061 497
rect 1119 297 1155 497
rect 1317 297 1353 497
rect 1411 297 1447 497
rect 1505 297 1541 497
rect 1599 297 1635 497
rect 1693 297 1729 497
rect 1787 297 1823 497
rect 1881 297 1917 497
rect 1975 297 2011 497
rect 2069 297 2105 497
rect 2163 297 2199 497
rect 2257 297 2293 497
rect 2351 297 2387 497
<< ndiff >>
rect 27 163 93 177
rect 27 129 39 163
rect 73 129 93 163
rect 27 95 93 129
rect 27 61 39 95
rect 73 61 93 95
rect 27 47 93 61
rect 123 163 177 177
rect 123 129 133 163
rect 167 129 177 163
rect 123 95 177 129
rect 123 61 133 95
rect 167 61 177 95
rect 123 47 177 61
rect 207 95 281 177
rect 207 61 227 95
rect 261 61 281 95
rect 207 47 281 61
rect 311 163 365 177
rect 311 129 321 163
rect 355 129 365 163
rect 311 95 365 129
rect 311 61 321 95
rect 355 61 365 95
rect 311 47 365 61
rect 395 95 469 177
rect 395 61 415 95
rect 449 61 469 95
rect 395 47 469 61
rect 499 163 553 177
rect 499 129 509 163
rect 543 129 553 163
rect 499 95 553 129
rect 499 61 509 95
rect 543 61 553 95
rect 499 47 553 61
rect 583 95 657 177
rect 583 61 603 95
rect 637 61 657 95
rect 583 47 657 61
rect 687 163 741 177
rect 687 129 697 163
rect 731 129 741 163
rect 687 95 741 129
rect 687 61 697 95
rect 731 61 741 95
rect 687 47 741 61
rect 771 95 845 177
rect 771 61 791 95
rect 825 61 845 95
rect 771 47 845 61
rect 875 163 929 177
rect 875 129 885 163
rect 919 129 929 163
rect 875 95 929 129
rect 875 61 885 95
rect 919 61 929 95
rect 875 47 929 61
rect 959 95 1033 177
rect 959 61 979 95
rect 1013 61 1033 95
rect 959 47 1033 61
rect 1063 163 1117 177
rect 1063 129 1073 163
rect 1107 129 1117 163
rect 1063 95 1117 129
rect 1063 61 1073 95
rect 1107 61 1117 95
rect 1063 47 1117 61
rect 1147 95 1325 177
rect 1147 61 1167 95
rect 1201 61 1271 95
rect 1305 61 1325 95
rect 1147 47 1325 61
rect 1355 163 1409 177
rect 1355 129 1365 163
rect 1399 129 1409 163
rect 1355 95 1409 129
rect 1355 61 1365 95
rect 1399 61 1409 95
rect 1355 47 1409 61
rect 1439 95 1513 177
rect 1439 61 1459 95
rect 1493 61 1513 95
rect 1439 47 1513 61
rect 1543 163 1597 177
rect 1543 129 1553 163
rect 1587 129 1597 163
rect 1543 95 1597 129
rect 1543 61 1553 95
rect 1587 61 1597 95
rect 1543 47 1597 61
rect 1627 95 1701 177
rect 1627 61 1647 95
rect 1681 61 1701 95
rect 1627 47 1701 61
rect 1731 163 1785 177
rect 1731 129 1741 163
rect 1775 129 1785 163
rect 1731 95 1785 129
rect 1731 61 1741 95
rect 1775 61 1785 95
rect 1731 47 1785 61
rect 1815 95 1889 177
rect 1815 61 1835 95
rect 1869 61 1889 95
rect 1815 47 1889 61
rect 1919 163 1973 177
rect 1919 129 1929 163
rect 1963 129 1973 163
rect 1919 95 1973 129
rect 1919 61 1929 95
rect 1963 61 1973 95
rect 1919 47 1973 61
rect 2003 95 2077 177
rect 2003 61 2023 95
rect 2057 61 2077 95
rect 2003 47 2077 61
rect 2107 163 2161 177
rect 2107 129 2117 163
rect 2151 129 2161 163
rect 2107 95 2161 129
rect 2107 61 2117 95
rect 2151 61 2161 95
rect 2107 47 2161 61
rect 2191 95 2265 177
rect 2191 61 2211 95
rect 2245 61 2265 95
rect 2191 47 2265 61
rect 2295 163 2349 177
rect 2295 129 2305 163
rect 2339 129 2349 163
rect 2295 95 2349 129
rect 2295 61 2305 95
rect 2339 61 2349 95
rect 2295 47 2349 61
rect 2379 163 2447 177
rect 2379 129 2401 163
rect 2435 129 2447 163
rect 2379 95 2447 129
rect 2379 61 2401 95
rect 2435 61 2447 95
rect 2379 47 2447 61
<< pdiff >>
rect 27 477 85 497
rect 27 443 39 477
rect 73 443 85 477
rect 27 409 85 443
rect 27 375 39 409
rect 73 375 85 409
rect 27 341 85 375
rect 27 307 39 341
rect 73 307 85 341
rect 27 297 85 307
rect 121 477 179 497
rect 121 443 133 477
rect 167 443 179 477
rect 121 409 179 443
rect 121 375 133 409
rect 167 375 179 409
rect 121 297 179 375
rect 215 477 273 497
rect 215 443 227 477
rect 261 443 273 477
rect 215 409 273 443
rect 215 375 227 409
rect 261 375 273 409
rect 215 341 273 375
rect 215 307 227 341
rect 261 307 273 341
rect 215 297 273 307
rect 309 477 367 497
rect 309 443 321 477
rect 355 443 367 477
rect 309 409 367 443
rect 309 375 321 409
rect 355 375 367 409
rect 309 297 367 375
rect 403 477 461 497
rect 403 443 415 477
rect 449 443 461 477
rect 403 409 461 443
rect 403 375 415 409
rect 449 375 461 409
rect 403 341 461 375
rect 403 307 415 341
rect 449 307 461 341
rect 403 297 461 307
rect 497 477 555 497
rect 497 443 509 477
rect 543 443 555 477
rect 497 409 555 443
rect 497 375 509 409
rect 543 375 555 409
rect 497 297 555 375
rect 591 477 649 497
rect 591 443 603 477
rect 637 443 649 477
rect 591 409 649 443
rect 591 375 603 409
rect 637 375 649 409
rect 591 341 649 375
rect 591 307 603 341
rect 637 307 649 341
rect 591 297 649 307
rect 685 409 743 497
rect 685 375 697 409
rect 731 375 743 409
rect 685 341 743 375
rect 685 307 697 341
rect 731 307 743 341
rect 685 297 743 307
rect 779 477 837 497
rect 779 443 791 477
rect 825 443 837 477
rect 779 409 837 443
rect 779 375 791 409
rect 825 375 837 409
rect 779 297 837 375
rect 873 409 931 497
rect 873 375 885 409
rect 919 375 931 409
rect 873 341 931 375
rect 873 307 885 341
rect 919 307 931 341
rect 873 297 931 307
rect 967 477 1025 497
rect 967 443 979 477
rect 1013 443 1025 477
rect 967 409 1025 443
rect 967 375 979 409
rect 1013 375 1025 409
rect 967 297 1025 375
rect 1061 409 1119 497
rect 1061 375 1073 409
rect 1107 375 1119 409
rect 1061 341 1119 375
rect 1061 307 1073 341
rect 1107 307 1119 341
rect 1061 297 1119 307
rect 1155 477 1209 497
rect 1155 443 1167 477
rect 1201 443 1209 477
rect 1155 409 1209 443
rect 1155 375 1167 409
rect 1201 375 1209 409
rect 1155 297 1209 375
rect 1263 477 1317 497
rect 1263 443 1271 477
rect 1305 443 1317 477
rect 1263 409 1317 443
rect 1263 375 1271 409
rect 1305 375 1317 409
rect 1263 297 1317 375
rect 1353 409 1411 497
rect 1353 375 1365 409
rect 1399 375 1411 409
rect 1353 341 1411 375
rect 1353 307 1365 341
rect 1399 307 1411 341
rect 1353 297 1411 307
rect 1447 477 1505 497
rect 1447 443 1459 477
rect 1493 443 1505 477
rect 1447 409 1505 443
rect 1447 375 1459 409
rect 1493 375 1505 409
rect 1447 297 1505 375
rect 1541 409 1599 497
rect 1541 375 1553 409
rect 1587 375 1599 409
rect 1541 341 1599 375
rect 1541 307 1553 341
rect 1587 307 1599 341
rect 1541 297 1599 307
rect 1635 477 1693 497
rect 1635 443 1647 477
rect 1681 443 1693 477
rect 1635 409 1693 443
rect 1635 375 1647 409
rect 1681 375 1693 409
rect 1635 297 1693 375
rect 1729 409 1787 497
rect 1729 375 1741 409
rect 1775 375 1787 409
rect 1729 341 1787 375
rect 1729 307 1741 341
rect 1775 307 1787 341
rect 1729 297 1787 307
rect 1823 477 1881 497
rect 1823 443 1835 477
rect 1869 443 1881 477
rect 1823 409 1881 443
rect 1823 375 1835 409
rect 1869 375 1881 409
rect 1823 341 1881 375
rect 1823 307 1835 341
rect 1869 307 1881 341
rect 1823 297 1881 307
rect 1917 409 1975 497
rect 1917 375 1929 409
rect 1963 375 1975 409
rect 1917 341 1975 375
rect 1917 307 1929 341
rect 1963 307 1975 341
rect 1917 297 1975 307
rect 2011 477 2069 497
rect 2011 443 2023 477
rect 2057 443 2069 477
rect 2011 409 2069 443
rect 2011 375 2023 409
rect 2057 375 2069 409
rect 2011 297 2069 375
rect 2105 409 2163 497
rect 2105 375 2117 409
rect 2151 375 2163 409
rect 2105 341 2163 375
rect 2105 307 2117 341
rect 2151 307 2163 341
rect 2105 297 2163 307
rect 2199 477 2257 497
rect 2199 443 2211 477
rect 2245 443 2257 477
rect 2199 409 2257 443
rect 2199 375 2211 409
rect 2245 375 2257 409
rect 2199 297 2257 375
rect 2293 409 2351 497
rect 2293 375 2305 409
rect 2339 375 2351 409
rect 2293 341 2351 375
rect 2293 307 2305 341
rect 2339 307 2351 341
rect 2293 297 2351 307
rect 2387 477 2447 497
rect 2387 443 2401 477
rect 2435 443 2447 477
rect 2387 409 2447 443
rect 2387 375 2401 409
rect 2435 375 2447 409
rect 2387 341 2447 375
rect 2387 307 2401 341
rect 2435 307 2447 341
rect 2387 297 2447 307
<< ndiffc >>
rect 39 129 73 163
rect 39 61 73 95
rect 133 129 167 163
rect 133 61 167 95
rect 227 61 261 95
rect 321 129 355 163
rect 321 61 355 95
rect 415 61 449 95
rect 509 129 543 163
rect 509 61 543 95
rect 603 61 637 95
rect 697 129 731 163
rect 697 61 731 95
rect 791 61 825 95
rect 885 129 919 163
rect 885 61 919 95
rect 979 61 1013 95
rect 1073 129 1107 163
rect 1073 61 1107 95
rect 1167 61 1201 95
rect 1271 61 1305 95
rect 1365 129 1399 163
rect 1365 61 1399 95
rect 1459 61 1493 95
rect 1553 129 1587 163
rect 1553 61 1587 95
rect 1647 61 1681 95
rect 1741 129 1775 163
rect 1741 61 1775 95
rect 1835 61 1869 95
rect 1929 129 1963 163
rect 1929 61 1963 95
rect 2023 61 2057 95
rect 2117 129 2151 163
rect 2117 61 2151 95
rect 2211 61 2245 95
rect 2305 129 2339 163
rect 2305 61 2339 95
rect 2401 129 2435 163
rect 2401 61 2435 95
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 133 443 167 477
rect 133 375 167 409
rect 227 443 261 477
rect 227 375 261 409
rect 227 307 261 341
rect 321 443 355 477
rect 321 375 355 409
rect 415 443 449 477
rect 415 375 449 409
rect 415 307 449 341
rect 509 443 543 477
rect 509 375 543 409
rect 603 443 637 477
rect 603 375 637 409
rect 603 307 637 341
rect 697 375 731 409
rect 697 307 731 341
rect 791 443 825 477
rect 791 375 825 409
rect 885 375 919 409
rect 885 307 919 341
rect 979 443 1013 477
rect 979 375 1013 409
rect 1073 375 1107 409
rect 1073 307 1107 341
rect 1167 443 1201 477
rect 1167 375 1201 409
rect 1271 443 1305 477
rect 1271 375 1305 409
rect 1365 375 1399 409
rect 1365 307 1399 341
rect 1459 443 1493 477
rect 1459 375 1493 409
rect 1553 375 1587 409
rect 1553 307 1587 341
rect 1647 443 1681 477
rect 1647 375 1681 409
rect 1741 375 1775 409
rect 1741 307 1775 341
rect 1835 443 1869 477
rect 1835 375 1869 409
rect 1835 307 1869 341
rect 1929 375 1963 409
rect 1929 307 1963 341
rect 2023 443 2057 477
rect 2023 375 2057 409
rect 2117 375 2151 409
rect 2117 307 2151 341
rect 2211 443 2245 477
rect 2211 375 2245 409
rect 2305 375 2339 409
rect 2305 307 2339 341
rect 2401 443 2435 477
rect 2401 375 2435 409
rect 2401 307 2435 341
<< poly >>
rect 85 497 121 523
rect 179 497 215 523
rect 273 497 309 523
rect 367 497 403 523
rect 461 497 497 523
rect 555 497 591 523
rect 649 497 685 523
rect 743 497 779 523
rect 837 497 873 523
rect 931 497 967 523
rect 1025 497 1061 523
rect 1119 497 1155 523
rect 1317 497 1353 523
rect 1411 497 1447 523
rect 1505 497 1541 523
rect 1599 497 1635 523
rect 1693 497 1729 523
rect 1787 497 1823 523
rect 1881 497 1917 523
rect 1975 497 2011 523
rect 2069 497 2105 523
rect 2163 497 2199 523
rect 2257 497 2293 523
rect 2351 497 2387 523
rect 85 282 121 297
rect 179 282 215 297
rect 273 282 309 297
rect 367 282 403 297
rect 461 282 497 297
rect 555 282 591 297
rect 649 282 685 297
rect 743 282 779 297
rect 837 282 873 297
rect 931 282 967 297
rect 1025 282 1061 297
rect 1119 282 1155 297
rect 1317 282 1353 297
rect 1411 282 1447 297
rect 1505 282 1541 297
rect 1599 282 1635 297
rect 1693 282 1729 297
rect 1787 282 1823 297
rect 1881 282 1917 297
rect 1975 282 2011 297
rect 2069 282 2105 297
rect 2163 282 2199 297
rect 2257 282 2293 297
rect 2351 282 2387 297
rect 83 265 123 282
rect 177 265 217 282
rect 271 265 311 282
rect 365 265 405 282
rect 459 265 499 282
rect 553 265 593 282
rect 83 249 593 265
rect 83 215 117 249
rect 151 215 185 249
rect 219 215 253 249
rect 287 215 321 249
rect 355 215 389 249
rect 423 215 457 249
rect 491 215 525 249
rect 559 215 593 249
rect 83 199 593 215
rect 647 265 687 282
rect 741 265 781 282
rect 835 265 875 282
rect 929 265 969 282
rect 1023 265 1063 282
rect 1117 265 1157 282
rect 647 249 1157 265
rect 647 215 681 249
rect 715 215 749 249
rect 783 215 817 249
rect 851 215 885 249
rect 919 215 953 249
rect 987 215 1021 249
rect 1055 215 1089 249
rect 1123 215 1157 249
rect 647 199 1157 215
rect 1315 265 1355 282
rect 1409 265 1449 282
rect 1503 265 1543 282
rect 1597 265 1637 282
rect 1691 265 1731 282
rect 1785 265 1825 282
rect 1315 249 1825 265
rect 1315 215 1349 249
rect 1383 215 1417 249
rect 1451 215 1485 249
rect 1519 215 1553 249
rect 1587 215 1621 249
rect 1655 215 1689 249
rect 1723 215 1757 249
rect 1791 215 1825 249
rect 1315 199 1825 215
rect 1879 265 1919 282
rect 1973 265 2013 282
rect 2067 265 2107 282
rect 2161 265 2201 282
rect 2255 265 2295 282
rect 2349 265 2389 282
rect 1879 249 2389 265
rect 1879 215 1895 249
rect 1929 215 1963 249
rect 1997 215 2031 249
rect 2065 215 2099 249
rect 2133 215 2167 249
rect 2201 215 2389 249
rect 1879 199 2389 215
rect 93 177 123 199
rect 177 177 207 199
rect 281 177 311 199
rect 365 177 395 199
rect 469 177 499 199
rect 553 177 583 199
rect 657 177 687 199
rect 741 177 771 199
rect 845 177 875 199
rect 929 177 959 199
rect 1033 177 1063 199
rect 1117 177 1147 199
rect 1325 177 1355 199
rect 1409 177 1439 199
rect 1513 177 1543 199
rect 1597 177 1627 199
rect 1701 177 1731 199
rect 1785 177 1815 199
rect 1889 177 1919 199
rect 1973 177 2003 199
rect 2077 177 2107 199
rect 2161 177 2191 199
rect 2265 177 2295 199
rect 2349 177 2379 199
rect 93 21 123 47
rect 177 21 207 47
rect 281 21 311 47
rect 365 21 395 47
rect 469 21 499 47
rect 553 21 583 47
rect 657 21 687 47
rect 741 21 771 47
rect 845 21 875 47
rect 929 21 959 47
rect 1033 21 1063 47
rect 1117 21 1147 47
rect 1325 21 1355 47
rect 1409 21 1439 47
rect 1513 21 1543 47
rect 1597 21 1627 47
rect 1701 21 1731 47
rect 1785 21 1815 47
rect 1889 21 1919 47
rect 1973 21 2003 47
rect 2077 21 2107 47
rect 2161 21 2191 47
rect 2265 21 2295 47
rect 2349 21 2379 47
<< polycont >>
rect 117 215 151 249
rect 185 215 219 249
rect 253 215 287 249
rect 321 215 355 249
rect 389 215 423 249
rect 457 215 491 249
rect 525 215 559 249
rect 681 215 715 249
rect 749 215 783 249
rect 817 215 851 249
rect 885 215 919 249
rect 953 215 987 249
rect 1021 215 1055 249
rect 1089 215 1123 249
rect 1349 215 1383 249
rect 1417 215 1451 249
rect 1485 215 1519 249
rect 1553 215 1587 249
rect 1621 215 1655 249
rect 1689 215 1723 249
rect 1757 215 1791 249
rect 1895 215 1929 249
rect 1963 215 1997 249
rect 2031 215 2065 249
rect 2099 215 2133 249
rect 2167 215 2201 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2484 561
rect 23 477 81 493
rect 23 443 39 477
rect 73 443 81 477
rect 23 409 81 443
rect 23 375 39 409
rect 73 375 81 409
rect 23 341 81 375
rect 125 477 175 527
rect 125 443 133 477
rect 167 443 175 477
rect 125 409 175 443
rect 125 375 133 409
rect 167 375 175 409
rect 125 359 175 375
rect 219 477 269 493
rect 219 443 227 477
rect 261 443 269 477
rect 219 409 269 443
rect 219 375 227 409
rect 261 375 269 409
rect 23 307 39 341
rect 73 325 81 341
rect 219 341 269 375
rect 313 477 363 527
rect 313 443 321 477
rect 355 443 363 477
rect 313 409 363 443
rect 313 375 321 409
rect 355 375 363 409
rect 313 359 363 375
rect 407 477 457 493
rect 407 443 415 477
rect 449 443 457 477
rect 407 409 457 443
rect 407 375 415 409
rect 449 375 457 409
rect 219 325 227 341
rect 73 307 227 325
rect 261 325 269 341
rect 407 341 457 375
rect 501 477 551 527
rect 501 443 509 477
rect 543 443 551 477
rect 501 409 551 443
rect 501 375 509 409
rect 543 375 551 409
rect 501 359 551 375
rect 595 477 1217 493
rect 595 443 603 477
rect 637 459 791 477
rect 637 443 645 459
rect 595 409 645 443
rect 783 443 791 459
rect 825 459 979 477
rect 825 443 833 459
rect 595 375 603 409
rect 637 375 645 409
rect 407 325 415 341
rect 261 307 415 325
rect 449 325 457 341
rect 595 341 645 375
rect 595 325 603 341
rect 449 307 603 325
rect 637 307 645 341
rect 23 291 645 307
rect 689 409 739 425
rect 689 375 697 409
rect 731 375 739 409
rect 689 341 739 375
rect 783 409 833 443
rect 971 443 979 459
rect 1013 459 1167 477
rect 1013 443 1021 459
rect 783 375 791 409
rect 825 375 833 409
rect 783 359 833 375
rect 877 409 927 425
rect 877 375 885 409
rect 919 375 927 409
rect 689 307 697 341
rect 731 325 739 341
rect 877 341 927 375
rect 971 409 1021 443
rect 1159 443 1167 459
rect 1201 443 1217 477
rect 971 375 979 409
rect 1013 375 1021 409
rect 971 359 1021 375
rect 1065 409 1115 425
rect 1065 375 1073 409
rect 1107 375 1115 409
rect 877 325 885 341
rect 731 307 885 325
rect 919 325 927 341
rect 1065 341 1115 375
rect 1159 409 1217 443
rect 1159 375 1167 409
rect 1201 375 1217 409
rect 1159 359 1217 375
rect 1255 477 2451 493
rect 1255 443 1271 477
rect 1305 459 1459 477
rect 1305 443 1313 459
rect 1255 409 1313 443
rect 1451 443 1459 459
rect 1493 459 1647 477
rect 1493 443 1501 459
rect 1255 375 1271 409
rect 1305 375 1313 409
rect 1255 359 1313 375
rect 1357 409 1407 425
rect 1357 375 1365 409
rect 1399 375 1407 409
rect 1065 325 1073 341
rect 919 307 1073 325
rect 1107 325 1115 341
rect 1357 341 1407 375
rect 1451 409 1501 443
rect 1639 443 1647 459
rect 1681 459 1835 477
rect 1681 443 1689 459
rect 1451 375 1459 409
rect 1493 375 1501 409
rect 1451 359 1501 375
rect 1545 409 1595 425
rect 1545 375 1553 409
rect 1587 375 1595 409
rect 1357 325 1365 341
rect 1107 307 1365 325
rect 1399 325 1407 341
rect 1545 341 1595 375
rect 1639 409 1689 443
rect 1827 443 1835 459
rect 1869 459 2023 477
rect 1869 443 1877 459
rect 1639 375 1647 409
rect 1681 375 1689 409
rect 1639 359 1689 375
rect 1733 409 1783 425
rect 1733 375 1741 409
rect 1775 375 1783 409
rect 1545 325 1553 341
rect 1399 307 1553 325
rect 1587 325 1595 341
rect 1733 341 1783 375
rect 1733 325 1741 341
rect 1587 307 1741 325
rect 1775 307 1783 341
rect 689 291 1783 307
rect 1827 409 1877 443
rect 2015 443 2023 459
rect 2057 459 2211 477
rect 2057 443 2065 459
rect 1827 375 1835 409
rect 1869 375 1877 409
rect 1827 341 1877 375
rect 1827 307 1835 341
rect 1869 307 1877 341
rect 1827 291 1877 307
rect 1921 409 1971 425
rect 1921 375 1929 409
rect 1963 375 1971 409
rect 1921 341 1971 375
rect 2015 409 2065 443
rect 2203 443 2211 459
rect 2245 459 2401 477
rect 2245 443 2253 459
rect 2015 375 2023 409
rect 2057 375 2065 409
rect 2015 359 2065 375
rect 2109 409 2159 425
rect 2109 375 2117 409
rect 2151 375 2159 409
rect 1921 307 1929 341
rect 1963 325 1971 341
rect 2109 341 2159 375
rect 2203 409 2253 443
rect 2435 443 2451 477
rect 2203 375 2211 409
rect 2245 375 2253 409
rect 2203 359 2253 375
rect 2289 409 2367 425
rect 2289 375 2305 409
rect 2339 375 2367 409
rect 2109 325 2117 341
rect 1963 307 2117 325
rect 2151 325 2159 341
rect 2289 341 2367 375
rect 2289 325 2305 341
rect 2151 307 2305 325
rect 2339 307 2367 341
rect 1921 291 2367 307
rect 2401 409 2451 443
rect 2435 375 2451 409
rect 2401 341 2451 375
rect 2435 307 2451 341
rect 2401 291 2451 307
rect 101 249 575 257
rect 101 215 117 249
rect 151 215 185 249
rect 219 215 253 249
rect 287 215 321 249
rect 355 215 389 249
rect 423 215 457 249
rect 491 215 525 249
rect 559 215 575 249
rect 665 249 1139 257
rect 665 215 681 249
rect 715 215 749 249
rect 783 215 817 249
rect 851 215 885 249
rect 919 215 953 249
rect 987 215 1021 249
rect 1055 215 1089 249
rect 1123 215 1139 249
rect 1333 249 1807 257
rect 1333 215 1349 249
rect 1383 215 1417 249
rect 1451 215 1485 249
rect 1519 215 1553 249
rect 1587 215 1621 249
rect 1655 215 1689 249
rect 1723 215 1757 249
rect 1791 215 1807 249
rect 1879 249 2217 257
rect 1879 215 1895 249
rect 1929 215 1963 249
rect 1997 215 2031 249
rect 2065 215 2099 249
rect 2133 215 2167 249
rect 2201 215 2217 249
rect 2289 181 2367 291
rect 23 163 83 181
rect 23 129 39 163
rect 73 129 83 163
rect 23 95 83 129
rect 23 61 39 95
rect 73 61 83 95
rect 23 17 83 61
rect 117 163 2367 181
rect 117 129 133 163
rect 167 145 321 163
rect 167 129 183 145
rect 117 95 183 129
rect 305 129 321 145
rect 355 145 509 163
rect 355 129 371 145
rect 117 61 133 95
rect 167 61 183 95
rect 117 51 183 61
rect 217 95 271 111
rect 217 61 227 95
rect 261 61 271 95
rect 217 17 271 61
rect 305 95 371 129
rect 493 129 509 145
rect 543 145 697 163
rect 543 129 559 145
rect 305 61 321 95
rect 355 61 371 95
rect 305 51 371 61
rect 405 95 459 111
rect 405 61 415 95
rect 449 61 459 95
rect 405 17 459 61
rect 493 95 559 129
rect 681 129 697 145
rect 731 145 885 163
rect 731 129 747 145
rect 493 61 509 95
rect 543 61 559 95
rect 493 51 559 61
rect 593 95 647 111
rect 593 61 603 95
rect 637 61 647 95
rect 593 17 647 61
rect 681 95 747 129
rect 869 129 885 145
rect 919 145 1073 163
rect 919 129 935 145
rect 681 61 697 95
rect 731 61 747 95
rect 681 51 747 61
rect 781 95 835 111
rect 781 61 791 95
rect 825 61 835 95
rect 781 17 835 61
rect 869 95 935 129
rect 1057 129 1073 145
rect 1107 145 1365 163
rect 1107 129 1123 145
rect 869 61 885 95
rect 919 61 935 95
rect 869 51 935 61
rect 969 95 1023 111
rect 969 61 979 95
rect 1013 61 1023 95
rect 969 17 1023 61
rect 1057 95 1123 129
rect 1349 129 1365 145
rect 1399 145 1553 163
rect 1399 129 1415 145
rect 1057 61 1073 95
rect 1107 61 1123 95
rect 1057 51 1123 61
rect 1157 95 1315 111
rect 1157 61 1167 95
rect 1201 61 1271 95
rect 1305 61 1315 95
rect 1157 17 1315 61
rect 1349 95 1415 129
rect 1537 129 1553 145
rect 1587 145 1741 163
rect 1587 129 1603 145
rect 1349 61 1365 95
rect 1399 61 1415 95
rect 1349 51 1415 61
rect 1449 95 1503 111
rect 1449 61 1459 95
rect 1493 61 1503 95
rect 1449 17 1503 61
rect 1537 95 1603 129
rect 1725 129 1741 145
rect 1775 145 1929 163
rect 1775 129 1791 145
rect 1537 61 1553 95
rect 1587 61 1603 95
rect 1537 51 1603 61
rect 1637 95 1691 111
rect 1637 61 1647 95
rect 1681 61 1691 95
rect 1637 17 1691 61
rect 1725 95 1791 129
rect 1913 129 1929 145
rect 1963 145 2117 163
rect 1963 129 1979 145
rect 1725 61 1741 95
rect 1775 61 1791 95
rect 1725 51 1791 61
rect 1825 95 1879 111
rect 1825 61 1835 95
rect 1869 61 1879 95
rect 1825 17 1879 61
rect 1913 95 1979 129
rect 2101 129 2117 145
rect 2151 145 2305 163
rect 2151 129 2167 145
rect 1913 61 1929 95
rect 1963 61 1979 95
rect 1913 51 1979 61
rect 2013 95 2067 111
rect 2013 61 2023 95
rect 2057 61 2067 95
rect 2013 17 2067 61
rect 2101 95 2167 129
rect 2289 129 2305 145
rect 2339 129 2367 163
rect 2101 61 2117 95
rect 2151 61 2167 95
rect 2101 51 2167 61
rect 2201 95 2255 111
rect 2201 61 2211 95
rect 2245 61 2255 95
rect 2201 17 2255 61
rect 2289 95 2367 129
rect 2289 61 2305 95
rect 2339 61 2367 95
rect 2289 51 2367 61
rect 2401 163 2451 181
rect 2435 129 2451 163
rect 2401 95 2451 129
rect 2435 61 2451 95
rect 2401 17 2451 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2484 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
<< metal1 >>
rect 0 561 2484 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2484 561
rect 0 496 2484 527
rect 0 17 2484 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2484 17
rect 0 -48 2484 -17
<< labels >>
flabel corelocali s 305 221 339 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 1593 221 1627 255 0 FreeSans 200 0 0 0 C
port 3 nsew
flabel corelocali s 2053 221 2087 255 0 FreeSans 200 0 0 0 D
port 4 nsew
flabel corelocali s 857 221 891 255 0 FreeSans 200 0 0 0 B
port 2 nsew
flabel corelocali s 2329 221 2363 255 0 FreeSans 200 0 0 0 Y
port 9 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
rlabel comment s 0 0 0 0 4 nor4_6
<< properties >>
string FIXED_BBOX 0 0 2484 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3497046
string GDS_START 3479092
<< end >>
