magic
tech sky130A
magscale 1 2
timestamp 1604502741
<< locali >>
rect 113 424 179 547
rect 585 424 651 547
rect 113 390 651 424
rect 585 364 651 390
rect 25 270 263 356
rect 297 270 363 356
rect 409 270 551 356
rect 585 236 619 364
rect 697 270 839 356
rect 889 270 1223 356
rect 109 202 619 236
rect 109 122 175 202
rect 309 122 375 202
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 23 581 253 615
rect 23 390 73 581
rect 219 492 253 581
rect 293 526 343 649
rect 383 492 449 596
rect 219 458 449 492
rect 495 581 921 615
rect 495 458 545 581
rect 691 390 725 581
rect 765 424 815 547
rect 855 458 921 581
rect 967 458 1033 649
rect 1067 424 1134 596
rect 765 390 1134 424
rect 1174 390 1224 649
rect 23 85 73 226
rect 661 202 1225 236
rect 209 85 275 165
rect 661 168 727 202
rect 409 134 727 168
rect 409 85 475 134
rect 23 51 475 85
rect 511 17 625 100
rect 661 70 727 134
rect 761 17 827 160
rect 861 70 927 202
rect 961 17 1125 161
rect 1159 70 1225 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
<< metal1 >>
rect 0 683 1248 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 0 617 1248 649
rect 0 17 1248 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
rect 0 -49 1248 -17
<< labels >>
rlabel locali s 889 270 1223 356 6 A1
port 1 nsew signal input
rlabel locali s 697 270 839 356 6 A2
port 2 nsew signal input
rlabel locali s 409 270 551 356 6 A3
port 3 nsew signal input
rlabel locali s 297 270 363 356 6 B1
port 4 nsew signal input
rlabel locali s 25 270 263 356 6 B2
port 5 nsew signal input
rlabel locali s 585 424 651 547 6 Y
port 6 nsew signal output
rlabel locali s 585 364 651 390 6 Y
port 6 nsew signal output
rlabel locali s 585 236 619 364 6 Y
port 6 nsew signal output
rlabel locali s 309 122 375 202 6 Y
port 6 nsew signal output
rlabel locali s 113 424 179 547 6 Y
port 6 nsew signal output
rlabel locali s 113 390 651 424 6 Y
port 6 nsew signal output
rlabel locali s 109 202 619 236 6 Y
port 6 nsew signal output
rlabel locali s 109 122 175 202 6 Y
port 6 nsew signal output
rlabel metal1 s 0 -49 1248 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 617 1248 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1248 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 638324
string GDS_START 627714
<< end >>
