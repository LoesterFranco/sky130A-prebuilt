magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 460 561
rect 18 333 85 490
rect 18 299 135 333
rect 206 323 257 490
rect 17 149 67 265
rect 101 165 135 299
rect 169 283 257 323
rect 169 199 215 283
rect 291 249 339 490
rect 391 367 443 527
rect 249 215 339 249
rect 101 131 341 165
rect 391 131 443 333
rect 101 129 172 131
rect 17 17 69 115
rect 119 77 172 129
rect 207 17 273 97
rect 307 77 341 131
rect 375 17 441 97
rect 0 -17 460 17
<< metal1 >>
rect 0 496 460 592
rect 0 -48 460 48
<< labels >>
rlabel locali s 391 131 443 333 6 A
port 1 nsew signal input
rlabel locali s 291 249 339 490 6 B
port 2 nsew signal input
rlabel locali s 249 215 339 249 6 B
port 2 nsew signal input
rlabel locali s 206 323 257 490 6 C
port 3 nsew signal input
rlabel locali s 169 283 257 323 6 C
port 3 nsew signal input
rlabel locali s 169 199 215 283 6 C
port 3 nsew signal input
rlabel locali s 17 149 67 265 6 D
port 4 nsew signal input
rlabel locali s 307 77 341 131 6 Y
port 5 nsew signal output
rlabel locali s 119 77 172 129 6 Y
port 5 nsew signal output
rlabel locali s 101 165 135 299 6 Y
port 5 nsew signal output
rlabel locali s 101 131 341 165 6 Y
port 5 nsew signal output
rlabel locali s 101 129 172 131 6 Y
port 5 nsew signal output
rlabel locali s 18 333 85 490 6 Y
port 5 nsew signal output
rlabel locali s 18 299 135 333 6 Y
port 5 nsew signal output
rlabel locali s 375 17 441 97 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 207 17 273 97 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 17 17 69 115 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 460 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 460 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 391 367 443 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 460 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 460 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 460 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1142854
string GDS_START 1138134
<< end >>
