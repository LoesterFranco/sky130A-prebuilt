magic
tech sky130A
magscale 1 2
timestamp 1601050088
<< locali >>
rect 377 446 433 547
rect 579 446 629 547
rect 377 412 629 446
rect 377 370 433 412
rect 377 350 411 370
rect 107 336 411 350
rect 37 316 411 336
rect 37 302 141 316
rect 37 282 71 302
rect 25 168 71 282
rect 217 268 359 282
rect 158 236 359 268
rect 729 236 795 310
rect 158 202 795 236
rect 950 236 1031 365
rect 25 134 762 168
rect 412 106 478 134
rect 712 102 762 134
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 23 370 73 649
rect 113 418 179 596
rect 219 452 253 649
rect 293 581 729 615
rect 293 418 343 581
rect 113 384 343 418
rect 473 480 539 581
rect 663 412 729 581
rect 763 412 829 649
rect 870 399 936 575
rect 976 399 1026 649
rect 870 378 916 399
rect 611 344 916 378
rect 611 336 645 344
rect 445 270 645 336
rect 882 202 916 344
rect 310 17 376 100
rect 514 17 676 100
rect 798 17 848 168
rect 882 69 1033 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 683 1056 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 0 617 1056 649
rect 0 17 1056 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -49 1056 -17
<< labels >>
rlabel locali s 729 236 795 310 6 A
port 1 nsew signal input
rlabel locali s 217 268 359 282 6 A
port 1 nsew signal input
rlabel locali s 158 236 359 268 6 A
port 1 nsew signal input
rlabel locali s 158 202 795 236 6 A
port 1 nsew signal input
rlabel locali s 950 236 1031 365 6 B_N
port 2 nsew signal input
rlabel locali s 712 102 762 134 6 Y
port 3 nsew signal output
rlabel locali s 579 446 629 547 6 Y
port 3 nsew signal output
rlabel locali s 412 106 478 134 6 Y
port 3 nsew signal output
rlabel locali s 377 446 433 547 6 Y
port 3 nsew signal output
rlabel locali s 377 412 629 446 6 Y
port 3 nsew signal output
rlabel locali s 377 370 433 412 6 Y
port 3 nsew signal output
rlabel locali s 377 350 411 370 6 Y
port 3 nsew signal output
rlabel locali s 107 336 411 350 6 Y
port 3 nsew signal output
rlabel locali s 37 316 411 336 6 Y
port 3 nsew signal output
rlabel locali s 37 302 141 316 6 Y
port 3 nsew signal output
rlabel locali s 37 282 71 302 6 Y
port 3 nsew signal output
rlabel locali s 25 168 71 282 6 Y
port 3 nsew signal output
rlabel locali s 25 134 762 168 6 Y
port 3 nsew signal output
rlabel metal1 s 0 -49 1056 49 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 617 1056 715 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1056 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1546732
string GDS_START 1538454
<< end >>
