magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1472 561
rect 119 289 257 527
rect 291 333 357 493
rect 391 367 425 527
rect 459 401 525 493
rect 559 435 593 527
rect 627 401 693 493
rect 459 333 693 401
rect 727 367 761 527
rect 795 333 861 493
rect 895 367 1033 527
rect 1067 333 1133 493
rect 1167 367 1201 527
rect 1235 333 1301 493
rect 291 289 1301 333
rect 1335 289 1401 527
rect 86 215 156 255
rect 559 215 620 289
rect 654 215 896 255
rect 958 215 1300 255
rect 559 181 593 215
rect 291 127 593 181
rect 119 17 169 109
rect 983 17 1033 109
rect 1167 17 1201 109
rect 1335 17 1401 181
rect 0 -17 1472 17
<< obsli1 >>
rect 17 289 85 493
rect 17 181 52 289
rect 201 215 525 255
rect 201 181 257 215
rect 17 143 257 181
rect 17 51 85 143
rect 627 143 1301 181
rect 627 127 945 143
rect 207 51 945 93
rect 1067 51 1133 143
rect 1235 51 1301 143
<< metal1 >>
rect 0 496 1472 592
rect 0 -48 1472 48
<< labels >>
rlabel locali s 86 215 156 255 6 A_N
port 1 nsew signal input
rlabel locali s 654 215 896 255 6 B
port 2 nsew signal input
rlabel locali s 958 215 1300 255 6 C
port 3 nsew signal input
rlabel locali s 1235 333 1301 493 6 Y
port 4 nsew signal output
rlabel locali s 1067 333 1133 493 6 Y
port 4 nsew signal output
rlabel locali s 795 333 861 493 6 Y
port 4 nsew signal output
rlabel locali s 627 401 693 493 6 Y
port 4 nsew signal output
rlabel locali s 559 215 620 289 6 Y
port 4 nsew signal output
rlabel locali s 559 181 593 215 6 Y
port 4 nsew signal output
rlabel locali s 459 401 525 493 6 Y
port 4 nsew signal output
rlabel locali s 459 333 693 401 6 Y
port 4 nsew signal output
rlabel locali s 291 333 357 493 6 Y
port 4 nsew signal output
rlabel locali s 291 289 1301 333 6 Y
port 4 nsew signal output
rlabel locali s 291 127 593 181 6 Y
port 4 nsew signal output
rlabel locali s 1335 17 1401 181 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 1167 17 1201 109 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 983 17 1033 109 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 119 17 169 109 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 1472 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1472 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 1335 289 1401 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 1167 367 1201 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 895 367 1033 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 727 367 761 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 559 435 593 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 391 367 425 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 119 289 257 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 1472 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 1472 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1472 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1836116
string GDS_START 1824330
<< end >>
