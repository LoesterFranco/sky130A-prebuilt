magic
tech sky130A
magscale 1 2
timestamp 1601050056
<< nwell >>
rect -38 332 1286 704
<< pwell >>
rect 0 0 1248 49
<< scpmos >>
rect 121 368 157 592
rect 211 368 247 592
rect 301 368 337 592
rect 391 368 427 592
rect 481 368 517 592
rect 571 368 607 592
rect 661 368 697 592
rect 751 368 787 592
rect 841 368 877 592
rect 931 368 967 592
rect 1021 368 1057 592
rect 1111 368 1147 592
<< nmoslvt >>
rect 137 74 167 222
rect 223 74 253 222
rect 309 74 339 222
rect 395 74 425 222
rect 481 74 511 222
rect 567 74 597 222
rect 653 74 683 222
rect 739 74 769 222
rect 941 74 971 222
rect 1027 74 1057 222
<< ndiff >>
rect 84 210 137 222
rect 84 176 92 210
rect 126 176 137 210
rect 84 120 137 176
rect 84 86 92 120
rect 126 86 137 120
rect 84 74 137 86
rect 167 136 223 222
rect 167 102 178 136
rect 212 102 223 136
rect 167 74 223 102
rect 253 210 309 222
rect 253 176 264 210
rect 298 176 309 210
rect 253 120 309 176
rect 253 86 264 120
rect 298 86 309 120
rect 253 74 309 86
rect 339 136 395 222
rect 339 102 350 136
rect 384 102 395 136
rect 339 74 395 102
rect 425 210 481 222
rect 425 176 436 210
rect 470 176 481 210
rect 425 120 481 176
rect 425 86 436 120
rect 470 86 481 120
rect 425 74 481 86
rect 511 189 567 222
rect 511 155 522 189
rect 556 155 567 189
rect 511 74 567 155
rect 597 123 653 222
rect 597 89 608 123
rect 642 89 653 123
rect 597 74 653 89
rect 683 210 739 222
rect 683 176 694 210
rect 728 176 739 210
rect 683 74 739 176
rect 769 123 826 222
rect 769 89 780 123
rect 814 89 826 123
rect 769 74 826 89
rect 888 210 941 222
rect 888 176 896 210
rect 930 176 941 210
rect 888 120 941 176
rect 888 86 896 120
rect 930 86 941 120
rect 888 74 941 86
rect 971 136 1027 222
rect 971 102 982 136
rect 1016 102 1027 136
rect 971 74 1027 102
rect 1057 210 1110 222
rect 1057 176 1068 210
rect 1102 176 1110 210
rect 1057 120 1110 176
rect 1057 86 1068 120
rect 1102 86 1110 120
rect 1057 74 1110 86
<< pdiff >>
rect 69 580 121 592
rect 69 546 77 580
rect 111 546 121 580
rect 69 497 121 546
rect 69 463 77 497
rect 111 463 121 497
rect 69 414 121 463
rect 69 380 77 414
rect 111 380 121 414
rect 69 368 121 380
rect 157 580 211 592
rect 157 546 167 580
rect 201 546 211 580
rect 157 508 211 546
rect 157 474 167 508
rect 201 474 211 508
rect 157 368 211 474
rect 247 580 301 592
rect 247 546 257 580
rect 291 546 301 580
rect 247 510 301 546
rect 247 476 257 510
rect 291 476 301 510
rect 247 440 301 476
rect 247 406 257 440
rect 291 406 301 440
rect 247 368 301 406
rect 337 580 391 592
rect 337 546 347 580
rect 381 546 391 580
rect 337 508 391 546
rect 337 474 347 508
rect 381 474 391 508
rect 337 368 391 474
rect 427 580 481 592
rect 427 546 437 580
rect 471 546 481 580
rect 427 510 481 546
rect 427 476 437 510
rect 471 476 481 510
rect 427 440 481 476
rect 427 406 437 440
rect 471 406 481 440
rect 427 368 481 406
rect 517 578 571 592
rect 517 544 527 578
rect 561 544 571 578
rect 517 368 571 544
rect 607 580 661 592
rect 607 546 617 580
rect 651 546 661 580
rect 607 508 661 546
rect 607 474 617 508
rect 651 474 661 508
rect 607 368 661 474
rect 697 578 751 592
rect 697 544 707 578
rect 741 544 751 578
rect 697 368 751 544
rect 787 580 841 592
rect 787 546 797 580
rect 831 546 841 580
rect 787 508 841 546
rect 787 474 797 508
rect 831 474 841 508
rect 787 368 841 474
rect 877 531 931 592
rect 877 497 887 531
rect 921 497 931 531
rect 877 440 931 497
rect 877 406 887 440
rect 921 406 931 440
rect 877 368 931 406
rect 967 580 1021 592
rect 967 546 977 580
rect 1011 546 1021 580
rect 967 508 1021 546
rect 967 474 977 508
rect 1011 474 1021 508
rect 967 368 1021 474
rect 1057 531 1111 592
rect 1057 497 1067 531
rect 1101 497 1111 531
rect 1057 440 1111 497
rect 1057 406 1067 440
rect 1101 406 1111 440
rect 1057 368 1111 406
rect 1147 580 1199 592
rect 1147 546 1157 580
rect 1191 546 1199 580
rect 1147 497 1199 546
rect 1147 463 1157 497
rect 1191 463 1199 497
rect 1147 414 1199 463
rect 1147 380 1157 414
rect 1191 380 1199 414
rect 1147 368 1199 380
<< ndiffc >>
rect 92 176 126 210
rect 92 86 126 120
rect 178 102 212 136
rect 264 176 298 210
rect 264 86 298 120
rect 350 102 384 136
rect 436 176 470 210
rect 436 86 470 120
rect 522 155 556 189
rect 608 89 642 123
rect 694 176 728 210
rect 780 89 814 123
rect 896 176 930 210
rect 896 86 930 120
rect 982 102 1016 136
rect 1068 176 1102 210
rect 1068 86 1102 120
<< pdiffc >>
rect 77 546 111 580
rect 77 463 111 497
rect 77 380 111 414
rect 167 546 201 580
rect 167 474 201 508
rect 257 546 291 580
rect 257 476 291 510
rect 257 406 291 440
rect 347 546 381 580
rect 347 474 381 508
rect 437 546 471 580
rect 437 476 471 510
rect 437 406 471 440
rect 527 544 561 578
rect 617 546 651 580
rect 617 474 651 508
rect 707 544 741 578
rect 797 546 831 580
rect 797 474 831 508
rect 887 497 921 531
rect 887 406 921 440
rect 977 546 1011 580
rect 977 474 1011 508
rect 1067 497 1101 531
rect 1067 406 1101 440
rect 1157 546 1191 580
rect 1157 463 1191 497
rect 1157 380 1191 414
<< poly >>
rect 121 592 157 618
rect 211 592 247 618
rect 301 592 337 618
rect 391 592 427 618
rect 481 592 517 618
rect 571 592 607 618
rect 661 592 697 618
rect 751 592 787 618
rect 841 592 877 618
rect 931 592 967 618
rect 1021 592 1057 618
rect 1111 592 1147 618
rect 121 336 157 368
rect 211 336 247 368
rect 301 336 337 368
rect 391 336 427 368
rect 121 320 427 336
rect 121 286 173 320
rect 207 286 241 320
rect 275 286 309 320
rect 343 286 377 320
rect 411 286 427 320
rect 121 270 427 286
rect 481 336 517 368
rect 571 336 607 368
rect 661 336 697 368
rect 751 336 787 368
rect 841 336 877 368
rect 931 336 967 368
rect 1021 336 1057 368
rect 1111 336 1147 368
rect 481 320 787 336
rect 481 286 601 320
rect 635 286 669 320
rect 703 286 737 320
rect 771 286 787 320
rect 481 270 787 286
rect 847 320 1147 336
rect 847 286 863 320
rect 897 286 931 320
rect 965 286 999 320
rect 1033 306 1147 320
rect 1033 286 1057 306
rect 847 270 1057 286
rect 137 222 167 270
rect 223 222 253 270
rect 309 222 339 270
rect 395 222 425 270
rect 481 222 511 270
rect 567 222 597 270
rect 653 222 683 270
rect 739 222 769 270
rect 941 222 971 270
rect 1027 222 1057 270
rect 137 48 167 74
rect 223 48 253 74
rect 309 48 339 74
rect 395 48 425 74
rect 481 48 511 74
rect 567 48 597 74
rect 653 48 683 74
rect 739 48 769 74
rect 941 48 971 74
rect 1027 48 1057 74
<< polycont >>
rect 173 286 207 320
rect 241 286 275 320
rect 309 286 343 320
rect 377 286 411 320
rect 601 286 635 320
rect 669 286 703 320
rect 737 286 771 320
rect 863 286 897 320
rect 931 286 965 320
rect 999 286 1033 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 61 580 111 596
rect 61 546 77 580
rect 61 497 111 546
rect 61 463 77 497
rect 61 424 111 463
rect 151 580 201 649
rect 151 546 167 580
rect 151 508 201 546
rect 151 474 167 508
rect 151 458 201 474
rect 241 580 307 596
rect 241 546 257 580
rect 291 546 307 580
rect 241 510 307 546
rect 241 476 257 510
rect 291 476 307 510
rect 241 440 307 476
rect 347 580 381 649
rect 347 508 381 546
rect 347 458 381 474
rect 421 580 471 596
rect 421 546 437 580
rect 421 510 471 546
rect 511 578 561 649
rect 511 544 527 578
rect 511 526 561 544
rect 601 580 667 596
rect 601 546 617 580
rect 651 546 667 580
rect 421 476 437 510
rect 601 508 667 546
rect 707 578 741 649
rect 707 526 741 544
rect 781 581 1207 615
rect 781 580 831 581
rect 781 546 797 580
rect 977 580 1011 581
rect 601 492 617 508
rect 471 476 617 492
rect 421 474 617 476
rect 651 492 667 508
rect 781 508 831 546
rect 781 492 797 508
rect 651 474 797 492
rect 421 458 831 474
rect 871 531 937 547
rect 871 497 887 531
rect 921 497 937 531
rect 241 424 257 440
rect 61 414 257 424
rect 61 380 77 414
rect 111 406 257 414
rect 291 424 307 440
rect 421 440 471 458
rect 421 424 437 440
rect 291 406 437 424
rect 871 440 937 497
rect 1157 580 1207 581
rect 977 508 1011 546
rect 977 458 1011 474
rect 1051 531 1117 547
rect 1051 497 1067 531
rect 1101 497 1117 531
rect 871 424 887 440
rect 111 390 471 406
rect 505 406 887 424
rect 921 424 937 440
rect 1051 440 1117 497
rect 1051 424 1067 440
rect 921 406 1067 424
rect 1101 406 1117 440
rect 505 390 1117 406
rect 1191 546 1207 580
rect 1157 497 1207 546
rect 1191 463 1207 497
rect 1157 414 1207 463
rect 61 364 111 380
rect 157 320 455 356
rect 157 286 173 320
rect 207 286 241 320
rect 275 286 309 320
rect 343 286 377 320
rect 411 286 455 320
rect 157 270 455 286
rect 505 236 551 390
rect 1191 380 1207 414
rect 1157 364 1207 380
rect 585 320 787 356
rect 585 286 601 320
rect 635 286 669 320
rect 703 286 737 320
rect 771 286 787 320
rect 585 270 787 286
rect 847 320 1049 356
rect 847 286 863 320
rect 897 286 931 320
rect 965 286 999 320
rect 1033 286 1049 320
rect 847 270 1049 286
rect 76 210 470 236
rect 76 176 92 210
rect 126 202 264 210
rect 76 120 126 176
rect 298 202 436 210
rect 76 86 92 120
rect 76 70 126 86
rect 162 136 228 168
rect 162 102 178 136
rect 212 102 228 136
rect 162 17 228 102
rect 264 120 298 176
rect 264 70 298 86
rect 334 136 400 168
rect 334 102 350 136
rect 384 102 400 136
rect 334 17 400 102
rect 436 120 470 176
rect 505 210 1118 236
rect 505 189 694 210
rect 505 155 522 189
rect 556 176 694 189
rect 728 176 896 210
rect 930 202 1068 210
rect 505 119 556 155
rect 592 123 658 142
rect 436 85 470 86
rect 592 89 608 123
rect 642 89 658 123
rect 592 85 658 89
rect 764 123 830 142
rect 764 89 780 123
rect 814 89 830 123
rect 764 85 830 89
rect 436 51 830 85
rect 880 120 930 176
rect 1102 176 1118 210
rect 880 86 896 120
rect 880 70 930 86
rect 966 136 1032 168
rect 966 102 982 136
rect 1016 102 1032 136
rect 966 17 1032 102
rect 1068 120 1118 176
rect 1102 86 1118 120
rect 1068 70 1118 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
<< metal1 >>
rect 0 683 1248 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 0 617 1248 649
rect 0 17 1248 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
rect 0 -49 1248 -17
<< labels >>
flabel pwell s 0 0 1248 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 1248 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
rlabel comment s 0 0 0 0 4 a21oi_4
flabel metal1 s 0 617 1248 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 1248 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 511 168 545 202 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 511 242 545 276 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 1248 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 4018290
string GDS_START 4008392
<< end >>
