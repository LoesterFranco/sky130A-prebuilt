magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1932 561
rect 103 451 169 527
rect 647 451 713 527
rect 30 199 99 323
rect 161 199 248 323
rect 103 17 169 93
rect 653 199 713 399
rect 1012 451 1078 527
rect 1196 451 1266 527
rect 960 211 1009 335
rect 1050 211 1116 335
rect 1211 199 1269 335
rect 560 17 618 161
rect 1030 17 1064 109
rect 1763 451 1829 527
rect 1202 17 1268 93
rect 1779 17 1813 109
rect 1863 51 1915 493
rect 0 -17 1932 17
<< obsli1 >>
rect 35 393 69 493
rect 203 459 509 493
rect 203 427 237 459
rect 307 393 341 425
rect 35 359 341 393
rect 375 391 441 425
rect 375 325 409 391
rect 475 359 509 459
rect 543 325 613 493
rect 765 459 967 493
rect 282 291 409 325
rect 282 187 316 291
rect 452 279 613 325
rect 452 257 524 279
rect 416 255 524 257
rect 416 221 490 255
rect 35 127 237 161
rect 35 52 69 127
rect 203 85 237 127
rect 282 153 306 187
rect 282 119 350 153
rect 384 85 418 152
rect 452 86 524 221
rect 765 357 799 459
rect 833 391 899 425
rect 833 357 865 391
rect 933 417 967 459
rect 1112 417 1146 493
rect 1300 427 1337 493
rect 933 383 1146 417
rect 833 323 899 357
rect 747 289 899 323
rect 747 184 781 289
rect 815 221 858 253
rect 815 219 881 221
rect 1303 255 1337 427
rect 1396 427 1438 493
rect 1472 459 1729 493
rect 1472 451 1538 459
rect 1303 221 1327 255
rect 747 169 810 184
rect 203 51 418 85
rect 676 85 710 159
rect 744 119 810 169
rect 844 177 878 185
rect 844 143 1148 177
rect 844 119 878 143
rect 925 85 996 93
rect 676 51 996 85
rect 1099 59 1148 143
rect 1303 131 1337 221
rect 1396 187 1430 427
rect 1569 397 1635 425
rect 1478 391 1635 397
rect 1478 357 1511 391
rect 1545 357 1635 391
rect 1478 351 1635 357
rect 1695 367 1729 459
rect 1396 153 1410 187
rect 1302 65 1337 131
rect 1478 117 1512 351
rect 1695 333 1825 367
rect 1638 221 1695 255
rect 1628 185 1676 187
rect 1628 153 1677 185
rect 1791 177 1825 333
rect 1642 119 1677 153
rect 1711 143 1825 177
rect 1406 83 1512 117
rect 1546 85 1580 117
rect 1711 85 1745 143
rect 1406 51 1440 83
rect 1546 51 1745 85
<< obsli1c >>
rect 490 221 524 255
rect 306 153 340 187
rect 865 357 899 391
rect 858 221 892 255
rect 1327 221 1361 255
rect 1511 357 1545 391
rect 1410 153 1444 187
rect 1695 221 1729 255
rect 1594 153 1628 187
<< metal1 >>
rect 0 496 1932 592
rect 0 -48 1932 48
<< obsm1 >>
rect 853 391 911 397
rect 853 357 865 391
rect 899 388 911 391
rect 1499 391 1557 397
rect 1499 388 1511 391
rect 899 360 1511 388
rect 899 357 911 360
rect 853 351 911 357
rect 1499 357 1511 360
rect 1545 357 1557 391
rect 1499 351 1557 357
rect 478 255 536 261
rect 478 221 490 255
rect 524 252 536 255
rect 846 255 904 261
rect 846 252 858 255
rect 524 224 858 252
rect 524 221 536 224
rect 478 215 536 221
rect 846 221 858 224
rect 892 221 904 255
rect 846 215 904 221
rect 1315 255 1373 261
rect 1315 221 1327 255
rect 1361 252 1373 255
rect 1683 255 1741 261
rect 1683 252 1695 255
rect 1361 224 1695 252
rect 1361 221 1373 224
rect 1315 215 1373 221
rect 1683 221 1695 224
rect 1729 221 1741 255
rect 1683 215 1741 221
rect 294 187 352 193
rect 294 153 306 187
rect 340 184 352 187
rect 1398 187 1456 193
rect 1398 184 1410 187
rect 340 156 1410 184
rect 340 153 352 156
rect 294 147 352 153
rect 1398 153 1410 156
rect 1444 184 1456 187
rect 1582 187 1640 193
rect 1582 184 1594 187
rect 1444 156 1594 184
rect 1444 153 1456 156
rect 1398 147 1456 153
rect 1582 153 1594 156
rect 1628 153 1640 187
rect 1582 147 1640 153
<< labels >>
rlabel locali s 161 199 248 323 6 A0
port 1 nsew signal input
rlabel locali s 30 199 99 323 6 A1
port 2 nsew signal input
rlabel locali s 1050 211 1116 335 6 A2
port 3 nsew signal input
rlabel locali s 960 211 1009 335 6 A3
port 4 nsew signal input
rlabel locali s 653 199 713 399 6 S0
port 5 nsew signal input
rlabel locali s 1211 199 1269 335 6 S1
port 6 nsew signal input
rlabel locali s 1863 51 1915 493 6 X
port 7 nsew signal output
rlabel locali s 1779 17 1813 109 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 1202 17 1268 93 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 1030 17 1064 109 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 560 17 618 161 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 103 17 169 93 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 0 -17 1932 17 8 VGND
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1932 48 8 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 1763 451 1829 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 1196 451 1266 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 1012 451 1078 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 647 451 713 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 103 451 169 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 0 527 1932 561 6 VPWR
port 9 nsew power bidirectional abutment
rlabel metal1 s 0 496 1932 592 6 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1932 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1749730
string GDS_START 1734254
<< end >>
