magic
tech sky130A
magscale 1 2
timestamp 1599588209
<< nwell >>
rect -38 332 1862 704
<< pwell >>
rect 0 0 1824 49
<< scpmos >>
rect 86 392 116 560
rect 210 392 240 560
rect 422 392 452 560
rect 536 392 566 592
rect 620 392 650 592
rect 727 508 757 592
rect 858 508 888 592
rect 1010 368 1040 592
rect 1110 368 1140 592
rect 1216 368 1246 592
rect 1306 368 1336 592
rect 1508 368 1538 568
rect 1618 368 1648 592
rect 1708 368 1738 592
<< nmoslvt >>
rect 84 112 114 222
rect 200 74 230 222
rect 420 82 450 230
rect 539 80 569 208
rect 611 80 641 208
rect 743 124 773 208
rect 821 124 851 208
rect 1019 74 1049 222
rect 1097 74 1127 222
rect 1205 74 1235 222
rect 1291 74 1321 222
rect 1510 94 1540 222
rect 1624 74 1654 222
rect 1710 74 1740 222
<< ndiff >>
rect 27 184 84 222
rect 27 150 39 184
rect 73 150 84 184
rect 27 112 84 150
rect 114 200 200 222
rect 114 166 141 200
rect 175 166 200 200
rect 114 120 200 166
rect 114 112 141 120
rect 129 86 141 112
rect 175 86 200 120
rect 129 74 200 86
rect 230 200 287 222
rect 230 166 241 200
rect 275 166 287 200
rect 230 120 287 166
rect 230 86 241 120
rect 275 86 287 120
rect 230 74 287 86
rect 363 218 420 230
rect 363 184 375 218
rect 409 184 420 218
rect 363 82 420 184
rect 450 208 500 230
rect 962 210 1019 222
rect 450 82 539 208
rect 465 48 477 82
rect 511 80 539 82
rect 569 80 611 208
rect 641 192 743 208
rect 641 158 675 192
rect 709 158 743 192
rect 641 124 743 158
rect 773 124 821 208
rect 851 183 908 208
rect 851 149 862 183
rect 896 149 908 183
rect 851 124 908 149
rect 962 176 974 210
rect 1008 176 1019 210
rect 641 80 691 124
rect 962 120 1019 176
rect 511 48 524 80
rect 465 36 524 48
rect 962 86 974 120
rect 1008 86 1019 120
rect 962 74 1019 86
rect 1049 74 1097 222
rect 1127 197 1205 222
rect 1127 163 1138 197
rect 1172 163 1205 197
rect 1127 120 1205 163
rect 1127 86 1138 120
rect 1172 86 1205 120
rect 1127 74 1205 86
rect 1235 210 1291 222
rect 1235 176 1246 210
rect 1280 176 1291 210
rect 1235 120 1291 176
rect 1235 86 1246 120
rect 1280 86 1291 120
rect 1235 74 1291 86
rect 1321 139 1392 222
rect 1321 105 1346 139
rect 1380 105 1392 139
rect 1321 74 1392 105
rect 1453 210 1510 222
rect 1453 176 1465 210
rect 1499 176 1510 210
rect 1453 140 1510 176
rect 1453 106 1465 140
rect 1499 106 1510 140
rect 1453 94 1510 106
rect 1540 210 1624 222
rect 1540 176 1565 210
rect 1599 176 1624 210
rect 1540 140 1624 176
rect 1540 106 1565 140
rect 1599 106 1624 140
rect 1540 94 1624 106
rect 1574 74 1624 94
rect 1654 210 1710 222
rect 1654 176 1665 210
rect 1699 176 1710 210
rect 1654 120 1710 176
rect 1654 86 1665 120
rect 1699 86 1710 120
rect 1654 74 1710 86
rect 1740 210 1797 222
rect 1740 176 1751 210
rect 1785 176 1797 210
rect 1740 120 1797 176
rect 1740 86 1751 120
rect 1785 86 1797 120
rect 1740 74 1797 86
<< pdiff >>
rect 134 590 192 602
rect 134 560 146 590
rect 27 548 86 560
rect 27 514 39 548
rect 73 514 86 548
rect 27 440 86 514
rect 27 406 39 440
rect 73 406 86 440
rect 27 392 86 406
rect 116 556 146 560
rect 180 560 192 590
rect 470 574 536 592
rect 470 560 485 574
rect 180 556 210 560
rect 116 392 210 556
rect 240 438 309 560
rect 240 404 258 438
rect 292 404 309 438
rect 240 392 309 404
rect 363 438 422 560
rect 363 404 375 438
rect 409 404 422 438
rect 363 392 422 404
rect 452 540 485 560
rect 519 540 536 574
rect 452 392 536 540
rect 566 392 620 592
rect 650 531 727 592
rect 650 497 663 531
rect 697 508 727 531
rect 757 508 858 592
rect 888 580 1010 592
rect 888 546 932 580
rect 966 546 1010 580
rect 888 508 1010 546
rect 697 497 709 508
rect 650 439 709 497
rect 650 405 663 439
rect 697 405 709 439
rect 650 392 709 405
rect 957 368 1010 508
rect 1040 580 1110 592
rect 1040 546 1063 580
rect 1097 546 1110 580
rect 1040 497 1110 546
rect 1040 463 1063 497
rect 1097 463 1110 497
rect 1040 414 1110 463
rect 1040 380 1063 414
rect 1097 380 1110 414
rect 1040 368 1110 380
rect 1140 582 1216 592
rect 1140 548 1163 582
rect 1197 548 1216 582
rect 1140 514 1216 548
rect 1140 480 1163 514
rect 1197 480 1216 514
rect 1140 446 1216 480
rect 1140 412 1163 446
rect 1197 412 1216 446
rect 1140 368 1216 412
rect 1246 580 1306 592
rect 1246 546 1259 580
rect 1293 546 1306 580
rect 1246 497 1306 546
rect 1246 463 1259 497
rect 1293 463 1306 497
rect 1246 414 1306 463
rect 1246 380 1259 414
rect 1293 380 1306 414
rect 1246 368 1306 380
rect 1336 580 1395 592
rect 1336 546 1349 580
rect 1383 546 1395 580
rect 1565 568 1618 592
rect 1336 478 1395 546
rect 1336 444 1349 478
rect 1383 444 1395 478
rect 1336 368 1395 444
rect 1449 556 1508 568
rect 1449 522 1461 556
rect 1495 522 1508 556
rect 1449 485 1508 522
rect 1449 451 1461 485
rect 1495 451 1508 485
rect 1449 414 1508 451
rect 1449 380 1461 414
rect 1495 380 1508 414
rect 1449 368 1508 380
rect 1538 556 1618 568
rect 1538 522 1561 556
rect 1595 522 1618 556
rect 1538 485 1618 522
rect 1538 451 1561 485
rect 1595 451 1618 485
rect 1538 414 1618 451
rect 1538 380 1561 414
rect 1595 380 1618 414
rect 1538 368 1618 380
rect 1648 580 1708 592
rect 1648 546 1661 580
rect 1695 546 1708 580
rect 1648 500 1708 546
rect 1648 466 1661 500
rect 1695 466 1708 500
rect 1648 414 1708 466
rect 1648 380 1661 414
rect 1695 380 1708 414
rect 1648 368 1708 380
rect 1738 580 1797 592
rect 1738 546 1751 580
rect 1785 546 1797 580
rect 1738 500 1797 546
rect 1738 466 1751 500
rect 1785 466 1797 500
rect 1738 414 1797 466
rect 1738 380 1751 414
rect 1785 380 1797 414
rect 1738 368 1797 380
<< ndiffc >>
rect 39 150 73 184
rect 141 166 175 200
rect 141 86 175 120
rect 241 166 275 200
rect 241 86 275 120
rect 375 184 409 218
rect 477 48 511 82
rect 675 158 709 192
rect 862 149 896 183
rect 974 176 1008 210
rect 974 86 1008 120
rect 1138 163 1172 197
rect 1138 86 1172 120
rect 1246 176 1280 210
rect 1246 86 1280 120
rect 1346 105 1380 139
rect 1465 176 1499 210
rect 1465 106 1499 140
rect 1565 176 1599 210
rect 1565 106 1599 140
rect 1665 176 1699 210
rect 1665 86 1699 120
rect 1751 176 1785 210
rect 1751 86 1785 120
<< pdiffc >>
rect 39 514 73 548
rect 39 406 73 440
rect 146 556 180 590
rect 258 404 292 438
rect 375 404 409 438
rect 485 540 519 574
rect 663 497 697 531
rect 932 546 966 580
rect 663 405 697 439
rect 1063 546 1097 580
rect 1063 463 1097 497
rect 1063 380 1097 414
rect 1163 548 1197 582
rect 1163 480 1197 514
rect 1163 412 1197 446
rect 1259 546 1293 580
rect 1259 463 1293 497
rect 1259 380 1293 414
rect 1349 546 1383 580
rect 1349 444 1383 478
rect 1461 522 1495 556
rect 1461 451 1495 485
rect 1461 380 1495 414
rect 1561 522 1595 556
rect 1561 451 1595 485
rect 1561 380 1595 414
rect 1661 546 1695 580
rect 1661 466 1695 500
rect 1661 380 1695 414
rect 1751 546 1785 580
rect 1751 466 1785 500
rect 1751 380 1785 414
<< poly >>
rect 536 592 566 618
rect 620 592 650 618
rect 727 592 757 618
rect 858 592 888 618
rect 1010 592 1040 618
rect 1110 592 1140 618
rect 1216 592 1246 618
rect 1306 592 1336 618
rect 86 560 116 586
rect 210 560 240 586
rect 422 560 452 586
rect 727 493 757 508
rect 858 493 888 508
rect 724 476 760 493
rect 724 460 807 476
rect 855 464 891 493
rect 724 426 757 460
rect 791 426 807 460
rect 724 410 807 426
rect 849 448 915 464
rect 849 414 865 448
rect 899 414 915 448
rect 849 398 915 414
rect 86 377 116 392
rect 210 377 240 392
rect 422 377 452 392
rect 536 377 566 392
rect 620 377 650 392
rect 83 356 119 377
rect 83 340 151 356
rect 83 306 101 340
rect 135 306 151 340
rect 207 310 243 377
rect 307 318 373 334
rect 83 290 151 306
rect 193 294 259 310
rect 84 222 114 290
rect 193 260 209 294
rect 243 260 259 294
rect 307 284 323 318
rect 357 298 373 318
rect 419 298 455 377
rect 533 360 569 377
rect 357 284 455 298
rect 497 344 569 360
rect 497 310 513 344
rect 547 310 569 344
rect 617 368 653 377
rect 617 338 773 368
rect 497 294 569 310
rect 307 268 455 284
rect 193 244 259 260
rect 420 245 455 268
rect 200 222 230 244
rect 420 230 450 245
rect 84 86 114 112
rect 539 208 569 294
rect 611 280 677 296
rect 611 246 627 280
rect 661 246 677 280
rect 611 230 677 246
rect 611 208 641 230
rect 743 208 773 338
rect 849 253 879 398
rect 1508 568 1538 594
rect 1618 592 1648 618
rect 1708 592 1738 618
rect 1010 353 1040 368
rect 1110 353 1140 368
rect 1216 353 1246 368
rect 1306 353 1336 368
rect 1508 353 1538 368
rect 1618 353 1648 368
rect 1708 353 1738 368
rect 1007 336 1043 353
rect 921 320 1043 336
rect 921 286 937 320
rect 971 300 1043 320
rect 1107 310 1143 353
rect 1213 326 1249 353
rect 1303 326 1339 353
rect 1505 326 1541 353
rect 1615 326 1651 353
rect 1705 326 1741 353
rect 1205 310 1541 326
rect 971 286 1049 300
rect 921 270 1049 286
rect 821 223 879 253
rect 821 208 851 223
rect 1019 222 1049 270
rect 1091 294 1157 310
rect 1091 260 1107 294
rect 1141 260 1157 294
rect 1091 244 1157 260
rect 1205 276 1221 310
rect 1255 276 1289 310
rect 1323 276 1541 310
rect 1205 260 1541 276
rect 1583 310 1741 326
rect 1583 276 1599 310
rect 1633 276 1741 310
rect 1583 260 1741 276
rect 1097 222 1127 244
rect 1205 222 1235 260
rect 1291 222 1321 260
rect 1510 222 1540 260
rect 1624 222 1654 260
rect 1710 222 1740 260
rect 200 48 230 74
rect 420 56 450 82
rect 743 102 773 124
rect 713 86 779 102
rect 821 98 851 124
rect 539 54 569 80
rect 611 54 641 80
rect 713 52 729 86
rect 763 52 779 86
rect 713 36 779 52
rect 1019 48 1049 74
rect 1097 48 1127 74
rect 1205 48 1235 74
rect 1291 48 1321 74
rect 1510 68 1540 94
rect 1624 48 1654 74
rect 1710 48 1740 74
<< polycont >>
rect 757 426 791 460
rect 865 414 899 448
rect 101 306 135 340
rect 209 260 243 294
rect 323 284 357 318
rect 513 310 547 344
rect 627 246 661 280
rect 937 286 971 320
rect 1107 260 1141 294
rect 1221 276 1255 310
rect 1289 276 1323 310
rect 1599 276 1633 310
rect 729 52 763 86
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 130 590 196 649
rect 17 548 89 564
rect 17 514 39 548
rect 73 514 89 548
rect 130 556 146 590
rect 180 556 196 590
rect 130 540 196 556
rect 466 574 539 649
rect 466 540 485 574
rect 519 540 539 574
rect 595 581 807 615
rect 17 506 89 514
rect 17 472 561 506
rect 17 440 89 472
rect 17 406 39 440
rect 73 406 89 440
rect 17 390 89 406
rect 237 404 258 438
rect 292 404 325 438
rect 17 226 51 390
rect 237 388 325 404
rect 359 404 375 438
rect 409 404 441 438
rect 359 388 441 404
rect 85 340 161 356
rect 85 306 101 340
rect 135 306 161 340
rect 291 334 325 388
rect 291 318 373 334
rect 85 290 161 306
rect 195 294 257 310
rect 195 260 209 294
rect 243 260 257 294
rect 195 236 257 260
rect 291 284 323 318
rect 357 284 373 318
rect 291 268 373 284
rect 17 184 89 226
rect 291 202 325 268
rect 407 260 441 388
rect 497 344 561 472
rect 497 310 513 344
rect 547 310 561 344
rect 497 294 561 310
rect 595 296 629 581
rect 663 531 697 547
rect 663 439 697 497
rect 741 460 807 581
rect 885 580 1013 649
rect 885 546 932 580
rect 966 546 1013 580
rect 885 530 1013 546
rect 1047 580 1113 596
rect 1047 546 1063 580
rect 1097 546 1113 580
rect 1047 497 1113 546
rect 1047 464 1063 497
rect 741 426 757 460
rect 791 426 807 460
rect 741 410 807 426
rect 849 463 1063 464
rect 1097 463 1113 497
rect 849 448 1113 463
rect 849 414 865 448
rect 899 414 1113 448
rect 663 364 697 405
rect 849 398 1063 414
rect 1019 380 1063 398
rect 1097 380 1113 414
rect 1147 582 1213 649
rect 1147 548 1163 582
rect 1197 548 1213 582
rect 1147 514 1213 548
rect 1147 480 1163 514
rect 1197 480 1213 514
rect 1147 446 1213 480
rect 1147 412 1163 446
rect 1197 412 1213 446
rect 1259 580 1293 596
rect 1259 497 1293 546
rect 1259 414 1293 463
rect 1333 580 1399 649
rect 1333 546 1349 580
rect 1383 546 1399 580
rect 1333 478 1399 546
rect 1333 444 1349 478
rect 1383 444 1399 478
rect 1333 428 1399 444
rect 1449 556 1511 572
rect 1449 522 1461 556
rect 1495 522 1511 556
rect 1449 485 1511 522
rect 1449 451 1461 485
rect 1495 451 1511 485
rect 1019 378 1113 380
rect 1449 414 1511 451
rect 1293 380 1415 394
rect 663 330 985 364
rect 595 280 677 296
rect 595 260 627 280
rect 407 246 627 260
rect 661 246 677 280
rect 407 234 677 246
rect 17 150 39 184
rect 73 150 89 184
rect 17 108 89 150
rect 125 200 191 202
rect 125 166 141 200
rect 175 166 191 200
rect 125 120 191 166
rect 125 86 141 120
rect 175 86 191 120
rect 125 17 191 86
rect 225 200 325 202
rect 225 166 241 200
rect 275 166 325 200
rect 359 226 677 234
rect 359 218 441 226
rect 359 184 375 218
rect 409 184 441 218
rect 714 192 748 330
rect 921 320 985 330
rect 921 286 937 320
rect 971 286 985 320
rect 921 270 985 286
rect 1019 344 1225 378
rect 1259 360 1415 380
rect 1019 226 1053 344
rect 1191 326 1225 344
rect 1191 310 1330 326
rect 1087 294 1157 310
rect 1087 260 1107 294
rect 1141 260 1157 294
rect 1191 276 1221 310
rect 1255 276 1289 310
rect 1323 276 1330 310
rect 1191 260 1330 276
rect 1087 236 1157 260
rect 1369 226 1415 360
rect 225 150 325 166
rect 636 158 675 192
rect 709 158 748 192
rect 846 183 912 212
rect 225 120 596 150
rect 225 86 241 120
rect 275 116 596 120
rect 275 86 325 116
rect 225 70 325 86
rect 562 102 596 116
rect 846 149 862 183
rect 896 149 912 183
rect 562 86 779 102
rect 461 48 477 82
rect 511 48 528 82
rect 562 52 729 86
rect 763 52 779 86
rect 562 51 779 52
rect 461 17 528 48
rect 846 17 912 149
rect 958 210 1053 226
rect 958 176 974 210
rect 1008 176 1053 210
rect 1230 210 1415 226
rect 958 120 1053 176
rect 958 86 974 120
rect 1008 86 1053 120
rect 958 70 1053 86
rect 1122 197 1188 202
rect 1122 163 1138 197
rect 1172 163 1188 197
rect 1122 120 1188 163
rect 1122 86 1138 120
rect 1172 86 1188 120
rect 1122 17 1188 86
rect 1230 176 1246 210
rect 1280 192 1415 210
rect 1449 380 1461 414
rect 1495 380 1511 414
rect 1449 326 1511 380
rect 1545 556 1611 649
rect 1545 522 1561 556
rect 1595 522 1611 556
rect 1545 485 1611 522
rect 1545 451 1561 485
rect 1595 451 1611 485
rect 1545 414 1611 451
rect 1545 380 1561 414
rect 1595 380 1611 414
rect 1545 364 1611 380
rect 1645 580 1717 596
rect 1645 546 1661 580
rect 1695 546 1717 580
rect 1645 500 1717 546
rect 1645 466 1661 500
rect 1695 466 1717 500
rect 1645 414 1717 466
rect 1645 380 1661 414
rect 1695 380 1717 414
rect 1645 364 1717 380
rect 1751 580 1801 649
rect 1785 546 1801 580
rect 1751 500 1801 546
rect 1785 466 1801 500
rect 1751 414 1801 466
rect 1785 380 1801 414
rect 1751 364 1801 380
rect 1449 310 1649 326
rect 1449 276 1599 310
rect 1633 276 1649 310
rect 1449 260 1649 276
rect 1449 226 1511 260
rect 1683 226 1717 364
rect 1449 210 1515 226
rect 1280 176 1296 192
rect 1230 120 1296 176
rect 1449 176 1465 210
rect 1499 176 1515 210
rect 1230 86 1246 120
rect 1280 86 1296 120
rect 1230 70 1296 86
rect 1330 139 1396 158
rect 1330 105 1346 139
rect 1380 105 1396 139
rect 1330 17 1396 105
rect 1449 140 1515 176
rect 1449 106 1465 140
rect 1499 106 1515 140
rect 1449 90 1515 106
rect 1549 210 1615 226
rect 1549 176 1565 210
rect 1599 176 1615 210
rect 1549 140 1615 176
rect 1549 106 1565 140
rect 1599 106 1615 140
rect 1549 17 1615 106
rect 1649 210 1717 226
rect 1649 176 1665 210
rect 1699 176 1717 210
rect 1649 120 1717 176
rect 1649 86 1665 120
rect 1699 86 1717 120
rect 1649 70 1717 86
rect 1751 210 1801 226
rect 1785 176 1801 210
rect 1751 120 1801 176
rect 1785 86 1801 120
rect 1751 17 1801 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
<< metal1 >>
rect 0 683 1824 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 0 617 1824 649
rect 0 17 1824 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
rect 0 -49 1824 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dlrbp_2
flabel pwell s 0 0 1824 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 0 617 1824 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 1824 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 1824 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 223 242 257 276 0 FreeSans 340 0 0 0 GATE
port 2 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 1 nsew
flabel corelocali s 1087 242 1121 276 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew
flabel corelocali s 1663 390 1697 424 0 FreeSans 340 0 0 0 Q_N
port 9 nsew
flabel corelocali s 1375 242 1409 276 0 FreeSans 340 0 0 0 Q
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 1824 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3128990
string GDS_START 3115200
<< end >>
