magic
tech sky130A
magscale 1 2
timestamp 1601050047
<< nwell >>
rect -38 332 1766 704
rect 300 311 1496 332
<< pwell >>
rect 0 0 1728 49
<< scpmos >>
rect 84 368 114 592
rect 187 368 217 568
rect 288 389 318 589
rect 389 347 419 547
rect 479 347 509 547
rect 576 347 606 547
rect 693 347 723 547
rect 794 347 824 547
rect 886 347 916 547
rect 987 347 1017 547
rect 1077 347 1107 547
rect 1196 347 1226 547
rect 1363 362 1393 562
rect 1614 368 1644 592
<< nmoslvt >>
rect 84 74 114 222
rect 207 75 237 203
rect 285 75 315 203
rect 363 75 393 203
rect 471 75 501 203
rect 573 75 603 203
rect 691 75 721 203
rect 777 75 807 203
rect 906 75 936 203
rect 984 75 1014 203
rect 1070 75 1100 203
rect 1282 75 1312 203
rect 1427 75 1457 203
rect 1617 74 1647 222
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 203 164 222
rect 114 82 207 203
rect 114 74 143 82
rect 129 48 143 74
rect 177 75 207 82
rect 237 75 285 203
rect 315 75 363 203
rect 393 127 471 203
rect 393 93 404 127
rect 438 93 471 127
rect 393 75 471 93
rect 501 134 573 203
rect 501 100 520 134
rect 554 100 573 134
rect 501 75 573 100
rect 603 82 691 203
rect 603 75 630 82
rect 177 48 192 75
rect 129 36 192 48
rect 618 48 630 75
rect 664 75 691 82
rect 721 134 777 203
rect 721 100 732 134
rect 766 100 777 134
rect 721 75 777 100
rect 807 126 906 203
rect 807 92 846 126
rect 880 92 906 126
rect 807 75 906 92
rect 936 75 984 203
rect 1014 137 1070 203
rect 1014 103 1025 137
rect 1059 103 1070 137
rect 1014 75 1070 103
rect 1100 85 1282 203
rect 1100 75 1127 85
rect 664 48 676 75
rect 1115 51 1127 75
rect 1161 51 1221 85
rect 1255 75 1282 85
rect 1312 78 1427 203
rect 1312 75 1366 78
rect 1255 51 1267 75
rect 618 36 676 48
rect 1115 39 1267 51
rect 1354 44 1366 75
rect 1400 75 1427 78
rect 1457 146 1510 203
rect 1457 112 1468 146
rect 1502 112 1510 146
rect 1457 75 1510 112
rect 1564 138 1617 222
rect 1564 104 1572 138
rect 1606 104 1617 138
rect 1400 44 1412 75
rect 1564 74 1617 104
rect 1647 210 1701 222
rect 1647 176 1658 210
rect 1692 176 1701 210
rect 1647 120 1701 176
rect 1647 86 1658 120
rect 1692 86 1701 120
rect 1647 74 1701 86
rect 1354 36 1412 44
<< pdiff >>
rect 27 580 84 592
rect 27 546 37 580
rect 71 546 84 580
rect 27 497 84 546
rect 27 463 37 497
rect 71 463 84 497
rect 27 414 84 463
rect 27 380 37 414
rect 71 380 84 414
rect 27 368 84 380
rect 114 580 169 592
rect 114 546 127 580
rect 161 568 169 580
rect 235 568 288 589
rect 161 546 187 568
rect 114 512 187 546
rect 114 478 127 512
rect 161 478 187 512
rect 114 444 187 478
rect 114 410 127 444
rect 161 410 187 444
rect 114 368 187 410
rect 217 389 288 568
rect 318 547 371 589
rect 624 576 675 588
rect 624 547 632 576
rect 318 389 389 547
rect 217 368 270 389
rect 336 347 389 389
rect 419 535 479 547
rect 419 501 432 535
rect 466 501 479 535
rect 419 467 479 501
rect 419 433 432 467
rect 466 433 479 467
rect 419 399 479 433
rect 419 365 432 399
rect 466 365 479 399
rect 419 347 479 365
rect 509 535 576 547
rect 509 501 522 535
rect 556 501 576 535
rect 509 443 576 501
rect 509 409 522 443
rect 556 409 576 443
rect 509 347 576 409
rect 606 542 632 547
rect 666 547 675 576
rect 1555 580 1614 592
rect 1244 547 1363 562
rect 666 542 693 547
rect 606 347 693 542
rect 723 508 794 547
rect 723 474 736 508
rect 770 474 794 508
rect 723 347 794 474
rect 824 511 886 547
rect 824 477 837 511
rect 871 477 886 511
rect 824 347 886 477
rect 916 347 987 547
rect 1017 535 1077 547
rect 1017 501 1030 535
rect 1064 501 1077 535
rect 1017 424 1077 501
rect 1017 390 1030 424
rect 1064 390 1077 424
rect 1017 347 1077 390
rect 1107 535 1196 547
rect 1107 501 1149 535
rect 1183 501 1196 535
rect 1107 451 1196 501
rect 1107 417 1149 451
rect 1183 417 1196 451
rect 1107 347 1196 417
rect 1226 537 1363 547
rect 1226 503 1240 537
rect 1274 503 1315 537
rect 1349 503 1363 537
rect 1226 362 1363 503
rect 1393 550 1460 562
rect 1393 516 1414 550
rect 1448 516 1460 550
rect 1393 440 1460 516
rect 1393 406 1414 440
rect 1448 406 1460 440
rect 1393 362 1460 406
rect 1555 546 1567 580
rect 1601 546 1614 580
rect 1555 497 1614 546
rect 1555 463 1567 497
rect 1601 463 1614 497
rect 1555 414 1614 463
rect 1555 380 1567 414
rect 1601 380 1614 414
rect 1555 368 1614 380
rect 1644 580 1701 592
rect 1644 546 1657 580
rect 1691 546 1701 580
rect 1644 497 1701 546
rect 1644 463 1657 497
rect 1691 463 1701 497
rect 1644 414 1701 463
rect 1644 380 1657 414
rect 1691 380 1701 414
rect 1644 368 1701 380
rect 1226 347 1279 362
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 143 48 177 82
rect 404 93 438 127
rect 520 100 554 134
rect 630 48 664 82
rect 732 100 766 134
rect 846 92 880 126
rect 1025 103 1059 137
rect 1127 51 1161 85
rect 1221 51 1255 85
rect 1366 44 1400 78
rect 1468 112 1502 146
rect 1572 104 1606 138
rect 1658 176 1692 210
rect 1658 86 1692 120
<< pdiffc >>
rect 37 546 71 580
rect 37 463 71 497
rect 37 380 71 414
rect 127 546 161 580
rect 127 478 161 512
rect 127 410 161 444
rect 432 501 466 535
rect 432 433 466 467
rect 432 365 466 399
rect 522 501 556 535
rect 522 409 556 443
rect 632 542 666 576
rect 736 474 770 508
rect 837 477 871 511
rect 1030 501 1064 535
rect 1030 390 1064 424
rect 1149 501 1183 535
rect 1149 417 1183 451
rect 1240 503 1274 537
rect 1315 503 1349 537
rect 1414 516 1448 550
rect 1414 406 1448 440
rect 1567 546 1601 580
rect 1567 463 1601 497
rect 1567 380 1601 414
rect 1657 546 1691 580
rect 1657 463 1691 497
rect 1657 380 1691 414
<< poly >>
rect 84 592 114 618
rect 285 615 1396 645
rect 285 604 321 615
rect 187 568 217 594
rect 288 589 318 604
rect 389 547 419 573
rect 479 547 509 573
rect 573 562 609 615
rect 576 547 606 562
rect 288 374 318 389
rect 84 353 114 368
rect 187 353 217 368
rect 81 326 117 353
rect 69 310 135 326
rect 184 310 220 353
rect 285 343 321 374
rect 693 547 723 573
rect 794 547 824 573
rect 886 547 916 573
rect 984 562 1020 615
rect 1360 577 1396 615
rect 1614 592 1644 618
rect 987 547 1017 562
rect 1077 547 1107 573
rect 1196 547 1226 573
rect 1363 562 1393 577
rect 1363 347 1393 362
rect 1614 353 1644 368
rect 69 276 85 310
rect 119 276 135 310
rect 69 260 135 276
rect 177 294 243 310
rect 177 260 193 294
rect 227 260 243 294
rect 84 222 114 260
rect 177 244 243 260
rect 207 203 237 244
rect 285 203 315 343
rect 389 332 419 347
rect 479 332 509 347
rect 576 332 606 347
rect 693 332 723 347
rect 794 332 824 347
rect 886 332 916 347
rect 987 332 1017 347
rect 1077 332 1107 347
rect 1196 332 1226 347
rect 386 315 422 332
rect 476 315 512 332
rect 357 299 423 315
rect 357 265 373 299
rect 407 265 423 299
rect 357 249 423 265
rect 465 299 531 315
rect 465 265 481 299
rect 515 265 531 299
rect 465 249 531 265
rect 363 203 393 249
rect 471 203 501 249
rect 573 218 609 332
rect 690 291 726 332
rect 791 315 827 332
rect 660 275 726 291
rect 660 241 676 275
rect 710 241 726 275
rect 768 299 834 315
rect 768 265 784 299
rect 818 265 834 299
rect 883 291 919 332
rect 768 249 834 265
rect 876 275 942 291
rect 660 225 726 241
rect 573 203 603 218
rect 691 203 721 225
rect 777 203 807 249
rect 876 241 892 275
rect 926 241 942 275
rect 876 225 942 241
rect 906 203 936 225
rect 984 218 1020 332
rect 1074 315 1110 332
rect 1193 315 1229 332
rect 1360 330 1396 347
rect 1062 299 1128 315
rect 1062 265 1078 299
rect 1112 265 1128 299
rect 1062 249 1128 265
rect 1176 299 1242 315
rect 1176 265 1192 299
rect 1226 265 1242 299
rect 1176 252 1242 265
rect 1360 314 1494 330
rect 1360 280 1376 314
rect 1410 280 1444 314
rect 1478 280 1494 314
rect 1611 310 1647 353
rect 1360 264 1494 280
rect 1542 294 1647 310
rect 984 203 1014 218
rect 1070 203 1100 249
rect 1176 222 1312 252
rect 1282 203 1312 222
rect 1427 203 1457 264
rect 1542 260 1558 294
rect 1592 260 1647 294
rect 1542 244 1647 260
rect 1617 222 1647 244
rect 84 48 114 74
rect 207 49 237 75
rect 285 49 315 75
rect 363 49 393 75
rect 471 49 501 75
rect 573 49 603 75
rect 691 49 721 75
rect 777 49 807 75
rect 906 49 936 75
rect 984 49 1014 75
rect 1070 49 1100 75
rect 1282 49 1312 75
rect 1427 49 1457 75
rect 1617 48 1647 74
<< polycont >>
rect 85 276 119 310
rect 193 260 227 294
rect 373 265 407 299
rect 481 265 515 299
rect 676 241 710 275
rect 784 265 818 299
rect 892 241 926 275
rect 1078 265 1112 299
rect 1192 265 1226 299
rect 1376 280 1410 314
rect 1444 280 1478 314
rect 1558 260 1592 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 17 580 71 596
rect 17 546 37 580
rect 17 497 71 546
rect 17 463 37 497
rect 17 414 71 463
rect 17 380 37 414
rect 111 580 177 649
rect 111 546 127 580
rect 161 546 177 580
rect 616 576 682 649
rect 111 512 177 546
rect 111 478 127 512
rect 161 478 177 512
rect 111 444 177 478
rect 111 410 127 444
rect 161 410 177 444
rect 416 535 482 551
rect 416 501 432 535
rect 466 501 482 535
rect 416 467 482 501
rect 416 433 432 467
rect 466 433 482 467
rect 416 424 482 433
rect 17 364 71 380
rect 211 399 482 424
rect 211 390 432 399
rect 211 376 245 390
rect 17 226 51 364
rect 107 342 245 376
rect 416 365 432 390
rect 466 365 482 399
rect 522 535 572 551
rect 556 501 572 535
rect 616 542 632 576
rect 666 542 682 576
rect 616 526 682 542
rect 522 492 572 501
rect 720 508 786 551
rect 720 492 736 508
rect 522 474 736 492
rect 770 474 786 508
rect 522 458 786 474
rect 821 511 887 649
rect 821 477 837 511
rect 871 477 887 511
rect 821 461 887 477
rect 1014 535 1099 551
rect 1014 501 1030 535
rect 1064 501 1099 535
rect 522 443 572 458
rect 556 409 572 443
rect 1014 424 1099 501
rect 522 393 572 409
rect 313 350 359 356
rect 107 326 141 342
rect 85 310 141 326
rect 119 276 141 310
rect 313 316 319 350
rect 353 316 359 350
rect 416 349 482 365
rect 606 390 1030 424
rect 1064 390 1099 424
rect 1133 535 1190 551
rect 1133 501 1149 535
rect 1183 501 1190 535
rect 1133 451 1190 501
rect 1224 537 1365 649
rect 1551 580 1617 649
rect 1224 503 1240 537
rect 1274 503 1315 537
rect 1349 503 1365 537
rect 1224 500 1365 503
rect 1400 550 1464 566
rect 1400 516 1414 550
rect 1448 516 1464 550
rect 1400 451 1464 516
rect 1133 417 1149 451
rect 1183 440 1464 451
rect 1183 417 1414 440
rect 1398 406 1414 417
rect 1448 406 1464 440
rect 1398 390 1464 406
rect 1551 546 1567 580
rect 1601 546 1617 580
rect 1551 497 1617 546
rect 1551 463 1567 497
rect 1601 463 1617 497
rect 1551 414 1617 463
rect 606 359 640 390
rect 313 315 359 316
rect 516 325 640 359
rect 1065 383 1099 390
rect 768 350 839 356
rect 516 315 550 325
rect 85 260 141 276
rect 17 210 73 226
rect 17 176 39 210
rect 17 120 73 176
rect 17 86 39 120
rect 107 150 141 260
rect 177 294 243 308
rect 177 260 193 294
rect 227 260 243 294
rect 177 244 243 260
rect 313 299 423 315
rect 313 265 373 299
rect 407 265 423 299
rect 313 252 423 265
rect 465 299 550 315
rect 465 265 481 299
rect 515 265 550 299
rect 768 316 799 350
rect 833 316 839 350
rect 768 299 839 316
rect 465 252 550 265
rect 660 275 726 291
rect 209 218 243 244
rect 660 241 676 275
rect 710 241 726 275
rect 768 265 784 299
rect 818 265 839 299
rect 985 350 1031 356
rect 985 316 991 350
rect 1025 316 1031 350
rect 1065 349 1310 383
rect 1551 380 1567 414
rect 1601 380 1617 414
rect 1551 364 1617 380
rect 1657 580 1708 596
rect 1691 546 1708 580
rect 1657 497 1708 546
rect 1691 463 1708 497
rect 1657 414 1708 463
rect 1691 380 1708 414
rect 985 315 1031 316
rect 985 299 1128 315
rect 768 252 839 265
rect 876 275 942 291
rect 660 218 726 241
rect 876 241 892 275
rect 926 241 942 275
rect 985 265 1078 299
rect 1112 265 1128 299
rect 985 255 1128 265
rect 1162 299 1242 315
rect 1162 265 1192 299
rect 1226 265 1242 299
rect 1162 264 1242 265
rect 876 221 942 241
rect 1162 221 1196 264
rect 1276 230 1310 349
rect 1360 314 1494 356
rect 1360 280 1376 314
rect 1410 280 1444 314
rect 1478 280 1494 314
rect 1360 264 1494 280
rect 1542 294 1608 310
rect 1542 260 1558 294
rect 1592 260 1608 294
rect 1542 230 1608 260
rect 876 218 1196 221
rect 209 187 1196 218
rect 1230 196 1608 230
rect 1657 226 1708 380
rect 1642 210 1708 226
rect 209 184 942 187
rect 1230 153 1264 196
rect 1642 176 1658 210
rect 1692 176 1708 210
rect 107 127 454 150
rect 107 116 404 127
rect 17 70 73 86
rect 388 93 404 116
rect 438 93 454 127
rect 125 48 143 82
rect 177 48 196 82
rect 388 71 454 93
rect 496 134 782 150
rect 496 100 520 134
rect 554 116 732 134
rect 554 100 578 116
rect 496 84 578 100
rect 716 100 732 116
rect 766 100 782 134
rect 716 84 782 100
rect 816 126 911 142
rect 816 92 846 126
rect 880 92 911 126
rect 125 17 196 48
rect 614 48 630 82
rect 664 48 680 82
rect 614 17 680 48
rect 816 17 911 92
rect 1009 137 1264 153
rect 1009 103 1025 137
rect 1059 119 1264 137
rect 1298 146 1518 162
rect 1298 128 1468 146
rect 1059 103 1075 119
rect 1009 87 1075 103
rect 1298 85 1332 128
rect 1452 112 1468 128
rect 1502 112 1518 146
rect 1452 96 1518 112
rect 1556 138 1606 154
rect 1556 104 1572 138
rect 1111 51 1127 85
rect 1161 51 1221 85
rect 1255 51 1332 85
rect 1366 78 1416 94
rect 1400 44 1416 78
rect 1366 17 1416 44
rect 1556 17 1606 104
rect 1642 120 1708 176
rect 1642 86 1658 120
rect 1692 86 1708 120
rect 1642 70 1708 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 319 316 353 350
rect 799 316 833 350
rect 991 316 1025 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
<< metal1 >>
rect 0 683 1728 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 0 617 1728 649
rect 307 350 365 356
rect 307 316 319 350
rect 353 347 365 350
rect 787 350 845 356
rect 787 347 799 350
rect 353 319 799 347
rect 353 316 365 319
rect 307 310 365 316
rect 787 316 799 319
rect 833 347 845 350
rect 979 350 1037 356
rect 979 347 991 350
rect 833 319 991 347
rect 833 316 845 319
rect 787 310 845 316
rect 979 316 991 319
rect 1025 316 1037 350
rect 979 310 1037 316
rect 0 17 1728 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
rect 0 -49 1728 -17
<< labels >>
rlabel comment s 0 0 0 0 4 fa_1
flabel pwell s 0 0 1728 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 1728 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 799 316 833 350 0 FreeSans 340 0 0 0 CIN
port 3 nsew
flabel metal1 s 0 617 1728 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 1728 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 895 242 929 276 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 1375 316 1409 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 1663 94 1697 128 0 FreeSans 340 0 0 0 COUT
port 8 nsew
flabel corelocali s 1663 168 1697 202 0 FreeSans 340 0 0 0 COUT
port 8 nsew
flabel corelocali s 1663 242 1697 276 0 FreeSans 340 0 0 0 COUT
port 8 nsew
flabel corelocali s 1663 316 1697 350 0 FreeSans 340 0 0 0 COUT
port 8 nsew
flabel corelocali s 1663 390 1697 424 0 FreeSans 340 0 0 0 COUT
port 8 nsew
flabel corelocali s 1663 464 1697 498 0 FreeSans 340 0 0 0 COUT
port 8 nsew
flabel corelocali s 1663 538 1697 572 0 FreeSans 340 0 0 0 COUT
port 8 nsew
flabel corelocali s 31 94 65 128 0 FreeSans 340 0 0 0 SUM
port 9 nsew
flabel corelocali s 31 168 65 202 0 FreeSans 340 0 0 0 SUM
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 1728 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 2467172
string GDS_START 2453134
<< end >>
