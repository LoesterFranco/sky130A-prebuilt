magic
tech sky130A
magscale 1 2
timestamp 1599588244
<< locali >>
rect 25 225 110 427
rect 161 310 257 419
rect 291 305 353 371
rect 686 236 752 334
rect 1419 581 1621 615
rect 1419 331 1453 581
rect 1587 467 1621 581
rect 1771 581 2053 615
rect 1771 467 1805 581
rect 1587 433 1805 467
rect 1409 282 1475 331
rect 2019 437 2053 581
rect 2019 403 2059 437
rect 2025 372 2059 403
rect 2211 372 2273 430
rect 2025 360 2273 372
rect 2025 338 2277 360
rect 2211 304 2277 338
rect 2774 344 2855 578
rect 2613 236 2672 310
rect 2821 210 2855 344
rect 2754 70 2855 210
rect 3079 70 3147 596
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3168 683
rect 23 495 89 596
rect 123 529 189 649
rect 223 581 455 615
rect 223 495 257 581
rect 23 461 257 495
rect 299 439 349 547
rect 389 504 455 581
rect 501 504 551 649
rect 591 470 657 596
rect 299 405 421 439
rect 387 271 421 405
rect 455 436 657 470
rect 455 366 556 436
rect 703 402 769 596
rect 809 436 843 649
rect 208 237 484 271
rect 28 17 94 191
rect 208 115 274 237
rect 366 17 416 203
rect 450 85 484 237
rect 522 207 556 366
rect 618 368 849 402
rect 883 368 981 596
rect 1015 407 1081 551
rect 1115 441 1225 507
rect 1015 373 1157 407
rect 522 119 572 207
rect 618 202 652 368
rect 815 334 849 368
rect 947 339 981 368
rect 815 268 913 334
rect 947 273 1089 339
rect 947 234 981 273
rect 1123 239 1157 373
rect 618 119 668 202
rect 872 200 981 234
rect 1033 205 1157 239
rect 1191 365 1225 441
rect 1319 415 1385 649
rect 1191 331 1375 365
rect 1487 399 1553 547
rect 1663 501 1737 649
rect 1875 422 1985 547
rect 1487 365 1803 399
rect 1033 166 1067 205
rect 1191 171 1225 331
rect 702 132 1067 166
rect 702 85 736 132
rect 450 51 736 85
rect 770 17 836 98
rect 1001 92 1067 132
rect 1101 137 1225 171
rect 1259 180 1307 297
rect 1341 248 1375 331
rect 1517 248 1583 317
rect 1341 214 1583 248
rect 1625 276 1703 317
rect 1625 242 1663 276
rect 1697 242 1703 276
rect 1625 236 1703 242
rect 1737 267 1803 365
rect 1851 301 1917 388
rect 1951 369 1985 422
rect 2087 532 2230 649
rect 2307 498 2357 596
rect 2093 464 2357 498
rect 2459 496 2525 649
rect 2668 496 2734 649
rect 2093 406 2159 464
rect 2307 462 2357 464
rect 2307 428 2740 462
rect 2307 394 2443 428
rect 1951 335 1991 369
rect 1957 304 1991 335
rect 1851 267 1923 301
rect 1737 180 1771 267
rect 1259 146 1771 180
rect 1101 92 1167 137
rect 1564 131 1630 146
rect 1298 17 1377 112
rect 1429 96 1528 112
rect 1666 96 1743 112
rect 1429 62 1743 96
rect 1805 17 1855 210
rect 1889 85 1923 267
rect 1957 270 2177 304
rect 2319 270 2375 310
rect 1957 119 1997 270
rect 2143 236 2375 270
rect 2031 85 2097 236
rect 2409 202 2443 394
rect 2545 344 2631 394
rect 2489 276 2579 344
rect 2706 310 2740 428
rect 2489 242 2527 276
rect 2561 242 2579 276
rect 2489 236 2579 242
rect 2706 244 2783 310
rect 2545 202 2579 236
rect 1889 51 2097 85
rect 2180 17 2230 202
rect 2266 85 2332 202
rect 2374 119 2443 202
rect 2477 85 2511 202
rect 2545 134 2623 202
rect 2266 51 2511 85
rect 2659 17 2718 200
rect 2889 337 2955 596
rect 2989 423 3041 649
rect 2889 271 2969 337
rect 2889 70 2943 271
rect 2979 17 3045 188
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3168 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 1663 242 1697 276
rect 2527 242 2561 276
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
<< metal1 >>
rect 0 683 3168 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3168 683
rect 0 617 3168 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 3168 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3168 17
rect 0 -49 3168 -17
<< obsm1 >>
rect 1651 276 1709 282
rect 1651 242 1663 276
rect 1697 273 1709 276
rect 2515 276 2573 282
rect 2515 273 2527 276
rect 1697 245 2527 273
rect 1697 242 1709 245
rect 1651 236 1709 242
rect 2515 242 2527 245
rect 2561 242 2573 276
rect 2515 236 2573 242
<< labels >>
rlabel locali s 291 305 353 371 6 D
port 1 nsew signal input
rlabel locali s 3079 70 3147 596 6 Q
port 2 nsew signal output
rlabel locali s 2821 210 2855 344 6 Q_N
port 3 nsew signal output
rlabel locali s 2774 344 2855 578 6 Q_N
port 3 nsew signal output
rlabel locali s 2754 70 2855 210 6 Q_N
port 3 nsew signal output
rlabel locali s 2613 236 2672 310 6 RESET_B
port 4 nsew signal input
rlabel locali s 25 225 110 427 6 SCD
port 5 nsew signal input
rlabel locali s 161 310 257 419 6 SCE
port 6 nsew signal input
rlabel locali s 2211 372 2273 430 6 SET_B
port 7 nsew signal input
rlabel locali s 2211 304 2277 338 6 SET_B
port 7 nsew signal input
rlabel locali s 2025 372 2059 403 6 SET_B
port 7 nsew signal input
rlabel locali s 2025 360 2273 372 6 SET_B
port 7 nsew signal input
rlabel locali s 2025 338 2277 360 6 SET_B
port 7 nsew signal input
rlabel locali s 2019 437 2053 581 6 SET_B
port 7 nsew signal input
rlabel locali s 2019 403 2059 437 6 SET_B
port 7 nsew signal input
rlabel locali s 1771 581 2053 615 6 SET_B
port 7 nsew signal input
rlabel locali s 1771 467 1805 581 6 SET_B
port 7 nsew signal input
rlabel locali s 1587 467 1621 581 6 SET_B
port 7 nsew signal input
rlabel locali s 1587 433 1805 467 6 SET_B
port 7 nsew signal input
rlabel locali s 1419 581 1621 615 6 SET_B
port 7 nsew signal input
rlabel locali s 1419 331 1453 581 6 SET_B
port 7 nsew signal input
rlabel locali s 1409 282 1475 331 6 SET_B
port 7 nsew signal input
rlabel locali s 686 236 752 334 6 CLK
port 8 nsew clock input
rlabel metal1 s 0 -49 3168 49 8 VGND
port 9 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 10 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 11 nsew power bidirectional
rlabel metal1 s 0 617 3168 715 6 VPWR
port 12 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 3168 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 989222
string GDS_START 966454
<< end >>
