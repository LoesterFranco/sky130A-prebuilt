magic
tech sky130A
magscale 1 2
timestamp 1604502697
<< nwell >>
rect -38 261 1050 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 83 47 113 177
rect 187 47 217 177
rect 271 47 301 177
rect 375 47 405 177
rect 571 47 601 177
rect 675 47 705 177
rect 759 47 789 177
rect 863 47 893 177
<< pmoshvt >>
rect 85 297 121 497
rect 179 297 215 497
rect 273 297 309 497
rect 367 297 403 497
rect 573 297 609 497
rect 667 297 703 497
rect 761 297 797 497
rect 855 297 891 497
<< ndiff >>
rect 27 163 83 177
rect 27 129 39 163
rect 73 129 83 163
rect 27 95 83 129
rect 27 61 39 95
rect 73 61 83 95
rect 27 47 83 61
rect 113 163 187 177
rect 113 129 133 163
rect 167 129 187 163
rect 113 47 187 129
rect 217 95 271 177
rect 217 61 227 95
rect 261 61 271 95
rect 217 47 271 61
rect 301 163 375 177
rect 301 129 321 163
rect 355 129 375 163
rect 301 47 375 129
rect 405 95 571 177
rect 405 61 415 95
rect 449 61 526 95
rect 560 61 571 95
rect 405 47 571 61
rect 601 95 675 177
rect 601 61 631 95
rect 665 61 675 95
rect 601 47 675 61
rect 705 163 759 177
rect 705 129 715 163
rect 749 129 759 163
rect 705 95 759 129
rect 705 61 715 95
rect 749 61 759 95
rect 705 47 759 61
rect 789 95 863 177
rect 789 61 809 95
rect 843 61 863 95
rect 789 47 863 61
rect 893 163 945 177
rect 893 129 903 163
rect 937 129 945 163
rect 893 95 945 129
rect 893 61 903 95
rect 937 61 945 95
rect 893 47 945 61
<< pdiff >>
rect 27 477 85 497
rect 27 443 39 477
rect 73 443 85 477
rect 27 409 85 443
rect 27 375 39 409
rect 73 375 85 409
rect 27 341 85 375
rect 27 307 39 341
rect 73 307 85 341
rect 27 297 85 307
rect 121 477 179 497
rect 121 443 133 477
rect 167 443 179 477
rect 121 409 179 443
rect 121 375 133 409
rect 167 375 179 409
rect 121 297 179 375
rect 215 477 273 497
rect 215 443 227 477
rect 261 443 273 477
rect 215 409 273 443
rect 215 375 227 409
rect 261 375 273 409
rect 215 341 273 375
rect 215 307 227 341
rect 261 307 273 341
rect 215 297 273 307
rect 309 409 367 497
rect 309 375 321 409
rect 355 375 367 409
rect 309 341 367 375
rect 309 307 321 341
rect 355 307 367 341
rect 309 297 367 307
rect 403 477 461 497
rect 403 443 415 477
rect 449 443 461 477
rect 403 409 461 443
rect 403 375 415 409
rect 449 375 461 409
rect 403 297 461 375
rect 515 477 573 497
rect 515 443 527 477
rect 561 443 573 477
rect 515 409 573 443
rect 515 375 527 409
rect 561 375 573 409
rect 515 297 573 375
rect 609 409 667 497
rect 609 375 621 409
rect 655 375 667 409
rect 609 341 667 375
rect 609 307 621 341
rect 655 307 667 341
rect 609 297 667 307
rect 703 477 761 497
rect 703 443 715 477
rect 749 443 761 477
rect 703 409 761 443
rect 703 375 715 409
rect 749 375 761 409
rect 703 341 761 375
rect 703 307 715 341
rect 749 307 761 341
rect 703 297 761 307
rect 797 477 855 497
rect 797 443 809 477
rect 843 443 855 477
rect 797 409 855 443
rect 797 375 809 409
rect 843 375 855 409
rect 797 297 855 375
rect 891 477 949 497
rect 891 443 903 477
rect 937 443 949 477
rect 891 409 949 443
rect 891 375 903 409
rect 937 375 949 409
rect 891 341 949 375
rect 891 307 903 341
rect 937 307 949 341
rect 891 297 949 307
<< ndiffc >>
rect 39 129 73 163
rect 39 61 73 95
rect 133 129 167 163
rect 227 61 261 95
rect 321 129 355 163
rect 415 61 449 95
rect 526 61 560 95
rect 631 61 665 95
rect 715 129 749 163
rect 715 61 749 95
rect 809 61 843 95
rect 903 129 937 163
rect 903 61 937 95
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 133 443 167 477
rect 133 375 167 409
rect 227 443 261 477
rect 227 375 261 409
rect 227 307 261 341
rect 321 375 355 409
rect 321 307 355 341
rect 415 443 449 477
rect 415 375 449 409
rect 527 443 561 477
rect 527 375 561 409
rect 621 375 655 409
rect 621 307 655 341
rect 715 443 749 477
rect 715 375 749 409
rect 715 307 749 341
rect 809 443 843 477
rect 809 375 843 409
rect 903 443 937 477
rect 903 375 937 409
rect 903 307 937 341
<< poly >>
rect 85 497 121 523
rect 179 497 215 523
rect 273 497 309 523
rect 367 497 403 523
rect 573 497 609 523
rect 667 497 703 523
rect 761 497 797 523
rect 855 497 891 523
rect 85 282 121 297
rect 179 282 215 297
rect 273 282 309 297
rect 367 282 403 297
rect 573 282 609 297
rect 667 282 703 297
rect 761 282 797 297
rect 855 282 891 297
rect 83 265 123 282
rect 177 265 217 282
rect 83 249 217 265
rect 83 215 95 249
rect 129 215 173 249
rect 207 215 217 249
rect 83 199 217 215
rect 83 177 113 199
rect 187 177 217 199
rect 271 265 311 282
rect 365 265 405 282
rect 271 249 405 265
rect 271 215 281 249
rect 315 215 359 249
rect 393 215 405 249
rect 271 199 405 215
rect 271 177 301 199
rect 375 177 405 199
rect 571 265 611 282
rect 665 265 705 282
rect 571 249 705 265
rect 571 215 583 249
rect 617 215 661 249
rect 695 215 705 249
rect 571 199 705 215
rect 571 177 601 199
rect 675 177 705 199
rect 759 265 799 282
rect 853 265 893 282
rect 759 249 893 265
rect 759 215 769 249
rect 803 215 847 249
rect 881 215 893 249
rect 759 199 893 215
rect 759 177 789 199
rect 863 177 893 199
rect 83 21 113 47
rect 187 21 217 47
rect 271 21 301 47
rect 375 21 405 47
rect 571 21 601 47
rect 675 21 705 47
rect 759 21 789 47
rect 863 21 893 47
<< polycont >>
rect 95 215 129 249
rect 173 215 207 249
rect 281 215 315 249
rect 359 215 393 249
rect 583 215 617 249
rect 661 215 695 249
rect 769 215 803 249
rect 847 215 881 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 30 477 81 493
rect 30 443 39 477
rect 73 443 81 477
rect 30 409 81 443
rect 30 375 39 409
rect 73 375 81 409
rect 30 341 81 375
rect 125 477 175 527
rect 125 443 133 477
rect 167 443 175 477
rect 125 409 175 443
rect 125 375 133 409
rect 167 375 175 409
rect 125 359 175 375
rect 219 477 457 493
rect 219 443 227 477
rect 261 459 415 477
rect 261 443 269 459
rect 219 409 269 443
rect 407 443 415 459
rect 449 443 457 477
rect 219 375 227 409
rect 261 375 269 409
rect 30 307 39 341
rect 73 325 81 341
rect 219 341 269 375
rect 219 325 227 341
rect 73 307 227 325
rect 261 307 269 341
rect 30 291 269 307
rect 313 409 363 425
rect 313 375 321 409
rect 355 375 363 409
rect 313 341 363 375
rect 407 409 457 443
rect 407 375 415 409
rect 449 375 457 409
rect 407 359 457 375
rect 519 477 757 493
rect 519 443 527 477
rect 561 459 715 477
rect 561 443 569 459
rect 519 409 569 443
rect 707 443 715 459
rect 749 443 757 477
rect 519 375 527 409
rect 561 375 569 409
rect 519 359 569 375
rect 613 409 663 425
rect 613 375 621 409
rect 655 375 663 409
rect 313 307 321 341
rect 355 325 363 341
rect 613 341 663 375
rect 613 325 621 341
rect 355 307 621 325
rect 655 307 663 341
rect 313 289 663 307
rect 707 409 757 443
rect 707 375 715 409
rect 749 375 757 409
rect 707 341 757 375
rect 801 477 851 527
rect 801 443 809 477
rect 843 443 851 477
rect 801 409 851 443
rect 801 375 809 409
rect 843 375 851 409
rect 801 359 851 375
rect 895 477 946 493
rect 895 443 903 477
rect 937 443 946 477
rect 895 409 946 443
rect 895 375 903 409
rect 937 375 946 409
rect 707 307 715 341
rect 749 325 757 341
rect 895 341 946 375
rect 895 325 903 341
rect 749 307 903 325
rect 937 307 946 341
rect 707 291 946 307
rect 40 249 223 257
rect 40 215 95 249
rect 129 215 173 249
rect 207 215 223 249
rect 265 249 425 255
rect 265 215 281 249
rect 315 215 359 249
rect 393 215 425 249
rect 481 181 529 289
rect 567 249 711 255
rect 567 215 583 249
rect 617 215 661 249
rect 695 215 711 249
rect 753 249 913 257
rect 753 215 769 249
rect 803 215 847 249
rect 881 215 913 249
rect 18 163 73 181
rect 18 129 39 163
rect 107 163 529 181
rect 107 129 133 163
rect 167 129 321 163
rect 355 129 529 163
rect 563 163 953 181
rect 563 145 715 163
rect 18 95 73 129
rect 563 95 597 145
rect 699 129 715 145
rect 749 145 903 163
rect 749 129 765 145
rect 18 61 39 95
rect 73 61 227 95
rect 261 61 415 95
rect 449 61 526 95
rect 560 61 597 95
rect 631 95 665 111
rect 631 17 665 61
rect 699 95 765 129
rect 877 129 903 145
rect 937 129 953 163
rect 699 61 715 95
rect 749 61 765 95
rect 699 51 765 61
rect 809 95 843 111
rect 809 17 843 61
rect 877 95 953 129
rect 877 61 903 95
rect 937 61 953 95
rect 877 51 953 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
flabel corelocali s 323 238 323 238 0 FreeSans 400 0 0 0 B2
port 4 nsew
flabel corelocali s 132 221 166 255 0 FreeSans 400 0 0 0 B1
port 3 nsew
flabel corelocali s 438 289 472 323 0 FreeSans 400 0 0 0 Y
port 9 nsew
flabel corelocali s 787 238 787 238 0 FreeSans 400 0 0 0 A1
port 1 nsew
flabel corelocali s 603 238 603 238 0 FreeSans 400 0 0 0 A2
port 2 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
rlabel comment s 0 0 0 0 4 o22ai_2
<< properties >>
string FIXED_BBOX 0 0 1012 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 863284
string GDS_START 855168
<< end >>
