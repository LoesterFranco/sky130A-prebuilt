magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 2822 704
rect 1491 305 1703 332
<< pwell >>
rect 0 0 2784 49
<< scnmos >>
rect 100 74 130 158
rect 208 74 238 158
rect 286 74 316 158
rect 372 74 402 158
rect 450 74 480 158
rect 656 74 686 222
rect 770 74 800 222
rect 968 81 998 165
rect 1120 81 1150 165
rect 1198 81 1228 165
rect 1396 118 1426 202
rect 1474 118 1504 202
rect 1656 74 1686 202
rect 1734 74 1764 202
rect 1880 74 1910 158
rect 1958 74 1988 158
rect 2140 74 2170 158
rect 2254 74 2284 158
rect 2535 112 2565 222
rect 2651 74 2681 222
<< pmoshvt >>
rect 85 464 115 592
rect 175 464 205 592
rect 259 464 289 592
rect 385 464 415 592
rect 469 464 499 592
rect 688 368 718 592
rect 778 368 808 592
rect 998 457 1028 541
rect 1098 457 1128 541
rect 1201 457 1231 541
rect 1348 457 1378 541
rect 1444 457 1474 541
rect 1580 341 1610 541
rect 1774 374 1804 458
rect 1886 374 1916 574
rect 2083 508 2113 592
rect 2173 508 2203 592
rect 2371 508 2401 592
rect 2569 403 2599 571
rect 2670 368 2700 592
<< ndiff >>
rect 599 188 656 222
rect 43 133 100 158
rect 43 99 55 133
rect 89 99 100 133
rect 43 74 100 99
rect 130 129 208 158
rect 130 95 155 129
rect 189 95 208 129
rect 130 74 208 95
rect 238 74 286 158
rect 316 133 372 158
rect 316 99 327 133
rect 361 99 372 133
rect 316 74 372 99
rect 402 74 450 158
rect 480 127 537 158
rect 480 93 491 127
rect 525 93 537 127
rect 480 74 537 93
rect 599 154 611 188
rect 645 154 656 188
rect 599 120 656 154
rect 599 86 611 120
rect 645 86 656 120
rect 599 74 656 86
rect 686 188 770 222
rect 686 154 711 188
rect 745 154 770 188
rect 686 120 770 154
rect 686 86 711 120
rect 745 86 770 120
rect 686 74 770 86
rect 800 210 857 222
rect 800 176 811 210
rect 845 176 857 210
rect 800 120 857 176
rect 1339 177 1396 202
rect 800 86 811 120
rect 845 86 857 120
rect 800 74 857 86
rect 911 153 968 165
rect 911 119 923 153
rect 957 119 968 153
rect 911 81 968 119
rect 998 140 1120 165
rect 998 106 1075 140
rect 1109 106 1120 140
rect 998 81 1120 106
rect 1150 81 1198 165
rect 1228 132 1285 165
rect 1228 98 1239 132
rect 1273 98 1285 132
rect 1339 143 1351 177
rect 1385 143 1396 177
rect 1339 118 1396 143
rect 1426 118 1474 202
rect 1504 188 1656 202
rect 1504 154 1515 188
rect 1549 154 1611 188
rect 1645 154 1656 188
rect 1504 120 1656 154
rect 1504 118 1531 120
rect 1228 81 1285 98
rect 1519 86 1531 118
rect 1565 86 1611 120
rect 1645 86 1656 120
rect 1519 74 1656 86
rect 1686 74 1734 202
rect 1764 188 1865 202
rect 1764 154 1797 188
rect 1831 158 1865 188
rect 2395 185 2535 222
rect 2395 158 2490 185
rect 1831 154 1880 158
rect 1764 120 1880 154
rect 1764 86 1797 120
rect 1831 86 1880 120
rect 1764 74 1880 86
rect 1910 74 1958 158
rect 1988 74 2140 158
rect 2170 133 2254 158
rect 2170 99 2181 133
rect 2215 99 2254 133
rect 2170 74 2254 99
rect 2284 133 2341 158
rect 2284 99 2295 133
rect 2329 99 2341 133
rect 2395 124 2407 158
rect 2441 151 2490 158
rect 2524 151 2535 185
rect 2441 124 2535 151
rect 2395 112 2535 124
rect 2565 194 2651 222
rect 2565 160 2592 194
rect 2626 160 2651 194
rect 2565 120 2651 160
rect 2565 112 2592 120
rect 2284 74 2341 99
rect 2580 86 2592 112
rect 2626 86 2651 120
rect 2580 74 2651 86
rect 2681 194 2738 222
rect 2681 160 2692 194
rect 2726 160 2738 194
rect 2681 120 2738 160
rect 2681 86 2692 120
rect 2726 86 2738 120
rect 2681 74 2738 86
<< pdiff >>
rect 517 616 575 628
rect 517 592 529 616
rect 27 580 85 592
rect 27 546 38 580
rect 72 546 85 580
rect 27 510 85 546
rect 27 476 38 510
rect 72 476 85 510
rect 27 464 85 476
rect 115 573 175 592
rect 115 539 128 573
rect 162 539 175 573
rect 115 464 175 539
rect 205 464 259 592
rect 289 566 385 592
rect 289 532 320 566
rect 354 532 385 566
rect 289 464 385 532
rect 415 464 469 592
rect 499 582 529 592
rect 563 582 575 616
rect 499 464 575 582
rect 629 414 688 592
rect 629 380 641 414
rect 675 380 688 414
rect 629 368 688 380
rect 718 573 778 592
rect 718 539 731 573
rect 765 539 778 573
rect 718 368 778 539
rect 808 573 867 592
rect 808 539 821 573
rect 855 539 867 573
rect 808 520 867 539
rect 808 368 861 520
rect 1249 587 1307 599
rect 1249 553 1261 587
rect 1295 553 1307 587
rect 1721 588 1779 600
rect 1249 541 1307 553
rect 1721 554 1733 588
rect 1767 554 1779 588
rect 1721 542 1779 554
rect 939 516 998 541
rect 939 482 951 516
rect 985 482 998 516
rect 939 457 998 482
rect 1028 516 1098 541
rect 1028 482 1051 516
rect 1085 482 1098 516
rect 1028 457 1098 482
rect 1128 457 1201 541
rect 1231 457 1348 541
rect 1378 516 1444 541
rect 1378 482 1397 516
rect 1431 482 1444 516
rect 1378 457 1444 482
rect 1474 520 1580 541
rect 1474 486 1533 520
rect 1567 486 1580 520
rect 1474 457 1580 486
rect 1527 341 1580 457
rect 1610 529 1667 541
rect 1610 495 1623 529
rect 1657 495 1667 529
rect 1610 434 1667 495
rect 1610 400 1623 434
rect 1657 400 1667 434
rect 1610 341 1667 400
rect 1721 458 1751 542
rect 1833 458 1886 574
rect 1721 374 1774 458
rect 1804 420 1886 458
rect 1804 386 1838 420
rect 1872 386 1886 420
rect 1804 374 1886 386
rect 1916 531 1972 574
rect 1916 497 1929 531
rect 1963 497 1972 531
rect 2026 571 2083 592
rect 2026 537 2036 571
rect 2070 537 2083 571
rect 2026 508 2083 537
rect 2113 571 2173 592
rect 2113 537 2126 571
rect 2160 537 2173 571
rect 2113 508 2173 537
rect 2203 567 2260 592
rect 2203 533 2216 567
rect 2250 533 2260 567
rect 2203 508 2260 533
rect 2314 567 2371 592
rect 2314 533 2324 567
rect 2358 533 2371 567
rect 2314 508 2371 533
rect 2401 571 2458 592
rect 2617 571 2670 592
rect 2401 537 2414 571
rect 2448 537 2458 571
rect 2401 508 2458 537
rect 2512 559 2569 571
rect 2512 525 2522 559
rect 2556 525 2569 559
rect 1916 442 1972 497
rect 1916 408 1929 442
rect 1963 408 1972 442
rect 1916 374 1972 408
rect 2512 449 2569 525
rect 2512 415 2522 449
rect 2556 415 2569 449
rect 2512 403 2569 415
rect 2599 559 2670 571
rect 2599 525 2622 559
rect 2656 525 2670 559
rect 2599 449 2670 525
rect 2599 415 2622 449
rect 2656 415 2670 449
rect 2599 403 2670 415
rect 2617 368 2670 403
rect 2700 580 2757 592
rect 2700 546 2713 580
rect 2747 546 2757 580
rect 2700 497 2757 546
rect 2700 463 2713 497
rect 2747 463 2757 497
rect 2700 414 2757 463
rect 2700 380 2713 414
rect 2747 380 2757 414
rect 2700 368 2757 380
<< ndiffc >>
rect 55 99 89 133
rect 155 95 189 129
rect 327 99 361 133
rect 491 93 525 127
rect 611 154 645 188
rect 611 86 645 120
rect 711 154 745 188
rect 711 86 745 120
rect 811 176 845 210
rect 811 86 845 120
rect 923 119 957 153
rect 1075 106 1109 140
rect 1239 98 1273 132
rect 1351 143 1385 177
rect 1515 154 1549 188
rect 1611 154 1645 188
rect 1531 86 1565 120
rect 1611 86 1645 120
rect 1797 154 1831 188
rect 1797 86 1831 120
rect 2181 99 2215 133
rect 2295 99 2329 133
rect 2407 124 2441 158
rect 2490 151 2524 185
rect 2592 160 2626 194
rect 2592 86 2626 120
rect 2692 160 2726 194
rect 2692 86 2726 120
<< pdiffc >>
rect 38 546 72 580
rect 38 476 72 510
rect 128 539 162 573
rect 320 532 354 566
rect 529 582 563 616
rect 641 380 675 414
rect 731 539 765 573
rect 821 539 855 573
rect 1261 553 1295 587
rect 1733 554 1767 588
rect 951 482 985 516
rect 1051 482 1085 516
rect 1397 482 1431 516
rect 1533 486 1567 520
rect 1623 495 1657 529
rect 1623 400 1657 434
rect 1838 386 1872 420
rect 1929 497 1963 531
rect 2036 537 2070 571
rect 2126 537 2160 571
rect 2216 533 2250 567
rect 2324 533 2358 567
rect 2414 537 2448 571
rect 2522 525 2556 559
rect 1929 408 1963 442
rect 2522 415 2556 449
rect 2622 525 2656 559
rect 2622 415 2656 449
rect 2713 546 2747 580
rect 2713 463 2747 497
rect 2713 380 2747 414
<< poly >>
rect 85 592 115 618
rect 175 592 205 618
rect 259 592 289 618
rect 385 592 415 618
rect 469 592 499 618
rect 688 592 718 618
rect 778 592 808 618
rect 894 615 1919 645
rect 85 449 115 464
rect 175 449 205 464
rect 259 449 289 464
rect 385 449 415 464
rect 469 449 499 464
rect 82 390 118 449
rect 172 390 208 449
rect 256 430 292 449
rect 382 432 418 449
rect 70 374 208 390
rect 70 340 86 374
rect 120 360 208 374
rect 250 414 316 430
rect 250 380 266 414
rect 300 380 316 414
rect 250 364 316 380
rect 358 416 424 432
rect 358 382 374 416
rect 408 382 424 416
rect 466 430 502 449
rect 466 414 569 430
rect 466 400 519 414
rect 358 366 424 382
rect 472 380 519 400
rect 553 380 569 414
rect 120 340 136 360
rect 70 306 136 340
rect 70 272 86 306
rect 120 272 136 306
rect 70 256 136 272
rect 100 158 130 256
rect 178 238 244 254
rect 178 204 194 238
rect 228 204 244 238
rect 178 188 244 204
rect 208 158 238 188
rect 286 158 316 364
rect 472 346 569 380
rect 894 492 924 615
rect 998 541 1028 567
rect 1095 556 1131 615
rect 1098 541 1128 556
rect 1201 541 1231 567
rect 1883 589 1919 615
rect 2083 592 2113 618
rect 2173 592 2203 618
rect 2371 592 2401 618
rect 1348 541 1378 567
rect 1444 541 1474 567
rect 1580 541 1610 567
rect 1886 574 1916 589
rect 876 462 924 492
rect 688 353 718 368
rect 778 353 808 368
rect 358 302 424 318
rect 358 268 374 302
rect 408 268 424 302
rect 358 252 424 268
rect 472 312 519 346
rect 553 312 569 346
rect 472 278 569 312
rect 685 310 721 353
rect 372 158 402 252
rect 472 244 519 278
rect 553 244 569 278
rect 655 294 721 310
rect 775 336 811 353
rect 876 336 906 462
rect 998 442 1028 457
rect 995 414 1031 442
rect 1098 431 1128 457
rect 1201 442 1231 457
rect 1348 442 1378 457
rect 1444 442 1474 457
rect 775 320 906 336
rect 775 300 793 320
rect 655 260 671 294
rect 705 260 721 294
rect 655 244 721 260
rect 770 286 793 300
rect 827 286 906 320
rect 770 270 906 286
rect 948 398 1031 414
rect 948 364 964 398
rect 998 364 1031 398
rect 1198 425 1234 442
rect 1198 409 1269 425
rect 948 353 1031 364
rect 1090 373 1156 389
rect 1090 353 1106 373
rect 948 339 1106 353
rect 1140 339 1156 373
rect 1198 375 1219 409
rect 1253 375 1269 409
rect 1198 359 1269 375
rect 1345 367 1381 442
rect 1441 367 1477 442
rect 948 330 1156 339
rect 948 296 964 330
rect 998 323 1156 330
rect 998 296 1031 323
rect 948 280 1031 296
rect 472 228 569 244
rect 472 204 502 228
rect 656 222 686 244
rect 770 222 800 270
rect 876 238 906 270
rect 450 174 502 204
rect 450 158 480 174
rect 876 208 998 238
rect 968 165 998 208
rect 1120 165 1150 323
rect 1239 253 1269 359
rect 1321 351 1387 367
rect 1321 317 1337 351
rect 1371 317 1387 351
rect 1321 301 1387 317
rect 1429 351 1504 367
rect 1429 317 1445 351
rect 1479 317 1504 351
rect 1774 458 1804 484
rect 2569 571 2599 597
rect 2670 592 2700 618
rect 2083 493 2113 508
rect 2173 493 2203 508
rect 2371 493 2401 508
rect 2080 488 2116 493
rect 2062 458 2116 488
rect 1774 359 1804 374
rect 1886 359 1916 374
rect 1580 326 1610 341
rect 1239 237 1305 253
rect 1239 217 1255 237
rect 1198 203 1255 217
rect 1289 203 1305 237
rect 1351 248 1381 301
rect 1429 296 1504 317
rect 1351 218 1426 248
rect 1198 187 1305 203
rect 1396 202 1426 218
rect 1474 202 1504 296
rect 1577 290 1613 326
rect 1771 290 1807 359
rect 1552 274 1686 290
rect 1552 240 1568 274
rect 1602 240 1636 274
rect 1670 240 1686 274
rect 1552 224 1686 240
rect 1656 202 1686 224
rect 1734 274 1807 290
rect 1734 240 1750 274
rect 1784 240 1807 274
rect 1734 224 1807 240
rect 1880 282 1919 359
rect 1734 202 1764 224
rect 1198 165 1228 187
rect 1396 92 1426 118
rect 1474 92 1504 118
rect 100 48 130 74
rect 208 48 238 74
rect 286 48 316 74
rect 372 48 402 74
rect 450 48 480 74
rect 656 48 686 74
rect 770 48 800 74
rect 968 55 998 81
rect 1120 55 1150 81
rect 1198 55 1228 81
rect 1880 158 1910 282
rect 2062 262 2092 458
rect 2170 410 2206 493
rect 2368 458 2404 493
rect 2374 410 2404 458
rect 1958 246 2092 262
rect 1958 212 1974 246
rect 2008 212 2042 246
rect 2076 212 2092 246
rect 1958 173 2092 212
rect 2140 394 2206 410
rect 2140 360 2156 394
rect 2190 360 2206 394
rect 2140 326 2206 360
rect 2140 292 2156 326
rect 2190 292 2206 326
rect 2140 276 2206 292
rect 2254 394 2404 410
rect 2254 360 2270 394
rect 2304 388 2404 394
rect 2569 388 2599 403
rect 2304 360 2602 388
rect 2254 358 2602 360
rect 2254 326 2320 358
rect 2254 292 2270 326
rect 2304 292 2320 326
rect 2254 276 2320 292
rect 1958 158 1988 173
rect 2140 158 2170 276
rect 2254 158 2284 276
rect 2535 222 2565 358
rect 2670 353 2700 368
rect 2667 310 2703 353
rect 2613 294 2703 310
rect 2613 260 2629 294
rect 2663 260 2703 294
rect 2613 244 2703 260
rect 2651 222 2681 244
rect 2535 86 2565 112
rect 1656 48 1686 74
rect 1734 48 1764 74
rect 1880 48 1910 74
rect 1958 48 1988 74
rect 2140 48 2170 74
rect 2254 48 2284 74
rect 2651 48 2681 74
<< polycont >>
rect 86 340 120 374
rect 266 380 300 414
rect 374 382 408 416
rect 519 380 553 414
rect 86 272 120 306
rect 194 204 228 238
rect 374 268 408 302
rect 519 312 553 346
rect 519 244 553 278
rect 671 260 705 294
rect 793 286 827 320
rect 964 364 998 398
rect 1106 339 1140 373
rect 1219 375 1253 409
rect 964 296 998 330
rect 1337 317 1371 351
rect 1445 317 1479 351
rect 1255 203 1289 237
rect 1568 240 1602 274
rect 1636 240 1670 274
rect 1750 240 1784 274
rect 1974 212 2008 246
rect 2042 212 2076 246
rect 2156 360 2190 394
rect 2156 292 2190 326
rect 2270 360 2304 394
rect 2270 292 2304 326
rect 2629 260 2663 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 17 580 72 596
rect 17 546 38 580
rect 17 510 72 546
rect 112 573 178 649
rect 513 616 579 649
rect 513 582 529 616
rect 563 582 579 616
rect 112 539 128 573
rect 162 539 178 573
rect 112 532 178 539
rect 286 566 477 582
rect 513 566 579 582
rect 715 573 781 649
rect 286 532 320 566
rect 354 532 477 566
rect 715 539 731 573
rect 765 539 781 573
rect 17 476 38 510
rect 443 498 681 532
rect 715 516 781 539
rect 821 579 1169 613
rect 821 573 855 579
rect 821 516 855 539
rect 889 516 1001 545
rect 72 476 409 498
rect 17 464 409 476
rect 17 460 72 464
rect 17 222 51 460
rect 217 414 316 430
rect 85 374 167 390
rect 85 340 86 374
rect 120 340 167 374
rect 217 380 266 414
rect 300 380 316 414
rect 217 364 316 380
rect 358 416 409 464
rect 358 382 374 416
rect 408 382 409 416
rect 358 366 409 382
rect 85 322 167 340
rect 85 306 409 322
rect 85 272 86 306
rect 120 302 409 306
rect 120 288 374 302
rect 120 272 136 288
rect 85 256 136 272
rect 358 268 374 288
rect 408 268 409 302
rect 178 238 244 254
rect 358 252 409 268
rect 178 222 194 238
rect 17 204 194 222
rect 228 204 244 238
rect 443 218 477 498
rect 647 482 681 498
rect 889 482 951 516
rect 985 482 1001 516
rect 647 448 1001 482
rect 1035 516 1101 545
rect 1035 482 1051 516
rect 1085 482 1101 516
rect 1035 453 1101 482
rect 1135 503 1169 579
rect 1245 587 1295 649
rect 1245 553 1261 587
rect 1245 537 1295 553
rect 1329 579 1499 613
rect 1329 503 1363 579
rect 1135 469 1363 503
rect 1397 516 1431 545
rect 511 414 561 430
rect 511 380 519 414
rect 553 380 561 414
rect 511 346 561 380
rect 511 312 519 346
rect 553 312 561 346
rect 511 278 561 312
rect 511 244 519 278
rect 553 244 561 278
rect 511 228 561 244
rect 595 380 641 414
rect 675 380 843 414
rect 595 364 843 380
rect 17 188 244 204
rect 17 133 105 188
rect 311 184 477 218
rect 595 202 629 364
rect 777 320 843 364
rect 663 294 743 310
rect 663 260 671 294
rect 705 260 743 294
rect 777 286 793 320
rect 827 286 843 320
rect 777 270 843 286
rect 663 236 743 260
rect 795 210 845 226
rect 595 188 661 202
rect 17 99 55 133
rect 89 99 105 133
rect 17 70 105 99
rect 139 129 205 154
rect 139 95 155 129
rect 189 95 205 129
rect 139 17 205 95
rect 311 133 377 184
rect 595 154 611 188
rect 645 154 661 188
rect 311 99 327 133
rect 361 99 377 133
rect 311 70 377 99
rect 475 127 541 150
rect 475 93 491 127
rect 525 93 541 127
rect 475 17 541 93
rect 595 120 661 154
rect 595 86 611 120
rect 645 86 661 120
rect 595 70 661 86
rect 695 188 761 202
rect 695 154 711 188
rect 745 154 761 188
rect 695 120 761 154
rect 695 86 711 120
rect 745 86 761 120
rect 695 17 761 86
rect 795 176 811 210
rect 795 120 845 176
rect 795 86 811 120
rect 889 119 923 448
rect 957 398 1001 414
rect 957 364 964 398
rect 998 364 1001 398
rect 957 330 1001 364
rect 957 296 964 330
rect 998 296 1001 330
rect 957 221 1001 296
rect 1035 289 1069 453
rect 1135 389 1169 469
rect 1397 435 1431 482
rect 1103 373 1169 389
rect 1103 339 1106 373
rect 1140 355 1169 373
rect 1203 409 1431 435
rect 1203 375 1219 409
rect 1253 401 1431 409
rect 1465 428 1499 579
rect 1533 520 1583 649
rect 1717 588 2086 615
rect 1717 554 1733 588
rect 1767 581 2086 588
rect 1767 554 1783 581
rect 1567 486 1583 520
rect 1533 462 1583 486
rect 1623 529 1673 545
rect 1717 538 1783 554
rect 2020 571 2086 581
rect 1657 504 1673 529
rect 1913 531 1979 547
rect 1913 504 1929 531
rect 1657 497 1929 504
rect 1963 497 1979 531
rect 2020 537 2036 571
rect 2070 537 2086 571
rect 2020 512 2086 537
rect 2126 571 2160 649
rect 2126 512 2160 537
rect 2200 567 2274 596
rect 2200 533 2216 567
rect 2250 533 2274 567
rect 1657 495 1979 497
rect 1623 470 1979 495
rect 2200 478 2274 533
rect 1623 434 1673 470
rect 1913 442 1979 470
rect 1253 375 1269 401
rect 1465 394 1589 428
rect 1203 359 1269 375
rect 1140 339 1146 355
rect 1103 323 1146 339
rect 1330 351 1387 367
rect 1330 321 1337 351
rect 1180 317 1337 321
rect 1371 317 1387 351
rect 1180 289 1387 317
rect 1429 351 1511 360
rect 1429 317 1445 351
rect 1479 350 1511 351
rect 1429 316 1471 317
rect 1505 316 1511 350
rect 1555 350 1589 394
rect 1657 400 1673 434
rect 1623 384 1673 400
rect 1818 420 1873 436
rect 1818 386 1838 420
rect 1872 386 1873 420
rect 1913 408 1929 442
rect 1963 408 1979 442
rect 1913 392 1979 408
rect 2013 444 2274 478
rect 2308 567 2374 596
rect 2308 533 2324 567
rect 2358 533 2374 567
rect 2308 478 2374 533
rect 2414 571 2464 649
rect 2448 537 2464 571
rect 2414 512 2464 537
rect 2506 559 2572 575
rect 2506 525 2522 559
rect 2556 525 2572 559
rect 2308 444 2388 478
rect 1818 358 1873 386
rect 2013 358 2047 444
rect 2240 410 2274 444
rect 1555 316 1768 350
rect 1818 324 2047 358
rect 2137 394 2206 410
rect 2137 360 2156 394
rect 2190 360 2206 394
rect 2137 350 2206 360
rect 1429 308 1511 316
rect 1035 287 1387 289
rect 1035 255 1214 287
rect 1330 274 1387 287
rect 1734 290 1768 316
rect 1552 274 1686 282
rect 957 187 1041 221
rect 957 119 973 153
rect 795 85 845 86
rect 1007 85 1041 187
rect 795 51 1041 85
rect 1075 140 1125 255
rect 1248 237 1296 253
rect 1330 240 1568 274
rect 1602 240 1636 274
rect 1670 240 1686 274
rect 1248 203 1255 237
rect 1289 206 1296 237
rect 1552 224 1686 240
rect 1734 274 1800 290
rect 1734 240 1750 274
rect 1784 240 1800 274
rect 1734 224 1800 240
rect 1289 203 1401 206
rect 1248 177 1401 203
rect 1839 188 1873 324
rect 2137 316 2143 350
rect 2177 326 2206 350
rect 2137 292 2156 316
rect 2190 292 2206 326
rect 2137 276 2206 292
rect 2240 394 2320 410
rect 2240 360 2270 394
rect 2304 360 2320 394
rect 2240 326 2320 360
rect 2240 292 2270 326
rect 2304 292 2320 326
rect 2240 276 2320 292
rect 1958 246 2092 262
rect 1958 212 1974 246
rect 2008 212 2042 246
rect 2076 242 2092 246
rect 2354 242 2388 444
rect 2076 212 2388 242
rect 1958 208 2388 212
rect 2506 449 2572 525
rect 2506 415 2522 449
rect 2556 415 2572 449
rect 2506 399 2572 415
rect 2606 559 2672 649
rect 2606 525 2622 559
rect 2656 525 2672 559
rect 2606 449 2672 525
rect 2606 415 2622 449
rect 2656 415 2672 449
rect 2606 399 2672 415
rect 2713 580 2763 596
rect 2747 546 2763 580
rect 2713 497 2763 546
rect 2747 463 2763 497
rect 2713 414 2763 463
rect 2506 310 2540 399
rect 2747 380 2763 414
rect 2506 294 2679 310
rect 2506 260 2629 294
rect 2663 260 2679 294
rect 2506 244 2679 260
rect 1958 196 2354 208
rect 2506 201 2540 244
rect 2713 210 2763 380
rect 1248 172 1351 177
rect 1109 106 1125 140
rect 1335 143 1351 172
rect 1385 143 1401 177
rect 1075 77 1125 106
rect 1223 132 1289 138
rect 1223 98 1239 132
rect 1273 98 1289 132
rect 1335 114 1401 143
rect 1491 154 1515 188
rect 1549 154 1611 188
rect 1645 154 1661 188
rect 1491 120 1661 154
rect 1223 17 1289 98
rect 1491 86 1531 120
rect 1565 86 1611 120
rect 1645 86 1661 120
rect 1491 17 1661 86
rect 1759 154 1797 188
rect 1831 154 1873 188
rect 1759 120 1873 154
rect 1759 86 1797 120
rect 1831 86 1873 120
rect 1759 70 1873 86
rect 2165 133 2231 162
rect 2165 99 2181 133
rect 2215 99 2231 133
rect 2165 17 2231 99
rect 2279 133 2354 196
rect 2474 185 2540 201
rect 2474 174 2490 185
rect 2279 99 2295 133
rect 2329 99 2354 133
rect 2391 158 2490 174
rect 2391 124 2407 158
rect 2441 151 2490 158
rect 2524 151 2540 185
rect 2441 124 2540 151
rect 2391 108 2540 124
rect 2576 194 2642 210
rect 2576 160 2592 194
rect 2626 160 2642 194
rect 2576 120 2642 160
rect 2279 70 2354 99
rect 2576 86 2592 120
rect 2626 86 2642 120
rect 2576 17 2642 86
rect 2676 194 2763 210
rect 2676 160 2692 194
rect 2726 160 2763 194
rect 2676 120 2763 160
rect 2676 86 2692 120
rect 2726 86 2763 120
rect 2676 70 2763 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 1471 317 1479 350
rect 1479 317 1505 350
rect 1471 316 1505 317
rect 2143 326 2177 350
rect 2143 316 2156 326
rect 2156 316 2177 326
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
<< metal1 >>
rect 0 683 2784 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 0 617 2784 649
rect 1459 350 1517 356
rect 1459 316 1471 350
rect 1505 347 1517 350
rect 2131 350 2189 356
rect 2131 347 2143 350
rect 1505 319 2143 347
rect 1505 316 1517 319
rect 1459 310 1517 316
rect 2131 316 2143 319
rect 2177 316 2189 350
rect 2131 310 2189 316
rect 0 17 2784 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
rect 0 -49 2784 -17
<< labels >>
rlabel comment s 0 0 0 0 4 sdfstp_1
flabel comment s 1253 276 1253 276 0 FreeSans 200 0 0 0 no_jumper_check
flabel comment s 1044 344 1044 344 0 FreeSans 200 0 0 0 no_jumper_check
flabel pwell s 0 0 2784 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 0 617 2784 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 2143 316 2177 350 0 FreeSans 340 0 0 0 SET_B
port 5 nsew
flabel metal1 s 0 617 2784 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 2784 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 2719 94 2753 128 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2719 168 2753 202 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2719 242 2753 276 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2719 316 2753 350 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2719 390 2753 424 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2719 464 2753 498 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2719 538 2753 572 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 511 242 545 276 0 FreeSans 340 0 0 0 SCD
port 3 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 SCD
port 3 nsew
flabel corelocali s 511 390 545 424 0 FreeSans 340 0 0 0 SCD
port 3 nsew
flabel corelocali s 703 242 737 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 SCE
port 4 nsew
flabel corelocali s 223 390 257 424 0 FreeSans 340 0 0 0 D
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 2784 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 362364
string GDS_START 341620
<< end >>
