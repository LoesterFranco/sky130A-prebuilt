magic
tech sky130A
magscale 1 2
timestamp 1599588209
<< nwell >>
rect -38 332 1958 704
<< pwell >>
rect 0 0 1920 49
<< scpmos >>
rect 127 376 157 576
rect 241 376 271 576
rect 420 376 450 576
rect 510 376 540 576
rect 632 368 662 592
rect 722 368 752 592
rect 812 368 842 592
rect 902 368 932 592
rect 1157 392 1187 592
rect 1247 392 1277 592
rect 1337 392 1367 592
rect 1427 392 1457 592
rect 1575 392 1605 592
rect 1673 392 1703 592
<< nmoslvt >>
rect 124 135 154 263
rect 210 135 240 263
rect 477 123 507 251
rect 563 123 593 251
rect 661 100 691 248
rect 747 100 777 248
rect 833 100 863 248
rect 919 100 949 248
rect 1097 120 1127 248
rect 1183 120 1213 248
rect 1316 123 1346 251
rect 1402 123 1432 251
rect 1598 76 1628 204
rect 1684 76 1714 204
<< ndiff >>
rect 71 183 124 263
rect 71 149 79 183
rect 113 149 124 183
rect 71 135 124 149
rect 154 250 210 263
rect 154 216 165 250
rect 199 216 210 250
rect 154 135 210 216
rect 240 224 293 263
rect 240 190 251 224
rect 285 190 293 224
rect 240 135 293 190
rect 424 191 477 251
rect 424 157 432 191
rect 466 157 477 191
rect 424 123 477 157
rect 507 228 563 251
rect 507 194 518 228
rect 552 194 563 228
rect 507 123 563 194
rect 593 248 643 251
rect 1263 248 1316 251
rect 593 149 661 248
rect 593 123 616 149
rect 608 115 616 123
rect 650 115 661 149
rect 608 100 661 115
rect 691 220 747 248
rect 691 186 702 220
rect 736 186 747 220
rect 691 146 747 186
rect 691 112 702 146
rect 736 112 747 146
rect 691 100 747 112
rect 777 149 833 248
rect 777 115 788 149
rect 822 115 833 149
rect 777 100 833 115
rect 863 220 919 248
rect 863 186 874 220
rect 908 186 919 220
rect 863 146 919 186
rect 863 112 874 146
rect 908 112 919 146
rect 863 100 919 112
rect 949 176 1097 248
rect 949 142 960 176
rect 994 142 1052 176
rect 1086 142 1097 176
rect 949 120 1097 142
rect 1127 236 1183 248
rect 1127 202 1138 236
rect 1172 202 1183 236
rect 1127 166 1183 202
rect 1127 132 1138 166
rect 1172 132 1183 166
rect 1127 120 1183 132
rect 1213 240 1316 248
rect 1213 206 1271 240
rect 1305 206 1316 240
rect 1213 169 1316 206
rect 1213 135 1242 169
rect 1276 135 1316 169
rect 1213 123 1316 135
rect 1346 228 1402 251
rect 1346 194 1357 228
rect 1391 194 1402 228
rect 1346 123 1402 194
rect 1432 202 1485 251
rect 1432 168 1443 202
rect 1477 168 1485 202
rect 1432 123 1485 168
rect 1213 120 1263 123
rect 949 100 1002 120
rect 1545 192 1598 204
rect 1545 158 1553 192
rect 1587 158 1598 192
rect 1545 122 1598 158
rect 1545 88 1553 122
rect 1587 88 1598 122
rect 1545 76 1598 88
rect 1628 169 1684 204
rect 1628 135 1639 169
rect 1673 135 1684 169
rect 1628 76 1684 135
rect 1714 192 1781 204
rect 1714 158 1730 192
rect 1764 158 1781 192
rect 1714 124 1781 158
rect 1714 90 1730 124
rect 1764 90 1781 124
rect 1714 76 1781 90
<< pdiff >>
rect 577 577 632 592
rect 577 576 585 577
rect 72 554 127 576
rect 72 520 80 554
rect 114 520 127 554
rect 72 486 127 520
rect 72 452 80 486
rect 114 452 127 486
rect 72 376 127 452
rect 157 568 241 576
rect 157 534 194 568
rect 228 534 241 568
rect 157 486 241 534
rect 157 452 194 486
rect 228 452 241 486
rect 157 376 241 452
rect 271 559 420 576
rect 271 525 295 559
rect 329 525 363 559
rect 397 525 420 559
rect 271 376 420 525
rect 450 568 510 576
rect 450 534 463 568
rect 497 534 510 568
rect 450 486 510 534
rect 450 452 463 486
rect 497 452 510 486
rect 450 376 510 452
rect 540 543 585 576
rect 619 543 632 577
rect 540 376 632 543
rect 577 368 632 376
rect 662 427 722 592
rect 662 393 675 427
rect 709 393 722 427
rect 662 368 722 393
rect 752 577 812 592
rect 752 543 765 577
rect 799 543 812 577
rect 752 368 812 543
rect 842 427 902 592
rect 842 393 855 427
rect 889 393 902 427
rect 842 368 902 393
rect 932 577 987 592
rect 932 543 945 577
rect 979 543 987 577
rect 932 368 987 543
rect 1102 577 1157 592
rect 1102 543 1110 577
rect 1144 543 1157 577
rect 1102 392 1157 543
rect 1187 438 1247 592
rect 1187 404 1200 438
rect 1234 404 1247 438
rect 1187 392 1247 404
rect 1277 577 1337 592
rect 1277 543 1290 577
rect 1324 543 1337 577
rect 1277 392 1337 543
rect 1367 531 1427 592
rect 1367 497 1380 531
rect 1414 497 1427 531
rect 1367 438 1427 497
rect 1367 404 1380 438
rect 1414 404 1427 438
rect 1367 392 1427 404
rect 1457 580 1575 592
rect 1457 546 1501 580
rect 1535 546 1575 580
rect 1457 493 1575 546
rect 1457 459 1501 493
rect 1535 459 1575 493
rect 1457 392 1575 459
rect 1605 540 1673 592
rect 1605 506 1622 540
rect 1656 506 1673 540
rect 1605 438 1673 506
rect 1605 404 1622 438
rect 1656 404 1673 438
rect 1605 392 1673 404
rect 1703 580 1758 592
rect 1703 546 1716 580
rect 1750 546 1758 580
rect 1703 509 1758 546
rect 1703 475 1716 509
rect 1750 475 1758 509
rect 1703 438 1758 475
rect 1703 404 1716 438
rect 1750 404 1758 438
rect 1703 392 1758 404
<< ndiffc >>
rect 79 149 113 183
rect 165 216 199 250
rect 251 190 285 224
rect 432 157 466 191
rect 518 194 552 228
rect 616 115 650 149
rect 702 186 736 220
rect 702 112 736 146
rect 788 115 822 149
rect 874 186 908 220
rect 874 112 908 146
rect 960 142 994 176
rect 1052 142 1086 176
rect 1138 202 1172 236
rect 1138 132 1172 166
rect 1271 206 1305 240
rect 1242 135 1276 169
rect 1357 194 1391 228
rect 1443 168 1477 202
rect 1553 158 1587 192
rect 1553 88 1587 122
rect 1639 135 1673 169
rect 1730 158 1764 192
rect 1730 90 1764 124
<< pdiffc >>
rect 80 520 114 554
rect 80 452 114 486
rect 194 534 228 568
rect 194 452 228 486
rect 295 525 329 559
rect 363 525 397 559
rect 463 534 497 568
rect 463 452 497 486
rect 585 543 619 577
rect 675 393 709 427
rect 765 543 799 577
rect 855 393 889 427
rect 945 543 979 577
rect 1110 543 1144 577
rect 1200 404 1234 438
rect 1290 543 1324 577
rect 1380 497 1414 531
rect 1380 404 1414 438
rect 1501 546 1535 580
rect 1501 459 1535 493
rect 1622 506 1656 540
rect 1622 404 1656 438
rect 1716 546 1750 580
rect 1716 475 1750 509
rect 1716 404 1750 438
<< poly >>
rect 127 576 157 602
rect 241 576 271 602
rect 420 576 450 602
rect 510 576 540 602
rect 632 592 662 618
rect 722 592 752 618
rect 812 592 842 618
rect 902 592 932 618
rect 1157 592 1187 618
rect 1247 592 1277 618
rect 1337 592 1367 618
rect 1427 592 1457 618
rect 1575 592 1605 618
rect 1673 592 1703 618
rect 127 361 157 376
rect 241 361 271 376
rect 420 361 450 376
rect 510 361 540 376
rect 1157 377 1187 392
rect 1247 377 1277 392
rect 1337 377 1367 392
rect 1427 377 1457 392
rect 1575 377 1605 392
rect 1673 377 1703 392
rect 124 278 160 361
rect 238 308 274 361
rect 210 278 274 308
rect 417 296 453 361
rect 507 296 543 361
rect 632 353 662 368
rect 722 353 752 368
rect 812 353 842 368
rect 902 353 932 368
rect 1154 360 1190 377
rect 632 338 665 353
rect 719 338 755 353
rect 809 338 845 353
rect 899 338 935 353
rect 635 320 935 338
rect 635 308 735 320
rect 124 263 154 278
rect 210 263 240 278
rect 417 266 593 296
rect 477 251 507 266
rect 563 251 593 266
rect 661 286 735 308
rect 769 286 803 320
rect 837 286 871 320
rect 905 300 935 320
rect 1081 344 1190 360
rect 1081 310 1097 344
rect 1131 318 1190 344
rect 1244 325 1280 377
rect 1334 355 1370 377
rect 1424 355 1460 377
rect 1334 325 1510 355
rect 1244 318 1274 325
rect 1131 310 1274 318
rect 905 286 949 300
rect 1081 288 1274 310
rect 661 270 949 286
rect 124 113 154 135
rect 210 113 240 135
rect 661 248 691 270
rect 747 248 777 270
rect 833 248 863 270
rect 919 248 949 270
rect 1097 248 1127 288
rect 1183 248 1213 288
rect 1316 251 1346 277
rect 1402 251 1432 325
rect 1480 296 1510 325
rect 1572 344 1608 377
rect 1670 344 1706 377
rect 1572 314 1856 344
rect 1598 310 1856 314
rect 1480 266 1530 296
rect 124 97 353 113
rect 477 101 507 123
rect 124 83 303 97
rect 287 63 303 83
rect 337 63 353 97
rect 287 47 353 63
rect 455 85 521 101
rect 563 97 593 123
rect 455 51 471 85
rect 505 51 521 85
rect 661 74 691 100
rect 747 74 777 100
rect 833 74 863 100
rect 919 74 949 100
rect 1097 94 1127 120
rect 1183 94 1213 120
rect 1316 101 1346 123
rect 1294 85 1360 101
rect 1402 97 1432 123
rect 455 35 521 51
rect 1294 51 1310 85
rect 1344 55 1360 85
rect 1500 55 1530 266
rect 1598 276 1738 310
rect 1772 276 1806 310
rect 1840 276 1856 310
rect 1598 204 1628 276
rect 1684 260 1856 276
rect 1684 204 1714 260
rect 1344 51 1530 55
rect 1294 25 1530 51
rect 1598 50 1628 76
rect 1684 50 1714 76
<< polycont >>
rect 735 286 769 320
rect 803 286 837 320
rect 871 286 905 320
rect 1097 310 1131 344
rect 303 63 337 97
rect 471 51 505 85
rect 1310 51 1344 85
rect 1738 276 1772 310
rect 1806 276 1840 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 64 554 130 649
rect 64 520 80 554
rect 114 520 130 554
rect 64 486 130 520
rect 64 452 80 486
rect 114 452 130 486
rect 178 568 244 580
rect 178 534 194 568
rect 228 534 244 568
rect 178 486 244 534
rect 279 559 413 649
rect 279 525 295 559
rect 329 525 363 559
rect 397 525 413 559
rect 279 520 413 525
rect 447 568 513 580
rect 447 534 463 568
rect 497 534 513 568
rect 569 577 635 649
rect 569 543 585 577
rect 619 543 635 577
rect 569 540 635 543
rect 749 577 815 649
rect 749 543 765 577
rect 799 543 815 577
rect 749 540 815 543
rect 929 577 995 649
rect 929 543 945 577
rect 979 543 995 577
rect 929 540 995 543
rect 1094 581 1766 615
rect 1094 577 1340 581
rect 1094 543 1110 577
rect 1144 543 1290 577
rect 1324 543 1340 577
rect 1485 580 1551 581
rect 1094 540 1340 543
rect 447 506 513 534
rect 1374 531 1430 547
rect 1374 506 1380 531
rect 447 497 1380 506
rect 1414 497 1430 531
rect 447 486 1430 497
rect 178 452 194 486
rect 228 452 463 486
rect 497 472 1430 486
rect 497 452 513 472
rect 1364 438 1430 472
rect 1485 546 1501 580
rect 1535 546 1551 580
rect 1716 580 1766 581
rect 1485 493 1551 546
rect 1485 459 1501 493
rect 1535 459 1551 493
rect 1485 456 1551 459
rect 1602 540 1676 547
rect 1602 506 1622 540
rect 1656 506 1676 540
rect 570 427 905 438
rect 570 418 675 427
rect 25 393 675 418
rect 709 393 855 427
rect 889 393 905 427
rect 25 384 905 393
rect 25 276 71 384
rect 25 242 31 276
rect 65 242 71 276
rect 25 236 71 242
rect 149 320 976 350
rect 149 316 735 320
rect 149 250 215 316
rect 719 286 735 316
rect 769 286 803 320
rect 837 286 871 320
rect 905 286 976 320
rect 1081 344 1147 430
rect 1081 310 1097 344
rect 1131 310 1147 344
rect 1081 294 1147 310
rect 1184 404 1200 438
rect 1234 404 1250 438
rect 1184 354 1250 404
rect 1364 404 1380 438
rect 1414 422 1430 438
rect 1602 438 1676 506
rect 1602 422 1622 438
rect 1414 404 1622 422
rect 1656 404 1676 438
rect 1364 388 1676 404
rect 1750 546 1766 580
rect 1716 509 1766 546
rect 1750 475 1766 509
rect 1716 438 1766 475
rect 1750 404 1766 438
rect 1716 388 1766 404
rect 1184 320 1689 354
rect 149 216 165 250
rect 199 216 215 250
rect 149 215 215 216
rect 251 248 552 282
rect 251 224 285 248
rect 63 183 113 202
rect 63 149 79 183
rect 502 228 552 248
rect 251 181 285 190
rect 113 149 285 181
rect 63 147 285 149
rect 63 131 113 147
rect 319 113 353 208
rect 287 97 353 113
rect 287 63 303 97
rect 337 63 353 97
rect 287 51 353 63
rect 387 191 466 214
rect 387 157 432 191
rect 502 194 518 228
rect 601 276 647 282
rect 601 242 607 276
rect 641 242 647 276
rect 719 270 976 286
rect 601 236 647 242
rect 942 260 976 270
rect 1184 260 1218 320
rect 942 236 1218 260
rect 601 220 908 236
rect 942 226 1138 236
rect 601 202 702 220
rect 502 168 552 194
rect 686 186 702 202
rect 736 202 874 220
rect 736 186 752 202
rect 387 135 466 157
rect 600 149 650 168
rect 387 17 421 135
rect 505 101 551 134
rect 455 85 551 101
rect 455 51 471 85
rect 505 51 551 85
rect 600 115 616 149
rect 600 17 650 115
rect 686 146 752 186
rect 858 186 874 202
rect 1122 202 1138 226
rect 1172 226 1218 236
rect 1255 240 1305 256
rect 1172 202 1188 226
rect 686 112 702 146
rect 736 112 752 146
rect 686 88 752 112
rect 788 149 822 168
rect 788 17 822 115
rect 858 146 908 186
rect 858 112 874 146
rect 858 96 908 112
rect 944 176 1088 192
rect 944 142 960 176
rect 994 142 1052 176
rect 1086 142 1088 176
rect 944 17 1088 142
rect 1122 166 1188 202
rect 1255 206 1271 240
rect 1255 192 1305 206
rect 1122 132 1138 166
rect 1172 132 1188 166
rect 1122 116 1188 132
rect 1226 169 1305 192
rect 1226 135 1242 169
rect 1276 135 1305 169
rect 1341 252 1587 286
rect 1341 228 1407 252
rect 1341 194 1357 228
rect 1391 194 1407 228
rect 1341 168 1407 194
rect 1443 202 1493 218
rect 1477 168 1493 202
rect 1226 17 1260 135
rect 1369 101 1409 134
rect 1294 85 1409 101
rect 1294 51 1310 85
rect 1344 51 1409 85
rect 1443 17 1493 168
rect 1537 192 1587 252
rect 1537 158 1553 192
rect 1537 122 1587 158
rect 1537 88 1553 122
rect 1623 169 1689 320
rect 1723 310 1899 350
rect 1723 276 1738 310
rect 1772 276 1806 310
rect 1840 276 1899 310
rect 1723 260 1899 276
rect 1819 242 1899 260
rect 1623 135 1639 169
rect 1673 135 1689 169
rect 1623 119 1689 135
rect 1725 192 1785 208
rect 1725 158 1730 192
rect 1764 158 1785 192
rect 1725 124 1785 158
rect 1537 85 1587 88
rect 1725 90 1730 124
rect 1764 90 1785 124
rect 1725 85 1785 90
rect 1537 51 1785 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 31 242 65 276
rect 607 242 641 276
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
<< metal1 >>
rect 0 683 1920 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 0 617 1920 649
rect 19 276 77 282
rect 19 242 31 276
rect 65 273 77 276
rect 595 276 653 282
rect 595 273 607 276
rect 65 245 607 273
rect 65 242 77 245
rect 19 236 77 242
rect 595 242 607 245
rect 641 242 653 276
rect 595 236 653 242
rect 0 17 1920 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
rect 0 -49 1920 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a221o_4
flabel pwell s 0 0 1920 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nwell s 0 617 1920 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 607 242 641 276 0 FreeSans 340 0 0 0 X
port 10 nsew
flabel metal1 s 0 617 1920 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 1920 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 1087 316 1121 350 0 FreeSans 340 0 0 0 C1
port 5 nsew
flabel corelocali s 1087 390 1121 424 0 FreeSans 340 0 0 0 C1
port 5 nsew
flabel corelocali s 1759 316 1793 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 1855 316 1889 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 511 94 545 128 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 1375 94 1409 128 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 319 94 353 128 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 319 168 353 202 0 FreeSans 340 0 0 0 A1
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 1920 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3527996
string GDS_START 3514544
<< end >>
