magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1656 561
rect 103 425 175 527
rect 17 199 66 323
rect 291 379 357 527
rect 459 379 525 527
rect 627 379 693 527
rect 795 379 861 527
rect 974 323 1040 425
rect 1142 323 1208 425
rect 1310 323 1376 425
rect 1478 323 1544 425
rect 974 289 1544 323
rect 974 170 1050 289
rect 1084 204 1639 255
rect 103 17 169 97
rect 275 17 341 97
rect 443 17 509 97
rect 611 17 677 97
rect 779 17 847 97
rect 974 127 1639 170
rect 0 -17 1656 17
<< obsli1 >>
rect 17 391 69 493
rect 17 357 175 391
rect 100 265 175 357
rect 215 345 257 493
rect 391 345 425 493
rect 559 345 593 493
rect 727 345 761 493
rect 895 459 1639 493
rect 895 345 940 459
rect 215 311 940 345
rect 1074 357 1108 459
rect 1242 357 1276 459
rect 1410 357 1444 459
rect 1578 289 1639 459
rect 100 199 940 265
rect 100 165 139 199
rect 17 131 139 165
rect 207 131 940 165
rect 17 51 69 131
rect 207 51 241 131
rect 375 51 409 131
rect 543 51 577 131
rect 711 51 745 131
rect 881 93 940 131
rect 881 51 1639 93
<< metal1 >>
rect 0 496 1656 592
rect 0 -48 1656 48
<< labels >>
rlabel locali s 1084 204 1639 255 6 A
port 1 nsew signal input
rlabel locali s 17 199 66 323 6 TE
port 2 nsew signal input
rlabel locali s 1478 323 1544 425 6 Z
port 3 nsew signal output
rlabel locali s 1310 323 1376 425 6 Z
port 3 nsew signal output
rlabel locali s 1142 323 1208 425 6 Z
port 3 nsew signal output
rlabel locali s 974 323 1040 425 6 Z
port 3 nsew signal output
rlabel locali s 974 289 1544 323 6 Z
port 3 nsew signal output
rlabel locali s 974 170 1050 289 6 Z
port 3 nsew signal output
rlabel locali s 974 127 1639 170 6 Z
port 3 nsew signal output
rlabel locali s 779 17 847 97 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 611 17 677 97 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 443 17 509 97 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 275 17 341 97 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 103 17 169 97 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 1656 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1656 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 795 379 861 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 627 379 693 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 459 379 525 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 291 379 357 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 103 425 175 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 1656 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 1656 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1656 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2006066
string GDS_START 1993444
<< end >>
