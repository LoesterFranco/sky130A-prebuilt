magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1932 561
rect 115 323 165 425
rect 283 323 333 425
rect 1235 443 1637 527
rect 1755 359 1789 527
rect 115 289 341 323
rect 719 289 1159 323
rect 301 255 341 289
rect 719 265 753 289
rect 18 215 267 255
rect 301 219 649 255
rect 301 181 341 219
rect 23 17 73 179
rect 107 145 341 181
rect 107 51 173 145
rect 207 17 241 111
rect 275 51 341 145
rect 375 129 581 185
rect 615 164 649 219
rect 683 199 753 265
rect 787 199 1057 255
rect 1093 215 1159 289
rect 1193 289 1653 323
rect 1193 215 1259 289
rect 1619 255 1653 289
rect 1295 215 1577 255
rect 1619 215 1915 255
rect 1102 164 1292 181
rect 615 147 1553 164
rect 615 129 1136 147
rect 1258 129 1553 147
rect 375 17 409 129
rect 547 119 581 129
rect 1167 17 1201 111
rect 1671 17 1705 111
rect 1839 17 1873 181
rect 0 -17 1932 17
<< obsli1 >>
rect 18 459 425 493
rect 18 289 81 459
rect 199 357 249 459
rect 375 323 425 459
rect 463 443 1201 493
rect 463 359 513 443
rect 1151 409 1201 443
rect 1671 409 1705 493
rect 547 367 1117 409
rect 547 323 606 367
rect 1151 357 1721 409
rect 1687 323 1721 357
rect 1831 323 1881 493
rect 375 289 606 323
rect 1687 289 1881 323
rect 1587 145 1805 181
rect 447 85 522 95
rect 607 85 1117 95
rect 447 51 1117 85
rect 1587 95 1637 145
rect 1235 51 1637 95
rect 1739 51 1805 145
<< metal1 >>
rect 0 496 1932 592
rect 0 -48 1932 48
<< labels >>
rlabel locali s 1295 215 1577 255 6 A1
port 1 nsew signal input
rlabel locali s 1619 255 1653 289 6 A2
port 2 nsew signal input
rlabel locali s 1619 215 1915 255 6 A2
port 2 nsew signal input
rlabel locali s 1193 289 1653 323 6 A2
port 2 nsew signal input
rlabel locali s 1193 215 1259 289 6 A2
port 2 nsew signal input
rlabel locali s 787 199 1057 255 6 B1
port 3 nsew signal input
rlabel locali s 1093 215 1159 289 6 B2
port 4 nsew signal input
rlabel locali s 719 289 1159 323 6 B2
port 4 nsew signal input
rlabel locali s 719 265 753 289 6 B2
port 4 nsew signal input
rlabel locali s 683 199 753 265 6 B2
port 4 nsew signal input
rlabel locali s 18 215 267 255 6 C1
port 5 nsew signal input
rlabel locali s 1258 129 1553 147 6 Y
port 6 nsew signal output
rlabel locali s 1102 164 1292 181 6 Y
port 6 nsew signal output
rlabel locali s 615 164 649 219 6 Y
port 6 nsew signal output
rlabel locali s 615 147 1553 164 6 Y
port 6 nsew signal output
rlabel locali s 615 129 1136 147 6 Y
port 6 nsew signal output
rlabel locali s 301 255 341 289 6 Y
port 6 nsew signal output
rlabel locali s 301 219 649 255 6 Y
port 6 nsew signal output
rlabel locali s 301 181 341 219 6 Y
port 6 nsew signal output
rlabel locali s 283 323 333 425 6 Y
port 6 nsew signal output
rlabel locali s 275 51 341 145 6 Y
port 6 nsew signal output
rlabel locali s 115 323 165 425 6 Y
port 6 nsew signal output
rlabel locali s 115 289 341 323 6 Y
port 6 nsew signal output
rlabel locali s 107 145 341 181 6 Y
port 6 nsew signal output
rlabel locali s 107 51 173 145 6 Y
port 6 nsew signal output
rlabel locali s 1839 17 1873 181 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1671 17 1705 111 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1167 17 1201 111 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 547 119 581 129 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 375 129 581 185 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 375 17 409 129 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 207 17 241 111 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 23 17 73 179 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 1932 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1932 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1755 359 1789 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1235 443 1637 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 1932 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 1932 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1932 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 4120944
string GDS_START 4107722
<< end >>
