magic
tech sky130A
magscale 1 2
timestamp 1599588209
<< nwell >>
rect -38 332 710 704
<< pwell >>
rect 0 0 672 49
<< scpmos >>
rect 86 368 116 592
rect 176 368 206 592
rect 266 368 296 592
rect 356 368 386 592
rect 556 464 586 592
<< nmoslvt >>
rect 93 74 123 222
rect 179 74 209 222
rect 265 74 295 222
rect 351 74 381 222
rect 555 140 585 224
<< ndiff >>
rect 36 202 93 222
rect 36 168 48 202
rect 82 168 93 202
rect 36 120 93 168
rect 36 86 48 120
rect 82 86 93 120
rect 36 74 93 86
rect 123 181 179 222
rect 123 147 134 181
rect 168 147 179 181
rect 123 74 179 147
rect 209 210 265 222
rect 209 176 220 210
rect 254 176 265 210
rect 209 120 265 176
rect 209 86 220 120
rect 254 86 265 120
rect 209 74 265 86
rect 295 188 351 222
rect 295 154 306 188
rect 340 154 351 188
rect 295 120 351 154
rect 295 86 306 120
rect 340 86 351 120
rect 295 74 351 86
rect 381 210 438 222
rect 381 176 392 210
rect 426 176 438 210
rect 381 120 438 176
rect 381 86 392 120
rect 426 86 438 120
rect 498 207 555 224
rect 498 173 510 207
rect 544 173 555 207
rect 498 140 555 173
rect 585 186 645 224
rect 585 152 597 186
rect 631 152 645 186
rect 585 140 645 152
rect 381 74 438 86
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 497 86 546
rect 27 463 39 497
rect 73 463 86 497
rect 27 414 86 463
rect 27 380 39 414
rect 73 380 86 414
rect 27 368 86 380
rect 116 531 176 592
rect 116 497 129 531
rect 163 497 176 531
rect 116 414 176 497
rect 116 380 129 414
rect 163 380 176 414
rect 116 368 176 380
rect 206 580 266 592
rect 206 546 219 580
rect 253 546 266 580
rect 206 497 266 546
rect 206 463 219 497
rect 253 463 266 497
rect 206 414 266 463
rect 206 380 219 414
rect 253 380 266 414
rect 206 368 266 380
rect 296 580 356 592
rect 296 546 309 580
rect 343 546 356 580
rect 296 497 356 546
rect 296 463 309 497
rect 343 463 356 497
rect 296 414 356 463
rect 296 380 309 414
rect 343 380 356 414
rect 296 368 356 380
rect 386 580 444 592
rect 386 546 399 580
rect 433 546 444 580
rect 386 497 444 546
rect 386 463 399 497
rect 433 463 444 497
rect 498 580 556 592
rect 498 546 509 580
rect 543 546 556 580
rect 498 510 556 546
rect 498 476 509 510
rect 543 476 556 510
rect 498 464 556 476
rect 586 580 645 592
rect 586 546 599 580
rect 633 546 645 580
rect 586 510 645 546
rect 586 476 599 510
rect 633 476 645 510
rect 586 464 645 476
rect 386 414 444 463
rect 386 380 399 414
rect 433 380 444 414
rect 386 368 444 380
<< ndiffc >>
rect 48 168 82 202
rect 48 86 82 120
rect 134 147 168 181
rect 220 176 254 210
rect 220 86 254 120
rect 306 154 340 188
rect 306 86 340 120
rect 392 176 426 210
rect 392 86 426 120
rect 510 173 544 207
rect 597 152 631 186
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 129 497 163 531
rect 129 380 163 414
rect 219 546 253 580
rect 219 463 253 497
rect 219 380 253 414
rect 309 546 343 580
rect 309 463 343 497
rect 309 380 343 414
rect 399 546 433 580
rect 399 463 433 497
rect 509 546 543 580
rect 509 476 543 510
rect 599 546 633 580
rect 599 476 633 510
rect 399 380 433 414
<< poly >>
rect 86 592 116 618
rect 176 592 206 618
rect 266 592 296 618
rect 356 592 386 618
rect 556 592 586 618
rect 556 449 586 464
rect 553 419 627 449
rect 86 353 116 368
rect 176 353 206 368
rect 266 353 296 368
rect 356 353 386 368
rect 483 361 549 377
rect 483 353 499 361
rect 83 310 119 353
rect 173 310 209 353
rect 263 327 499 353
rect 533 327 549 361
rect 263 323 549 327
rect 483 311 549 323
rect 21 294 209 310
rect 21 260 37 294
rect 71 260 209 294
rect 597 269 627 419
rect 21 244 209 260
rect 93 222 123 244
rect 179 222 209 244
rect 265 237 483 267
rect 265 222 295 237
rect 351 222 381 237
rect 453 118 483 237
rect 555 239 627 269
rect 555 224 585 239
rect 555 118 585 140
rect 453 102 585 118
rect 453 88 512 102
rect 93 48 123 74
rect 179 48 209 74
rect 265 48 295 74
rect 351 48 381 74
rect 496 68 512 88
rect 546 68 585 102
rect 496 52 585 68
<< polycont >>
rect 499 327 533 361
rect 37 260 71 294
rect 512 68 546 102
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 23 581 253 615
rect 23 580 73 581
rect 23 546 39 580
rect 219 580 253 581
rect 23 497 73 546
rect 23 463 39 497
rect 23 414 73 463
rect 23 380 39 414
rect 23 364 73 380
rect 121 531 184 547
rect 121 497 129 531
rect 163 497 184 531
rect 121 414 184 497
rect 121 380 129 414
rect 163 380 184 414
rect 21 294 87 310
rect 21 260 37 294
rect 71 260 87 294
rect 21 236 87 260
rect 121 236 184 380
rect 219 497 253 546
rect 219 414 253 463
rect 219 330 253 380
rect 293 580 343 649
rect 293 546 309 580
rect 293 497 343 546
rect 293 463 309 497
rect 293 414 343 463
rect 293 380 309 414
rect 293 364 343 380
rect 383 580 433 596
rect 383 546 399 580
rect 383 497 433 546
rect 383 463 399 497
rect 383 414 433 463
rect 383 380 399 414
rect 383 330 433 380
rect 219 296 433 330
rect 483 580 549 596
rect 483 546 509 580
rect 543 546 549 580
rect 483 510 549 546
rect 483 476 509 510
rect 543 476 549 510
rect 483 361 549 476
rect 583 580 649 649
rect 583 546 599 580
rect 633 546 649 580
rect 583 510 649 546
rect 583 476 599 510
rect 633 476 649 510
rect 583 460 649 476
rect 483 327 499 361
rect 533 327 549 361
rect 32 168 48 202
rect 82 168 98 202
rect 32 120 98 168
rect 134 181 184 236
rect 168 147 184 181
rect 134 125 184 147
rect 220 228 442 262
rect 220 210 254 228
rect 390 210 442 228
rect 32 86 48 120
rect 82 86 98 120
rect 32 85 98 86
rect 220 120 254 176
rect 220 85 254 86
rect 32 51 254 85
rect 290 188 356 194
rect 290 154 306 188
rect 340 154 356 188
rect 290 120 356 154
rect 290 86 306 120
rect 340 86 356 120
rect 290 17 356 86
rect 390 176 392 210
rect 426 176 442 210
rect 390 120 442 176
rect 483 228 549 327
rect 483 207 560 228
rect 483 173 510 207
rect 544 173 560 207
rect 483 168 560 173
rect 596 186 649 202
rect 596 152 597 186
rect 631 152 649 186
rect 390 86 392 120
rect 426 86 442 120
rect 390 70 442 86
rect 496 102 562 134
rect 496 68 512 102
rect 546 68 562 102
rect 496 52 562 68
rect 596 17 649 152
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel comment s 0 0 0 0 4 einvp_2
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 127 242 161 276 0 FreeSans 340 0 0 0 Z
port 7 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 Z
port 7 nsew
flabel corelocali s 127 390 161 424 0 FreeSans 340 0 0 0 Z
port 7 nsew
flabel corelocali s 127 464 161 498 0 FreeSans 340 0 0 0 Z
port 7 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 511 94 545 128 0 FreeSans 340 0 0 0 TE
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 672 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 2443580
string GDS_START 2436858
<< end >>
