magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 998 704
<< pwell >>
rect 0 0 960 49
<< scnmos >>
rect 137 112 167 222
rect 264 74 294 222
rect 364 74 394 222
rect 533 74 563 222
rect 633 74 663 222
rect 846 112 876 222
<< pmoshvt >>
rect 86 368 116 536
rect 283 368 313 592
rect 367 368 397 592
rect 500 368 530 592
rect 614 368 644 592
rect 844 424 874 592
<< ndiff >>
rect 27 186 137 222
rect 27 152 92 186
rect 126 152 137 186
rect 27 112 137 152
rect 167 210 264 222
rect 167 176 205 210
rect 239 176 264 210
rect 167 120 264 176
rect 167 112 205 120
rect 193 86 205 112
rect 239 86 264 120
rect 193 74 264 86
rect 294 210 364 222
rect 294 176 305 210
rect 339 176 364 210
rect 294 120 364 176
rect 294 86 305 120
rect 339 86 364 120
rect 294 74 364 86
rect 394 120 533 222
rect 394 86 405 120
rect 439 86 488 120
rect 522 86 533 120
rect 394 74 533 86
rect 563 194 633 222
rect 563 160 588 194
rect 622 160 633 194
rect 563 120 633 160
rect 563 86 588 120
rect 622 86 633 120
rect 563 74 633 86
rect 663 184 846 222
rect 663 150 697 184
rect 731 150 785 184
rect 819 150 846 184
rect 663 116 846 150
rect 663 82 697 116
rect 731 82 785 116
rect 819 112 846 116
rect 876 184 933 222
rect 876 150 887 184
rect 921 150 933 184
rect 876 112 933 150
rect 819 82 831 112
rect 663 74 831 82
<< pdiff >>
rect 134 614 265 626
rect 134 580 146 614
rect 180 580 219 614
rect 253 592 265 614
rect 253 580 283 592
rect 134 536 283 580
rect 27 524 86 536
rect 27 490 39 524
rect 73 490 86 524
rect 27 414 86 490
rect 27 380 39 414
rect 73 380 86 414
rect 27 368 86 380
rect 116 368 283 536
rect 313 368 367 592
rect 397 368 500 592
rect 530 368 614 592
rect 644 462 703 592
rect 644 428 657 462
rect 691 428 703 462
rect 644 368 703 428
rect 789 580 844 592
rect 789 546 797 580
rect 831 546 844 580
rect 789 470 844 546
rect 789 436 797 470
rect 831 436 844 470
rect 789 424 844 436
rect 874 580 933 592
rect 874 546 887 580
rect 921 546 933 580
rect 874 470 933 546
rect 874 436 887 470
rect 921 436 933 470
rect 874 424 933 436
<< ndiffc >>
rect 92 152 126 186
rect 205 176 239 210
rect 205 86 239 120
rect 305 176 339 210
rect 305 86 339 120
rect 405 86 439 120
rect 488 86 522 120
rect 588 160 622 194
rect 588 86 622 120
rect 697 150 731 184
rect 785 150 819 184
rect 697 82 731 116
rect 785 82 819 116
rect 887 150 921 184
<< pdiffc >>
rect 146 580 180 614
rect 219 580 253 614
rect 39 490 73 524
rect 39 380 73 414
rect 657 428 691 462
rect 797 546 831 580
rect 797 436 831 470
rect 887 546 921 580
rect 887 436 921 470
<< poly >>
rect 283 592 313 618
rect 367 592 397 618
rect 500 592 530 618
rect 611 607 748 637
rect 614 592 644 607
rect 86 536 116 562
rect 86 353 116 368
rect 283 353 313 368
rect 367 353 397 368
rect 500 353 530 368
rect 614 353 644 368
rect 83 322 119 353
rect 280 336 316 353
rect 83 310 167 322
rect 21 294 167 310
rect 21 260 37 294
rect 71 260 167 294
rect 215 320 316 336
rect 215 286 231 320
rect 265 286 316 320
rect 215 270 316 286
rect 364 336 400 353
rect 497 336 533 353
rect 364 320 449 336
rect 364 286 399 320
rect 433 286 449 320
rect 364 270 449 286
rect 497 320 563 336
rect 497 286 513 320
rect 547 286 563 320
rect 497 270 563 286
rect 21 244 167 260
rect 137 222 167 244
rect 264 222 294 270
rect 364 222 394 270
rect 533 222 563 270
rect 611 310 647 353
rect 718 310 748 607
rect 844 592 874 618
rect 844 409 874 424
rect 841 356 877 409
rect 611 294 748 310
rect 611 260 630 294
rect 664 260 698 294
rect 732 260 748 294
rect 803 340 876 356
rect 803 306 819 340
rect 853 306 876 340
rect 803 290 876 306
rect 611 244 748 260
rect 633 222 663 244
rect 846 222 876 290
rect 137 86 167 112
rect 846 86 876 112
rect 264 48 294 74
rect 364 48 394 74
rect 533 48 563 74
rect 633 48 663 74
<< polycont >>
rect 37 260 71 294
rect 231 286 265 320
rect 399 286 433 320
rect 513 286 547 320
rect 630 260 664 294
rect 698 260 732 294
rect 819 306 853 340
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 130 614 269 649
rect 130 580 146 614
rect 180 580 219 614
rect 253 580 269 614
rect 793 580 837 649
rect 793 546 797 580
rect 831 546 837 580
rect 23 524 759 546
rect 23 490 39 524
rect 73 512 759 524
rect 73 490 155 512
rect 23 414 155 490
rect 315 462 691 478
rect 23 380 39 414
rect 73 380 155 414
rect 23 364 155 380
rect 21 294 87 310
rect 21 260 37 294
rect 71 260 87 294
rect 21 236 87 260
rect 121 202 155 364
rect 215 320 281 430
rect 215 286 231 320
rect 265 286 281 320
rect 215 270 281 286
rect 315 428 657 462
rect 315 412 691 428
rect 315 226 349 412
rect 725 378 759 512
rect 793 470 837 546
rect 793 436 797 470
rect 831 436 837 470
rect 793 420 837 436
rect 871 580 937 596
rect 871 546 887 580
rect 921 546 937 580
rect 871 470 937 546
rect 871 436 887 470
rect 921 436 937 470
rect 871 420 937 436
rect 383 320 455 356
rect 383 286 399 320
rect 433 286 455 320
rect 383 270 455 286
rect 497 344 759 378
rect 497 320 563 344
rect 497 286 513 320
rect 547 286 563 320
rect 793 340 869 356
rect 497 270 563 286
rect 614 294 748 310
rect 614 260 630 294
rect 664 260 698 294
rect 732 260 748 294
rect 793 306 819 340
rect 853 306 869 340
rect 793 290 869 306
rect 614 252 748 260
rect 903 252 937 420
rect 614 244 937 252
rect 23 186 155 202
rect 23 152 92 186
rect 126 152 155 186
rect 23 136 155 152
rect 189 210 255 226
rect 189 176 205 210
rect 239 176 255 210
rect 189 120 255 176
rect 189 86 205 120
rect 239 86 255 120
rect 189 17 255 86
rect 289 210 355 226
rect 714 218 937 244
rect 289 176 305 210
rect 339 194 647 210
rect 339 176 588 194
rect 289 120 355 176
rect 572 160 588 176
rect 622 160 647 194
rect 871 184 937 218
rect 289 86 305 120
rect 339 86 355 120
rect 289 70 355 86
rect 389 120 538 136
rect 389 86 405 120
rect 439 86 488 120
rect 522 86 538 120
rect 389 17 538 86
rect 572 120 647 160
rect 572 86 588 120
rect 622 86 647 120
rect 572 70 647 86
rect 681 150 697 184
rect 731 150 785 184
rect 819 150 835 184
rect 681 116 835 150
rect 681 82 697 116
rect 731 82 785 116
rect 819 82 835 116
rect 871 150 887 184
rect 921 150 937 184
rect 871 108 937 150
rect 681 17 835 82
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
rlabel comment s 0 0 0 0 4 nor4bb_1
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 D_N
port 4 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 C_N
port 3 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 223 390 257 424 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 607 94 641 128 0 FreeSans 340 0 0 0 Y
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 960 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1183406
string GDS_START 1175944
<< end >>
