magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 236 333 312 493
rect 426 333 535 493
rect 236 299 535 333
rect 85 199 165 265
rect 203 199 267 265
rect 304 199 359 265
rect 482 97 535 299
rect 426 51 535 97
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 17 319 102 385
rect 17 165 51 319
rect 152 299 202 527
rect 358 367 392 527
rect 400 165 444 265
rect 17 131 444 165
rect 17 89 102 131
rect 152 17 218 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
rlabel locali s 85 199 165 265 6 A_N
port 1 nsew signal input
rlabel locali s 304 199 359 265 6 B
port 2 nsew signal input
rlabel locali s 203 199 267 265 6 C
port 3 nsew signal input
rlabel locali s 482 97 535 299 6 Y
port 4 nsew signal output
rlabel locali s 426 333 535 493 6 Y
port 4 nsew signal output
rlabel locali s 426 51 535 97 6 Y
port 4 nsew signal output
rlabel locali s 236 333 312 493 6 Y
port 4 nsew signal output
rlabel locali s 236 299 535 333 6 Y
port 4 nsew signal output
rlabel metal1 s 0 -48 552 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 552 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 552 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2267644
string GDS_START 2261998
<< end >>
