magic
tech sky130A
magscale 1 2
timestamp 1604502729
<< locali >>
rect 25 290 95 356
rect 323 282 389 547
rect 323 230 455 282
rect 497 264 563 356
rect 653 244 743 310
rect 697 236 743 244
rect 254 196 580 230
rect 254 70 288 196
rect 514 154 580 196
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 39 390 89 649
rect 129 388 195 596
rect 161 330 195 388
rect 233 581 463 615
rect 233 364 283 581
rect 161 264 279 330
rect 423 424 463 581
rect 503 458 569 649
rect 609 424 643 596
rect 423 390 643 424
rect 683 412 753 649
rect 423 364 463 390
rect 609 378 643 390
rect 793 378 843 596
rect 161 256 195 264
rect 54 222 195 256
rect 609 344 843 378
rect 54 90 104 222
rect 152 17 218 188
rect 324 17 390 162
rect 616 202 650 210
rect 788 202 838 226
rect 616 168 838 202
rect 616 120 650 168
rect 428 70 650 120
rect 686 17 752 134
rect 788 70 838 168
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel locali s 497 264 563 356 6 A1
port 1 nsew signal input
rlabel locali s 697 236 743 244 6 A2
port 2 nsew signal input
rlabel locali s 653 244 743 310 6 A2
port 2 nsew signal input
rlabel locali s 25 290 95 356 6 B1_N
port 3 nsew signal input
rlabel locali s 514 154 580 196 6 Y
port 4 nsew signal output
rlabel locali s 323 282 389 547 6 Y
port 4 nsew signal output
rlabel locali s 323 230 455 282 6 Y
port 4 nsew signal output
rlabel locali s 254 196 580 230 6 Y
port 4 nsew signal output
rlabel locali s 254 70 288 196 6 Y
port 4 nsew signal output
rlabel metal1 s 0 -49 864 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 617 864 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 4105984
string GDS_START 4097992
<< end >>
