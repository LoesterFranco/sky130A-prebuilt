magic
tech sky130A
magscale 1 2
timestamp 1604502710
<< nwell >>
rect -38 332 2054 704
<< pwell >>
rect 0 0 2016 49
<< scpmos >>
rect 84 368 120 592
rect 183 368 219 592
rect 283 368 319 592
rect 373 368 409 592
rect 463 368 499 592
rect 573 368 609 592
rect 663 368 699 592
rect 764 368 800 592
rect 854 368 890 592
rect 956 368 992 592
rect 1046 368 1082 592
rect 1146 368 1182 592
rect 1236 368 1272 592
rect 1336 368 1372 592
rect 1426 368 1462 592
rect 1526 368 1562 592
rect 1626 368 1662 592
rect 1716 368 1752 592
rect 1806 368 1842 592
rect 1896 368 1932 592
<< nmoslvt >>
rect 84 74 114 222
rect 184 74 214 222
rect 382 74 412 222
rect 482 74 512 222
rect 636 74 666 222
rect 722 74 752 222
rect 822 74 852 222
rect 922 74 952 222
rect 1008 74 1038 222
rect 1094 74 1124 222
rect 1292 74 1322 222
rect 1378 74 1408 222
rect 1464 74 1494 222
rect 1550 74 1580 222
rect 1636 74 1666 222
rect 1722 74 1752 222
rect 1808 74 1838 222
rect 1902 74 1932 222
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 210 184 222
rect 114 176 125 210
rect 159 176 184 210
rect 114 120 184 176
rect 114 86 125 120
rect 159 86 184 120
rect 114 74 184 86
rect 214 152 271 222
rect 214 118 225 152
rect 259 118 271 152
rect 214 74 271 118
rect 325 148 382 222
rect 325 114 337 148
rect 371 114 382 148
rect 325 74 382 114
rect 412 169 482 222
rect 412 135 437 169
rect 471 135 482 169
rect 412 74 482 135
rect 512 210 636 222
rect 512 176 523 210
rect 557 176 591 210
rect 625 176 636 210
rect 512 120 636 176
rect 512 86 523 120
rect 557 86 591 120
rect 625 86 636 120
rect 512 74 636 86
rect 666 174 722 222
rect 666 140 677 174
rect 711 140 722 174
rect 666 74 722 140
rect 752 210 822 222
rect 752 176 777 210
rect 811 176 822 210
rect 752 120 822 176
rect 752 86 777 120
rect 811 86 822 120
rect 752 74 822 86
rect 852 207 922 222
rect 852 173 877 207
rect 911 173 922 207
rect 852 74 922 173
rect 952 120 1008 222
rect 952 86 963 120
rect 997 86 1008 120
rect 952 74 1008 86
rect 1038 207 1094 222
rect 1038 173 1049 207
rect 1083 173 1094 207
rect 1038 74 1094 173
rect 1124 120 1181 222
rect 1124 86 1135 120
rect 1169 86 1181 120
rect 1124 74 1181 86
rect 1235 122 1292 222
rect 1235 88 1247 122
rect 1281 88 1292 122
rect 1235 74 1292 88
rect 1322 209 1378 222
rect 1322 175 1333 209
rect 1367 175 1378 209
rect 1322 74 1378 175
rect 1408 120 1464 222
rect 1408 86 1419 120
rect 1453 86 1464 120
rect 1408 74 1464 86
rect 1494 207 1550 222
rect 1494 173 1505 207
rect 1539 173 1550 207
rect 1494 74 1550 173
rect 1580 210 1636 222
rect 1580 176 1591 210
rect 1625 176 1636 210
rect 1580 120 1636 176
rect 1580 86 1591 120
rect 1625 86 1636 120
rect 1580 74 1636 86
rect 1666 152 1722 222
rect 1666 118 1677 152
rect 1711 118 1722 152
rect 1666 74 1722 118
rect 1752 210 1808 222
rect 1752 176 1763 210
rect 1797 176 1808 210
rect 1752 120 1808 176
rect 1752 86 1763 120
rect 1797 86 1808 120
rect 1752 74 1808 86
rect 1838 152 1902 222
rect 1838 118 1849 152
rect 1883 118 1902 152
rect 1838 74 1902 118
rect 1932 210 1989 222
rect 1932 176 1943 210
rect 1977 176 1989 210
rect 1932 120 1989 176
rect 1932 86 1943 120
rect 1977 86 1989 120
rect 1932 74 1989 86
<< pdiff >>
rect 27 580 84 592
rect 27 546 39 580
rect 73 546 84 580
rect 27 501 84 546
rect 27 467 39 501
rect 73 467 84 501
rect 27 424 84 467
rect 27 390 39 424
rect 73 390 84 424
rect 27 368 84 390
rect 120 539 183 592
rect 120 505 139 539
rect 173 505 183 539
rect 120 432 183 505
rect 120 398 139 432
rect 173 398 183 432
rect 120 368 183 398
rect 219 580 283 592
rect 219 546 239 580
rect 273 546 283 580
rect 219 498 283 546
rect 219 464 239 498
rect 273 464 283 498
rect 219 368 283 464
rect 319 531 373 592
rect 319 497 329 531
rect 363 497 373 531
rect 319 414 373 497
rect 319 380 329 414
rect 363 380 373 414
rect 319 368 373 380
rect 409 580 463 592
rect 409 546 419 580
rect 453 546 463 580
rect 409 492 463 546
rect 409 458 419 492
rect 453 458 463 492
rect 409 368 463 458
rect 499 564 573 592
rect 499 530 519 564
rect 553 530 573 564
rect 499 368 573 530
rect 609 580 663 592
rect 609 546 619 580
rect 653 546 663 580
rect 609 492 663 546
rect 609 458 619 492
rect 653 458 663 492
rect 609 368 663 458
rect 699 576 764 592
rect 699 542 709 576
rect 743 542 764 576
rect 699 368 764 542
rect 800 580 854 592
rect 800 546 810 580
rect 844 546 854 580
rect 800 504 854 546
rect 800 470 810 504
rect 844 470 854 504
rect 800 424 854 470
rect 800 390 810 424
rect 844 390 854 424
rect 800 368 854 390
rect 890 578 956 592
rect 890 544 900 578
rect 934 544 956 578
rect 890 508 956 544
rect 890 474 900 508
rect 934 474 956 508
rect 890 368 956 474
rect 992 580 1046 592
rect 992 546 1002 580
rect 1036 546 1046 580
rect 992 497 1046 546
rect 992 463 1002 497
rect 1036 463 1046 497
rect 992 414 1046 463
rect 992 380 1002 414
rect 1036 380 1046 414
rect 992 368 1046 380
rect 1082 580 1146 592
rect 1082 546 1092 580
rect 1126 546 1146 580
rect 1082 508 1146 546
rect 1082 474 1092 508
rect 1126 474 1146 508
rect 1082 368 1146 474
rect 1182 580 1236 592
rect 1182 546 1192 580
rect 1226 546 1236 580
rect 1182 502 1236 546
rect 1182 468 1192 502
rect 1226 468 1236 502
rect 1182 424 1236 468
rect 1182 390 1192 424
rect 1226 390 1236 424
rect 1182 368 1236 390
rect 1272 580 1336 592
rect 1272 546 1282 580
rect 1316 546 1336 580
rect 1272 508 1336 546
rect 1272 474 1282 508
rect 1316 474 1336 508
rect 1272 368 1336 474
rect 1372 580 1426 592
rect 1372 546 1382 580
rect 1416 546 1426 580
rect 1372 502 1426 546
rect 1372 468 1382 502
rect 1416 468 1426 502
rect 1372 424 1426 468
rect 1372 390 1382 424
rect 1416 390 1426 424
rect 1372 368 1426 390
rect 1462 580 1526 592
rect 1462 546 1472 580
rect 1506 546 1526 580
rect 1462 508 1526 546
rect 1462 474 1472 508
rect 1506 474 1526 508
rect 1462 368 1526 474
rect 1562 580 1626 592
rect 1562 546 1572 580
rect 1606 546 1626 580
rect 1562 502 1626 546
rect 1562 468 1572 502
rect 1606 468 1626 502
rect 1562 424 1626 468
rect 1562 390 1572 424
rect 1606 390 1626 424
rect 1562 368 1626 390
rect 1662 580 1716 592
rect 1662 546 1672 580
rect 1706 546 1716 580
rect 1662 508 1716 546
rect 1662 474 1672 508
rect 1706 474 1716 508
rect 1662 368 1716 474
rect 1752 580 1806 592
rect 1752 546 1762 580
rect 1796 546 1806 580
rect 1752 502 1806 546
rect 1752 468 1762 502
rect 1796 468 1806 502
rect 1752 424 1806 468
rect 1752 390 1762 424
rect 1796 390 1806 424
rect 1752 368 1806 390
rect 1842 580 1896 592
rect 1842 546 1852 580
rect 1886 546 1896 580
rect 1842 508 1896 546
rect 1842 474 1852 508
rect 1886 474 1896 508
rect 1842 368 1896 474
rect 1932 580 1988 592
rect 1932 546 1942 580
rect 1976 546 1988 580
rect 1932 502 1988 546
rect 1932 468 1942 502
rect 1976 468 1988 502
rect 1932 424 1988 468
rect 1932 390 1942 424
rect 1976 390 1988 424
rect 1932 368 1988 390
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 125 176 159 210
rect 125 86 159 120
rect 225 118 259 152
rect 337 114 371 148
rect 437 135 471 169
rect 523 176 557 210
rect 591 176 625 210
rect 523 86 557 120
rect 591 86 625 120
rect 677 140 711 174
rect 777 176 811 210
rect 777 86 811 120
rect 877 173 911 207
rect 963 86 997 120
rect 1049 173 1083 207
rect 1135 86 1169 120
rect 1247 88 1281 122
rect 1333 175 1367 209
rect 1419 86 1453 120
rect 1505 173 1539 207
rect 1591 176 1625 210
rect 1591 86 1625 120
rect 1677 118 1711 152
rect 1763 176 1797 210
rect 1763 86 1797 120
rect 1849 118 1883 152
rect 1943 176 1977 210
rect 1943 86 1977 120
<< pdiffc >>
rect 39 546 73 580
rect 39 467 73 501
rect 39 390 73 424
rect 139 505 173 539
rect 139 398 173 432
rect 239 546 273 580
rect 239 464 273 498
rect 329 497 363 531
rect 329 380 363 414
rect 419 546 453 580
rect 419 458 453 492
rect 519 530 553 564
rect 619 546 653 580
rect 619 458 653 492
rect 709 542 743 576
rect 810 546 844 580
rect 810 470 844 504
rect 810 390 844 424
rect 900 544 934 578
rect 900 474 934 508
rect 1002 546 1036 580
rect 1002 463 1036 497
rect 1002 380 1036 414
rect 1092 546 1126 580
rect 1092 474 1126 508
rect 1192 546 1226 580
rect 1192 468 1226 502
rect 1192 390 1226 424
rect 1282 546 1316 580
rect 1282 474 1316 508
rect 1382 546 1416 580
rect 1382 468 1416 502
rect 1382 390 1416 424
rect 1472 546 1506 580
rect 1472 474 1506 508
rect 1572 546 1606 580
rect 1572 468 1606 502
rect 1572 390 1606 424
rect 1672 546 1706 580
rect 1672 474 1706 508
rect 1762 546 1796 580
rect 1762 468 1796 502
rect 1762 390 1796 424
rect 1852 546 1886 580
rect 1852 474 1886 508
rect 1942 546 1976 580
rect 1942 468 1976 502
rect 1942 390 1976 424
<< poly >>
rect 84 592 120 618
rect 183 592 219 618
rect 283 592 319 618
rect 373 592 409 618
rect 463 592 499 618
rect 573 592 609 618
rect 663 592 699 618
rect 764 592 800 618
rect 854 592 890 618
rect 956 592 992 618
rect 1046 592 1082 618
rect 1146 592 1182 618
rect 1236 592 1272 618
rect 1336 592 1372 618
rect 1426 592 1462 618
rect 1526 592 1562 618
rect 1626 592 1662 618
rect 1716 592 1752 618
rect 1806 592 1842 618
rect 1896 592 1932 618
rect 84 343 120 368
rect 183 343 219 368
rect 283 343 319 368
rect 373 343 409 368
rect 463 349 499 368
rect 573 349 609 368
rect 663 349 699 368
rect 764 349 800 368
rect 84 320 409 343
rect 84 286 100 320
rect 134 286 168 320
rect 202 286 236 320
rect 270 313 409 320
rect 457 320 800 349
rect 270 286 319 313
rect 84 270 319 286
rect 457 286 473 320
rect 507 286 541 320
rect 575 286 609 320
rect 643 319 800 320
rect 854 330 890 368
rect 956 330 992 368
rect 1046 330 1082 368
rect 1146 330 1182 368
rect 643 286 752 319
rect 457 271 752 286
rect 854 314 1182 330
rect 854 280 870 314
rect 904 280 938 314
rect 972 280 1006 314
rect 1040 280 1074 314
rect 1108 300 1182 314
rect 1236 336 1272 368
rect 1336 336 1372 368
rect 1426 336 1462 368
rect 1526 336 1562 368
rect 1626 336 1662 368
rect 1716 336 1752 368
rect 1806 336 1842 368
rect 1896 336 1932 368
rect 1236 320 1580 336
rect 1108 280 1124 300
rect 854 271 1124 280
rect 84 222 114 270
rect 184 222 214 270
rect 382 241 752 271
rect 382 222 412 241
rect 482 222 512 241
rect 636 222 666 241
rect 722 222 752 241
rect 822 241 1124 271
rect 1236 286 1252 320
rect 1286 286 1320 320
rect 1354 286 1388 320
rect 1422 286 1456 320
rect 1490 286 1524 320
rect 1558 286 1580 320
rect 1236 270 1580 286
rect 1626 320 1932 336
rect 1626 286 1673 320
rect 1707 286 1741 320
rect 1775 286 1809 320
rect 1843 286 1877 320
rect 1911 286 1932 320
rect 1626 270 1932 286
rect 822 222 852 241
rect 922 222 952 241
rect 1008 222 1038 241
rect 1094 222 1124 241
rect 1292 222 1322 270
rect 1378 222 1408 270
rect 1464 222 1494 270
rect 1550 222 1580 270
rect 1636 222 1666 270
rect 1722 222 1752 270
rect 1808 222 1838 270
rect 1902 222 1932 270
rect 84 48 114 74
rect 184 48 214 74
rect 382 48 412 74
rect 482 48 512 74
rect 636 48 666 74
rect 722 48 752 74
rect 822 48 852 74
rect 922 48 952 74
rect 1008 48 1038 74
rect 1094 48 1124 74
rect 1292 48 1322 74
rect 1378 48 1408 74
rect 1464 48 1494 74
rect 1550 48 1580 74
rect 1636 48 1666 74
rect 1722 48 1752 74
rect 1808 48 1838 74
rect 1902 48 1932 74
<< polycont >>
rect 100 286 134 320
rect 168 286 202 320
rect 236 286 270 320
rect 473 286 507 320
rect 541 286 575 320
rect 609 286 643 320
rect 870 280 904 314
rect 938 280 972 314
rect 1006 280 1040 314
rect 1074 280 1108 314
rect 1252 286 1286 320
rect 1320 286 1354 320
rect 1388 286 1422 320
rect 1456 286 1490 320
rect 1524 286 1558 320
rect 1673 286 1707 320
rect 1741 286 1775 320
rect 1809 286 1843 320
rect 1877 286 1911 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 23 581 469 615
rect 23 580 89 581
rect 23 546 39 580
rect 73 546 89 580
rect 223 580 289 581
rect 23 501 89 546
rect 23 467 39 501
rect 73 467 89 501
rect 23 424 89 467
rect 23 390 39 424
rect 73 390 89 424
rect 123 539 189 547
rect 123 505 139 539
rect 173 505 189 539
rect 123 432 189 505
rect 223 546 239 580
rect 273 546 289 580
rect 403 580 469 581
rect 223 498 289 546
rect 223 464 239 498
rect 273 464 289 498
rect 223 458 289 464
rect 329 531 363 547
rect 123 398 139 432
rect 173 424 189 432
rect 329 424 363 497
rect 403 546 419 580
rect 453 546 469 580
rect 403 492 469 546
rect 503 564 569 649
rect 503 530 519 564
rect 553 530 569 564
rect 503 526 569 530
rect 603 580 669 596
rect 603 546 619 580
rect 653 546 669 580
rect 603 492 669 546
rect 709 576 759 649
rect 743 542 759 576
rect 709 526 759 542
rect 794 580 860 596
rect 794 546 810 580
rect 844 546 860 580
rect 794 504 860 546
rect 794 492 810 504
rect 403 458 419 492
rect 453 458 619 492
rect 653 470 810 492
rect 844 470 860 504
rect 653 458 860 470
rect 900 578 950 649
rect 934 544 950 578
rect 900 508 950 544
rect 934 474 950 508
rect 900 458 950 474
rect 986 580 1052 596
rect 986 546 1002 580
rect 1036 546 1052 580
rect 986 497 1052 546
rect 986 463 1002 497
rect 1036 463 1052 497
rect 794 424 860 458
rect 986 424 1052 463
rect 1092 580 1142 649
rect 1126 546 1142 580
rect 1092 508 1142 546
rect 1126 474 1142 508
rect 1092 458 1142 474
rect 1176 580 1242 596
rect 1176 546 1192 580
rect 1226 546 1242 580
rect 1176 502 1242 546
rect 1176 468 1192 502
rect 1226 468 1242 502
rect 1176 424 1242 468
rect 1282 580 1332 649
rect 1316 546 1332 580
rect 1282 508 1332 546
rect 1316 474 1332 508
rect 1282 458 1332 474
rect 1366 580 1432 596
rect 1366 546 1382 580
rect 1416 546 1432 580
rect 1366 502 1432 546
rect 1366 468 1382 502
rect 1416 468 1432 502
rect 1366 424 1432 468
rect 1472 580 1522 649
rect 1506 546 1522 580
rect 1472 508 1522 546
rect 1506 474 1522 508
rect 1472 458 1522 474
rect 1556 580 1622 596
rect 1556 546 1572 580
rect 1606 546 1622 580
rect 1556 502 1622 546
rect 1556 468 1572 502
rect 1606 468 1622 502
rect 1556 424 1622 468
rect 1656 580 1706 649
rect 1656 546 1672 580
rect 1656 508 1706 546
rect 1656 474 1672 508
rect 1656 458 1706 474
rect 1746 580 1812 596
rect 1746 546 1762 580
rect 1796 546 1812 580
rect 1746 502 1812 546
rect 1746 468 1762 502
rect 1796 468 1812 502
rect 1746 424 1812 468
rect 1852 580 1886 649
rect 1852 508 1886 546
rect 1852 458 1886 474
rect 1926 580 1992 596
rect 1926 546 1942 580
rect 1976 546 1992 580
rect 1926 502 1992 546
rect 1926 468 1942 502
rect 1976 468 1992 502
rect 1926 424 1992 468
rect 173 414 743 424
rect 173 398 329 414
rect 123 390 329 398
rect 363 390 743 414
rect 794 390 810 424
rect 844 414 1192 424
rect 844 390 1002 414
rect 363 380 421 390
rect 329 364 421 380
rect 25 320 286 356
rect 25 286 100 320
rect 134 286 168 320
rect 202 286 236 320
rect 270 286 286 320
rect 25 270 286 286
rect 363 236 421 364
rect 457 320 659 356
rect 457 286 473 320
rect 507 286 541 320
rect 575 286 609 320
rect 643 286 659 320
rect 457 270 659 286
rect 693 310 743 390
rect 986 380 1002 390
rect 1036 390 1192 414
rect 1226 390 1382 424
rect 1416 390 1572 424
rect 1606 390 1762 424
rect 1796 390 1942 424
rect 1976 390 1992 424
rect 1036 380 1052 390
rect 986 364 1052 380
rect 793 330 935 356
rect 793 314 1124 330
rect 23 210 73 226
rect 23 176 39 210
rect 23 120 73 176
rect 23 86 39 120
rect 23 17 73 86
rect 109 210 487 236
rect 109 176 125 210
rect 159 202 487 210
rect 159 176 175 202
rect 109 120 175 176
rect 421 169 487 202
rect 109 86 125 120
rect 159 86 175 120
rect 109 70 175 86
rect 209 152 275 168
rect 209 118 225 152
rect 259 118 275 152
rect 209 17 275 118
rect 321 148 387 168
rect 321 114 337 148
rect 371 114 387 148
rect 421 135 437 169
rect 471 135 487 169
rect 421 119 487 135
rect 521 210 627 226
rect 521 176 523 210
rect 557 176 591 210
rect 625 176 627 210
rect 693 200 727 310
rect 793 280 870 314
rect 904 280 938 314
rect 972 280 1006 314
rect 1040 280 1074 314
rect 1108 280 1124 314
rect 793 264 1124 280
rect 1177 320 1607 356
rect 1177 286 1252 320
rect 1286 286 1320 320
rect 1354 286 1388 320
rect 1422 286 1456 320
rect 1490 286 1524 320
rect 1558 286 1607 320
rect 1177 270 1607 286
rect 1657 320 1991 356
rect 1657 286 1673 320
rect 1707 286 1741 320
rect 1775 286 1809 320
rect 1843 286 1877 320
rect 1911 286 1991 320
rect 1657 270 1991 286
rect 521 120 627 176
rect 321 85 387 114
rect 521 86 523 120
rect 557 86 591 120
rect 625 86 627 120
rect 661 174 727 200
rect 661 140 677 174
rect 711 140 727 174
rect 661 119 727 140
rect 761 210 827 226
rect 761 176 777 210
rect 811 176 827 210
rect 761 124 827 176
rect 861 209 1555 226
rect 861 207 1333 209
rect 861 173 877 207
rect 911 173 1049 207
rect 1083 175 1333 207
rect 1367 207 1555 209
rect 1367 175 1505 207
rect 1083 173 1505 175
rect 1539 173 1555 207
rect 861 158 1555 173
rect 1489 154 1555 158
rect 1591 210 1993 236
rect 1625 202 1763 210
rect 761 120 1185 124
rect 521 85 627 86
rect 761 86 777 120
rect 811 86 963 120
rect 997 86 1135 120
rect 1169 86 1185 120
rect 761 85 1185 86
rect 321 51 1185 85
rect 1231 122 1297 124
rect 1231 88 1247 122
rect 1281 120 1297 122
rect 1591 120 1625 176
rect 1797 202 1943 210
rect 1281 88 1419 120
rect 1231 86 1419 88
rect 1453 86 1591 120
rect 1231 70 1625 86
rect 1661 152 1727 168
rect 1661 118 1677 152
rect 1711 118 1727 152
rect 1661 17 1727 118
rect 1763 120 1797 176
rect 1977 176 1993 210
rect 1763 70 1797 86
rect 1833 152 1899 168
rect 1833 118 1849 152
rect 1883 118 1899 152
rect 1833 17 1899 118
rect 1943 120 1993 176
rect 1977 86 1993 120
rect 1943 70 1993 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
flabel pwell s 0 0 2016 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 0 617 2016 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
rlabel comment s 0 0 0 0 4 a41oi_4
flabel metal1 s 0 617 2016 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 2016 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 1183 316 1217 350 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 1279 316 1313 350 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 1375 316 1409 350 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 1471 316 1505 350 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 1567 316 1601 350 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 1663 316 1697 350 0 FreeSans 340 0 0 0 A4
port 4 nsew
flabel corelocali s 1759 316 1793 350 0 FreeSans 340 0 0 0 A4
port 4 nsew
flabel corelocali s 1855 316 1889 350 0 FreeSans 340 0 0 0 A4
port 4 nsew
flabel corelocali s 1951 316 1985 350 0 FreeSans 340 0 0 0 A4
port 4 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 B1
port 5 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 B1
port 5 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 B1
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 2016 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3104364
string GDS_START 3088464
<< end >>
