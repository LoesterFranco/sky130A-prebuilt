magic
tech sky130A
magscale 1 2
timestamp 1604502693
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 79 47 109 177
rect 174 47 204 177
rect 266 47 296 177
rect 431 47 461 177
rect 515 47 545 177
<< pmoshvt >>
rect 79 297 109 497
rect 151 297 181 497
rect 303 297 333 497
rect 431 297 461 497
rect 515 297 545 497
<< ndiff >>
rect 27 93 79 177
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 165 174 177
rect 109 131 119 165
rect 153 131 174 165
rect 109 47 174 131
rect 204 161 266 177
rect 204 127 219 161
rect 253 127 266 161
rect 204 93 266 127
rect 204 59 219 93
rect 253 59 266 93
rect 204 47 266 59
rect 296 93 431 177
rect 296 59 319 93
rect 353 59 387 93
rect 421 59 431 93
rect 296 47 431 59
rect 461 125 515 177
rect 461 91 471 125
rect 505 91 515 125
rect 461 47 515 91
rect 545 161 617 177
rect 545 127 555 161
rect 589 127 617 161
rect 545 93 617 127
rect 545 59 555 93
rect 589 59 617 93
rect 545 47 617 59
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 297 151 497
rect 181 485 303 497
rect 181 383 191 485
rect 293 383 303 485
rect 181 297 303 383
rect 333 297 431 497
rect 461 297 515 497
rect 545 485 601 497
rect 545 451 555 485
rect 589 451 601 485
rect 545 417 601 451
rect 545 383 555 417
rect 589 383 601 417
rect 545 349 601 383
rect 545 315 555 349
rect 589 315 601 349
rect 545 297 601 315
<< ndiffc >>
rect 35 59 69 93
rect 119 131 153 165
rect 219 127 253 161
rect 219 59 253 93
rect 319 59 353 93
rect 387 59 421 93
rect 471 91 505 125
rect 555 127 589 161
rect 555 59 589 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 191 383 293 485
rect 555 451 589 485
rect 555 383 589 417
rect 555 315 589 349
<< poly >>
rect 79 497 109 523
rect 151 497 181 523
rect 303 497 333 523
rect 431 497 461 523
rect 515 497 545 523
rect 79 265 109 297
rect 22 249 109 265
rect 22 215 38 249
rect 72 215 109 249
rect 22 199 109 215
rect 151 265 181 297
rect 303 265 333 297
rect 431 265 461 297
rect 151 249 224 265
rect 151 215 174 249
rect 208 215 224 249
rect 151 213 224 215
rect 158 199 224 213
rect 266 249 333 265
rect 266 215 282 249
rect 316 215 333 249
rect 266 213 333 215
rect 395 249 461 265
rect 395 215 411 249
rect 445 215 461 249
rect 266 199 332 213
rect 395 199 461 215
rect 79 177 109 199
rect 174 177 204 199
rect 266 177 296 199
rect 431 177 461 199
rect 515 265 545 297
rect 515 249 581 265
rect 515 215 531 249
rect 565 215 581 249
rect 515 199 581 215
rect 515 177 545 199
rect 79 21 109 47
rect 174 21 204 47
rect 266 21 296 47
rect 431 21 461 47
rect 515 21 545 47
<< polycont >>
rect 38 215 72 249
rect 174 215 208 249
rect 282 215 316 249
rect 411 215 445 249
rect 531 215 565 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 18 485 72 527
rect 18 451 35 485
rect 69 451 72 485
rect 18 417 72 451
rect 18 383 35 417
rect 69 383 72 417
rect 18 349 72 383
rect 18 315 35 349
rect 69 315 72 349
rect 18 299 72 315
rect 106 485 309 493
rect 106 383 191 485
rect 293 383 309 485
rect 106 357 309 383
rect 18 249 72 265
rect 18 215 38 249
rect 18 199 72 215
rect 18 137 69 199
rect 106 165 140 357
rect 174 249 248 323
rect 208 215 248 249
rect 174 199 248 215
rect 282 249 340 323
rect 316 215 340 249
rect 282 199 340 215
rect 386 249 445 493
rect 539 485 627 527
rect 539 451 555 485
rect 589 451 627 485
rect 539 417 627 451
rect 539 383 555 417
rect 589 383 627 417
rect 539 349 627 383
rect 539 315 555 349
rect 589 315 627 349
rect 539 299 627 315
rect 386 215 411 249
rect 386 199 445 215
rect 515 249 627 265
rect 515 215 531 249
rect 565 215 627 249
rect 515 199 627 215
rect 103 131 119 165
rect 153 131 169 165
rect 203 161 505 165
rect 203 127 219 161
rect 253 131 505 161
rect 253 127 269 131
rect 203 97 269 127
rect 471 125 505 131
rect 18 93 269 97
rect 18 59 35 93
rect 69 59 219 93
rect 253 59 269 93
rect 18 51 269 59
rect 303 93 437 97
rect 303 59 319 93
rect 353 59 387 93
rect 421 59 437 93
rect 471 75 505 91
rect 539 161 627 165
rect 539 127 555 161
rect 589 127 627 161
rect 539 93 627 127
rect 303 17 437 59
rect 539 59 555 93
rect 589 59 627 93
rect 539 17 627 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel corelocali s 398 425 432 459 0 FreeSans 250 0 0 0 A2
port 2 nsew
flabel corelocali s 398 357 432 391 0 FreeSans 250 0 0 0 A2
port 2 nsew
flabel corelocali s 398 289 432 323 0 FreeSans 250 0 0 0 A2
port 2 nsew
flabel corelocali s 214 357 248 391 0 FreeSans 250 0 0 0 Y
port 10 nsew
flabel corelocali s 214 425 248 459 0 FreeSans 250 0 0 0 Y
port 10 nsew
flabel corelocali s 122 357 156 391 0 FreeSans 250 0 0 0 Y
port 10 nsew
flabel corelocali s 122 425 156 459 0 FreeSans 250 0 0 0 Y
port 10 nsew
flabel corelocali s 582 221 616 255 0 FreeSans 250 0 0 0 A1
port 1 nsew
flabel corelocali s 398 221 432 255 0 FreeSans 250 0 0 0 A2
port 2 nsew
flabel corelocali s 306 221 340 255 0 FreeSans 250 0 0 0 A3
port 3 nsew
flabel corelocali s 214 221 248 255 0 FreeSans 250 0 0 0 B2
port 5 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 250 0 0 0 B1
port 4 nsew
flabel corelocali s 30 153 64 187 0 FreeSans 250 0 0 0 B1
port 4 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew
rlabel comment s 0 0 0 0 4 o32ai_1
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 912600
string GDS_START 905924
string path 0.000 0.000 3.220 0.000 
<< end >>
