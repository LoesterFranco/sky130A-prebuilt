magic
tech sky130A
magscale 1 2
timestamp 1604502701
<< nwell >>
rect -38 332 2246 704
<< pwell >>
rect 0 0 2208 49
<< scpmos >>
rect 108 464 138 592
rect 208 464 238 592
rect 292 464 322 592
rect 382 464 412 592
rect 490 464 520 592
rect 632 368 662 592
rect 870 368 900 592
rect 1072 508 1102 592
rect 1172 508 1202 592
rect 1252 508 1282 592
rect 1376 424 1406 592
rect 1517 424 1547 592
rect 1658 508 1688 592
rect 1742 508 1772 592
rect 1891 424 1921 592
rect 2093 368 2123 592
<< nmoslvt >>
rect 92 74 122 158
rect 193 74 223 158
rect 271 74 301 158
rect 420 74 450 158
rect 498 74 528 158
rect 600 74 630 222
rect 798 74 828 222
rect 988 100 1018 184
rect 1124 100 1154 184
rect 1239 100 1269 184
rect 1403 74 1433 184
rect 1490 74 1520 184
rect 1658 100 1688 184
rect 1736 100 1766 184
rect 1905 74 1935 184
rect 2096 78 2126 226
<< ndiff >>
rect 543 158 600 222
rect 35 130 92 158
rect 35 96 47 130
rect 81 96 92 130
rect 35 74 92 96
rect 122 130 193 158
rect 122 96 133 130
rect 167 96 193 130
rect 122 74 193 96
rect 223 74 271 158
rect 301 130 420 158
rect 301 96 346 130
rect 380 96 420 130
rect 301 74 420 96
rect 450 74 498 158
rect 528 142 600 158
rect 528 108 555 142
rect 589 108 600 142
rect 528 74 600 108
rect 630 192 687 222
rect 630 158 641 192
rect 675 158 687 192
rect 630 120 687 158
rect 630 86 641 120
rect 675 86 687 120
rect 630 74 687 86
rect 741 122 798 222
rect 741 88 753 122
rect 787 88 798 122
rect 741 74 798 88
rect 828 210 881 222
rect 828 176 839 210
rect 873 176 881 210
rect 2042 214 2096 226
rect 828 120 881 176
rect 828 86 839 120
rect 873 86 881 120
rect 935 170 988 184
rect 935 136 943 170
rect 977 136 988 170
rect 935 100 988 136
rect 1018 170 1124 184
rect 1018 136 1079 170
rect 1113 136 1124 170
rect 1018 100 1124 136
rect 1154 100 1239 184
rect 1269 100 1403 184
rect 828 74 881 86
rect 1284 88 1403 100
rect 1284 54 1293 88
rect 1327 74 1403 88
rect 1433 154 1490 184
rect 1433 120 1445 154
rect 1479 120 1490 154
rect 1433 74 1490 120
rect 1520 159 1658 184
rect 1520 125 1613 159
rect 1647 125 1658 159
rect 1520 100 1658 125
rect 1688 100 1736 184
rect 1766 146 1905 184
rect 1766 112 1777 146
rect 1811 112 1846 146
rect 1880 112 1905 146
rect 1766 100 1905 112
rect 1520 74 1570 100
rect 1855 74 1905 100
rect 1935 146 1988 184
rect 1935 112 1946 146
rect 1980 112 1988 146
rect 1935 74 1988 112
rect 2042 180 2051 214
rect 2085 180 2096 214
rect 2042 124 2096 180
rect 2042 90 2051 124
rect 2085 90 2096 124
rect 2042 78 2096 90
rect 2126 214 2181 226
rect 2126 180 2137 214
rect 2171 180 2181 214
rect 2126 124 2181 180
rect 2126 90 2137 124
rect 2171 90 2181 124
rect 2126 78 2181 90
rect 1327 54 1339 74
rect 1284 42 1339 54
<< pdiff >>
rect 1300 622 1358 634
rect 1300 592 1312 622
rect 49 580 108 592
rect 49 546 61 580
rect 95 546 108 580
rect 49 510 108 546
rect 49 476 61 510
rect 95 476 108 510
rect 49 464 108 476
rect 138 580 208 592
rect 138 546 161 580
rect 195 546 208 580
rect 138 510 208 546
rect 138 476 161 510
rect 195 476 208 510
rect 138 464 208 476
rect 238 464 292 592
rect 322 580 382 592
rect 322 546 335 580
rect 369 546 382 580
rect 322 512 382 546
rect 322 478 335 512
rect 369 478 382 512
rect 322 464 382 478
rect 412 464 490 592
rect 520 580 632 592
rect 520 546 567 580
rect 601 546 632 580
rect 520 464 632 546
rect 579 368 632 464
rect 662 421 721 592
rect 662 387 675 421
rect 709 387 721 421
rect 662 368 721 387
rect 775 580 870 592
rect 775 546 805 580
rect 839 546 870 580
rect 775 368 870 546
rect 900 421 959 592
rect 1013 578 1072 592
rect 1013 544 1025 578
rect 1059 544 1072 578
rect 1013 508 1072 544
rect 1102 567 1172 592
rect 1102 533 1125 567
rect 1159 533 1172 567
rect 1102 508 1172 533
rect 1202 508 1252 592
rect 1282 588 1312 592
rect 1346 592 1358 622
rect 1346 588 1376 592
rect 1282 508 1376 588
rect 900 387 913 421
rect 947 387 959 421
rect 900 368 959 387
rect 1323 424 1376 508
rect 1406 470 1517 592
rect 1406 436 1422 470
rect 1456 436 1517 470
rect 1406 424 1517 436
rect 1547 580 1658 592
rect 1547 546 1577 580
rect 1611 546 1658 580
rect 1547 508 1658 546
rect 1688 508 1742 592
rect 1772 580 1891 592
rect 1772 546 1809 580
rect 1843 546 1891 580
rect 1772 508 1891 546
rect 1547 470 1623 508
rect 1547 436 1577 470
rect 1611 436 1623 470
rect 1547 424 1623 436
rect 1838 424 1891 508
rect 1921 580 1980 592
rect 1921 546 1934 580
rect 1968 546 1980 580
rect 1921 470 1980 546
rect 1921 436 1934 470
rect 1968 436 1980 470
rect 1921 424 1980 436
rect 2034 580 2093 592
rect 2034 546 2046 580
rect 2080 546 2093 580
rect 2034 497 2093 546
rect 2034 463 2046 497
rect 2080 463 2093 497
rect 2034 414 2093 463
rect 2034 380 2046 414
rect 2080 380 2093 414
rect 2034 368 2093 380
rect 2123 580 2181 592
rect 2123 546 2136 580
rect 2170 546 2181 580
rect 2123 497 2181 546
rect 2123 463 2136 497
rect 2170 463 2181 497
rect 2123 414 2181 463
rect 2123 380 2136 414
rect 2170 380 2181 414
rect 2123 368 2181 380
<< ndiffc >>
rect 47 96 81 130
rect 133 96 167 130
rect 346 96 380 130
rect 555 108 589 142
rect 641 158 675 192
rect 641 86 675 120
rect 753 88 787 122
rect 839 176 873 210
rect 839 86 873 120
rect 943 136 977 170
rect 1079 136 1113 170
rect 1293 54 1327 88
rect 1445 120 1479 154
rect 1613 125 1647 159
rect 1777 112 1811 146
rect 1846 112 1880 146
rect 1946 112 1980 146
rect 2051 180 2085 214
rect 2051 90 2085 124
rect 2137 180 2171 214
rect 2137 90 2171 124
<< pdiffc >>
rect 61 546 95 580
rect 61 476 95 510
rect 161 546 195 580
rect 161 476 195 510
rect 335 546 369 580
rect 335 478 369 512
rect 567 546 601 580
rect 675 387 709 421
rect 805 546 839 580
rect 1025 544 1059 578
rect 1125 533 1159 567
rect 1312 588 1346 622
rect 913 387 947 421
rect 1422 436 1456 470
rect 1577 546 1611 580
rect 1809 546 1843 580
rect 1577 436 1611 470
rect 1934 546 1968 580
rect 1934 436 1968 470
rect 2046 546 2080 580
rect 2046 463 2080 497
rect 2046 380 2080 414
rect 2136 546 2170 580
rect 2136 463 2170 497
rect 2136 380 2170 414
<< poly >>
rect 108 592 138 618
rect 208 592 238 618
rect 292 592 322 618
rect 382 592 412 618
rect 490 592 520 618
rect 632 592 662 618
rect 870 592 900 618
rect 1072 592 1102 618
rect 1172 592 1202 618
rect 1252 592 1282 618
rect 108 449 138 464
rect 208 449 238 464
rect 292 449 322 464
rect 382 449 412 464
rect 490 449 520 464
rect 21 419 241 449
rect 21 257 51 419
rect 99 355 165 371
rect 289 357 325 449
rect 379 428 415 449
rect 487 428 523 449
rect 373 412 439 428
rect 373 378 389 412
rect 423 378 439 412
rect 99 321 115 355
rect 149 335 165 355
rect 265 341 331 357
rect 149 321 223 335
rect 99 305 223 321
rect 21 241 151 257
rect 21 227 101 241
rect 85 207 101 227
rect 135 207 151 241
rect 85 191 151 207
rect 92 158 122 191
rect 193 158 223 305
rect 265 307 281 341
rect 315 307 331 341
rect 265 291 331 307
rect 373 344 439 378
rect 373 310 389 344
rect 423 310 439 344
rect 373 294 439 310
rect 481 412 547 428
rect 481 378 497 412
rect 531 378 547 412
rect 481 344 547 378
rect 1376 592 1406 618
rect 1517 592 1547 618
rect 1658 592 1688 618
rect 1742 592 1772 618
rect 1891 592 1921 618
rect 2093 592 2123 618
rect 1072 493 1102 508
rect 1172 493 1202 508
rect 1252 493 1282 508
rect 1069 476 1105 493
rect 991 460 1105 476
rect 991 426 1007 460
rect 1041 446 1105 460
rect 1041 426 1057 446
rect 1169 440 1205 493
rect 1249 463 1285 493
rect 991 410 1057 426
rect 1147 424 1213 440
rect 1147 390 1163 424
rect 1197 390 1213 424
rect 1147 368 1213 390
rect 632 353 662 368
rect 870 353 900 368
rect 481 310 497 344
rect 531 310 547 344
rect 481 294 547 310
rect 629 310 665 353
rect 867 326 903 353
rect 988 338 1213 368
rect 988 326 1018 338
rect 758 310 1018 326
rect 629 294 716 310
rect 271 158 301 291
rect 384 230 450 246
rect 384 196 400 230
rect 434 196 450 230
rect 384 180 450 196
rect 420 158 450 180
rect 498 158 528 294
rect 629 274 666 294
rect 600 260 666 274
rect 700 260 716 294
rect 758 276 774 310
rect 808 296 1018 310
rect 808 276 828 296
rect 758 260 828 276
rect 600 244 716 260
rect 600 222 630 244
rect 798 222 828 260
rect 988 184 1018 296
rect 1255 272 1285 463
rect 1658 493 1688 508
rect 1742 493 1772 508
rect 1376 409 1406 424
rect 1517 409 1547 424
rect 1655 415 1691 493
rect 1739 463 1805 493
rect 1373 386 1409 409
rect 1514 386 1550 409
rect 1661 399 1727 415
rect 1329 370 1433 386
rect 1329 336 1345 370
rect 1379 336 1433 370
rect 1329 320 1433 336
rect 1514 370 1580 386
rect 1514 336 1530 370
rect 1564 350 1580 370
rect 1661 365 1677 399
rect 1711 365 1727 399
rect 1564 336 1619 350
rect 1514 320 1619 336
rect 1124 256 1197 272
rect 1124 222 1147 256
rect 1181 222 1197 256
rect 1124 206 1197 222
rect 1239 256 1305 272
rect 1239 222 1255 256
rect 1289 222 1305 256
rect 1239 206 1305 222
rect 1124 184 1154 206
rect 1239 184 1269 206
rect 1403 184 1433 320
rect 1481 256 1547 272
rect 1481 222 1497 256
rect 1531 222 1547 256
rect 1481 206 1547 222
rect 1589 233 1619 320
rect 1661 331 1727 365
rect 1661 297 1677 331
rect 1711 297 1727 331
rect 1661 281 1727 297
rect 1775 272 1805 463
rect 1891 409 1921 424
rect 1888 386 1924 409
rect 1853 370 1935 386
rect 1853 336 1869 370
rect 1903 336 1935 370
rect 2093 353 2123 368
rect 1853 320 1935 336
rect 2090 330 2126 353
rect 1775 256 1863 272
rect 1775 233 1813 256
rect 1490 184 1520 206
rect 1589 203 1688 233
rect 1658 184 1688 203
rect 1736 222 1813 233
rect 1847 222 1863 256
rect 1736 203 1863 222
rect 1736 184 1766 203
rect 1905 184 1935 320
rect 1983 314 2126 330
rect 1983 280 1999 314
rect 2033 280 2126 314
rect 1983 264 2126 280
rect 2096 226 2126 264
rect 988 74 1018 100
rect 1124 74 1154 100
rect 1239 74 1269 100
rect 92 48 122 74
rect 193 48 223 74
rect 271 48 301 74
rect 420 48 450 74
rect 498 48 528 74
rect 600 48 630 74
rect 798 48 828 74
rect 1658 74 1688 100
rect 1736 74 1766 100
rect 1403 48 1433 74
rect 1490 48 1520 74
rect 1905 48 1935 74
rect 2096 52 2126 78
<< polycont >>
rect 389 378 423 412
rect 115 321 149 355
rect 101 207 135 241
rect 281 307 315 341
rect 389 310 423 344
rect 497 378 531 412
rect 1007 426 1041 460
rect 1163 390 1197 424
rect 497 310 531 344
rect 400 196 434 230
rect 666 260 700 294
rect 774 276 808 310
rect 1345 336 1379 370
rect 1530 336 1564 370
rect 1677 365 1711 399
rect 1147 222 1181 256
rect 1255 222 1289 256
rect 1497 222 1531 256
rect 1677 297 1711 331
rect 1869 336 1903 370
rect 1813 222 1847 256
rect 1999 280 2033 314
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 17 580 111 596
rect 17 546 61 580
rect 95 546 111 580
rect 17 510 111 546
rect 17 476 61 510
rect 95 476 111 510
rect 17 425 111 476
rect 145 580 211 649
rect 145 546 161 580
rect 195 546 211 580
rect 145 510 211 546
rect 145 476 161 510
rect 195 476 211 510
rect 145 460 211 476
rect 319 580 385 596
rect 319 546 335 580
rect 369 546 385 580
rect 319 512 385 546
rect 534 580 635 649
rect 534 546 567 580
rect 601 546 635 580
rect 771 580 873 649
rect 1296 622 1362 649
rect 771 546 805 580
rect 839 546 873 580
rect 907 578 1075 596
rect 534 530 635 546
rect 907 544 1025 578
rect 1059 544 1075 578
rect 907 542 1075 544
rect 1109 567 1175 596
rect 1296 588 1312 622
rect 1346 588 1362 622
rect 1296 572 1362 588
rect 1577 580 1627 596
rect 907 512 941 542
rect 319 478 335 512
rect 369 496 385 512
rect 669 496 941 512
rect 1109 533 1125 567
rect 1159 533 1175 567
rect 1611 546 1627 580
rect 1109 508 1175 533
rect 369 478 941 496
rect 319 462 879 478
rect 373 425 439 428
rect 17 412 439 425
rect 17 391 389 412
rect 17 355 165 391
rect 373 378 389 391
rect 423 378 439 412
rect 17 321 115 355
rect 149 321 165 355
rect 17 305 165 321
rect 217 341 331 357
rect 217 307 281 341
rect 315 307 331 341
rect 17 157 51 305
rect 217 291 331 307
rect 373 344 439 378
rect 373 310 389 344
rect 423 310 439 344
rect 373 294 439 310
rect 481 412 548 428
rect 481 378 497 412
rect 531 378 548 412
rect 481 344 548 378
rect 481 310 497 344
rect 531 310 548 344
rect 481 294 548 310
rect 582 260 616 462
rect 659 421 811 428
rect 659 387 675 421
rect 709 387 811 421
rect 659 364 811 387
rect 771 310 811 364
rect 85 241 450 257
rect 85 207 101 241
rect 135 230 450 241
rect 135 207 400 230
rect 85 196 400 207
rect 434 196 450 230
rect 85 191 450 196
rect 217 180 450 191
rect 484 226 616 260
rect 650 294 737 310
rect 650 260 666 294
rect 700 260 737 294
rect 650 236 737 260
rect 771 276 774 310
rect 808 276 811 310
rect 845 330 879 462
rect 991 460 1045 476
rect 991 444 1007 460
rect 913 426 1007 444
rect 1041 426 1045 460
rect 913 421 1045 426
rect 947 410 1045 421
rect 947 387 963 410
rect 913 364 963 387
rect 845 296 957 330
rect 771 260 811 276
rect 217 162 263 180
rect 17 130 81 157
rect 17 96 47 130
rect 17 70 81 96
rect 117 130 183 157
rect 484 146 518 226
rect 771 192 805 260
rect 625 158 641 192
rect 675 158 805 192
rect 839 210 889 226
rect 873 176 889 210
rect 117 96 133 130
rect 167 96 183 130
rect 117 17 183 96
rect 297 130 518 146
rect 297 96 346 130
rect 380 96 518 130
rect 297 80 518 96
rect 555 142 589 158
rect 555 17 589 108
rect 625 120 691 158
rect 625 86 641 120
rect 675 86 691 120
rect 625 70 691 86
rect 737 122 803 124
rect 737 88 753 122
rect 787 88 803 122
rect 737 17 803 88
rect 839 120 889 176
rect 873 86 889 120
rect 923 188 957 296
rect 923 170 977 188
rect 923 136 943 170
rect 923 119 977 136
rect 839 85 889 86
rect 1011 85 1045 410
rect 1079 474 1175 508
rect 1209 504 1543 538
rect 1079 340 1113 474
rect 1209 440 1243 504
rect 1147 424 1243 440
rect 1147 390 1163 424
rect 1197 390 1243 424
rect 1403 436 1422 470
rect 1456 436 1475 470
rect 1403 420 1475 436
rect 1147 374 1243 390
rect 1329 370 1395 386
rect 1329 340 1345 370
rect 1079 336 1345 340
rect 1379 336 1395 370
rect 1079 306 1395 336
rect 1079 170 1113 306
rect 1429 272 1463 420
rect 1509 386 1543 504
rect 1577 483 1627 546
rect 1769 580 1884 649
rect 1769 546 1809 580
rect 1843 546 1884 580
rect 1769 530 1884 546
rect 1918 580 1987 596
rect 1918 546 1934 580
rect 1968 546 1987 580
rect 1577 470 1779 483
rect 1611 449 1779 470
rect 1611 436 1627 449
rect 1577 420 1627 436
rect 1661 399 1711 415
rect 1509 370 1580 386
rect 1509 336 1530 370
rect 1564 336 1580 370
rect 1509 320 1580 336
rect 1661 365 1677 399
rect 1661 331 1711 365
rect 1661 298 1677 331
rect 1614 297 1677 298
rect 1614 272 1711 297
rect 1079 119 1113 136
rect 1147 256 1197 272
rect 1181 222 1197 256
rect 1147 172 1197 222
rect 1239 256 1463 272
rect 1239 222 1255 256
rect 1289 222 1463 256
rect 1239 206 1463 222
rect 1497 264 1711 272
rect 1745 386 1779 449
rect 1918 470 1987 546
rect 1918 436 1934 470
rect 1968 436 1987 470
rect 1918 420 1987 436
rect 1745 370 1919 386
rect 1745 336 1869 370
rect 1903 336 1919 370
rect 1745 320 1919 336
rect 1953 330 1987 420
rect 2030 580 2080 649
rect 2030 546 2046 580
rect 2030 497 2080 546
rect 2030 463 2046 497
rect 2030 414 2080 463
rect 2030 380 2046 414
rect 2030 364 2080 380
rect 2120 580 2187 596
rect 2120 546 2136 580
rect 2170 546 2187 580
rect 2120 497 2187 546
rect 2120 463 2136 497
rect 2170 463 2187 497
rect 2120 414 2187 463
rect 2120 380 2136 414
rect 2170 380 2187 414
rect 1497 256 1648 264
rect 1531 238 1648 256
rect 1531 222 1563 238
rect 1745 230 1779 320
rect 1953 314 2049 330
rect 1953 280 1999 314
rect 2033 280 2049 314
rect 1953 272 2049 280
rect 1497 206 1563 222
rect 1429 172 1463 206
rect 1147 138 1395 172
rect 1147 85 1181 138
rect 839 51 1181 85
rect 1277 88 1327 104
rect 1277 54 1293 88
rect 1277 17 1327 54
rect 1361 85 1395 138
rect 1429 154 1495 172
rect 1429 120 1445 154
rect 1479 120 1495 154
rect 1429 119 1495 120
rect 1529 85 1563 206
rect 1682 196 1779 230
rect 1813 264 2049 272
rect 1813 256 1996 264
rect 1847 222 1996 256
rect 1813 206 1996 222
rect 1682 188 1716 196
rect 1597 159 1716 188
rect 1597 125 1613 159
rect 1647 154 1716 159
rect 1647 125 1663 154
rect 1597 96 1663 125
rect 1761 146 1896 162
rect 1761 112 1777 146
rect 1811 112 1846 146
rect 1880 112 1896 146
rect 1361 51 1563 85
rect 1761 17 1896 112
rect 1930 146 1996 206
rect 1930 112 1946 146
rect 1980 112 1996 146
rect 1930 70 1996 112
rect 2035 214 2085 230
rect 2035 180 2051 214
rect 2035 124 2085 180
rect 2035 90 2051 124
rect 2035 17 2085 90
rect 2120 214 2187 380
rect 2120 180 2137 214
rect 2171 180 2187 214
rect 2120 124 2187 180
rect 2120 90 2137 124
rect 2171 90 2187 124
rect 2120 74 2187 90
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
<< metal1 >>
rect 0 683 2208 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 0 617 2208 649
rect 0 17 2208 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
rect 0 -49 2208 -17
<< labels >>
rlabel comment s 0 0 0 0 4 sdfxtp_1
flabel comment s 980 313 980 313 0 FreeSans 200 0 0 0 no_jumper_check
flabel pwell s 0 0 2208 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 2208 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 2208 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 2208 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 223 168 257 202 0 FreeSans 340 0 0 0 SCE
port 4 nsew
flabel corelocali s 2143 94 2177 128 0 FreeSans 340 0 0 0 Q
port 9 nsew
flabel corelocali s 2143 168 2177 202 0 FreeSans 340 0 0 0 Q
port 9 nsew
flabel corelocali s 2143 242 2177 276 0 FreeSans 340 0 0 0 Q
port 9 nsew
flabel corelocali s 2143 316 2177 350 0 FreeSans 340 0 0 0 Q
port 9 nsew
flabel corelocali s 2143 390 2177 424 0 FreeSans 340 0 0 0 Q
port 9 nsew
flabel corelocali s 2143 464 2177 498 0 FreeSans 340 0 0 0 Q
port 9 nsew
flabel corelocali s 2143 538 2177 572 0 FreeSans 340 0 0 0 Q
port 9 nsew
flabel corelocali s 703 242 737 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 SCD
port 3 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 D
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 2208 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 297098
string GDS_START 280448
<< end >>
