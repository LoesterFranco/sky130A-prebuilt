magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 2300 561
rect 106 427 172 527
rect 28 195 98 325
rect 293 397 346 493
rect 297 214 346 397
rect 464 408 498 527
rect 573 357 624 493
rect 860 455 926 527
rect 547 271 624 357
rect 103 17 169 93
rect 375 17 441 112
rect 479 17 545 165
rect 804 142 879 340
rect 1282 471 1348 527
rect 1475 435 1549 527
rect 1872 439 1922 527
rect 804 57 855 142
rect 889 17 955 108
rect 1301 153 1407 209
rect 1383 17 1449 109
rect 2024 451 2090 527
rect 2144 299 2194 527
rect 2228 292 2280 465
rect 2230 289 2280 292
rect 1905 213 2023 255
rect 1817 17 1851 105
rect 1965 127 2023 213
rect 2238 159 2280 289
rect 2144 17 2178 109
rect 2228 53 2280 159
rect 0 -17 2300 17
<< obsli1 >>
rect 18 393 69 493
rect 18 391 173 393
rect 18 359 135 391
rect 132 357 135 359
rect 169 357 173 391
rect 132 265 173 357
rect 207 380 241 493
rect 380 411 430 480
rect 207 346 263 380
rect 132 199 195 265
rect 229 255 263 346
rect 132 161 167 199
rect 19 127 167 161
rect 229 135 263 221
rect 396 291 430 411
rect 692 421 726 493
rect 981 437 1055 487
rect 981 421 1015 437
rect 1094 427 1167 493
rect 396 252 494 291
rect 658 387 1015 421
rect 411 237 494 252
rect 658 237 692 387
rect 411 199 617 237
rect 411 180 445 199
rect 19 69 69 127
rect 203 69 263 135
rect 307 146 445 180
rect 307 79 341 146
rect 583 85 617 199
rect 651 203 692 237
rect 651 135 685 203
rect 736 85 770 337
rect 583 51 770 85
rect 913 179 947 387
rect 1049 357 1065 391
rect 1049 315 1099 357
rect 981 255 1015 279
rect 981 213 1015 221
rect 1065 207 1099 315
rect 1133 277 1167 427
rect 1201 421 1235 475
rect 1399 421 1433 475
rect 1201 387 1433 421
rect 1594 401 1628 493
rect 1664 425 1838 493
rect 1803 423 1838 425
rect 1803 407 1842 423
rect 1491 367 1628 401
rect 1491 353 1543 367
rect 1257 319 1543 353
rect 1662 357 1689 391
rect 1723 387 1768 391
rect 1723 357 1774 387
rect 1662 333 1774 357
rect 1133 243 1475 277
rect 913 143 1029 179
rect 995 101 1029 143
rect 1065 141 1195 207
rect 995 67 1063 101
rect 1233 95 1267 243
rect 1441 201 1475 243
rect 1509 167 1543 319
rect 1097 61 1267 95
rect 1491 89 1543 167
rect 1577 331 1774 333
rect 1808 349 1842 407
rect 1956 417 1990 475
rect 1956 383 2109 417
rect 1577 299 1704 331
rect 1808 315 2041 349
rect 1577 141 1619 299
rect 1808 297 1842 315
rect 1681 255 1715 265
rect 1681 184 1715 221
rect 1749 263 1842 297
rect 2075 265 2109 383
rect 1749 107 1783 263
rect 2075 259 2204 265
rect 1825 173 1859 229
rect 1825 139 1931 173
rect 1491 55 1557 89
rect 1601 51 1783 107
rect 1897 93 1931 139
rect 2069 199 2204 259
rect 2069 93 2103 199
rect 1897 59 2103 93
<< obsli1c >>
rect 135 357 169 391
rect 229 221 263 255
rect 1065 357 1099 391
rect 981 221 1015 255
rect 1689 357 1723 391
rect 1681 221 1715 255
<< metal1 >>
rect 0 496 2300 592
rect 1926 193 1984 261
rect 1289 184 1419 193
rect 1926 184 2035 193
rect 1289 156 2035 184
rect 1289 147 1419 156
rect 1977 147 2035 156
rect 0 -48 2300 48
<< obsm1 >>
rect 123 391 183 397
rect 123 357 135 391
rect 169 388 183 391
rect 1053 391 1111 397
rect 1053 388 1065 391
rect 169 360 1065 388
rect 169 357 183 360
rect 123 351 183 357
rect 1053 357 1065 360
rect 1099 388 1111 391
rect 1677 391 1735 397
rect 1677 388 1689 391
rect 1099 360 1689 388
rect 1099 357 1111 360
rect 1053 351 1111 357
rect 1677 357 1689 360
rect 1723 357 1735 391
rect 1677 351 1735 357
rect 217 255 275 261
rect 217 221 229 255
rect 263 252 275 255
rect 969 255 1027 261
rect 969 252 981 255
rect 263 224 981 252
rect 263 221 275 224
rect 217 215 275 221
rect 969 221 981 224
rect 1015 252 1027 255
rect 1669 255 1727 261
rect 1669 252 1681 255
rect 1015 224 1681 252
rect 1015 221 1027 224
rect 969 215 1027 221
rect 1669 221 1681 224
rect 1715 221 1727 255
rect 1669 215 1727 221
<< labels >>
rlabel locali s 573 357 624 493 6 D
port 1 nsew signal input
rlabel locali s 547 271 624 357 6 D
port 1 nsew signal input
rlabel locali s 2238 159 2280 289 6 Q
port 2 nsew signal output
rlabel locali s 2230 289 2280 292 6 Q
port 2 nsew signal output
rlabel locali s 2228 292 2280 465 6 Q
port 2 nsew signal output
rlabel locali s 2228 53 2280 159 6 Q
port 2 nsew signal output
rlabel locali s 1301 153 1407 209 6 RESET_B
port 3 nsew signal input
rlabel locali s 1965 127 2023 213 6 RESET_B
port 3 nsew signal input
rlabel locali s 1905 213 2023 255 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 1977 147 2035 156 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 1926 193 1984 261 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 1926 184 2035 193 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 1289 184 1419 193 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 1289 156 2035 184 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 1289 147 1419 156 6 RESET_B
port 3 nsew signal input
rlabel locali s 804 142 879 340 6 SCD
port 4 nsew signal input
rlabel locali s 804 57 855 142 6 SCD
port 4 nsew signal input
rlabel locali s 297 214 346 397 6 SCE
port 5 nsew signal input
rlabel locali s 293 397 346 493 6 SCE
port 5 nsew signal input
rlabel locali s 28 195 98 325 6 CLK_N
port 6 nsew clock input
rlabel locali s 2144 17 2178 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1817 17 1851 105 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1383 17 1449 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 889 17 955 108 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 479 17 545 165 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 375 17 441 112 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 103 17 169 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 2300 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 2300 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 2144 299 2194 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 2024 451 2090 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1872 439 1922 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1475 435 1549 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1282 471 1348 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 860 455 926 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 464 408 498 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 106 427 172 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 2300 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 2300 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2300 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 176854
string GDS_START 158022
<< end >>
