magic
tech sky130A
magscale 1 2
timestamp 1604502729
<< locali >>
rect 17 364 91 596
rect 17 226 51 364
rect 193 270 263 356
rect 301 260 367 356
rect 409 270 475 356
rect 509 270 583 356
rect 17 70 89 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 125 458 218 649
rect 439 424 505 576
rect 547 458 610 649
rect 125 390 651 424
rect 125 330 159 390
rect 85 264 159 330
rect 617 226 651 390
rect 123 17 189 226
rect 225 192 549 226
rect 225 90 292 192
rect 353 17 426 156
rect 483 90 549 192
rect 583 90 651 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel locali s 193 270 263 356 6 A1
port 1 nsew signal input
rlabel locali s 301 260 367 356 6 A2
port 2 nsew signal input
rlabel locali s 409 270 475 356 6 A3
port 3 nsew signal input
rlabel locali s 509 270 583 356 6 B1
port 4 nsew signal input
rlabel locali s 17 364 91 596 6 X
port 5 nsew signal output
rlabel locali s 17 226 51 364 6 X
port 5 nsew signal output
rlabel locali s 17 70 89 226 6 X
port 5 nsew signal output
rlabel metal1 s 0 -49 672 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 672 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1369902
string GDS_START 1363536
<< end >>
