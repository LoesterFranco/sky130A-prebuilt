magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 736 561
rect 17 433 85 485
rect 119 435 169 527
rect 17 112 69 433
rect 383 435 433 527
rect 569 435 619 527
rect 201 215 267 327
rect 307 265 367 324
rect 307 199 383 265
rect 17 60 85 112
rect 119 17 185 113
rect 445 120 489 265
rect 541 199 617 325
rect 663 199 714 325
rect 340 83 530 120
rect 576 79 617 199
rect 651 17 719 162
rect 0 -17 736 17
<< obsli1 >>
rect 207 399 273 485
rect 103 365 273 399
rect 307 393 341 493
rect 475 393 509 493
rect 667 393 701 493
rect 103 181 137 365
rect 307 359 701 393
rect 103 162 267 181
rect 103 147 306 162
rect 223 60 306 147
<< metal1 >>
rect 0 496 736 592
rect 0 -48 736 48
<< labels >>
rlabel locali s 307 265 367 324 6 A1
port 1 nsew signal input
rlabel locali s 307 199 383 265 6 A1
port 1 nsew signal input
rlabel locali s 445 120 489 265 6 A2
port 2 nsew signal input
rlabel locali s 340 83 530 120 6 A2
port 2 nsew signal input
rlabel locali s 576 79 617 199 6 A3
port 3 nsew signal input
rlabel locali s 541 199 617 325 6 A3
port 3 nsew signal input
rlabel locali s 663 199 714 325 6 A4
port 4 nsew signal input
rlabel locali s 201 215 267 327 6 B1
port 5 nsew signal input
rlabel locali s 17 433 85 485 6 X
port 6 nsew signal output
rlabel locali s 17 112 69 433 6 X
port 6 nsew signal output
rlabel locali s 17 60 85 112 6 X
port 6 nsew signal output
rlabel locali s 651 17 719 162 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 119 17 185 113 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 736 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 736 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 569 435 619 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 383 435 433 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 119 435 169 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 736 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 736 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3682810
string GDS_START 3674928
<< end >>
