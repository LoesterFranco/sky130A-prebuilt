magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 1785 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 89 47 119 177
rect 183 47 213 177
rect 277 47 307 177
rect 371 47 401 177
rect 455 47 485 177
rect 549 47 579 177
rect 643 47 673 177
rect 747 47 777 177
rect 945 47 975 177
rect 1039 47 1069 177
rect 1133 47 1163 177
rect 1227 47 1257 177
rect 1323 47 1353 177
rect 1417 47 1447 177
rect 1511 47 1541 177
rect 1605 47 1635 177
<< pmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 457 297 493 497
rect 551 297 587 497
rect 645 297 681 497
rect 739 297 775 497
rect 937 297 973 497
rect 1031 297 1067 497
rect 1125 297 1161 497
rect 1219 297 1255 497
rect 1325 297 1361 497
rect 1419 297 1455 497
rect 1513 297 1549 497
rect 1607 297 1643 497
<< ndiff >>
rect 27 142 89 177
rect 27 108 35 142
rect 69 108 89 142
rect 27 47 89 108
rect 119 97 183 177
rect 119 63 129 97
rect 163 63 183 97
rect 119 47 183 63
rect 213 142 277 177
rect 213 108 223 142
rect 257 108 277 142
rect 213 47 277 108
rect 307 97 371 177
rect 307 63 317 97
rect 351 63 371 97
rect 307 47 371 63
rect 401 142 455 177
rect 401 108 411 142
rect 445 108 455 142
rect 401 47 455 108
rect 485 165 549 177
rect 485 131 505 165
rect 539 131 549 165
rect 485 47 549 131
rect 579 97 643 177
rect 579 63 599 97
rect 633 63 643 97
rect 579 47 643 63
rect 673 165 747 177
rect 673 131 693 165
rect 727 131 747 165
rect 673 47 747 131
rect 777 97 829 177
rect 777 63 787 97
rect 821 63 829 97
rect 777 47 829 63
rect 883 97 945 177
rect 883 63 891 97
rect 925 63 945 97
rect 883 47 945 63
rect 975 165 1039 177
rect 975 131 985 165
rect 1019 131 1039 165
rect 975 47 1039 131
rect 1069 97 1133 177
rect 1069 63 1079 97
rect 1113 63 1133 97
rect 1069 47 1133 63
rect 1163 165 1227 177
rect 1163 131 1173 165
rect 1207 131 1227 165
rect 1163 47 1227 131
rect 1257 97 1323 177
rect 1257 63 1274 97
rect 1308 63 1323 97
rect 1257 47 1323 63
rect 1353 165 1417 177
rect 1353 131 1373 165
rect 1407 131 1417 165
rect 1353 47 1417 131
rect 1447 97 1511 177
rect 1447 63 1467 97
rect 1501 63 1511 97
rect 1447 47 1511 63
rect 1541 165 1605 177
rect 1541 131 1561 165
rect 1595 131 1605 165
rect 1541 47 1605 131
rect 1635 165 1697 177
rect 1635 131 1655 165
rect 1689 131 1697 165
rect 1635 97 1697 131
rect 1635 63 1655 97
rect 1689 63 1697 97
rect 1635 47 1697 63
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 485 175 497
rect 117 451 129 485
rect 163 451 175 485
rect 117 417 175 451
rect 117 383 129 417
rect 163 383 175 417
rect 117 349 175 383
rect 117 315 129 349
rect 163 315 175 349
rect 117 297 175 315
rect 211 485 269 497
rect 211 451 223 485
rect 257 451 269 485
rect 211 417 269 451
rect 211 383 223 417
rect 257 383 269 417
rect 211 297 269 383
rect 305 485 363 497
rect 305 451 317 485
rect 351 451 363 485
rect 305 417 363 451
rect 305 383 317 417
rect 351 383 363 417
rect 305 349 363 383
rect 305 315 317 349
rect 351 315 363 349
rect 305 297 363 315
rect 399 485 457 497
rect 399 451 411 485
rect 445 451 457 485
rect 399 417 457 451
rect 399 383 411 417
rect 445 383 457 417
rect 399 297 457 383
rect 493 485 551 497
rect 493 451 505 485
rect 539 451 551 485
rect 493 417 551 451
rect 493 383 505 417
rect 539 383 551 417
rect 493 349 551 383
rect 493 315 505 349
rect 539 315 551 349
rect 493 297 551 315
rect 587 485 645 497
rect 587 451 599 485
rect 633 451 645 485
rect 587 417 645 451
rect 587 383 599 417
rect 633 383 645 417
rect 587 297 645 383
rect 681 485 739 497
rect 681 451 693 485
rect 727 451 739 485
rect 681 417 739 451
rect 681 383 693 417
rect 727 383 739 417
rect 681 349 739 383
rect 681 315 693 349
rect 727 315 739 349
rect 681 297 739 315
rect 775 485 937 497
rect 775 451 787 485
rect 821 451 891 485
rect 925 451 937 485
rect 775 417 937 451
rect 775 383 787 417
rect 821 383 891 417
rect 925 383 937 417
rect 775 297 937 383
rect 973 485 1031 497
rect 973 451 985 485
rect 1019 451 1031 485
rect 973 417 1031 451
rect 973 383 985 417
rect 1019 383 1031 417
rect 973 349 1031 383
rect 973 315 985 349
rect 1019 315 1031 349
rect 973 297 1031 315
rect 1067 485 1125 497
rect 1067 451 1079 485
rect 1113 451 1125 485
rect 1067 417 1125 451
rect 1067 383 1079 417
rect 1113 383 1125 417
rect 1067 297 1125 383
rect 1161 485 1219 497
rect 1161 451 1173 485
rect 1207 451 1219 485
rect 1161 417 1219 451
rect 1161 383 1173 417
rect 1207 383 1219 417
rect 1161 349 1219 383
rect 1161 315 1173 349
rect 1207 315 1219 349
rect 1161 297 1219 315
rect 1255 485 1325 497
rect 1255 451 1274 485
rect 1308 451 1325 485
rect 1255 417 1325 451
rect 1255 383 1274 417
rect 1308 383 1325 417
rect 1255 297 1325 383
rect 1361 485 1419 497
rect 1361 451 1373 485
rect 1407 451 1419 485
rect 1361 417 1419 451
rect 1361 383 1373 417
rect 1407 383 1419 417
rect 1361 349 1419 383
rect 1361 315 1373 349
rect 1407 315 1419 349
rect 1361 297 1419 315
rect 1455 485 1513 497
rect 1455 451 1467 485
rect 1501 451 1513 485
rect 1455 417 1513 451
rect 1455 383 1467 417
rect 1501 383 1513 417
rect 1455 297 1513 383
rect 1549 485 1607 497
rect 1549 451 1561 485
rect 1595 451 1607 485
rect 1549 417 1607 451
rect 1549 383 1561 417
rect 1595 383 1607 417
rect 1549 349 1607 383
rect 1549 315 1561 349
rect 1595 315 1607 349
rect 1549 297 1607 315
rect 1643 485 1697 497
rect 1643 451 1655 485
rect 1689 451 1697 485
rect 1643 417 1697 451
rect 1643 383 1655 417
rect 1689 383 1697 417
rect 1643 349 1697 383
rect 1643 315 1655 349
rect 1689 315 1697 349
rect 1643 297 1697 315
<< ndiffc >>
rect 35 108 69 142
rect 129 63 163 97
rect 223 108 257 142
rect 317 63 351 97
rect 411 108 445 142
rect 505 131 539 165
rect 599 63 633 97
rect 693 131 727 165
rect 787 63 821 97
rect 891 63 925 97
rect 985 131 1019 165
rect 1079 63 1113 97
rect 1173 131 1207 165
rect 1274 63 1308 97
rect 1373 131 1407 165
rect 1467 63 1501 97
rect 1561 131 1595 165
rect 1655 131 1689 165
rect 1655 63 1689 97
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 451 163 485
rect 129 383 163 417
rect 129 315 163 349
rect 223 451 257 485
rect 223 383 257 417
rect 317 451 351 485
rect 317 383 351 417
rect 317 315 351 349
rect 411 451 445 485
rect 411 383 445 417
rect 505 451 539 485
rect 505 383 539 417
rect 505 315 539 349
rect 599 451 633 485
rect 599 383 633 417
rect 693 451 727 485
rect 693 383 727 417
rect 693 315 727 349
rect 787 451 821 485
rect 891 451 925 485
rect 787 383 821 417
rect 891 383 925 417
rect 985 451 1019 485
rect 985 383 1019 417
rect 985 315 1019 349
rect 1079 451 1113 485
rect 1079 383 1113 417
rect 1173 451 1207 485
rect 1173 383 1207 417
rect 1173 315 1207 349
rect 1274 451 1308 485
rect 1274 383 1308 417
rect 1373 451 1407 485
rect 1373 383 1407 417
rect 1373 315 1407 349
rect 1467 451 1501 485
rect 1467 383 1501 417
rect 1561 451 1595 485
rect 1561 383 1595 417
rect 1561 315 1595 349
rect 1655 451 1689 485
rect 1655 383 1689 417
rect 1655 315 1689 349
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 457 497 493 523
rect 551 497 587 523
rect 645 497 681 523
rect 739 497 775 523
rect 937 497 973 523
rect 1031 497 1067 523
rect 1125 497 1161 523
rect 1219 497 1255 523
rect 1325 497 1361 523
rect 1419 497 1455 523
rect 1513 497 1549 523
rect 1607 497 1643 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 457 282 493 297
rect 551 282 587 297
rect 645 282 681 297
rect 739 282 775 297
rect 937 282 973 297
rect 1031 282 1067 297
rect 1125 282 1161 297
rect 1219 282 1255 297
rect 1325 282 1361 297
rect 1419 282 1455 297
rect 1513 282 1549 297
rect 1607 282 1643 297
rect 79 261 119 282
rect 21 259 119 261
rect 173 259 213 282
rect 267 259 307 282
rect 361 259 401 282
rect 21 249 401 259
rect 21 215 38 249
rect 72 215 129 249
rect 163 215 223 249
rect 257 215 317 249
rect 351 215 401 249
rect 21 205 401 215
rect 89 177 119 205
rect 183 177 213 205
rect 277 177 307 205
rect 371 177 401 205
rect 455 259 495 282
rect 549 259 589 282
rect 643 259 683 282
rect 737 259 777 282
rect 935 259 975 282
rect 1029 259 1069 282
rect 1123 259 1163 282
rect 1217 259 1257 282
rect 455 249 777 259
rect 455 215 504 249
rect 538 215 599 249
rect 633 215 693 249
rect 727 215 777 249
rect 455 205 777 215
rect 869 249 1257 259
rect 869 215 885 249
rect 919 215 985 249
rect 1019 215 1079 249
rect 1113 215 1173 249
rect 1207 215 1257 249
rect 869 205 1257 215
rect 455 177 485 205
rect 549 177 579 205
rect 643 177 673 205
rect 747 177 777 205
rect 945 177 975 205
rect 1039 177 1069 205
rect 1133 177 1163 205
rect 1227 177 1257 205
rect 1323 259 1363 282
rect 1417 259 1457 282
rect 1511 259 1551 282
rect 1605 261 1645 282
rect 1605 259 1702 261
rect 1323 249 1702 259
rect 1323 215 1439 249
rect 1473 215 1533 249
rect 1567 215 1652 249
rect 1686 215 1702 249
rect 1323 205 1702 215
rect 1323 177 1353 205
rect 1417 177 1447 205
rect 1511 177 1541 205
rect 1605 177 1635 205
rect 89 21 119 47
rect 183 21 213 47
rect 277 21 307 47
rect 371 21 401 47
rect 455 21 485 47
rect 549 21 579 47
rect 643 21 673 47
rect 747 21 777 47
rect 945 21 975 47
rect 1039 21 1069 47
rect 1133 21 1163 47
rect 1227 21 1257 47
rect 1323 21 1353 47
rect 1417 21 1447 47
rect 1511 21 1541 47
rect 1605 21 1635 47
<< polycont >>
rect 38 215 72 249
rect 129 215 163 249
rect 223 215 257 249
rect 317 215 351 249
rect 504 215 538 249
rect 599 215 633 249
rect 693 215 727 249
rect 885 215 919 249
rect 985 215 1019 249
rect 1079 215 1113 249
rect 1173 215 1207 249
rect 1439 215 1473 249
rect 1533 215 1567 249
rect 1652 215 1686 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 18 485 69 527
rect 18 451 35 485
rect 18 417 69 451
rect 18 383 35 417
rect 18 349 69 383
rect 18 315 35 349
rect 18 289 69 315
rect 103 485 179 493
rect 103 451 129 485
rect 163 451 179 485
rect 103 417 179 451
rect 103 383 129 417
rect 163 383 179 417
rect 103 349 179 383
rect 223 485 257 527
rect 223 417 257 451
rect 223 367 257 383
rect 291 485 367 493
rect 291 451 317 485
rect 351 451 367 485
rect 291 417 367 451
rect 291 383 317 417
rect 351 383 367 417
rect 103 315 129 349
rect 163 333 179 349
rect 291 349 367 383
rect 411 485 445 527
rect 411 417 445 451
rect 411 367 445 383
rect 479 485 555 493
rect 479 451 505 485
rect 539 451 555 485
rect 479 417 555 451
rect 479 383 505 417
rect 539 383 555 417
rect 291 333 317 349
rect 163 315 317 333
rect 351 333 367 349
rect 479 349 555 383
rect 599 485 633 527
rect 599 417 633 451
rect 599 367 633 383
rect 667 485 743 493
rect 667 451 693 485
rect 727 451 743 485
rect 667 417 743 451
rect 667 383 693 417
rect 727 383 743 417
rect 479 333 505 349
rect 351 315 505 333
rect 539 333 555 349
rect 667 349 743 383
rect 787 485 925 527
rect 821 451 891 485
rect 787 417 925 451
rect 821 383 891 417
rect 787 367 925 383
rect 959 485 1035 493
rect 959 451 985 485
rect 1019 451 1035 485
rect 959 417 1035 451
rect 959 383 985 417
rect 1019 383 1035 417
rect 667 333 693 349
rect 539 315 693 333
rect 727 333 743 349
rect 959 349 1035 383
rect 1079 485 1113 527
rect 1079 417 1113 451
rect 1079 367 1113 383
rect 1147 485 1223 493
rect 1147 451 1173 485
rect 1207 451 1223 485
rect 1147 417 1223 451
rect 1147 383 1173 417
rect 1207 383 1223 417
rect 959 333 985 349
rect 727 315 985 333
rect 1019 333 1035 349
rect 1147 349 1223 383
rect 1274 485 1308 527
rect 1274 417 1308 451
rect 1274 367 1308 383
rect 1347 485 1423 493
rect 1347 451 1373 485
rect 1407 451 1423 485
rect 1347 417 1423 451
rect 1347 383 1373 417
rect 1407 383 1423 417
rect 1147 333 1173 349
rect 1019 315 1173 333
rect 1207 333 1223 349
rect 1347 349 1423 383
rect 1467 485 1501 527
rect 1467 417 1501 451
rect 1467 367 1501 383
rect 1535 485 1611 493
rect 1535 451 1561 485
rect 1595 451 1611 485
rect 1535 417 1611 451
rect 1535 383 1561 417
rect 1595 383 1611 417
rect 1347 333 1373 349
rect 1207 315 1373 333
rect 1407 333 1423 349
rect 1535 349 1611 383
rect 1535 333 1561 349
rect 1407 315 1561 333
rect 1595 315 1611 349
rect 103 289 1611 315
rect 1655 485 1707 527
rect 1689 451 1707 485
rect 1655 417 1707 451
rect 1689 383 1707 417
rect 1655 349 1707 383
rect 1689 315 1707 349
rect 1655 289 1707 315
rect 21 249 367 255
rect 21 215 38 249
rect 72 215 129 249
rect 163 215 223 249
rect 257 215 317 249
rect 351 215 367 249
rect 438 249 805 255
rect 438 215 504 249
rect 538 215 599 249
rect 633 215 693 249
rect 727 215 805 249
rect 850 249 1223 255
rect 850 215 885 249
rect 919 215 985 249
rect 1019 215 1079 249
rect 1113 215 1173 249
rect 1207 215 1223 249
rect 1309 181 1365 289
rect 1423 249 1702 255
rect 1423 215 1439 249
rect 1473 215 1533 249
rect 1567 215 1652 249
rect 1686 215 1702 249
rect 18 142 445 181
rect 18 108 35 142
rect 69 131 223 142
rect 18 51 69 108
rect 257 131 411 142
rect 103 63 129 97
rect 163 63 179 97
rect 103 17 179 63
rect 223 51 257 108
rect 479 165 1223 181
rect 479 131 505 165
rect 539 131 693 165
rect 727 131 985 165
rect 1019 131 1173 165
rect 1207 131 1223 165
rect 1309 165 1611 181
rect 1309 131 1373 165
rect 1407 131 1561 165
rect 1595 131 1611 165
rect 1655 165 1706 181
rect 1689 131 1706 165
rect 411 97 445 108
rect 1655 97 1706 131
rect 291 63 317 97
rect 351 63 367 97
rect 291 17 367 63
rect 411 63 599 97
rect 633 63 787 97
rect 821 63 837 97
rect 411 51 837 63
rect 875 63 891 97
rect 925 63 1079 97
rect 1113 63 1274 97
rect 1308 63 1467 97
rect 1501 63 1655 97
rect 1689 63 1706 97
rect 875 51 1706 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
<< metal1 >>
rect 0 561 1748 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 0 496 1748 527
rect 0 17 1748 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
rect 0 -48 1748 -17
<< labels >>
flabel corelocali s 1660 221 1694 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 1558 221 1592 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 1446 221 1480 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 200 0 0 0 D
port 4 nsew
flabel corelocali s 132 221 166 255 0 FreeSans 200 0 0 0 D
port 4 nsew
flabel corelocali s 231 238 231 238 0 FreeSans 200 0 0 0 D
port 4 nsew
flabel corelocali s 302 221 336 255 0 FreeSans 200 0 0 0 D
port 4 nsew
flabel corelocali s 438 221 472 255 0 FreeSans 200 0 0 0 C
port 3 nsew
flabel corelocali s 540 221 574 255 0 FreeSans 200 0 0 0 C
port 3 nsew
flabel corelocali s 744 221 778 255 0 FreeSans 200 0 0 0 C
port 3 nsew
flabel corelocali s 652 221 686 255 0 FreeSans 200 0 0 0 C
port 3 nsew
flabel corelocali s 1146 221 1181 255 0 FreeSans 200 0 0 0 B
port 2 nsew
flabel corelocali s 850 221 884 255 0 FreeSans 200 0 0 0 B
port 2 nsew
flabel corelocali s 942 221 976 255 0 FreeSans 200 0 0 0 B
port 2 nsew
flabel corelocali s 1044 221 1078 255 0 FreeSans 200 0 0 0 B
port 2 nsew
flabel corelocali s 1320 221 1354 255 0 FreeSans 200 0 0 0 Y
port 9 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
rlabel comment s 0 0 0 0 4 nand4_4
<< properties >>
string FIXED_BBOX 0 0 1748 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2315866
string GDS_START 2302012
<< end >>
