magic
tech sky130A
magscale 1 2
timestamp 1601050082
<< locali >>
rect 25 290 167 356
rect 201 290 267 356
rect 1481 430 1515 596
rect 993 290 1223 356
rect 1273 270 1375 356
rect 1481 364 1799 430
rect 1753 230 1799 364
rect 1448 196 1799 230
rect 1448 70 1514 196
rect 1648 154 1799 196
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 23 424 89 596
rect 123 458 189 649
rect 223 492 289 596
rect 378 526 445 649
rect 223 458 452 492
rect 23 390 335 424
rect 301 256 335 390
rect 386 290 452 458
rect 486 353 552 592
rect 593 387 659 649
rect 693 353 759 592
rect 793 387 859 649
rect 893 424 959 592
rect 993 458 1233 649
rect 1267 424 1333 572
rect 1375 458 1441 649
rect 1555 464 1621 649
rect 1735 464 1801 649
rect 893 390 1447 424
rect 893 353 959 390
rect 486 319 959 353
rect 508 272 552 319
rect 23 222 374 256
rect 23 70 73 222
rect 109 17 175 188
rect 209 117 306 188
rect 340 185 374 222
rect 408 219 474 256
rect 508 219 574 272
rect 610 251 832 285
rect 1413 330 1447 390
rect 440 185 474 219
rect 610 185 644 251
rect 766 219 832 251
rect 878 256 944 269
rect 1413 264 1713 330
rect 878 236 1130 256
rect 878 222 1312 236
rect 878 219 944 222
rect 340 151 406 185
rect 440 151 644 185
rect 680 185 730 217
rect 1080 202 1312 222
rect 978 185 1044 188
rect 680 151 1044 185
rect 372 117 406 151
rect 978 133 1044 151
rect 1080 133 1130 202
rect 209 51 338 117
rect 372 51 721 117
rect 1176 17 1226 168
rect 1262 90 1312 202
rect 1348 17 1414 226
rect 1548 17 1614 162
rect 1734 17 1801 120
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
<< metal1 >>
rect 0 683 1824 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 0 617 1824 649
rect 0 17 1824 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
rect 0 -49 1824 -17
<< labels >>
rlabel locali s 201 290 267 356 6 A_N
port 1 nsew signal input
rlabel locali s 25 290 167 356 6 B_N
port 2 nsew signal input
rlabel locali s 993 290 1223 356 6 C
port 3 nsew signal input
rlabel locali s 1273 270 1375 356 6 D
port 4 nsew signal input
rlabel locali s 1753 230 1799 364 6 X
port 5 nsew signal output
rlabel locali s 1648 154 1799 196 6 X
port 5 nsew signal output
rlabel locali s 1481 430 1515 596 6 X
port 5 nsew signal output
rlabel locali s 1481 364 1799 430 6 X
port 5 nsew signal output
rlabel locali s 1448 196 1799 230 6 X
port 5 nsew signal output
rlabel locali s 1448 70 1514 196 6 X
port 5 nsew signal output
rlabel metal1 s 0 -49 1824 49 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1824 715 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1824 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3160286
string GDS_START 3145826
<< end >>
