magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1932 561
rect 57 298 91 527
rect 125 265 191 485
rect 225 299 259 527
rect 293 288 349 493
rect 383 443 450 527
rect 921 447 987 527
rect 1755 455 1822 527
rect 293 265 342 288
rect 125 199 342 265
rect 57 17 91 147
rect 125 75 175 199
rect 293 185 342 199
rect 225 17 259 147
rect 293 70 345 185
rect 379 17 429 105
rect 599 215 712 265
rect 971 17 1005 173
rect 1521 289 1637 323
rect 1521 199 1555 289
rect 1685 215 1767 265
rect 1771 17 1805 113
rect 0 -17 1932 17
<< obsli1 >>
rect 486 447 780 481
rect 1054 455 1673 489
rect 486 409 520 447
rect 1054 413 1088 455
rect 383 375 520 409
rect 588 379 1088 413
rect 383 265 417 375
rect 463 307 780 341
rect 376 199 417 265
rect 382 173 417 199
rect 382 139 497 173
rect 463 85 497 139
rect 531 119 565 307
rect 746 265 780 307
rect 814 323 891 339
rect 814 305 857 323
rect 835 289 857 305
rect 835 275 891 289
rect 746 199 801 265
rect 625 159 701 181
rect 835 159 869 275
rect 925 241 959 379
rect 1005 289 1089 343
rect 625 125 869 159
rect 903 207 959 241
rect 903 91 937 207
rect 1041 187 1089 289
rect 690 85 777 91
rect 463 51 777 85
rect 811 57 937 91
rect 1075 153 1089 187
rect 1041 83 1089 153
rect 1125 119 1159 421
rect 1193 178 1227 455
rect 1856 421 1915 493
rect 1263 323 1346 409
rect 1453 387 1915 421
rect 1263 289 1317 323
rect 1351 289 1419 323
rect 1266 199 1351 254
rect 1309 187 1351 199
rect 1193 165 1235 178
rect 1193 144 1275 165
rect 1201 131 1275 144
rect 1125 85 1133 119
rect 1167 85 1207 97
rect 1125 53 1207 85
rect 1241 64 1275 131
rect 1309 153 1317 187
rect 1309 126 1351 153
rect 1385 85 1419 289
rect 1453 119 1487 387
rect 1818 375 1915 387
rect 1671 299 1835 341
rect 1801 265 1835 299
rect 1589 189 1651 255
rect 1801 199 1847 265
rect 1589 187 1630 189
rect 1589 153 1593 187
rect 1627 153 1630 187
rect 1801 181 1835 199
rect 1589 146 1630 153
rect 1687 150 1835 181
rect 1679 147 1835 150
rect 1679 119 1737 147
rect 1521 85 1614 93
rect 1385 51 1614 85
rect 1679 85 1685 119
rect 1719 85 1737 119
rect 1881 117 1915 375
rect 1679 59 1737 85
rect 1855 51 1915 117
<< obsli1c >>
rect 857 289 891 323
rect 1041 153 1075 187
rect 1317 289 1351 323
rect 1133 85 1167 119
rect 1317 153 1351 187
rect 1593 153 1627 187
rect 1685 85 1719 119
<< metal1 >>
rect 0 496 1932 592
rect 0 -48 1932 48
<< obsm1 >>
rect 845 323 903 329
rect 845 289 857 323
rect 891 320 903 323
rect 1305 323 1363 329
rect 1305 320 1317 323
rect 891 292 1317 320
rect 891 289 903 292
rect 845 283 903 289
rect 1305 289 1317 292
rect 1351 289 1363 323
rect 1305 283 1363 289
rect 1029 187 1087 193
rect 1029 153 1041 187
rect 1075 184 1087 187
rect 1305 187 1363 193
rect 1305 184 1317 187
rect 1075 156 1317 184
rect 1075 153 1087 156
rect 1029 147 1087 153
rect 1305 153 1317 156
rect 1351 184 1363 187
rect 1581 187 1639 193
rect 1581 184 1593 187
rect 1351 156 1593 184
rect 1351 153 1363 156
rect 1305 147 1363 153
rect 1581 153 1593 156
rect 1627 153 1639 187
rect 1581 147 1639 153
rect 1121 119 1179 125
rect 1121 85 1133 119
rect 1167 116 1179 119
rect 1673 119 1731 125
rect 1673 116 1685 119
rect 1167 88 1685 116
rect 1167 85 1179 88
rect 1121 79 1179 85
rect 1673 85 1685 88
rect 1719 85 1731 119
rect 1673 79 1731 85
<< labels >>
rlabel locali s 1685 215 1767 265 6 A
port 1 nsew signal input
rlabel locali s 1521 289 1637 323 6 B
port 2 nsew signal input
rlabel locali s 1521 199 1555 289 6 B
port 2 nsew signal input
rlabel locali s 599 215 712 265 6 C
port 3 nsew signal input
rlabel locali s 293 288 349 493 6 X
port 4 nsew signal output
rlabel locali s 293 265 342 288 6 X
port 4 nsew signal output
rlabel locali s 293 185 342 199 6 X
port 4 nsew signal output
rlabel locali s 293 70 345 185 6 X
port 4 nsew signal output
rlabel locali s 125 265 191 485 6 X
port 4 nsew signal output
rlabel locali s 125 199 342 265 6 X
port 4 nsew signal output
rlabel locali s 125 75 175 199 6 X
port 4 nsew signal output
rlabel locali s 1771 17 1805 113 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 971 17 1005 173 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 379 17 429 105 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 225 17 259 147 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 57 17 91 147 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 1932 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1932 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 1755 455 1822 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 921 447 987 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 383 443 450 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 225 299 259 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 57 298 91 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 1932 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 1932 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1932 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 580264
string GDS_START 567078
<< end >>
