magic
tech sky130A
magscale 1 2
timestamp 1599588244
<< locali >>
rect 25 290 110 356
rect 462 284 551 356
rect 585 284 651 356
rect 767 368 839 596
rect 805 234 839 368
rect 763 184 839 234
rect 965 236 1031 318
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 42 424 108 564
rect 156 458 222 649
rect 286 424 352 596
rect 413 458 479 649
rect 522 424 588 596
rect 640 458 706 649
rect 42 390 187 424
rect 153 334 187 390
rect 286 390 733 424
rect 286 388 352 390
rect 153 268 252 334
rect 153 256 187 268
rect 23 222 187 256
rect 286 234 320 388
rect 23 70 73 222
rect 109 17 175 188
rect 221 78 320 234
rect 354 234 420 318
rect 699 334 733 390
rect 873 420 923 649
rect 964 386 1033 540
rect 699 268 771 334
rect 354 200 729 234
rect 595 17 661 166
rect 695 150 729 200
rect 873 352 1033 386
rect 873 150 907 352
rect 967 150 1033 202
rect 695 116 1033 150
rect 865 17 931 82
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 683 1056 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 0 617 1056 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 1056 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -49 1056 -17
<< labels >>
rlabel locali s 25 290 110 356 6 A_N
port 1 nsew signal input
rlabel locali s 965 236 1031 318 6 B_N
port 2 nsew signal input
rlabel locali s 462 284 551 356 6 C
port 3 nsew signal input
rlabel locali s 585 284 651 356 6 D
port 4 nsew signal input
rlabel locali s 805 234 839 368 6 X
port 5 nsew signal output
rlabel locali s 767 368 839 596 6 X
port 5 nsew signal output
rlabel locali s 763 184 839 234 6 X
port 5 nsew signal output
rlabel metal1 s 0 -49 1056 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 7 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 617 1056 715 6 VPWR
port 9 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1056 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3240880
string GDS_START 3232492
<< end >>
