magic
tech sky130A
magscale 1 2
timestamp 1599588209
<< nwell >>
rect -38 332 230 704
<< pwell >>
rect 0 0 192 49
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 192 683
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 192 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 31 -17 65 17
rect 127 -17 161 17
<< metal1 >>
rect 0 683 192 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 192 683
rect 0 617 192 649
rect 0 17 192 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 192 17
rect 0 -49 192 -17
<< labels >>
flabel pwell s 0 0 192 49 0 FreeSans 200 0 0 0 VNB
port 2 nsew
flabel nwell s 0 617 192 666 0 FreeSans 200 0 0 0 VPB
port 3 nsew
rlabel comment s 0 0 0 0 4 fill_2
flabel metal1 s 0 617 192 666 0 FreeSans 200 0 0 0 VPWR
port 4 nsew
flabel metal1 s 0 0 192 49 0 FreeSans 200 0 0 0 VGND
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 192 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1802856
string GDS_START 1801436
<< end >>
