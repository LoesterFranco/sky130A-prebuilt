magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 828 561
rect 23 268 73 467
rect 179 387 269 527
rect 382 387 448 527
rect 490 352 528 493
rect 562 387 628 527
rect 662 353 700 493
rect 734 387 800 527
rect 662 352 811 353
rect 490 307 811 352
rect 23 199 175 268
rect 213 149 271 268
rect 305 199 380 265
rect 755 169 811 307
rect 490 123 811 169
rect 490 103 528 123
rect 381 17 447 89
rect 562 17 628 89
rect 662 51 700 123
rect 734 17 800 89
rect 0 -17 828 17
<< obsli1 >>
rect 109 350 145 493
rect 304 350 340 493
rect 109 316 456 350
rect 414 271 456 316
rect 93 113 160 161
rect 414 204 721 271
rect 414 161 456 204
rect 307 123 456 161
rect 307 113 345 123
rect 93 75 345 113
rect 93 51 160 75
<< metal1 >>
rect 0 496 828 592
rect 0 -48 828 48
<< labels >>
rlabel locali s 23 268 73 467 6 A
port 1 nsew signal input
rlabel locali s 23 199 175 268 6 A
port 1 nsew signal input
rlabel locali s 213 149 271 268 6 B
port 2 nsew signal input
rlabel locali s 305 199 380 265 6 C
port 3 nsew signal input
rlabel locali s 755 169 811 307 6 X
port 4 nsew signal output
rlabel locali s 662 353 700 493 6 X
port 4 nsew signal output
rlabel locali s 662 352 811 353 6 X
port 4 nsew signal output
rlabel locali s 662 51 700 123 6 X
port 4 nsew signal output
rlabel locali s 490 352 528 493 6 X
port 4 nsew signal output
rlabel locali s 490 307 811 352 6 X
port 4 nsew signal output
rlabel locali s 490 123 811 169 6 X
port 4 nsew signal output
rlabel locali s 490 103 528 123 6 X
port 4 nsew signal output
rlabel locali s 734 17 800 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 562 17 628 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 381 17 447 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 828 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 828 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 734 387 800 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 562 387 628 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 382 387 448 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 179 387 269 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 828 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 828 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3807562
string GDS_START 3800726
<< end >>
