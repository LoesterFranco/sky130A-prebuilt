magic
tech sky130A
magscale 1 2
timestamp 1599588232
<< locali >>
rect 21 260 87 356
rect 121 326 167 578
rect 225 394 291 596
rect 441 394 554 596
rect 225 360 554 394
rect 121 310 233 326
rect 133 260 233 310
rect 281 260 359 326
rect 313 88 359 260
rect 395 236 461 310
rect 519 202 554 360
rect 409 88 554 202
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 23 390 73 649
rect 341 428 407 649
rect 27 192 279 226
rect 27 70 93 192
rect 127 17 193 156
rect 229 70 279 192
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
rlabel locali s 21 260 87 356 6 A1
port 1 nsew signal input
rlabel locali s 133 260 233 310 6 A2
port 2 nsew signal input
rlabel locali s 121 326 167 578 6 A2
port 2 nsew signal input
rlabel locali s 121 310 233 326 6 A2
port 2 nsew signal input
rlabel locali s 313 88 359 260 6 B1
port 3 nsew signal input
rlabel locali s 281 260 359 326 6 B1
port 3 nsew signal input
rlabel locali s 395 236 461 310 6 C1
port 4 nsew signal input
rlabel locali s 519 202 554 360 6 Y
port 5 nsew signal output
rlabel locali s 441 394 554 596 6 Y
port 5 nsew signal output
rlabel locali s 409 88 554 202 6 Y
port 5 nsew signal output
rlabel locali s 225 394 291 596 6 Y
port 5 nsew signal output
rlabel locali s 225 360 554 394 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -49 576 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 7 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 617 576 715 6 VPWR
port 9 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 576 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1784214
string GDS_START 1777886
<< end >>
