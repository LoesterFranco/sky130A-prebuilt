magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 975 325 1025 493
rect 1163 325 1213 493
rect 1455 325 1505 425
rect 1643 325 1693 425
rect 975 291 1693 325
rect 85 215 405 257
rect 459 215 781 257
rect 1295 181 1361 291
rect 1413 215 1735 257
rect 1769 215 2188 257
rect 973 129 1361 181
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 31 359 81 527
rect 125 325 175 493
rect 219 359 269 527
rect 313 325 363 493
rect 407 359 457 527
rect 501 325 551 493
rect 595 359 645 527
rect 689 325 739 493
rect 783 359 931 527
rect 1069 359 1119 527
rect 1257 359 1307 527
rect 1355 459 1787 493
rect 1355 359 1411 459
rect 1549 359 1599 459
rect 17 291 863 325
rect 1737 325 1787 459
rect 1831 359 1881 527
rect 1925 325 1975 493
rect 2019 359 2069 527
rect 2113 325 2175 493
rect 1737 291 2175 325
rect 17 181 51 291
rect 829 257 863 291
rect 829 215 1261 257
rect 17 129 371 181
rect 415 145 841 181
rect 415 95 465 145
rect 20 51 465 95
rect 509 17 543 111
rect 577 51 653 145
rect 697 17 731 111
rect 765 51 841 145
rect 892 95 929 167
rect 1395 147 2171 181
rect 1395 95 1429 147
rect 1531 145 2171 147
rect 892 51 1429 95
rect 1463 17 1497 111
rect 1531 51 1607 145
rect 1651 17 1685 111
rect 1719 51 1795 145
rect 1839 17 1873 111
rect 1907 51 1983 145
rect 2027 17 2061 111
rect 2095 51 2171 145
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
<< metal1 >>
rect 0 561 2208 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 0 496 2208 527
rect 0 17 2208 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
rect 0 -48 2208 -17
<< labels >>
rlabel locali s 459 215 781 257 6 A1_N
port 1 nsew signal input
rlabel locali s 85 215 405 257 6 A2_N
port 2 nsew signal input
rlabel locali s 1769 215 2188 257 6 B1
port 3 nsew signal input
rlabel locali s 1413 215 1735 257 6 B2
port 4 nsew signal input
rlabel locali s 1643 325 1693 425 6 Y
port 5 nsew signal output
rlabel locali s 1455 325 1505 425 6 Y
port 5 nsew signal output
rlabel locali s 1295 181 1361 291 6 Y
port 5 nsew signal output
rlabel locali s 1163 325 1213 493 6 Y
port 5 nsew signal output
rlabel locali s 975 325 1025 493 6 Y
port 5 nsew signal output
rlabel locali s 975 291 1693 325 6 Y
port 5 nsew signal output
rlabel locali s 973 129 1361 181 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -48 2208 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 2208 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2208 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 686526
string GDS_START 670836
<< end >>
