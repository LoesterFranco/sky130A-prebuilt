magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 17 823 136 889
rect 931 823 1209 877
rect 1275 823 1553 877
rect 17 199 136 265
rect 2348 823 2467 889
rect 2501 823 2620 889
rect 3415 823 3693 877
rect 3759 823 4037 877
rect 931 211 1209 265
rect 1275 211 1553 265
rect 2348 199 2467 265
rect 2501 199 2620 265
rect 4832 823 4951 889
rect 3415 211 3693 265
rect 3759 211 4037 265
rect 4832 199 4951 265
<< obsli1 >>
rect 0 1071 29 1105
rect 63 1071 121 1105
rect 155 1071 213 1105
rect 247 1071 305 1105
rect 339 1071 397 1105
rect 431 1071 489 1105
rect 523 1071 581 1105
rect 615 1071 673 1105
rect 707 1071 765 1105
rect 799 1071 857 1105
rect 891 1071 949 1105
rect 983 1071 1041 1105
rect 1075 1071 1133 1105
rect 1167 1071 1225 1105
rect 1259 1071 1317 1105
rect 1351 1071 1409 1105
rect 1443 1071 1501 1105
rect 1535 1071 1593 1105
rect 1627 1071 1685 1105
rect 1719 1071 1777 1105
rect 1811 1071 1869 1105
rect 1903 1071 1961 1105
rect 1995 1071 2053 1105
rect 2087 1071 2145 1105
rect 2179 1071 2237 1105
rect 2271 1071 2329 1105
rect 2363 1071 2421 1105
rect 2455 1071 2513 1105
rect 2547 1071 2605 1105
rect 2639 1071 2697 1105
rect 2731 1071 2789 1105
rect 2823 1071 2881 1105
rect 2915 1071 2973 1105
rect 3007 1071 3065 1105
rect 3099 1071 3157 1105
rect 3191 1071 3249 1105
rect 3283 1071 3341 1105
rect 3375 1071 3433 1105
rect 3467 1071 3525 1105
rect 3559 1071 3617 1105
rect 3651 1071 3709 1105
rect 3743 1071 3801 1105
rect 3835 1071 3893 1105
rect 3927 1071 3985 1105
rect 4019 1071 4077 1105
rect 4111 1071 4169 1105
rect 4203 1071 4261 1105
rect 4295 1071 4353 1105
rect 4387 1071 4445 1105
rect 4479 1071 4537 1105
rect 4571 1071 4629 1105
rect 4663 1071 4721 1105
rect 4755 1071 4813 1105
rect 4847 1071 4905 1105
rect 4939 1071 4968 1105
rect 54 966 112 1071
rect 154 923 204 1032
rect 238 966 296 1071
rect 397 1003 803 1037
rect 397 934 447 1003
rect 170 875 204 923
rect 481 875 547 969
rect 581 934 615 1003
rect 649 911 715 969
rect 749 945 803 1003
rect 837 979 887 1071
rect 921 945 987 1037
rect 1021 979 1075 1071
rect 1109 945 1175 1037
rect 749 911 1175 945
rect 1209 911 1275 1071
rect 1309 945 1375 1037
rect 1409 979 1463 1071
rect 1497 945 1563 1037
rect 1597 979 1647 1071
rect 1681 1003 2087 1037
rect 1681 945 1735 1003
rect 1309 911 1735 945
rect 1769 911 1835 969
rect 1869 934 1903 1003
rect 649 875 695 911
rect 170 809 407 875
rect 441 815 695 875
rect 1789 875 1835 911
rect 1937 875 2003 969
rect 2037 934 2087 1003
rect 2188 966 2246 1071
rect 2280 923 2330 1032
rect 2372 966 2430 1071
rect 2538 966 2596 1071
rect 2638 923 2688 1032
rect 2722 966 2780 1071
rect 2881 1003 3287 1037
rect 2881 934 2931 1003
rect 2280 875 2314 923
rect 170 767 204 809
rect 44 561 104 767
rect 138 595 204 767
rect 243 561 298 767
rect 347 660 407 775
rect 347 626 361 660
rect 395 626 407 660
rect 347 595 407 626
rect 441 731 507 815
rect 441 697 457 731
rect 491 697 507 731
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 407 561
rect 44 321 104 527
rect 138 321 204 493
rect 243 321 298 527
rect 347 462 407 493
rect 347 428 361 462
rect 395 428 407 462
rect 170 279 204 321
rect 347 313 407 428
rect 441 391 507 697
rect 541 660 595 781
rect 541 626 551 660
rect 585 626 595 660
rect 541 595 595 626
rect 629 731 695 815
rect 1789 815 2043 875
rect 629 697 645 731
rect 679 697 695 731
rect 441 357 457 391
rect 491 357 507 391
rect 170 213 407 279
rect 441 273 507 357
rect 541 462 595 493
rect 541 428 551 462
rect 585 428 595 462
rect 541 307 595 428
rect 629 391 695 697
rect 729 755 1175 789
rect 729 660 789 755
rect 729 626 741 660
rect 775 626 789 660
rect 729 595 789 626
rect 833 561 887 721
rect 921 660 987 755
rect 921 626 937 660
rect 971 626 987 660
rect 921 595 987 626
rect 1021 561 1075 721
rect 1109 660 1175 755
rect 1109 626 1125 660
rect 1159 626 1175 660
rect 1109 595 1175 626
rect 1209 561 1275 789
rect 1309 755 1755 789
rect 1309 660 1375 755
rect 1309 626 1325 660
rect 1359 626 1375 660
rect 1309 595 1375 626
rect 1409 561 1463 721
rect 1497 660 1563 755
rect 1497 626 1513 660
rect 1547 626 1563 660
rect 1497 595 1563 626
rect 1597 561 1651 721
rect 1695 660 1755 755
rect 1695 626 1709 660
rect 1743 626 1755 660
rect 1695 595 1755 626
rect 1789 731 1855 815
rect 1789 697 1805 731
rect 1839 697 1855 731
rect 729 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1755 561
rect 629 357 645 391
rect 679 357 695 391
rect 629 273 695 357
rect 729 462 789 493
rect 729 428 741 462
rect 775 428 789 462
rect 729 333 789 428
rect 833 367 887 527
rect 921 462 987 493
rect 921 428 937 462
rect 971 428 987 462
rect 921 333 987 428
rect 1021 367 1075 527
rect 1109 462 1175 493
rect 1109 428 1125 462
rect 1159 428 1175 462
rect 1109 333 1175 428
rect 729 299 1175 333
rect 1209 299 1275 527
rect 1309 462 1375 493
rect 1309 428 1325 462
rect 1359 428 1375 462
rect 1309 333 1375 428
rect 1409 367 1463 527
rect 1497 462 1563 493
rect 1497 428 1513 462
rect 1547 428 1563 462
rect 1497 333 1563 428
rect 1597 367 1651 527
rect 1695 462 1755 493
rect 1695 428 1709 462
rect 1743 428 1755 462
rect 1695 333 1755 428
rect 1309 299 1755 333
rect 1789 391 1855 697
rect 1889 660 1943 781
rect 1889 626 1899 660
rect 1933 626 1943 660
rect 1889 595 1943 626
rect 1977 731 2043 815
rect 2077 809 2314 875
rect 2654 875 2688 923
rect 2965 875 3031 969
rect 3065 934 3099 1003
rect 3133 911 3199 969
rect 3233 945 3287 1003
rect 3321 979 3371 1071
rect 3405 945 3471 1037
rect 3505 979 3559 1071
rect 3593 945 3659 1037
rect 3233 911 3659 945
rect 3693 911 3759 1071
rect 3793 945 3859 1037
rect 3893 979 3947 1071
rect 3981 945 4047 1037
rect 4081 979 4131 1071
rect 4165 1003 4571 1037
rect 4165 945 4219 1003
rect 3793 911 4219 945
rect 4253 911 4319 969
rect 4353 934 4387 1003
rect 3133 875 3179 911
rect 1977 697 1993 731
rect 2027 697 2043 731
rect 1789 357 1805 391
rect 1839 357 1855 391
rect 441 213 695 273
rect 1789 273 1855 357
rect 1889 462 1943 493
rect 1889 428 1899 462
rect 1933 428 1943 462
rect 1889 307 1943 428
rect 1977 391 2043 697
rect 2077 660 2137 775
rect 2280 767 2314 809
rect 2654 809 2891 875
rect 2925 815 3179 875
rect 4273 875 4319 911
rect 4421 875 4487 969
rect 4521 934 4571 1003
rect 4672 966 4730 1071
rect 4764 923 4814 1032
rect 4856 966 4914 1071
rect 4764 875 4798 923
rect 2654 767 2688 809
rect 2077 626 2089 660
rect 2123 626 2137 660
rect 2077 595 2137 626
rect 2186 561 2241 767
rect 2280 595 2346 767
rect 2380 561 2440 767
rect 2528 561 2588 767
rect 2622 595 2688 767
rect 2727 561 2782 767
rect 2831 660 2891 775
rect 2831 626 2845 660
rect 2879 626 2891 660
rect 2831 595 2891 626
rect 2925 731 2991 815
rect 2925 697 2941 731
rect 2975 697 2991 731
rect 2077 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2891 561
rect 1977 357 1993 391
rect 2027 357 2043 391
rect 1977 273 2043 357
rect 2077 462 2137 493
rect 2077 428 2089 462
rect 2123 428 2137 462
rect 2077 313 2137 428
rect 2186 321 2241 527
rect 2280 321 2346 493
rect 2380 321 2440 527
rect 2528 321 2588 527
rect 2622 321 2688 493
rect 2727 321 2782 527
rect 2831 462 2891 493
rect 2831 428 2845 462
rect 2879 428 2891 462
rect 2280 279 2314 321
rect 170 165 204 213
rect 54 17 112 122
rect 154 56 204 165
rect 238 17 296 122
rect 397 85 447 154
rect 481 119 547 213
rect 649 177 695 213
rect 1789 213 2043 273
rect 2077 213 2314 279
rect 2654 279 2688 321
rect 2831 313 2891 428
rect 2925 391 2991 697
rect 3025 660 3079 781
rect 3025 626 3035 660
rect 3069 626 3079 660
rect 3025 595 3079 626
rect 3113 731 3179 815
rect 4273 815 4527 875
rect 3113 697 3129 731
rect 3163 697 3179 731
rect 2925 357 2941 391
rect 2975 357 2991 391
rect 1789 177 1835 213
rect 581 85 615 154
rect 649 119 715 177
rect 749 143 1175 177
rect 749 85 803 143
rect 397 51 803 85
rect 837 17 887 109
rect 921 51 987 143
rect 1021 17 1075 109
rect 1109 51 1175 143
rect 1209 17 1275 177
rect 1309 143 1735 177
rect 1309 51 1375 143
rect 1409 17 1463 109
rect 1497 51 1563 143
rect 1597 17 1647 109
rect 1681 85 1735 143
rect 1769 119 1835 177
rect 1869 85 1903 154
rect 1937 119 2003 213
rect 2280 165 2314 213
rect 2654 213 2891 279
rect 2925 273 2991 357
rect 3025 462 3079 493
rect 3025 428 3035 462
rect 3069 428 3079 462
rect 3025 307 3079 428
rect 3113 391 3179 697
rect 3213 755 3659 789
rect 3213 660 3273 755
rect 3213 626 3225 660
rect 3259 626 3273 660
rect 3213 595 3273 626
rect 3317 561 3371 721
rect 3405 660 3471 755
rect 3405 626 3421 660
rect 3455 626 3471 660
rect 3405 595 3471 626
rect 3505 561 3559 721
rect 3593 660 3659 755
rect 3593 626 3609 660
rect 3643 626 3659 660
rect 3593 595 3659 626
rect 3693 561 3759 789
rect 3793 755 4239 789
rect 3793 660 3859 755
rect 3793 626 3809 660
rect 3843 626 3859 660
rect 3793 595 3859 626
rect 3893 561 3947 721
rect 3981 660 4047 755
rect 3981 626 3997 660
rect 4031 626 4047 660
rect 3981 595 4047 626
rect 4081 561 4135 721
rect 4179 660 4239 755
rect 4179 626 4193 660
rect 4227 626 4239 660
rect 4179 595 4239 626
rect 4273 731 4339 815
rect 4273 697 4289 731
rect 4323 697 4339 731
rect 3213 527 3249 561
rect 3283 527 3341 561
rect 3375 527 3433 561
rect 3467 527 3525 561
rect 3559 527 3617 561
rect 3651 527 3709 561
rect 3743 527 3801 561
rect 3835 527 3893 561
rect 3927 527 3985 561
rect 4019 527 4077 561
rect 4111 527 4169 561
rect 4203 527 4239 561
rect 3113 357 3129 391
rect 3163 357 3179 391
rect 3113 273 3179 357
rect 3213 462 3273 493
rect 3213 428 3225 462
rect 3259 428 3273 462
rect 3213 333 3273 428
rect 3317 367 3371 527
rect 3405 462 3471 493
rect 3405 428 3421 462
rect 3455 428 3471 462
rect 3405 333 3471 428
rect 3505 367 3559 527
rect 3593 462 3659 493
rect 3593 428 3609 462
rect 3643 428 3659 462
rect 3593 333 3659 428
rect 3213 299 3659 333
rect 3693 299 3759 527
rect 3793 462 3859 493
rect 3793 428 3809 462
rect 3843 428 3859 462
rect 3793 333 3859 428
rect 3893 367 3947 527
rect 3981 462 4047 493
rect 3981 428 3997 462
rect 4031 428 4047 462
rect 3981 333 4047 428
rect 4081 367 4135 527
rect 4179 462 4239 493
rect 4179 428 4193 462
rect 4227 428 4239 462
rect 4179 333 4239 428
rect 3793 299 4239 333
rect 4273 391 4339 697
rect 4373 660 4427 781
rect 4373 626 4383 660
rect 4417 626 4427 660
rect 4373 595 4427 626
rect 4461 731 4527 815
rect 4561 809 4798 875
rect 4461 697 4477 731
rect 4511 697 4527 731
rect 4273 357 4289 391
rect 4323 357 4339 391
rect 2925 213 3179 273
rect 4273 273 4339 357
rect 4373 462 4427 493
rect 4373 428 4383 462
rect 4417 428 4427 462
rect 4373 307 4427 428
rect 4461 391 4527 697
rect 4561 660 4621 775
rect 4764 767 4798 809
rect 4561 626 4573 660
rect 4607 626 4621 660
rect 4561 595 4621 626
rect 4670 561 4725 767
rect 4764 595 4830 767
rect 4864 561 4924 767
rect 4561 527 4629 561
rect 4663 527 4721 561
rect 4755 527 4813 561
rect 4847 527 4905 561
rect 4939 527 4968 561
rect 4461 357 4477 391
rect 4511 357 4527 391
rect 4461 273 4527 357
rect 4561 462 4621 493
rect 4561 428 4573 462
rect 4607 428 4621 462
rect 4561 313 4621 428
rect 4670 321 4725 527
rect 4764 321 4830 493
rect 4864 321 4924 527
rect 4764 279 4798 321
rect 2654 165 2688 213
rect 2037 85 2087 154
rect 1681 51 2087 85
rect 2188 17 2246 122
rect 2280 56 2330 165
rect 2372 17 2430 122
rect 2538 17 2596 122
rect 2638 56 2688 165
rect 2722 17 2780 122
rect 2881 85 2931 154
rect 2965 119 3031 213
rect 3133 177 3179 213
rect 4273 213 4527 273
rect 4561 213 4798 279
rect 4273 177 4319 213
rect 3065 85 3099 154
rect 3133 119 3199 177
rect 3233 143 3659 177
rect 3233 85 3287 143
rect 2881 51 3287 85
rect 3321 17 3371 109
rect 3405 51 3471 143
rect 3505 17 3559 109
rect 3593 51 3659 143
rect 3693 17 3759 177
rect 3793 143 4219 177
rect 3793 51 3859 143
rect 3893 17 3947 109
rect 3981 51 4047 143
rect 4081 17 4131 109
rect 4165 85 4219 143
rect 4253 119 4319 177
rect 4353 85 4387 154
rect 4421 119 4487 213
rect 4764 165 4798 213
rect 4521 85 4571 154
rect 4165 51 4571 85
rect 4672 17 4730 122
rect 4764 56 4814 165
rect 4856 17 4914 122
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3341 17
rect 3375 -17 3433 17
rect 3467 -17 3525 17
rect 3559 -17 3617 17
rect 3651 -17 3709 17
rect 3743 -17 3801 17
rect 3835 -17 3893 17
rect 3927 -17 3985 17
rect 4019 -17 4077 17
rect 4111 -17 4169 17
rect 4203 -17 4261 17
rect 4295 -17 4353 17
rect 4387 -17 4445 17
rect 4479 -17 4537 17
rect 4571 -17 4629 17
rect 4663 -17 4721 17
rect 4755 -17 4813 17
rect 4847 -17 4905 17
rect 4939 -17 4968 17
<< obsli1c >>
rect 29 1071 63 1105
rect 121 1071 155 1105
rect 213 1071 247 1105
rect 305 1071 339 1105
rect 397 1071 431 1105
rect 489 1071 523 1105
rect 581 1071 615 1105
rect 673 1071 707 1105
rect 765 1071 799 1105
rect 857 1071 891 1105
rect 949 1071 983 1105
rect 1041 1071 1075 1105
rect 1133 1071 1167 1105
rect 1225 1071 1259 1105
rect 1317 1071 1351 1105
rect 1409 1071 1443 1105
rect 1501 1071 1535 1105
rect 1593 1071 1627 1105
rect 1685 1071 1719 1105
rect 1777 1071 1811 1105
rect 1869 1071 1903 1105
rect 1961 1071 1995 1105
rect 2053 1071 2087 1105
rect 2145 1071 2179 1105
rect 2237 1071 2271 1105
rect 2329 1071 2363 1105
rect 2421 1071 2455 1105
rect 2513 1071 2547 1105
rect 2605 1071 2639 1105
rect 2697 1071 2731 1105
rect 2789 1071 2823 1105
rect 2881 1071 2915 1105
rect 2973 1071 3007 1105
rect 3065 1071 3099 1105
rect 3157 1071 3191 1105
rect 3249 1071 3283 1105
rect 3341 1071 3375 1105
rect 3433 1071 3467 1105
rect 3525 1071 3559 1105
rect 3617 1071 3651 1105
rect 3709 1071 3743 1105
rect 3801 1071 3835 1105
rect 3893 1071 3927 1105
rect 3985 1071 4019 1105
rect 4077 1071 4111 1105
rect 4169 1071 4203 1105
rect 4261 1071 4295 1105
rect 4353 1071 4387 1105
rect 4445 1071 4479 1105
rect 4537 1071 4571 1105
rect 4629 1071 4663 1105
rect 4721 1071 4755 1105
rect 4813 1071 4847 1105
rect 4905 1071 4939 1105
rect 361 626 395 660
rect 457 697 491 731
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 361 428 395 462
rect 551 626 585 660
rect 645 697 679 731
rect 457 357 491 391
rect 551 428 585 462
rect 741 626 775 660
rect 937 626 971 660
rect 1125 626 1159 660
rect 1325 626 1359 660
rect 1513 626 1547 660
rect 1709 626 1743 660
rect 1805 697 1839 731
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 645 357 679 391
rect 741 428 775 462
rect 937 428 971 462
rect 1125 428 1159 462
rect 1325 428 1359 462
rect 1513 428 1547 462
rect 1709 428 1743 462
rect 1899 626 1933 660
rect 1993 697 2027 731
rect 1805 357 1839 391
rect 1899 428 1933 462
rect 2089 626 2123 660
rect 2845 626 2879 660
rect 2941 697 2975 731
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 1993 357 2027 391
rect 2089 428 2123 462
rect 2845 428 2879 462
rect 3035 626 3069 660
rect 3129 697 3163 731
rect 2941 357 2975 391
rect 3035 428 3069 462
rect 3225 626 3259 660
rect 3421 626 3455 660
rect 3609 626 3643 660
rect 3809 626 3843 660
rect 3997 626 4031 660
rect 4193 626 4227 660
rect 4289 697 4323 731
rect 3249 527 3283 561
rect 3341 527 3375 561
rect 3433 527 3467 561
rect 3525 527 3559 561
rect 3617 527 3651 561
rect 3709 527 3743 561
rect 3801 527 3835 561
rect 3893 527 3927 561
rect 3985 527 4019 561
rect 4077 527 4111 561
rect 4169 527 4203 561
rect 3129 357 3163 391
rect 3225 428 3259 462
rect 3421 428 3455 462
rect 3609 428 3643 462
rect 3809 428 3843 462
rect 3997 428 4031 462
rect 4193 428 4227 462
rect 4383 626 4417 660
rect 4477 697 4511 731
rect 4289 357 4323 391
rect 4383 428 4417 462
rect 4573 626 4607 660
rect 4629 527 4663 561
rect 4721 527 4755 561
rect 4813 527 4847 561
rect 4905 527 4939 561
rect 4477 357 4511 391
rect 4573 428 4607 462
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
rect 2881 -17 2915 17
rect 2973 -17 3007 17
rect 3065 -17 3099 17
rect 3157 -17 3191 17
rect 3249 -17 3283 17
rect 3341 -17 3375 17
rect 3433 -17 3467 17
rect 3525 -17 3559 17
rect 3617 -17 3651 17
rect 3709 -17 3743 17
rect 3801 -17 3835 17
rect 3893 -17 3927 17
rect 3985 -17 4019 17
rect 4077 -17 4111 17
rect 4169 -17 4203 17
rect 4261 -17 4295 17
rect 4353 -17 4387 17
rect 4445 -17 4479 17
rect 4537 -17 4571 17
rect 4629 -17 4663 17
rect 4721 -17 4755 17
rect 4813 -17 4847 17
rect 4905 -17 4939 17
<< metal1 >>
rect 0 1105 4968 1136
rect 0 1071 29 1105
rect 63 1071 121 1105
rect 155 1071 213 1105
rect 247 1071 305 1105
rect 339 1071 397 1105
rect 431 1071 489 1105
rect 523 1071 581 1105
rect 615 1071 673 1105
rect 707 1071 765 1105
rect 799 1071 857 1105
rect 891 1071 949 1105
rect 983 1071 1041 1105
rect 1075 1071 1133 1105
rect 1167 1071 1225 1105
rect 1259 1071 1317 1105
rect 1351 1071 1409 1105
rect 1443 1071 1501 1105
rect 1535 1071 1593 1105
rect 1627 1071 1685 1105
rect 1719 1071 1777 1105
rect 1811 1071 1869 1105
rect 1903 1071 1961 1105
rect 1995 1071 2053 1105
rect 2087 1071 2145 1105
rect 2179 1071 2237 1105
rect 2271 1071 2329 1105
rect 2363 1071 2421 1105
rect 2455 1071 2513 1105
rect 2547 1071 2605 1105
rect 2639 1071 2697 1105
rect 2731 1071 2789 1105
rect 2823 1071 2881 1105
rect 2915 1071 2973 1105
rect 3007 1071 3065 1105
rect 3099 1071 3157 1105
rect 3191 1071 3249 1105
rect 3283 1071 3341 1105
rect 3375 1071 3433 1105
rect 3467 1071 3525 1105
rect 3559 1071 3617 1105
rect 3651 1071 3709 1105
rect 3743 1071 3801 1105
rect 3835 1071 3893 1105
rect 3927 1071 3985 1105
rect 4019 1071 4077 1105
rect 4111 1071 4169 1105
rect 4203 1071 4261 1105
rect 4295 1071 4353 1105
rect 4387 1071 4445 1105
rect 4479 1071 4537 1105
rect 4571 1071 4629 1105
rect 4663 1071 4721 1105
rect 4755 1071 4813 1105
rect 4847 1071 4905 1105
rect 4939 1071 4968 1105
rect 0 1040 4968 1071
rect 445 731 503 737
rect 445 697 457 731
rect 491 728 503 731
rect 633 731 691 737
rect 633 728 645 731
rect 491 700 645 728
rect 491 697 503 700
rect 445 691 503 697
rect 633 697 645 700
rect 679 728 691 731
rect 1793 731 1851 737
rect 1793 728 1805 731
rect 679 700 1805 728
rect 679 697 691 700
rect 633 691 691 697
rect 1793 697 1805 700
rect 1839 728 1851 731
rect 1981 731 2039 737
rect 1981 728 1993 731
rect 1839 700 1993 728
rect 1839 697 1851 700
rect 1793 691 1851 697
rect 1981 697 1993 700
rect 2027 728 2039 731
rect 2929 731 2987 737
rect 2929 728 2941 731
rect 2027 700 2941 728
rect 2027 697 2039 700
rect 1981 691 2039 697
rect 2929 697 2941 700
rect 2975 728 2987 731
rect 3117 731 3175 737
rect 3117 728 3129 731
rect 2975 700 3129 728
rect 2975 697 2987 700
rect 2929 691 2987 697
rect 3117 697 3129 700
rect 3163 728 3175 731
rect 4277 731 4335 737
rect 4277 728 4289 731
rect 3163 700 4289 728
rect 3163 697 3175 700
rect 3117 691 3175 697
rect 4277 697 4289 700
rect 4323 728 4335 731
rect 4465 731 4523 737
rect 4465 728 4477 731
rect 4323 700 4477 728
rect 4323 697 4335 700
rect 4277 691 4335 697
rect 4465 697 4477 700
rect 4511 697 4523 731
rect 4465 691 4523 697
rect 0 561 4968 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 3249 561
rect 3283 527 3341 561
rect 3375 527 3433 561
rect 3467 527 3525 561
rect 3559 527 3617 561
rect 3651 527 3709 561
rect 3743 527 3801 561
rect 3835 527 3893 561
rect 3927 527 3985 561
rect 4019 527 4077 561
rect 4111 527 4169 561
rect 4203 527 4629 561
rect 4663 527 4721 561
rect 4755 527 4813 561
rect 4847 527 4905 561
rect 4939 527 4968 561
rect 0 496 4968 527
rect 445 391 503 397
rect 445 357 457 391
rect 491 388 503 391
rect 633 391 691 397
rect 633 388 645 391
rect 491 360 645 388
rect 491 357 503 360
rect 445 351 503 357
rect 633 357 645 360
rect 679 388 691 391
rect 1793 391 1851 397
rect 1793 388 1805 391
rect 679 360 1805 388
rect 679 357 691 360
rect 633 351 691 357
rect 1793 357 1805 360
rect 1839 388 1851 391
rect 1981 391 2039 397
rect 1981 388 1993 391
rect 1839 360 1993 388
rect 1839 357 1851 360
rect 1793 351 1851 357
rect 1981 357 1993 360
rect 2027 388 2039 391
rect 2929 391 2987 397
rect 2929 388 2941 391
rect 2027 360 2941 388
rect 2027 357 2039 360
rect 1981 351 2039 357
rect 2929 357 2941 360
rect 2975 388 2987 391
rect 3117 391 3175 397
rect 3117 388 3129 391
rect 2975 360 3129 388
rect 2975 357 2987 360
rect 2929 351 2987 357
rect 3117 357 3129 360
rect 3163 388 3175 391
rect 4277 391 4335 397
rect 4277 388 4289 391
rect 3163 360 4289 388
rect 3163 357 3175 360
rect 3117 351 3175 357
rect 4277 357 4289 360
rect 4323 388 4335 391
rect 4465 391 4523 397
rect 4465 388 4477 391
rect 4323 360 4477 388
rect 4323 357 4335 360
rect 4277 351 4335 357
rect 4465 357 4477 360
rect 4511 357 4523 391
rect 4465 351 4523 357
rect 0 17 4968 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3341 17
rect 3375 -17 3433 17
rect 3467 -17 3525 17
rect 3559 -17 3617 17
rect 3651 -17 3709 17
rect 3743 -17 3801 17
rect 3835 -17 3893 17
rect 3927 -17 3985 17
rect 4019 -17 4077 17
rect 4111 -17 4169 17
rect 4203 -17 4261 17
rect 4295 -17 4353 17
rect 4387 -17 4445 17
rect 4479 -17 4537 17
rect 4571 -17 4629 17
rect 4663 -17 4721 17
rect 4755 -17 4813 17
rect 4847 -17 4905 17
rect 4939 -17 4968 17
rect 0 -48 4968 -17
<< obsm1 >>
rect 349 660 407 666
rect 349 626 361 660
rect 395 657 407 660
rect 539 660 597 666
rect 539 657 551 660
rect 395 629 551 657
rect 395 626 407 629
rect 349 620 407 626
rect 539 626 551 629
rect 585 657 597 660
rect 729 660 787 666
rect 729 657 741 660
rect 585 629 741 657
rect 585 626 597 629
rect 539 620 597 626
rect 729 626 741 629
rect 775 657 787 660
rect 925 660 983 666
rect 925 657 937 660
rect 775 629 937 657
rect 775 626 787 629
rect 729 620 787 626
rect 925 626 937 629
rect 971 657 983 660
rect 1113 660 1171 666
rect 1113 657 1125 660
rect 971 629 1125 657
rect 971 626 983 629
rect 925 620 983 626
rect 1113 626 1125 629
rect 1159 626 1171 660
rect 1113 620 1171 626
rect 1313 660 1371 666
rect 1313 626 1325 660
rect 1359 657 1371 660
rect 1501 660 1559 666
rect 1501 657 1513 660
rect 1359 629 1513 657
rect 1359 626 1371 629
rect 1313 620 1371 626
rect 1501 626 1513 629
rect 1547 657 1559 660
rect 1697 660 1755 666
rect 1697 657 1709 660
rect 1547 629 1709 657
rect 1547 626 1559 629
rect 1501 620 1559 626
rect 1697 626 1709 629
rect 1743 657 1755 660
rect 1887 660 1945 666
rect 1887 657 1899 660
rect 1743 629 1899 657
rect 1743 626 1755 629
rect 1697 620 1755 626
rect 1887 626 1899 629
rect 1933 657 1945 660
rect 2077 660 2135 666
rect 2077 657 2089 660
rect 1933 629 2089 657
rect 1933 626 1945 629
rect 1887 620 1945 626
rect 2077 626 2089 629
rect 2123 626 2135 660
rect 2077 620 2135 626
rect 2833 660 2891 666
rect 2833 626 2845 660
rect 2879 657 2891 660
rect 3023 660 3081 666
rect 3023 657 3035 660
rect 2879 629 3035 657
rect 2879 626 2891 629
rect 2833 620 2891 626
rect 3023 626 3035 629
rect 3069 657 3081 660
rect 3213 660 3271 666
rect 3213 657 3225 660
rect 3069 629 3225 657
rect 3069 626 3081 629
rect 3023 620 3081 626
rect 3213 626 3225 629
rect 3259 657 3271 660
rect 3409 660 3467 666
rect 3409 657 3421 660
rect 3259 629 3421 657
rect 3259 626 3271 629
rect 3213 620 3271 626
rect 3409 626 3421 629
rect 3455 657 3467 660
rect 3597 660 3655 666
rect 3597 657 3609 660
rect 3455 629 3609 657
rect 3455 626 3467 629
rect 3409 620 3467 626
rect 3597 626 3609 629
rect 3643 626 3655 660
rect 3597 620 3655 626
rect 3797 660 3855 666
rect 3797 626 3809 660
rect 3843 657 3855 660
rect 3985 660 4043 666
rect 3985 657 3997 660
rect 3843 629 3997 657
rect 3843 626 3855 629
rect 3797 620 3855 626
rect 3985 626 3997 629
rect 4031 657 4043 660
rect 4181 660 4239 666
rect 4181 657 4193 660
rect 4031 629 4193 657
rect 4031 626 4043 629
rect 3985 620 4043 626
rect 4181 626 4193 629
rect 4227 657 4239 660
rect 4371 660 4429 666
rect 4371 657 4383 660
rect 4227 629 4383 657
rect 4227 626 4239 629
rect 4181 620 4239 626
rect 4371 626 4383 629
rect 4417 657 4429 660
rect 4561 660 4619 666
rect 4561 657 4573 660
rect 4417 629 4573 657
rect 4417 626 4429 629
rect 4371 620 4429 626
rect 4561 626 4573 629
rect 4607 626 4619 660
rect 4561 620 4619 626
rect 349 462 407 468
rect 349 428 361 462
rect 395 459 407 462
rect 539 462 597 468
rect 539 459 551 462
rect 395 431 551 459
rect 395 428 407 431
rect 349 422 407 428
rect 539 428 551 431
rect 585 459 597 462
rect 729 462 787 468
rect 729 459 741 462
rect 585 431 741 459
rect 585 428 597 431
rect 539 422 597 428
rect 729 428 741 431
rect 775 459 787 462
rect 925 462 983 468
rect 925 459 937 462
rect 775 431 937 459
rect 775 428 787 431
rect 729 422 787 428
rect 925 428 937 431
rect 971 459 983 462
rect 1113 462 1171 468
rect 1113 459 1125 462
rect 971 431 1125 459
rect 971 428 983 431
rect 925 422 983 428
rect 1113 428 1125 431
rect 1159 428 1171 462
rect 1113 422 1171 428
rect 1313 462 1371 468
rect 1313 428 1325 462
rect 1359 459 1371 462
rect 1501 462 1559 468
rect 1501 459 1513 462
rect 1359 431 1513 459
rect 1359 428 1371 431
rect 1313 422 1371 428
rect 1501 428 1513 431
rect 1547 459 1559 462
rect 1697 462 1755 468
rect 1697 459 1709 462
rect 1547 431 1709 459
rect 1547 428 1559 431
rect 1501 422 1559 428
rect 1697 428 1709 431
rect 1743 459 1755 462
rect 1887 462 1945 468
rect 1887 459 1899 462
rect 1743 431 1899 459
rect 1743 428 1755 431
rect 1697 422 1755 428
rect 1887 428 1899 431
rect 1933 459 1945 462
rect 2077 462 2135 468
rect 2077 459 2089 462
rect 1933 431 2089 459
rect 1933 428 1945 431
rect 1887 422 1945 428
rect 2077 428 2089 431
rect 2123 428 2135 462
rect 2077 422 2135 428
rect 2833 462 2891 468
rect 2833 428 2845 462
rect 2879 459 2891 462
rect 3023 462 3081 468
rect 3023 459 3035 462
rect 2879 431 3035 459
rect 2879 428 2891 431
rect 2833 422 2891 428
rect 3023 428 3035 431
rect 3069 459 3081 462
rect 3213 462 3271 468
rect 3213 459 3225 462
rect 3069 431 3225 459
rect 3069 428 3081 431
rect 3023 422 3081 428
rect 3213 428 3225 431
rect 3259 459 3271 462
rect 3409 462 3467 468
rect 3409 459 3421 462
rect 3259 431 3421 459
rect 3259 428 3271 431
rect 3213 422 3271 428
rect 3409 428 3421 431
rect 3455 459 3467 462
rect 3597 462 3655 468
rect 3597 459 3609 462
rect 3455 431 3609 459
rect 3455 428 3467 431
rect 3409 422 3467 428
rect 3597 428 3609 431
rect 3643 428 3655 462
rect 3597 422 3655 428
rect 3797 462 3855 468
rect 3797 428 3809 462
rect 3843 459 3855 462
rect 3985 462 4043 468
rect 3985 459 3997 462
rect 3843 431 3997 459
rect 3843 428 3855 431
rect 3797 422 3855 428
rect 3985 428 3997 431
rect 4031 459 4043 462
rect 4181 462 4239 468
rect 4181 459 4193 462
rect 4031 431 4193 459
rect 4031 428 4043 431
rect 3985 422 4043 428
rect 4181 428 4193 431
rect 4227 459 4239 462
rect 4371 462 4429 468
rect 4371 459 4383 462
rect 4227 431 4383 459
rect 4227 428 4239 431
rect 4181 422 4239 428
rect 4371 428 4383 431
rect 4417 459 4429 462
rect 4561 462 4619 468
rect 4561 459 4573 462
rect 4417 431 4573 459
rect 4417 428 4429 431
rect 4371 422 4429 428
rect 4561 428 4573 431
rect 4607 428 4619 462
rect 4561 422 4619 428
<< labels >>
rlabel locali s 931 211 1209 265 6 D[0]
port 1 nsew signal input
rlabel locali s 931 823 1209 877 6 D[1]
port 2 nsew signal input
rlabel locali s 1275 211 1553 265 6 D[2]
port 3 nsew signal input
rlabel locali s 1275 823 1553 877 6 D[3]
port 4 nsew signal input
rlabel locali s 3415 211 3693 265 6 D[4]
port 5 nsew signal input
rlabel locali s 3415 823 3693 877 6 D[5]
port 6 nsew signal input
rlabel locali s 3759 211 4037 265 6 D[6]
port 7 nsew signal input
rlabel locali s 3759 823 4037 877 6 D[7]
port 8 nsew signal input
rlabel locali s 17 199 136 265 6 S[0]
port 9 nsew signal input
rlabel locali s 17 823 136 889 6 S[1]
port 10 nsew signal input
rlabel locali s 2348 199 2467 265 6 S[2]
port 11 nsew signal input
rlabel locali s 2348 823 2467 889 6 S[3]
port 12 nsew signal input
rlabel locali s 2501 199 2620 265 6 S[4]
port 13 nsew signal input
rlabel locali s 2501 823 2620 889 6 S[5]
port 14 nsew signal input
rlabel locali s 4832 199 4951 265 6 S[6]
port 15 nsew signal input
rlabel locali s 4832 823 4951 889 6 S[7]
port 16 nsew signal input
rlabel metal1 s 4465 728 4523 737 6 Z
port 17 nsew signal output
rlabel metal1 s 4465 691 4523 700 6 Z
port 17 nsew signal output
rlabel metal1 s 4465 388 4523 397 6 Z
port 17 nsew signal output
rlabel metal1 s 4465 351 4523 360 6 Z
port 17 nsew signal output
rlabel metal1 s 4277 728 4335 737 6 Z
port 17 nsew signal output
rlabel metal1 s 4277 691 4335 700 6 Z
port 17 nsew signal output
rlabel metal1 s 4277 388 4335 397 6 Z
port 17 nsew signal output
rlabel metal1 s 4277 351 4335 360 6 Z
port 17 nsew signal output
rlabel metal1 s 3117 728 3175 737 6 Z
port 17 nsew signal output
rlabel metal1 s 3117 691 3175 700 6 Z
port 17 nsew signal output
rlabel metal1 s 3117 388 3175 397 6 Z
port 17 nsew signal output
rlabel metal1 s 3117 351 3175 360 6 Z
port 17 nsew signal output
rlabel metal1 s 2929 728 2987 737 6 Z
port 17 nsew signal output
rlabel metal1 s 2929 691 2987 700 6 Z
port 17 nsew signal output
rlabel metal1 s 2929 388 2987 397 6 Z
port 17 nsew signal output
rlabel metal1 s 2929 351 2987 360 6 Z
port 17 nsew signal output
rlabel metal1 s 1981 728 2039 737 6 Z
port 17 nsew signal output
rlabel metal1 s 1981 691 2039 700 6 Z
port 17 nsew signal output
rlabel metal1 s 1981 388 2039 397 6 Z
port 17 nsew signal output
rlabel metal1 s 1981 351 2039 360 6 Z
port 17 nsew signal output
rlabel metal1 s 1793 728 1851 737 6 Z
port 17 nsew signal output
rlabel metal1 s 1793 691 1851 700 6 Z
port 17 nsew signal output
rlabel metal1 s 1793 388 1851 397 6 Z
port 17 nsew signal output
rlabel metal1 s 1793 351 1851 360 6 Z
port 17 nsew signal output
rlabel metal1 s 633 728 691 737 6 Z
port 17 nsew signal output
rlabel metal1 s 633 691 691 700 6 Z
port 17 nsew signal output
rlabel metal1 s 633 388 691 397 6 Z
port 17 nsew signal output
rlabel metal1 s 633 351 691 360 6 Z
port 17 nsew signal output
rlabel metal1 s 445 728 503 737 6 Z
port 17 nsew signal output
rlabel metal1 s 445 700 4523 728 6 Z
port 17 nsew signal output
rlabel metal1 s 445 691 503 700 6 Z
port 17 nsew signal output
rlabel metal1 s 445 388 503 397 6 Z
port 17 nsew signal output
rlabel metal1 s 445 360 4523 388 6 Z
port 17 nsew signal output
rlabel metal1 s 445 351 503 360 6 Z
port 17 nsew signal output
rlabel metal1 s 0 1040 4968 1136 6 VGND
port 18 nsew ground bidirectional
rlabel metal1 s 0 -48 4968 48 8 VGND
port 18 nsew ground bidirectional
rlabel metal1 s 0 496 4968 592 6 VPWR
port 19 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 4968 1088
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2964294
string GDS_START 2893498
<< end >>
