magic
tech sky130A
magscale 1 2
timestamp 1601050056
<< nwell >>
rect -38 332 1862 704
<< pwell >>
rect 0 0 1824 49
<< scpmos >>
rect 83 368 119 536
rect 173 368 209 536
rect 263 368 299 536
rect 353 368 389 536
rect 479 368 515 592
rect 569 368 605 592
rect 1006 368 1042 592
rect 1131 368 1167 592
rect 1221 368 1257 592
rect 1345 368 1381 592
rect 1435 368 1471 592
rect 1525 368 1561 592
rect 1615 368 1651 592
rect 1705 368 1741 592
<< nmoslvt >>
rect 84 74 114 202
rect 184 74 214 202
rect 270 74 300 202
rect 370 74 400 202
rect 568 74 598 222
rect 668 74 698 222
rect 787 74 817 222
rect 873 74 903 222
rect 973 74 1003 222
rect 1091 74 1121 222
rect 1177 74 1207 222
rect 1295 74 1325 222
rect 1381 74 1411 222
rect 1506 74 1536 222
rect 1592 74 1622 222
rect 1710 74 1740 222
<< ndiff >>
rect 27 190 84 202
rect 27 156 39 190
rect 73 156 84 190
rect 27 120 84 156
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 133 184 202
rect 114 99 125 133
rect 159 99 184 133
rect 114 74 184 99
rect 214 190 270 202
rect 214 156 225 190
rect 259 156 270 190
rect 214 120 270 156
rect 214 86 225 120
rect 259 86 270 120
rect 214 74 270 86
rect 300 189 370 202
rect 300 155 325 189
rect 359 155 370 189
rect 300 74 370 155
rect 400 120 457 202
rect 400 86 411 120
rect 445 86 457 120
rect 400 74 457 86
rect 511 136 568 222
rect 511 102 523 136
rect 557 102 568 136
rect 511 74 568 102
rect 598 189 668 222
rect 598 155 623 189
rect 657 155 668 189
rect 598 74 668 155
rect 698 136 787 222
rect 698 102 723 136
rect 757 102 787 136
rect 698 74 787 102
rect 817 189 873 222
rect 817 155 828 189
rect 862 155 873 189
rect 817 74 873 155
rect 903 136 973 222
rect 903 102 928 136
rect 962 102 973 136
rect 903 74 973 102
rect 1003 84 1091 222
rect 1003 74 1030 84
rect 1018 50 1030 74
rect 1064 74 1091 84
rect 1121 136 1177 222
rect 1121 102 1132 136
rect 1166 102 1177 136
rect 1121 74 1177 102
rect 1207 84 1295 222
rect 1207 74 1234 84
rect 1064 50 1076 74
rect 1018 38 1076 50
rect 1222 50 1234 74
rect 1268 74 1295 84
rect 1325 136 1381 222
rect 1325 102 1336 136
rect 1370 102 1381 136
rect 1325 74 1381 102
rect 1411 84 1506 222
rect 1411 74 1441 84
rect 1268 50 1280 74
rect 1222 38 1280 50
rect 1426 50 1441 74
rect 1475 74 1506 84
rect 1536 136 1592 222
rect 1536 102 1547 136
rect 1581 102 1592 136
rect 1536 74 1592 102
rect 1622 84 1710 222
rect 1622 74 1649 84
rect 1475 50 1491 74
rect 1426 38 1491 50
rect 1637 50 1649 74
rect 1683 74 1710 84
rect 1740 210 1797 222
rect 1740 176 1751 210
rect 1785 176 1797 210
rect 1740 120 1797 176
rect 1740 86 1751 120
rect 1785 86 1797 120
rect 1740 74 1797 86
rect 1683 50 1695 74
rect 1637 38 1695 50
<< pdiff >>
rect 404 627 464 639
rect 404 593 417 627
rect 451 593 464 627
rect 620 627 678 639
rect 404 592 464 593
rect 620 593 632 627
rect 666 593 678 627
rect 1057 627 1116 639
rect 620 592 678 593
rect 1057 593 1069 627
rect 1103 593 1116 627
rect 1272 627 1330 639
rect 1057 592 1116 593
rect 1272 593 1284 627
rect 1318 593 1330 627
rect 1272 592 1330 593
rect 404 536 479 592
rect 27 524 83 536
rect 27 490 39 524
rect 73 490 83 524
rect 27 414 83 490
rect 27 380 39 414
rect 73 380 83 414
rect 27 368 83 380
rect 119 524 173 536
rect 119 490 129 524
rect 163 490 173 524
rect 119 414 173 490
rect 119 380 129 414
rect 163 380 173 414
rect 119 368 173 380
rect 209 516 263 536
rect 209 482 219 516
rect 253 482 263 516
rect 209 368 263 482
rect 299 524 353 536
rect 299 490 309 524
rect 343 490 353 524
rect 299 440 353 490
rect 299 406 309 440
rect 343 406 353 440
rect 299 368 353 406
rect 389 368 479 536
rect 515 491 569 592
rect 515 457 525 491
rect 559 457 569 491
rect 515 368 569 457
rect 605 368 678 592
rect 950 577 1006 592
rect 950 543 962 577
rect 996 543 1006 577
rect 950 368 1006 543
rect 1042 368 1131 592
rect 1167 577 1221 592
rect 1167 543 1177 577
rect 1211 543 1221 577
rect 1167 368 1221 543
rect 1257 368 1345 592
rect 1381 577 1435 592
rect 1381 543 1391 577
rect 1425 543 1435 577
rect 1381 368 1435 543
rect 1471 531 1525 592
rect 1471 497 1481 531
rect 1515 497 1525 531
rect 1471 437 1525 497
rect 1471 403 1481 437
rect 1515 403 1525 437
rect 1471 368 1525 403
rect 1561 580 1615 592
rect 1561 546 1571 580
rect 1605 546 1615 580
rect 1561 505 1615 546
rect 1561 471 1571 505
rect 1605 471 1615 505
rect 1561 368 1615 471
rect 1651 531 1705 592
rect 1651 497 1661 531
rect 1695 497 1705 531
rect 1651 437 1705 497
rect 1651 403 1661 437
rect 1695 403 1705 437
rect 1651 368 1705 403
rect 1741 580 1797 592
rect 1741 546 1751 580
rect 1785 546 1797 580
rect 1741 508 1797 546
rect 1741 474 1751 508
rect 1785 474 1797 508
rect 1741 437 1797 474
rect 1741 403 1751 437
rect 1785 403 1797 437
rect 1741 368 1797 403
<< ndiffc >>
rect 39 156 73 190
rect 39 86 73 120
rect 125 99 159 133
rect 225 156 259 190
rect 225 86 259 120
rect 325 155 359 189
rect 411 86 445 120
rect 523 102 557 136
rect 623 155 657 189
rect 723 102 757 136
rect 828 155 862 189
rect 928 102 962 136
rect 1030 50 1064 84
rect 1132 102 1166 136
rect 1234 50 1268 84
rect 1336 102 1370 136
rect 1441 50 1475 84
rect 1547 102 1581 136
rect 1649 50 1683 84
rect 1751 176 1785 210
rect 1751 86 1785 120
<< pdiffc >>
rect 417 593 451 627
rect 632 593 666 627
rect 1069 593 1103 627
rect 1284 593 1318 627
rect 39 490 73 524
rect 39 380 73 414
rect 129 490 163 524
rect 129 380 163 414
rect 219 482 253 516
rect 309 490 343 524
rect 309 406 343 440
rect 525 457 559 491
rect 962 543 996 577
rect 1177 543 1211 577
rect 1391 543 1425 577
rect 1481 497 1515 531
rect 1481 403 1515 437
rect 1571 546 1605 580
rect 1571 471 1605 505
rect 1661 497 1695 531
rect 1661 403 1695 437
rect 1751 546 1785 580
rect 1751 474 1785 508
rect 1751 403 1785 437
<< poly >>
rect 479 592 515 618
rect 569 592 605 618
rect 1006 592 1042 618
rect 1131 592 1167 618
rect 1221 592 1257 618
rect 1345 592 1381 618
rect 1435 592 1471 618
rect 1525 592 1561 618
rect 1615 592 1651 618
rect 1705 592 1741 618
rect 83 536 119 562
rect 173 536 209 562
rect 263 536 299 562
rect 353 536 389 562
rect 716 575 918 591
rect 716 541 732 575
rect 766 541 800 575
rect 834 541 868 575
rect 902 541 918 575
rect 716 525 918 541
rect 83 330 119 368
rect 173 330 209 368
rect 83 314 209 330
rect 83 280 125 314
rect 159 294 209 314
rect 263 336 299 368
rect 353 336 389 368
rect 479 336 515 368
rect 569 336 605 368
rect 787 336 817 525
rect 1006 336 1042 368
rect 1131 336 1167 368
rect 263 320 431 336
rect 159 280 214 294
rect 83 264 214 280
rect 263 286 313 320
rect 347 286 381 320
rect 415 286 431 320
rect 263 270 431 286
rect 479 320 817 336
rect 479 286 495 320
rect 529 286 563 320
rect 597 286 631 320
rect 665 286 699 320
rect 733 286 767 320
rect 801 300 817 320
rect 965 320 1167 336
rect 801 286 903 300
rect 479 270 903 286
rect 965 286 981 320
rect 1015 286 1049 320
rect 1083 286 1117 320
rect 1151 315 1167 320
rect 1221 345 1257 368
rect 1345 345 1381 368
rect 1221 315 1381 345
rect 1435 336 1471 368
rect 1525 336 1561 368
rect 1615 336 1651 368
rect 1429 320 1651 336
rect 1151 286 1325 315
rect 965 285 1325 286
rect 965 270 1207 285
rect 84 202 114 264
rect 184 202 214 264
rect 270 202 300 270
rect 370 202 400 270
rect 568 222 598 270
rect 668 222 698 270
rect 787 222 817 270
rect 873 222 903 270
rect 973 222 1003 270
rect 1091 222 1121 270
rect 1177 222 1207 270
rect 1295 222 1325 285
rect 1429 286 1445 320
rect 1479 286 1513 320
rect 1547 286 1581 320
rect 1615 300 1651 320
rect 1705 300 1741 368
rect 1615 286 1741 300
rect 1429 270 1741 286
rect 1429 267 1459 270
rect 1381 237 1459 267
rect 1381 222 1411 237
rect 1506 222 1536 270
rect 1592 222 1622 270
rect 1710 222 1740 270
rect 84 48 114 74
rect 184 48 214 74
rect 270 48 300 74
rect 370 48 400 74
rect 568 48 598 74
rect 668 48 698 74
rect 787 48 817 74
rect 873 48 903 74
rect 973 48 1003 74
rect 1091 48 1121 74
rect 1177 48 1207 74
rect 1295 48 1325 74
rect 1381 48 1411 74
rect 1506 48 1536 74
rect 1592 48 1622 74
rect 1710 48 1740 74
<< polycont >>
rect 732 541 766 575
rect 800 541 834 575
rect 868 541 902 575
rect 125 280 159 314
rect 313 286 347 320
rect 381 286 415 320
rect 495 286 529 320
rect 563 286 597 320
rect 631 286 665 320
rect 699 286 733 320
rect 767 286 801 320
rect 981 286 1015 320
rect 1049 286 1083 320
rect 1117 286 1151 320
rect 1445 286 1479 320
rect 1513 286 1547 320
rect 1581 286 1615 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 23 524 73 649
rect 23 490 39 524
rect 23 414 73 490
rect 23 380 39 414
rect 23 364 73 380
rect 113 524 179 540
rect 113 490 129 524
rect 163 490 179 524
rect 113 424 179 490
rect 219 516 253 649
rect 400 627 468 649
rect 400 593 417 627
rect 451 593 468 627
rect 616 627 682 649
rect 616 593 632 627
rect 666 593 682 627
rect 1053 627 1120 649
rect 716 575 918 591
rect 716 559 732 575
rect 219 458 253 482
rect 293 541 732 559
rect 766 541 800 575
rect 834 541 868 575
rect 902 541 918 575
rect 293 525 918 541
rect 962 577 1012 596
rect 1053 593 1069 627
rect 1103 593 1120 627
rect 1268 627 1334 649
rect 996 559 1012 577
rect 1161 577 1227 596
rect 1268 593 1284 627
rect 1318 593 1334 627
rect 1161 559 1177 577
rect 996 543 1177 559
rect 1211 559 1227 577
rect 1375 581 1801 615
rect 1375 577 1425 581
rect 1375 559 1391 577
rect 1211 543 1391 559
rect 1571 580 1605 581
rect 962 525 1425 543
rect 1465 531 1531 547
rect 293 524 359 525
rect 293 490 309 524
rect 343 490 359 524
rect 1465 497 1481 531
rect 1515 497 1531 531
rect 1465 491 1531 497
rect 293 440 359 490
rect 509 457 525 491
rect 559 457 1531 491
rect 293 424 309 440
rect 113 414 309 424
rect 113 380 129 414
rect 163 406 309 414
rect 343 406 359 440
rect 1465 437 1531 457
rect 1751 580 1801 581
rect 1571 505 1605 546
rect 1571 455 1605 471
rect 1645 531 1711 547
rect 1645 497 1661 531
rect 1695 497 1711 531
rect 163 390 359 406
rect 163 380 179 390
rect 113 364 179 380
rect 397 389 1307 423
rect 217 350 263 356
rect 217 330 223 350
rect 109 316 223 330
rect 257 316 263 350
rect 397 336 431 389
rect 889 350 1167 355
rect 109 314 263 316
rect 109 280 125 314
rect 159 280 263 314
rect 109 264 263 280
rect 297 320 431 336
rect 297 286 313 320
rect 347 286 381 320
rect 415 286 431 320
rect 297 270 431 286
rect 479 320 817 336
rect 479 286 495 320
rect 529 286 563 320
rect 597 286 631 320
rect 665 286 699 320
rect 733 286 767 320
rect 801 286 817 320
rect 479 270 817 286
rect 889 316 895 350
rect 929 320 1167 350
rect 929 316 981 320
rect 889 286 981 316
rect 1015 286 1049 320
rect 1083 286 1117 320
rect 1151 286 1167 320
rect 889 270 1167 286
rect 1273 353 1307 389
rect 1465 403 1481 437
rect 1515 421 1531 437
rect 1645 437 1711 497
rect 1645 421 1661 437
rect 1515 403 1661 421
rect 1695 403 1711 437
rect 1465 387 1711 403
rect 1785 546 1801 580
rect 1751 508 1801 546
rect 1785 474 1801 508
rect 1751 437 1801 474
rect 1785 403 1801 437
rect 1751 387 1801 403
rect 1273 320 1631 353
rect 1273 286 1445 320
rect 1479 286 1513 320
rect 1547 286 1581 320
rect 1615 286 1631 320
rect 1273 270 1631 286
rect 479 236 513 270
rect 1665 236 1699 387
rect 23 196 275 230
rect 23 190 73 196
rect 23 156 39 190
rect 209 190 275 196
rect 23 120 73 156
rect 23 86 39 120
rect 23 70 73 86
rect 109 133 175 162
rect 109 99 125 133
rect 159 99 175 133
rect 109 17 175 99
rect 209 156 225 190
rect 259 156 275 190
rect 209 120 275 156
rect 309 202 513 236
rect 607 202 1699 236
rect 1735 210 1801 226
rect 309 189 375 202
rect 309 155 325 189
rect 359 155 375 189
rect 607 189 673 202
rect 309 154 375 155
rect 507 136 573 168
rect 209 86 225 120
rect 259 86 411 120
rect 445 86 461 120
rect 209 70 461 86
rect 507 102 523 136
rect 557 102 573 136
rect 607 155 623 189
rect 657 155 673 189
rect 812 189 878 202
rect 607 119 673 155
rect 707 136 773 168
rect 507 85 573 102
rect 707 102 723 136
rect 757 102 773 136
rect 812 155 828 189
rect 862 155 878 189
rect 1735 176 1751 210
rect 1785 176 1801 210
rect 1735 168 1801 176
rect 812 119 878 155
rect 912 136 1801 168
rect 707 85 773 102
rect 912 102 928 136
rect 962 134 1132 136
rect 962 102 978 134
rect 912 85 978 102
rect 1116 102 1132 134
rect 1166 134 1336 136
rect 1166 102 1182 134
rect 507 51 978 85
rect 1014 84 1080 100
rect 1014 50 1030 84
rect 1064 50 1080 84
rect 1116 70 1182 102
rect 1320 102 1336 134
rect 1370 134 1547 136
rect 1370 102 1386 134
rect 1218 84 1284 100
rect 1014 17 1080 50
rect 1218 50 1234 84
rect 1268 50 1284 84
rect 1320 70 1386 102
rect 1531 102 1547 134
rect 1581 134 1801 136
rect 1581 102 1597 134
rect 1422 84 1495 100
rect 1218 17 1284 50
rect 1422 50 1441 84
rect 1475 50 1495 84
rect 1531 70 1597 102
rect 1735 120 1801 134
rect 1633 84 1699 100
rect 1422 17 1495 50
rect 1633 50 1649 84
rect 1683 50 1699 84
rect 1735 86 1751 120
rect 1785 86 1801 120
rect 1735 70 1801 86
rect 1633 17 1699 50
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 223 316 257 350
rect 895 316 929 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
<< metal1 >>
rect 0 683 1824 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 0 617 1824 649
rect 211 350 269 356
rect 211 316 223 350
rect 257 347 269 350
rect 883 350 941 356
rect 883 347 895 350
rect 257 319 895 347
rect 257 316 269 319
rect 211 310 269 316
rect 883 316 895 319
rect 929 316 941 350
rect 883 310 941 316
rect 0 17 1824 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
rect 0 -49 1824 -17
<< labels >>
flabel pwell s 0 0 1824 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 0 617 1824 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
rlabel comment s 0 0 0 0 4 xnor2_4
flabel comment s 797 440 797 440 0 FreeSans 200 0 0 0 no_jumper_check
flabel metal1 s 0 617 1824 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 1824 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 1471 390 1505 424 0 FreeSans 340 0 0 0 Y
port 7 nsew
flabel corelocali s 1279 316 1313 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 1375 316 1409 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 1471 316 1505 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 1567 316 1601 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 A
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 1824 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 440604
string GDS_START 428126
<< end >>
