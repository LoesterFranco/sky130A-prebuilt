magic
tech sky130A
magscale 1 2
timestamp 1604502710
<< nwell >>
rect -38 335 2918 704
rect -38 332 732 335
rect 1210 332 2918 335
rect 1624 311 1956 332
<< pwell >>
rect 0 0 2880 49
<< scpmos >>
rect 83 464 119 592
rect 307 483 343 611
rect 389 483 425 611
rect 481 483 517 611
rect 589 483 625 611
rect 683 483 719 611
rect 911 387 947 611
rect 1001 387 1037 611
rect 1209 457 1245 541
rect 1303 457 1339 541
rect 1383 457 1419 541
rect 1508 457 1544 541
rect 1710 347 1746 547
rect 1834 366 1870 566
rect 2004 508 2040 592
rect 2082 508 2118 592
rect 2252 508 2288 592
rect 2342 508 2378 592
rect 2459 392 2495 592
rect 2661 368 2697 592
rect 2751 368 2787 592
<< nmoslvt >>
rect 84 74 114 158
rect 282 81 312 165
rect 360 81 390 165
rect 517 81 547 165
rect 595 81 625 165
rect 688 81 718 165
rect 893 119 923 267
rect 1007 119 1037 267
rect 1205 119 1235 203
rect 1324 119 1354 203
rect 1402 119 1432 203
rect 1480 119 1510 203
rect 1693 74 1723 222
rect 1794 74 1824 222
rect 2048 74 2078 158
rect 2126 74 2156 158
rect 2212 74 2242 158
rect 2284 74 2314 158
rect 2482 74 2512 202
rect 2680 74 2710 222
rect 2766 74 2796 222
<< ndiff >>
rect 843 234 893 267
rect 837 169 893 234
rect 27 133 84 158
rect 27 99 39 133
rect 73 99 84 133
rect 27 74 84 99
rect 114 128 171 158
rect 114 94 125 128
rect 159 94 171 128
rect 114 74 171 94
rect 225 127 282 165
rect 225 93 237 127
rect 271 93 282 127
rect 225 81 282 93
rect 312 81 360 165
rect 390 153 517 165
rect 390 119 471 153
rect 505 119 517 153
rect 390 81 517 119
rect 547 81 595 165
rect 625 140 688 165
rect 625 106 643 140
rect 677 106 688 140
rect 625 81 688 106
rect 718 140 783 165
rect 718 106 741 140
rect 775 106 783 140
rect 837 135 845 169
rect 879 135 893 169
rect 837 119 893 135
rect 923 134 1007 267
rect 923 119 948 134
rect 718 81 783 106
rect 938 100 948 119
rect 982 119 1007 134
rect 1037 239 1091 267
rect 1037 205 1047 239
rect 1081 205 1091 239
rect 1037 165 1091 205
rect 1525 203 1693 222
rect 1037 131 1047 165
rect 1081 131 1091 165
rect 1037 119 1091 131
rect 1145 180 1205 203
rect 1145 146 1160 180
rect 1194 146 1205 180
rect 1145 119 1205 146
rect 1235 179 1324 203
rect 1235 145 1279 179
rect 1313 145 1324 179
rect 1235 119 1324 145
rect 1354 119 1402 203
rect 1432 119 1480 203
rect 1510 119 1693 203
rect 982 100 992 119
rect 938 84 992 100
rect 1525 82 1693 119
rect 1525 48 1551 82
rect 1585 74 1693 82
rect 1723 189 1794 222
rect 1723 155 1734 189
rect 1768 155 1794 189
rect 1723 74 1794 155
rect 1824 158 1874 222
rect 2623 210 2680 222
rect 1824 146 2048 158
rect 1824 112 1902 146
rect 1936 112 2003 146
rect 2037 112 2048 146
rect 1824 74 2048 112
rect 2078 74 2126 158
rect 2156 133 2212 158
rect 2156 99 2167 133
rect 2201 99 2212 133
rect 2156 74 2212 99
rect 2242 74 2284 158
rect 2314 133 2371 158
rect 2314 99 2325 133
rect 2359 99 2371 133
rect 2314 74 2371 99
rect 2425 120 2482 202
rect 2425 86 2437 120
rect 2471 86 2482 120
rect 2425 74 2482 86
rect 2512 190 2569 202
rect 2512 156 2523 190
rect 2557 156 2569 190
rect 2512 120 2569 156
rect 2512 86 2523 120
rect 2557 86 2569 120
rect 2512 74 2569 86
rect 2623 176 2635 210
rect 2669 176 2680 210
rect 2623 120 2680 176
rect 2623 86 2635 120
rect 2669 86 2680 120
rect 2623 74 2680 86
rect 2710 210 2766 222
rect 2710 176 2721 210
rect 2755 176 2766 210
rect 2710 120 2766 176
rect 2710 86 2721 120
rect 2755 86 2766 120
rect 2710 74 2766 86
rect 2796 210 2853 222
rect 2796 176 2807 210
rect 2841 176 2853 210
rect 2796 120 2853 176
rect 2796 86 2807 120
rect 2841 86 2853 120
rect 2796 74 2853 86
rect 1585 48 1612 74
rect 1525 36 1612 48
<< pdiff >>
rect 189 599 307 611
rect 189 592 263 599
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 510 83 546
rect 27 476 39 510
rect 73 476 83 510
rect 27 464 83 476
rect 119 580 263 592
rect 119 546 139 580
rect 173 565 263 580
rect 297 565 307 599
rect 173 546 307 565
rect 119 529 307 546
rect 119 510 263 529
rect 119 476 139 510
rect 173 495 263 510
rect 297 495 307 529
rect 173 483 307 495
rect 343 483 389 611
rect 425 599 481 611
rect 425 565 437 599
rect 471 565 481 599
rect 425 529 481 565
rect 425 495 437 529
rect 471 495 481 529
rect 425 483 481 495
rect 517 483 589 611
rect 625 575 683 611
rect 625 541 635 575
rect 669 541 683 575
rect 625 483 683 541
rect 719 599 795 611
rect 719 565 749 599
rect 783 565 795 599
rect 719 529 795 565
rect 719 495 749 529
rect 783 495 795 529
rect 719 483 795 495
rect 173 476 270 483
rect 119 464 270 476
rect 855 439 911 611
rect 855 405 867 439
rect 901 405 911 439
rect 855 387 911 405
rect 947 593 1001 611
rect 947 559 957 593
rect 991 559 1001 593
rect 947 387 1001 559
rect 1037 439 1089 611
rect 1037 405 1047 439
rect 1081 405 1089 439
rect 1037 387 1089 405
rect 1434 582 1493 594
rect 1434 548 1446 582
rect 1480 548 1493 582
rect 1434 541 1493 548
rect 1948 566 2004 592
rect 1761 547 1834 566
rect 1153 516 1209 541
rect 1153 482 1165 516
rect 1199 482 1209 516
rect 1153 457 1209 482
rect 1245 529 1303 541
rect 1245 495 1255 529
rect 1289 495 1303 529
rect 1245 457 1303 495
rect 1339 457 1383 541
rect 1419 457 1508 541
rect 1544 521 1600 541
rect 1544 487 1554 521
rect 1588 487 1600 521
rect 1544 457 1600 487
rect 1654 524 1710 547
rect 1654 490 1666 524
rect 1700 490 1710 524
rect 1654 468 1710 490
rect 1660 347 1710 468
rect 1746 535 1834 547
rect 1746 501 1773 535
rect 1807 501 1834 535
rect 1746 464 1834 501
rect 1746 430 1773 464
rect 1807 430 1834 464
rect 1746 393 1834 430
rect 1746 359 1773 393
rect 1807 366 1834 393
rect 1870 554 2004 566
rect 1870 520 1880 554
rect 1914 520 1960 554
rect 1994 520 2004 554
rect 1870 508 2004 520
rect 2040 508 2082 592
rect 2118 580 2252 592
rect 2118 546 2128 580
rect 2162 546 2198 580
rect 2232 546 2252 580
rect 2118 508 2252 546
rect 2288 567 2342 592
rect 2288 533 2298 567
rect 2332 533 2342 567
rect 2288 508 2342 533
rect 2378 580 2459 592
rect 2378 546 2405 580
rect 2439 546 2459 580
rect 2378 509 2459 546
rect 2378 508 2405 509
rect 1870 486 1925 508
rect 1870 452 1880 486
rect 1914 452 1925 486
rect 1870 418 1925 452
rect 1870 384 1880 418
rect 1914 384 1925 418
rect 1870 366 1925 384
rect 1807 359 1819 366
rect 1746 347 1819 359
rect 2393 475 2405 508
rect 2439 475 2459 509
rect 2393 438 2459 475
rect 2393 404 2405 438
rect 2439 404 2459 438
rect 2393 392 2459 404
rect 2495 580 2551 592
rect 2495 546 2505 580
rect 2539 546 2551 580
rect 2495 509 2551 546
rect 2495 475 2505 509
rect 2539 475 2551 509
rect 2495 438 2551 475
rect 2495 404 2505 438
rect 2539 404 2551 438
rect 2495 392 2551 404
rect 2605 580 2661 592
rect 2605 546 2617 580
rect 2651 546 2661 580
rect 2605 497 2661 546
rect 2605 463 2617 497
rect 2651 463 2661 497
rect 2605 414 2661 463
rect 2605 380 2617 414
rect 2651 380 2661 414
rect 2605 368 2661 380
rect 2697 580 2751 592
rect 2697 546 2707 580
rect 2741 546 2751 580
rect 2697 497 2751 546
rect 2697 463 2707 497
rect 2741 463 2751 497
rect 2697 414 2751 463
rect 2697 380 2707 414
rect 2741 380 2751 414
rect 2697 368 2751 380
rect 2787 580 2853 592
rect 2787 546 2807 580
rect 2841 546 2853 580
rect 2787 497 2853 546
rect 2787 463 2807 497
rect 2841 463 2853 497
rect 2787 414 2853 463
rect 2787 380 2807 414
rect 2841 380 2853 414
rect 2787 368 2853 380
<< ndiffc >>
rect 39 99 73 133
rect 125 94 159 128
rect 237 93 271 127
rect 471 119 505 153
rect 643 106 677 140
rect 741 106 775 140
rect 845 135 879 169
rect 948 100 982 134
rect 1047 205 1081 239
rect 1047 131 1081 165
rect 1160 146 1194 180
rect 1279 145 1313 179
rect 1551 48 1585 82
rect 1734 155 1768 189
rect 1902 112 1936 146
rect 2003 112 2037 146
rect 2167 99 2201 133
rect 2325 99 2359 133
rect 2437 86 2471 120
rect 2523 156 2557 190
rect 2523 86 2557 120
rect 2635 176 2669 210
rect 2635 86 2669 120
rect 2721 176 2755 210
rect 2721 86 2755 120
rect 2807 176 2841 210
rect 2807 86 2841 120
<< pdiffc >>
rect 39 546 73 580
rect 39 476 73 510
rect 139 546 173 580
rect 263 565 297 599
rect 139 476 173 510
rect 263 495 297 529
rect 437 565 471 599
rect 437 495 471 529
rect 635 541 669 575
rect 749 565 783 599
rect 749 495 783 529
rect 867 405 901 439
rect 957 559 991 593
rect 1047 405 1081 439
rect 1446 548 1480 582
rect 1165 482 1199 516
rect 1255 495 1289 529
rect 1554 487 1588 521
rect 1666 490 1700 524
rect 1773 501 1807 535
rect 1773 430 1807 464
rect 1773 359 1807 393
rect 1880 520 1914 554
rect 1960 520 1994 554
rect 2128 546 2162 580
rect 2198 546 2232 580
rect 2298 533 2332 567
rect 2405 546 2439 580
rect 1880 452 1914 486
rect 1880 384 1914 418
rect 2405 475 2439 509
rect 2405 404 2439 438
rect 2505 546 2539 580
rect 2505 475 2539 509
rect 2505 404 2539 438
rect 2617 546 2651 580
rect 2617 463 2651 497
rect 2617 380 2651 414
rect 2707 546 2741 580
rect 2707 463 2741 497
rect 2707 380 2741 414
rect 2807 546 2841 580
rect 2807 463 2841 497
rect 2807 380 2841 414
<< poly >>
rect 83 592 119 618
rect 307 611 343 637
rect 389 611 425 637
rect 481 611 517 637
rect 589 611 625 637
rect 683 611 719 637
rect 911 611 947 637
rect 1001 611 1037 637
rect 1106 615 1870 645
rect 83 367 119 464
rect 307 367 343 483
rect 83 351 343 367
rect 83 317 137 351
rect 171 317 205 351
rect 239 317 273 351
rect 307 317 343 351
rect 83 301 343 317
rect 84 158 114 301
rect 389 253 425 483
rect 481 432 517 483
rect 467 416 533 432
rect 589 430 625 483
rect 683 432 719 483
rect 467 382 483 416
rect 517 382 533 416
rect 467 366 533 382
rect 575 414 641 430
rect 575 380 591 414
rect 625 380 641 414
rect 575 346 641 380
rect 162 237 228 253
rect 162 203 178 237
rect 212 217 228 237
rect 354 237 425 253
rect 467 302 533 318
rect 467 268 483 302
rect 517 268 533 302
rect 575 312 591 346
rect 625 312 641 346
rect 575 296 641 312
rect 683 416 823 432
rect 683 382 773 416
rect 807 382 823 416
rect 1106 439 1138 615
rect 1209 541 1245 567
rect 1303 541 1339 615
rect 1383 541 1419 567
rect 1508 541 1544 567
rect 1710 547 1746 573
rect 1834 566 1870 615
rect 2004 592 2040 618
rect 2082 592 2118 618
rect 2252 592 2288 618
rect 2342 592 2378 618
rect 2459 592 2495 618
rect 2661 592 2697 618
rect 2751 592 2787 618
rect 683 366 823 382
rect 467 252 533 268
rect 212 203 312 217
rect 162 187 312 203
rect 354 203 370 237
rect 404 203 425 237
rect 354 187 425 203
rect 503 210 533 252
rect 282 165 312 187
rect 360 165 390 187
rect 503 180 547 210
rect 517 165 547 180
rect 595 165 625 296
rect 683 215 713 366
rect 911 355 947 387
rect 1001 372 1037 387
rect 879 339 947 355
rect 879 322 895 339
rect 755 306 895 322
rect 755 272 771 306
rect 805 305 895 306
rect 929 305 947 339
rect 805 282 947 305
rect 993 339 1059 372
rect 993 305 1009 339
rect 1043 312 1059 339
rect 1106 312 1136 439
rect 1209 393 1245 457
rect 1303 431 1339 457
rect 1383 415 1419 457
rect 1508 425 1544 457
rect 1383 399 1466 415
rect 1180 377 1246 393
rect 1180 343 1196 377
rect 1230 357 1246 377
rect 1383 365 1416 399
rect 1450 365 1466 399
rect 1230 343 1332 357
rect 1383 349 1466 365
rect 1508 409 1628 425
rect 1508 375 1578 409
rect 1612 375 1628 409
rect 1508 359 1628 375
rect 1180 316 1332 343
rect 1043 305 1136 312
rect 993 282 1136 305
rect 805 272 821 282
rect 755 256 821 272
rect 893 267 923 282
rect 1007 267 1037 282
rect 683 180 718 215
rect 688 165 718 180
rect 893 93 923 119
rect 1106 248 1136 282
rect 1294 301 1332 316
rect 1294 271 1354 301
rect 1106 218 1235 248
rect 1205 203 1235 218
rect 1324 203 1354 271
rect 1402 203 1432 349
rect 1514 267 1544 359
rect 2004 466 2040 508
rect 1957 450 2040 466
rect 1957 416 1973 450
rect 2007 416 2040 450
rect 2082 476 2118 508
rect 2082 460 2170 476
rect 2082 446 2120 460
rect 1957 400 2040 416
rect 2088 426 2120 446
rect 2154 426 2170 460
rect 2252 447 2288 508
rect 2088 392 2170 426
rect 2222 431 2288 447
rect 2222 411 2238 431
rect 1710 315 1746 347
rect 1834 345 1870 366
rect 2088 358 2120 392
rect 2154 358 2170 392
rect 1834 315 2040 345
rect 1480 237 1544 267
rect 1618 299 1746 315
rect 1618 265 1634 299
rect 1668 285 1746 299
rect 1668 265 1723 285
rect 1618 249 1723 265
rect 1480 203 1510 237
rect 1693 222 1723 249
rect 1794 251 1962 267
rect 1794 237 1912 251
rect 1794 222 1824 237
rect 1007 93 1037 119
rect 1205 93 1235 119
rect 1324 93 1354 119
rect 1402 93 1432 119
rect 84 48 114 74
rect 282 55 312 81
rect 360 55 390 81
rect 517 55 547 81
rect 595 55 625 81
rect 688 51 718 81
rect 1480 51 1510 119
rect 688 21 1510 51
rect 1896 217 1912 237
rect 1946 217 1962 251
rect 1896 201 1962 217
rect 2010 226 2040 315
rect 2088 324 2170 358
rect 2088 290 2120 324
rect 2154 290 2170 324
rect 2088 274 2170 290
rect 2212 397 2238 411
rect 2272 397 2288 431
rect 2212 381 2288 397
rect 2010 196 2078 226
rect 2048 158 2078 196
rect 2126 158 2156 274
rect 2212 158 2242 381
rect 2342 333 2378 508
rect 2348 285 2378 333
rect 2459 285 2495 392
rect 2661 326 2697 368
rect 2751 326 2787 368
rect 2312 269 2495 285
rect 2312 249 2328 269
rect 2284 235 2328 249
rect 2362 249 2495 269
rect 2605 310 2787 326
rect 2605 276 2621 310
rect 2655 290 2787 310
rect 2655 276 2796 290
rect 2605 260 2796 276
rect 2362 235 2512 249
rect 2284 219 2512 235
rect 2680 222 2710 260
rect 2766 222 2796 260
rect 2284 158 2314 219
rect 2482 202 2512 219
rect 1693 48 1723 74
rect 1794 48 1824 74
rect 2048 48 2078 74
rect 2126 48 2156 74
rect 2212 48 2242 74
rect 2284 48 2314 74
rect 2482 48 2512 74
rect 2680 48 2710 74
rect 2766 48 2796 74
<< polycont >>
rect 137 317 171 351
rect 205 317 239 351
rect 273 317 307 351
rect 483 382 517 416
rect 591 380 625 414
rect 178 203 212 237
rect 483 268 517 302
rect 591 312 625 346
rect 773 382 807 416
rect 370 203 404 237
rect 771 272 805 306
rect 895 305 929 339
rect 1009 305 1043 339
rect 1196 343 1230 377
rect 1416 365 1450 399
rect 1578 375 1612 409
rect 1973 416 2007 450
rect 2120 426 2154 460
rect 2120 358 2154 392
rect 1634 265 1668 299
rect 1912 217 1946 251
rect 2120 290 2154 324
rect 2238 397 2272 431
rect 2328 235 2362 269
rect 2621 276 2655 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2880 683
rect 123 599 313 649
rect 23 580 89 596
rect 23 546 39 580
rect 73 546 89 580
rect 23 510 89 546
rect 23 476 39 510
rect 73 476 89 510
rect 23 435 89 476
rect 123 580 263 599
rect 123 546 139 580
rect 173 565 263 580
rect 297 565 313 599
rect 173 546 313 565
rect 123 529 313 546
rect 123 510 263 529
rect 123 476 139 510
rect 173 495 263 510
rect 297 495 313 529
rect 173 476 313 495
rect 123 469 313 476
rect 421 599 487 615
rect 421 565 437 599
rect 471 565 487 599
rect 421 529 487 565
rect 619 575 685 649
rect 619 541 635 575
rect 669 541 685 575
rect 619 537 685 541
rect 723 599 799 615
rect 723 565 749 599
rect 783 565 799 599
rect 421 495 437 529
rect 471 503 487 529
rect 723 529 799 565
rect 941 593 1007 649
rect 941 559 957 593
rect 991 559 1007 593
rect 1430 582 1497 649
rect 1430 548 1446 582
rect 1480 548 1497 582
rect 723 503 749 529
rect 471 495 749 503
rect 783 525 799 529
rect 1149 525 1199 545
rect 783 516 1199 525
rect 783 495 1165 516
rect 421 489 1165 495
rect 421 469 799 489
rect 689 466 799 469
rect 1149 482 1165 489
rect 1239 529 1374 545
rect 1430 532 1497 548
rect 1239 495 1255 529
rect 1289 498 1374 529
rect 1538 521 1604 545
rect 1538 498 1554 521
rect 1289 495 1554 498
rect 23 416 541 435
rect 23 401 483 416
rect 23 253 57 401
rect 475 382 483 401
rect 517 382 541 416
rect 121 351 359 367
rect 475 366 541 382
rect 589 414 655 430
rect 589 380 591 414
rect 625 380 655 414
rect 121 317 137 351
rect 171 317 205 351
rect 239 317 273 351
rect 307 332 359 351
rect 589 346 655 380
rect 307 317 541 332
rect 121 302 541 317
rect 121 298 483 302
rect 475 268 483 298
rect 517 268 541 302
rect 589 312 591 346
rect 625 312 655 346
rect 589 296 655 312
rect 23 237 228 253
rect 23 203 178 237
rect 212 203 228 237
rect 23 187 228 203
rect 313 237 420 253
rect 475 252 541 268
rect 689 262 723 466
rect 1149 461 1199 482
rect 1340 487 1554 495
rect 1588 487 1604 521
rect 1340 464 1604 487
rect 1650 524 1716 649
rect 2112 580 2248 649
rect 1864 554 2078 570
rect 1650 490 1666 524
rect 1700 490 1716 524
rect 1650 464 1716 490
rect 1750 535 1823 551
rect 1750 501 1773 535
rect 1807 501 1823 535
rect 1750 464 1823 501
rect 867 439 917 455
rect 757 424 833 432
rect 757 416 799 424
rect 757 382 773 416
rect 807 382 833 390
rect 901 423 917 439
rect 1031 439 1115 455
rect 901 405 997 423
rect 867 389 997 405
rect 1031 405 1047 439
rect 1081 405 1115 439
rect 1149 427 1306 461
rect 1031 393 1115 405
rect 1031 389 1233 393
rect 757 366 833 382
rect 963 355 997 389
rect 1077 377 1233 389
rect 879 339 929 355
rect 879 330 895 339
rect 313 203 370 237
rect 404 203 420 237
rect 23 133 73 187
rect 313 162 420 203
rect 575 228 723 262
rect 757 306 895 330
rect 757 272 771 306
rect 805 305 895 306
rect 805 272 929 305
rect 757 252 929 272
rect 963 339 1043 355
rect 963 305 1009 339
rect 963 289 1043 305
rect 1077 343 1196 377
rect 1230 343 1233 377
rect 1077 327 1233 343
rect 575 169 609 228
rect 757 203 844 252
rect 963 218 997 289
rect 1077 244 1124 327
rect 1272 293 1306 427
rect 878 184 997 218
rect 1031 239 1124 244
rect 1031 205 1047 239
rect 1081 205 1124 239
rect 1031 197 1124 205
rect 1158 259 1306 293
rect 1031 184 1084 197
rect 878 169 914 184
rect 454 153 609 169
rect 23 99 39 133
rect 23 70 73 99
rect 109 128 175 153
rect 109 94 125 128
rect 159 94 175 128
rect 109 17 175 94
rect 221 127 287 128
rect 221 93 237 127
rect 271 93 287 127
rect 454 119 471 153
rect 505 119 609 153
rect 643 140 683 156
rect 221 85 287 93
rect 677 106 683 140
rect 643 85 683 106
rect 221 51 683 85
rect 733 140 793 156
rect 733 106 741 140
rect 775 106 793 140
rect 829 135 845 169
rect 879 135 914 169
rect 1034 165 1084 184
rect 829 119 914 135
rect 948 134 1000 150
rect 733 17 793 106
rect 982 100 1000 134
rect 948 17 1000 100
rect 1034 131 1047 165
rect 1081 131 1084 165
rect 1034 93 1084 131
rect 1158 180 1223 259
rect 1340 225 1374 464
rect 1158 146 1160 180
rect 1194 146 1223 180
rect 1158 130 1223 146
rect 1263 191 1374 225
rect 1408 399 1463 415
rect 1408 365 1416 399
rect 1450 365 1463 399
rect 1408 218 1463 365
rect 1497 315 1531 464
rect 1750 430 1773 464
rect 1807 430 1823 464
rect 1565 424 1703 430
rect 1565 409 1663 424
rect 1565 375 1578 409
rect 1612 390 1663 409
rect 1697 390 1703 424
rect 1612 375 1703 390
rect 1565 359 1703 375
rect 1750 393 1823 430
rect 1750 359 1773 393
rect 1807 359 1823 393
rect 1864 520 1880 554
rect 1914 520 1960 554
rect 1994 520 2078 554
rect 2112 546 2128 580
rect 2162 546 2198 580
rect 2232 546 2248 580
rect 2282 567 2348 596
rect 1864 504 2078 520
rect 2282 533 2298 567
rect 2332 533 2348 567
rect 2282 512 2348 533
rect 1864 486 1920 504
rect 1864 452 1880 486
rect 1914 452 1920 486
rect 1864 418 1920 452
rect 1864 384 1880 418
rect 1914 384 1920 418
rect 1864 368 1920 384
rect 1957 450 2010 466
rect 1957 416 1973 450
rect 2007 416 2010 450
rect 1750 343 1823 359
rect 1497 299 1684 315
rect 1497 265 1634 299
rect 1668 265 1684 299
rect 1497 252 1684 265
rect 1750 226 1784 343
rect 1957 267 2010 416
rect 1718 218 1784 226
rect 1263 179 1329 191
rect 1408 189 1784 218
rect 1408 184 1734 189
rect 1263 145 1279 179
rect 1313 145 1329 179
rect 1718 155 1734 184
rect 1768 155 1784 189
rect 1263 129 1329 145
rect 1403 116 1684 150
rect 1718 119 1784 155
rect 1818 251 2010 267
rect 1818 217 1912 251
rect 1946 217 2010 251
rect 1818 201 2010 217
rect 2044 240 2078 504
rect 2112 478 2348 512
rect 2389 580 2455 649
rect 2389 546 2405 580
rect 2439 546 2455 580
rect 2389 509 2455 546
rect 2112 460 2170 478
rect 2112 426 2120 460
rect 2154 426 2170 460
rect 2389 475 2405 509
rect 2439 475 2455 509
rect 2112 392 2170 426
rect 2112 358 2120 392
rect 2154 358 2170 392
rect 2222 431 2288 444
rect 2222 397 2238 431
rect 2272 424 2288 431
rect 2222 390 2239 397
rect 2273 390 2288 424
rect 2222 384 2288 390
rect 2389 438 2455 475
rect 2389 404 2405 438
rect 2439 404 2455 438
rect 2389 388 2455 404
rect 2489 580 2555 596
rect 2489 546 2505 580
rect 2539 546 2555 580
rect 2489 509 2555 546
rect 2489 475 2505 509
rect 2539 475 2555 509
rect 2489 438 2555 475
rect 2489 404 2505 438
rect 2539 404 2555 438
rect 2489 388 2555 404
rect 2112 350 2170 358
rect 2112 324 2446 350
rect 2112 290 2120 324
rect 2154 316 2446 324
rect 2154 290 2170 316
rect 2112 274 2170 290
rect 2204 269 2378 282
rect 2204 240 2328 269
rect 2044 235 2328 240
rect 2362 235 2378 269
rect 2044 222 2378 235
rect 2044 206 2238 222
rect 1403 93 1451 116
rect 1034 53 1451 93
rect 1650 85 1684 116
rect 1818 85 1852 201
rect 2044 162 2078 206
rect 2412 188 2446 316
rect 1886 146 2078 162
rect 1886 112 1902 146
rect 1936 112 2003 146
rect 2037 112 2078 146
rect 1886 96 2078 112
rect 2151 133 2217 162
rect 2151 99 2167 133
rect 2201 99 2217 133
rect 1521 48 1551 82
rect 1585 48 1616 82
rect 1650 51 1852 85
rect 1521 17 1616 48
rect 2151 17 2217 99
rect 2309 154 2446 188
rect 2521 326 2555 388
rect 2601 580 2667 649
rect 2601 546 2617 580
rect 2651 546 2667 580
rect 2601 497 2667 546
rect 2601 463 2617 497
rect 2651 463 2667 497
rect 2601 414 2667 463
rect 2601 380 2617 414
rect 2651 380 2667 414
rect 2601 364 2667 380
rect 2705 580 2757 596
rect 2705 546 2707 580
rect 2741 546 2757 580
rect 2705 497 2757 546
rect 2705 463 2707 497
rect 2741 463 2757 497
rect 2705 414 2757 463
rect 2705 380 2707 414
rect 2741 380 2757 414
rect 2521 310 2671 326
rect 2521 276 2621 310
rect 2655 276 2671 310
rect 2521 260 2671 276
rect 2705 282 2757 380
rect 2791 580 2857 649
rect 2791 546 2807 580
rect 2841 546 2857 580
rect 2791 497 2857 546
rect 2791 463 2807 497
rect 2841 463 2857 497
rect 2791 414 2857 463
rect 2791 380 2807 414
rect 2841 380 2857 414
rect 2791 364 2857 380
rect 2521 190 2573 260
rect 2521 156 2523 190
rect 2557 156 2573 190
rect 2309 133 2375 154
rect 2309 99 2325 133
rect 2359 99 2375 133
rect 2521 120 2573 156
rect 2309 70 2375 99
rect 2421 86 2437 120
rect 2471 86 2487 120
rect 2421 17 2487 86
rect 2521 86 2523 120
rect 2557 86 2573 120
rect 2521 70 2573 86
rect 2619 210 2669 226
rect 2619 176 2635 210
rect 2619 120 2669 176
rect 2619 86 2635 120
rect 2619 17 2669 86
rect 2705 210 2771 282
rect 2705 176 2721 210
rect 2755 176 2771 210
rect 2705 120 2771 176
rect 2705 86 2721 120
rect 2755 86 2771 120
rect 2705 70 2771 86
rect 2807 210 2857 226
rect 2841 176 2857 210
rect 2807 120 2857 176
rect 2841 86 2857 120
rect 2807 17 2857 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2880 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 799 416 833 424
rect 799 390 807 416
rect 807 390 833 416
rect 1663 390 1697 424
rect 2239 397 2272 424
rect 2272 397 2273 424
rect 2239 390 2273 397
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
<< metal1 >>
rect 0 683 2880 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2880 683
rect 0 617 2880 649
rect 787 424 845 430
rect 787 390 799 424
rect 833 421 845 424
rect 1651 424 1709 430
rect 1651 421 1663 424
rect 833 393 1663 421
rect 833 390 845 393
rect 787 384 845 390
rect 1651 390 1663 393
rect 1697 421 1709 424
rect 2227 424 2285 430
rect 2227 421 2239 424
rect 1697 393 2239 421
rect 1697 390 1709 393
rect 1651 384 1709 390
rect 2227 390 2239 393
rect 2273 390 2285 424
rect 2227 384 2285 390
rect 0 17 2880 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2880 17
rect 0 -49 2880 -17
<< labels >>
flabel pwell s 0 0 2880 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 0 617 2880 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
rlabel comment s 0 0 0 0 4 sdfrtp_2
flabel comment s 1481 630 1481 630 0 FreeSans 300 0 0 0 no_jumper_check
flabel comment s 1107 36 1107 36 0 FreeSans 300 0 0 0 no_jumper_check
flabel metal1 s 2239 390 2273 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew
flabel metal1 s 0 617 2880 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 2880 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 319 168 353 202 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 SCD
port 4 nsew
flabel corelocali s 607 390 641 424 0 FreeSans 340 0 0 0 SCD
port 4 nsew
flabel corelocali s 799 242 833 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 2719 94 2753 128 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2719 168 2753 202 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2719 242 2753 276 0 FreeSans 340 0 0 0 Q
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 2880 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 210386
string GDS_START 189392
<< end >>
