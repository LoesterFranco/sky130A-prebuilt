magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1104 561
rect 17 309 1086 493
rect 17 171 533 275
rect 567 205 1086 309
rect 17 17 1086 171
rect 0 -17 1104 17
<< metal1 >>
rect 0 496 1104 592
rect 14 428 1090 468
rect 17 416 1087 428
rect 0 -48 1104 48
<< labels >>
rlabel locali s 567 205 1086 309 6 KAPWR
port 1 nsew power bidirectional abutment
rlabel locali s 17 309 1086 493 6 KAPWR
port 1 nsew power bidirectional abutment
rlabel metal1 s 17 416 1087 428 6 KAPWR
port 1 nsew power bidirectional abutment
rlabel metal1 s 14 428 1090 468 6 KAPWR
port 1 nsew power bidirectional abutment
rlabel locali s 17 171 533 275 6 VGND
port 2 nsew ground bidirectional abutment
rlabel locali s 17 17 1086 171 6 VGND
port 2 nsew ground bidirectional abutment
rlabel locali s 0 -17 1104 17 8 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1104 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel locali s 0 527 1104 561 6 VPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 0 496 1104 592 6 VPWR
port 3 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1104 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2277740
string GDS_START 2272624
<< end >>
