magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 2024 561
rect 103 333 169 417
rect 271 333 340 417
rect 442 435 508 527
rect 610 435 676 527
rect 882 333 948 417
rect 1050 333 1116 417
rect 103 299 1116 333
rect 1574 367 1624 527
rect 1758 367 1792 527
rect 1926 299 2007 527
rect 22 215 337 255
rect 371 181 407 299
rect 441 215 708 255
rect 754 215 1076 255
rect 1218 215 1452 255
rect 1658 215 2007 255
rect 103 131 676 181
rect 794 17 828 109
rect 962 17 1028 109
rect 1234 17 1268 109
rect 1402 17 1436 109
rect 1674 17 1708 109
rect 1842 17 1894 109
rect 0 -17 2024 17
<< obsli1 >>
rect 18 451 408 493
rect 18 299 69 451
rect 203 367 237 451
rect 374 401 408 451
rect 542 401 576 485
rect 710 401 760 493
rect 374 367 760 401
rect 798 451 1536 493
rect 798 367 848 451
rect 982 367 1016 451
rect 1150 367 1184 451
rect 1218 333 1284 417
rect 1318 367 1352 451
rect 1386 333 1452 417
rect 1486 367 1536 451
rect 1658 333 1724 493
rect 1826 333 1892 493
rect 1218 299 1892 333
rect 18 93 69 181
rect 710 147 2007 181
rect 710 93 760 147
rect 18 51 760 93
rect 862 51 928 147
rect 1062 51 1196 147
rect 1302 51 1368 147
rect 1470 51 1608 147
rect 1742 51 1808 147
rect 1929 51 2007 147
<< metal1 >>
rect 0 496 2024 592
rect 0 -48 2024 48
<< labels >>
rlabel locali s 1658 215 2007 255 6 A1
port 1 nsew signal input
rlabel locali s 1218 215 1452 255 6 A2
port 2 nsew signal input
rlabel locali s 754 215 1076 255 6 A3
port 3 nsew signal input
rlabel locali s 441 215 708 255 6 B1
port 4 nsew signal input
rlabel locali s 22 215 337 255 6 B2
port 5 nsew signal input
rlabel locali s 1050 333 1116 417 6 Y
port 6 nsew signal output
rlabel locali s 882 333 948 417 6 Y
port 6 nsew signal output
rlabel locali s 371 181 407 299 6 Y
port 6 nsew signal output
rlabel locali s 271 333 340 417 6 Y
port 6 nsew signal output
rlabel locali s 103 333 169 417 6 Y
port 6 nsew signal output
rlabel locali s 103 299 1116 333 6 Y
port 6 nsew signal output
rlabel locali s 103 131 676 181 6 Y
port 6 nsew signal output
rlabel locali s 1842 17 1894 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1674 17 1708 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1402 17 1436 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1234 17 1268 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 962 17 1028 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 794 17 828 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 2024 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 2024 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1926 299 2007 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1758 367 1792 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1574 367 1624 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 610 435 676 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 442 435 508 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 2024 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 2024 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2024 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 895886
string GDS_START 879908
<< end >>
