magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 113 333 189 493
rect 301 337 377 493
rect 301 333 533 337
rect 113 299 533 333
rect 21 215 377 265
rect 479 181 533 299
rect 113 145 533 181
rect 113 51 189 145
rect 301 51 377 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 26 299 79 527
rect 233 367 267 527
rect 421 435 463 527
rect 26 17 79 109
rect 233 17 267 109
rect 421 17 471 110
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
rlabel locali s 21 215 377 265 6 A
port 1 nsew signal input
rlabel locali s 479 181 533 299 6 Y
port 2 nsew signal output
rlabel locali s 301 337 377 493 6 Y
port 2 nsew signal output
rlabel locali s 301 333 533 337 6 Y
port 2 nsew signal output
rlabel locali s 301 51 377 145 6 Y
port 2 nsew signal output
rlabel locali s 113 333 189 493 6 Y
port 2 nsew signal output
rlabel locali s 113 299 533 333 6 Y
port 2 nsew signal output
rlabel locali s 113 145 533 181 6 Y
port 2 nsew signal output
rlabel locali s 113 51 189 145 6 Y
port 2 nsew signal output
rlabel metal1 s 0 -48 552 48 8 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 496 552 592 6 VPWR
port 4 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 552 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2107354
string GDS_START 2102076
<< end >>
