magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 368 561
rect 18 299 82 527
rect 118 265 157 475
rect 193 357 259 493
rect 299 367 350 527
rect 193 301 263 357
rect 30 199 82 265
rect 118 199 195 265
rect 229 225 263 301
rect 301 259 350 331
rect 229 191 333 225
rect 115 17 181 89
rect 299 78 333 191
rect 0 -17 368 17
<< obsli1 >>
rect 18 123 261 157
rect 18 53 76 123
rect 215 62 261 123
<< metal1 >>
rect 0 496 368 592
rect 0 -48 368 48
<< labels >>
rlabel locali s 30 199 82 265 6 A1
port 1 nsew signal input
rlabel locali s 118 265 157 475 6 A2
port 2 nsew signal input
rlabel locali s 118 199 195 265 6 A2
port 2 nsew signal input
rlabel locali s 301 259 350 331 6 B1
port 3 nsew signal input
rlabel locali s 299 78 333 191 6 Y
port 4 nsew signal output
rlabel locali s 229 225 263 301 6 Y
port 4 nsew signal output
rlabel locali s 229 191 333 225 6 Y
port 4 nsew signal output
rlabel locali s 193 357 259 493 6 Y
port 4 nsew signal output
rlabel locali s 193 301 263 357 6 Y
port 4 nsew signal output
rlabel locali s 115 17 181 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 368 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 368 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 299 367 350 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 18 299 82 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 368 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 368 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 368 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1334808
string GDS_START 1330090
<< end >>
