magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 21 236 87 313
rect 189 300 263 366
rect 1254 70 1321 596
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 24 381 90 591
rect 124 415 190 649
rect 231 522 331 591
rect 472 556 541 649
rect 575 581 836 615
rect 575 522 609 581
rect 231 488 609 522
rect 231 415 331 488
rect 24 347 155 381
rect 121 202 155 347
rect 297 354 331 415
rect 365 388 445 454
rect 666 413 768 547
rect 411 379 445 388
rect 297 266 377 354
rect 23 166 155 202
rect 227 200 377 266
rect 23 132 263 166
rect 297 152 377 200
rect 411 345 700 379
rect 23 111 89 132
rect 125 17 191 98
rect 229 85 263 132
rect 411 119 461 345
rect 495 245 594 311
rect 636 294 700 345
rect 495 85 529 245
rect 229 51 529 85
rect 563 17 629 211
rect 663 117 697 294
rect 734 211 768 413
rect 802 357 836 581
rect 894 505 1013 649
rect 1053 471 1131 596
rect 870 405 1131 471
rect 1053 388 1131 405
rect 802 291 868 357
rect 902 261 1063 327
rect 1097 326 1131 388
rect 1165 364 1215 649
rect 902 211 936 261
rect 1097 260 1177 326
rect 1097 227 1131 260
rect 731 161 936 211
rect 663 51 871 117
rect 970 17 1020 227
rect 1056 91 1131 227
rect 1168 17 1218 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
<< metal1 >>
rect 0 683 1344 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 0 617 1344 649
rect 0 17 1344 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
rect 0 -49 1344 -17
<< labels >>
rlabel locali s 21 236 87 313 6 D
port 1 nsew signal input
rlabel locali s 1254 70 1321 596 6 Q
port 2 nsew signal output
rlabel locali s 189 300 263 366 6 GATE_N
port 3 nsew clock input
rlabel metal1 s 0 -49 1344 49 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 617 1344 715 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1344 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 2319528
string GDS_START 2308360
<< end >>
