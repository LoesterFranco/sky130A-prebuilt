magic
tech sky130A
magscale 1 2
timestamp 1601050047
<< nwell >>
rect -38 332 902 704
<< pwell >>
rect 0 0 864 49
<< scpmos >>
rect 124 392 154 592
rect 225 368 255 592
rect 324 368 354 592
rect 424 368 454 592
rect 514 368 544 592
rect 646 368 676 592
rect 748 368 778 592
<< nmoslvt >>
rect 81 94 111 222
rect 176 74 206 222
rect 262 74 292 222
rect 469 100 499 248
rect 555 100 585 248
rect 667 100 697 248
rect 753 100 783 248
<< ndiff >>
rect 27 210 81 222
rect 27 176 36 210
rect 70 176 81 210
rect 27 140 81 176
rect 27 106 36 140
rect 70 106 81 140
rect 27 94 81 106
rect 111 162 176 222
rect 111 128 122 162
rect 156 128 176 162
rect 111 94 176 128
rect 126 74 176 94
rect 206 184 262 222
rect 206 150 217 184
rect 251 150 262 184
rect 206 116 262 150
rect 206 82 217 116
rect 251 82 262 116
rect 206 74 262 82
rect 292 128 342 222
rect 292 116 349 128
rect 292 82 303 116
rect 337 82 349 116
rect 419 112 469 248
rect 292 74 349 82
rect 403 100 469 112
rect 499 236 555 248
rect 499 202 510 236
rect 544 202 555 236
rect 499 100 555 202
rect 585 100 667 248
rect 697 236 753 248
rect 697 202 708 236
rect 742 202 753 236
rect 697 168 753 202
rect 697 134 708 168
rect 742 134 753 168
rect 697 100 753 134
rect 783 220 837 248
rect 783 186 794 220
rect 828 186 837 220
rect 783 146 837 186
rect 783 112 794 146
rect 828 112 837 146
rect 783 100 837 112
rect 403 66 411 100
rect 445 66 454 100
rect 403 54 454 66
rect 600 66 609 100
rect 643 66 652 100
rect 600 54 652 66
<< pdiff >>
rect 65 580 124 592
rect 65 546 77 580
rect 111 546 124 580
rect 65 510 124 546
rect 65 476 77 510
rect 111 476 124 510
rect 65 440 124 476
rect 65 406 77 440
rect 111 406 124 440
rect 65 392 124 406
rect 154 580 225 592
rect 154 546 173 580
rect 207 546 225 580
rect 154 508 225 546
rect 154 474 173 508
rect 207 474 225 508
rect 154 392 225 474
rect 172 368 225 392
rect 255 580 324 592
rect 255 546 272 580
rect 306 546 324 580
rect 255 503 324 546
rect 255 469 272 503
rect 306 469 324 503
rect 255 424 324 469
rect 255 390 272 424
rect 306 390 324 424
rect 255 368 324 390
rect 354 580 424 592
rect 354 546 377 580
rect 411 546 424 580
rect 354 499 424 546
rect 354 465 377 499
rect 411 465 424 499
rect 354 368 424 465
rect 454 580 514 592
rect 454 546 467 580
rect 501 546 514 580
rect 454 503 514 546
rect 454 469 467 503
rect 501 469 514 503
rect 454 424 514 469
rect 454 390 467 424
rect 501 390 514 424
rect 454 368 514 390
rect 544 580 646 592
rect 544 546 574 580
rect 608 546 646 580
rect 544 499 646 546
rect 544 465 574 499
rect 608 465 646 499
rect 544 368 646 465
rect 676 580 748 592
rect 676 546 689 580
rect 723 546 748 580
rect 676 503 748 546
rect 676 469 689 503
rect 723 469 748 503
rect 676 424 748 469
rect 676 390 689 424
rect 723 390 748 424
rect 676 368 748 390
rect 778 580 837 592
rect 778 546 791 580
rect 825 546 837 580
rect 778 503 837 546
rect 778 469 791 503
rect 825 469 837 503
rect 778 424 837 469
rect 778 390 791 424
rect 825 390 837 424
rect 778 368 837 390
<< ndiffc >>
rect 36 176 70 210
rect 36 106 70 140
rect 122 128 156 162
rect 217 150 251 184
rect 217 82 251 116
rect 303 82 337 116
rect 510 202 544 236
rect 708 202 742 236
rect 708 134 742 168
rect 794 186 828 220
rect 794 112 828 146
rect 411 66 445 100
rect 609 66 643 100
<< pdiffc >>
rect 77 546 111 580
rect 77 476 111 510
rect 77 406 111 440
rect 173 546 207 580
rect 173 474 207 508
rect 272 546 306 580
rect 272 469 306 503
rect 272 390 306 424
rect 377 546 411 580
rect 377 465 411 499
rect 467 546 501 580
rect 467 469 501 503
rect 467 390 501 424
rect 574 546 608 580
rect 574 465 608 499
rect 689 546 723 580
rect 689 469 723 503
rect 689 390 723 424
rect 791 546 825 580
rect 791 469 825 503
rect 791 390 825 424
<< poly >>
rect 124 592 154 618
rect 225 592 255 618
rect 324 592 354 618
rect 424 592 454 618
rect 514 592 544 618
rect 646 592 676 618
rect 748 592 778 618
rect 124 377 154 392
rect 121 356 157 377
rect 44 340 157 356
rect 225 353 255 368
rect 324 353 354 368
rect 424 353 454 368
rect 514 353 544 368
rect 646 353 676 368
rect 748 353 778 368
rect 44 306 60 340
rect 94 326 157 340
rect 222 336 258 353
rect 321 336 357 353
rect 421 336 457 353
rect 511 336 547 353
rect 646 336 679 353
rect 745 336 781 353
rect 94 306 111 326
rect 44 290 111 306
rect 81 222 111 290
rect 222 320 357 336
rect 222 286 238 320
rect 272 286 306 320
rect 340 286 357 320
rect 222 267 357 286
rect 405 320 585 336
rect 405 286 421 320
rect 455 286 585 320
rect 405 280 585 286
rect 405 270 499 280
rect 176 237 357 267
rect 469 248 499 270
rect 555 248 585 280
rect 649 320 783 336
rect 649 286 665 320
rect 699 286 733 320
rect 767 286 783 320
rect 649 270 783 286
rect 667 248 697 270
rect 753 248 783 270
rect 176 222 206 237
rect 262 222 292 237
rect 81 68 111 94
rect 176 48 206 74
rect 262 48 292 74
rect 469 74 499 100
rect 555 74 585 100
rect 667 74 697 100
rect 753 74 783 100
<< polycont >>
rect 60 306 94 340
rect 238 286 272 320
rect 306 286 340 320
rect 421 286 455 320
rect 665 286 699 320
rect 733 286 767 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 61 580 127 596
rect 61 546 77 580
rect 111 546 127 580
rect 61 510 127 546
rect 61 476 77 510
rect 111 476 127 510
rect 61 440 127 476
rect 166 580 215 649
rect 166 546 173 580
rect 207 546 215 580
rect 166 508 215 546
rect 166 474 173 508
rect 207 474 215 508
rect 166 458 215 474
rect 252 580 327 596
rect 252 546 272 580
rect 306 546 327 580
rect 252 503 327 546
rect 252 469 272 503
rect 306 469 327 503
rect 61 406 77 440
rect 111 424 127 440
rect 252 424 327 469
rect 361 580 427 649
rect 361 546 377 580
rect 411 546 427 580
rect 361 499 427 546
rect 361 465 377 499
rect 411 465 427 499
rect 361 458 427 465
rect 467 580 517 596
rect 501 546 517 580
rect 467 503 517 546
rect 501 469 517 503
rect 467 424 517 469
rect 558 580 624 649
rect 558 546 574 580
rect 608 546 624 580
rect 558 499 624 546
rect 558 465 574 499
rect 608 465 624 499
rect 558 458 624 465
rect 673 580 739 596
rect 673 546 689 580
rect 723 546 739 580
rect 673 503 739 546
rect 673 469 689 503
rect 723 469 739 503
rect 673 424 739 469
rect 111 406 178 424
rect 61 390 178 406
rect 252 390 272 424
rect 306 390 467 424
rect 501 390 689 424
rect 723 390 739 424
rect 775 580 841 649
rect 775 546 791 580
rect 825 546 841 580
rect 775 503 841 546
rect 775 469 791 503
rect 825 469 841 503
rect 775 424 841 469
rect 775 390 791 424
rect 825 390 841 424
rect 25 340 110 356
rect 25 306 60 340
rect 94 306 110 340
rect 25 290 110 306
rect 144 252 178 390
rect 217 320 359 356
rect 217 286 238 320
rect 272 286 306 320
rect 340 286 359 320
rect 405 320 471 336
rect 405 286 421 320
rect 455 286 471 320
rect 405 270 471 286
rect 405 252 439 270
rect 20 218 439 252
rect 505 236 560 390
rect 601 320 839 356
rect 601 286 665 320
rect 699 286 733 320
rect 767 286 839 320
rect 601 270 839 286
rect 20 210 70 218
rect 20 176 36 210
rect 494 202 510 236
rect 544 202 560 236
rect 594 202 708 236
rect 742 202 758 236
rect 20 140 70 176
rect 20 106 36 140
rect 20 90 70 106
rect 106 162 164 182
rect 106 128 122 162
rect 156 128 164 162
rect 106 17 164 128
rect 201 150 217 184
rect 251 168 421 184
rect 594 168 758 202
rect 251 150 708 168
rect 201 116 251 150
rect 387 134 708 150
rect 742 134 758 168
rect 792 220 844 236
rect 792 186 794 220
rect 828 186 844 220
rect 792 146 844 186
rect 201 82 217 116
rect 201 66 251 82
rect 287 82 303 116
rect 337 82 353 116
rect 792 112 794 146
rect 828 112 844 146
rect 792 100 844 112
rect 287 17 353 82
rect 395 66 411 100
rect 445 66 609 100
rect 643 66 844 100
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel comment s 0 0 0 0 4 nand3b_2
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 B
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 864 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 2083096
string GDS_START 2074966
<< end >>
