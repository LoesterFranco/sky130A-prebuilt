magic
tech sky130A
magscale 1 2
timestamp 1601050047
<< nwell >>
rect -38 332 1382 704
<< pwell >>
rect 0 0 1344 49
<< scpmos >>
rect 86 392 116 592
rect 176 392 206 592
rect 266 392 296 592
rect 359 392 389 592
rect 459 392 489 592
rect 549 392 579 592
rect 726 392 756 592
rect 826 392 856 592
rect 938 368 968 592
rect 1038 368 1068 592
rect 1128 368 1158 592
rect 1218 368 1248 592
<< nmoslvt >>
rect 89 119 119 247
rect 175 119 205 247
rect 261 119 291 247
rect 347 119 377 247
rect 433 119 463 247
rect 519 119 549 247
rect 637 119 667 247
rect 723 119 753 247
rect 935 74 965 222
rect 1027 74 1057 222
rect 1127 74 1157 222
rect 1213 74 1243 222
<< ndiff >>
rect 32 235 89 247
rect 32 201 44 235
rect 78 201 89 235
rect 32 165 89 201
rect 32 131 44 165
rect 78 131 89 165
rect 32 119 89 131
rect 119 166 175 247
rect 119 132 130 166
rect 164 132 175 166
rect 119 119 175 132
rect 205 235 261 247
rect 205 201 216 235
rect 250 201 261 235
rect 205 119 261 201
rect 291 166 347 247
rect 291 132 302 166
rect 336 132 347 166
rect 291 119 347 132
rect 377 235 433 247
rect 377 201 388 235
rect 422 201 433 235
rect 377 165 433 201
rect 377 131 388 165
rect 422 131 433 165
rect 377 119 433 131
rect 463 170 519 247
rect 463 136 474 170
rect 508 136 519 170
rect 463 119 519 136
rect 549 124 637 247
rect 549 119 576 124
rect 564 90 576 119
rect 610 119 637 124
rect 667 165 723 247
rect 667 131 678 165
rect 712 131 723 165
rect 667 119 723 131
rect 753 234 810 247
rect 753 200 764 234
rect 798 200 810 234
rect 753 187 810 200
rect 753 119 803 187
rect 610 90 622 119
rect 564 78 622 90
rect 870 210 935 222
rect 870 176 882 210
rect 916 176 935 210
rect 870 120 935 176
rect 870 86 882 120
rect 916 86 935 120
rect 870 74 935 86
rect 965 210 1027 222
rect 965 176 982 210
rect 1016 176 1027 210
rect 965 120 1027 176
rect 965 86 982 120
rect 1016 86 1027 120
rect 965 74 1027 86
rect 1057 142 1127 222
rect 1057 108 1068 142
rect 1102 108 1127 142
rect 1057 74 1127 108
rect 1157 210 1213 222
rect 1157 176 1168 210
rect 1202 176 1213 210
rect 1157 120 1213 176
rect 1157 86 1168 120
rect 1202 86 1213 120
rect 1157 74 1213 86
rect 1243 120 1301 222
rect 1243 86 1254 120
rect 1288 86 1301 120
rect 1243 74 1301 86
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 509 86 546
rect 27 475 39 509
rect 73 475 86 509
rect 27 440 86 475
rect 27 406 39 440
rect 73 406 86 440
rect 27 392 86 406
rect 116 440 176 592
rect 116 406 129 440
rect 163 406 176 440
rect 116 392 176 406
rect 206 584 266 592
rect 206 550 219 584
rect 253 550 266 584
rect 206 516 266 550
rect 206 482 219 516
rect 253 482 266 516
rect 206 392 266 482
rect 296 580 359 592
rect 296 546 312 580
rect 346 546 359 580
rect 296 509 359 546
rect 296 475 312 509
rect 346 475 359 509
rect 296 438 359 475
rect 296 404 312 438
rect 346 404 359 438
rect 296 392 359 404
rect 389 580 459 592
rect 389 546 402 580
rect 436 546 459 580
rect 389 509 459 546
rect 389 475 402 509
rect 436 475 459 509
rect 389 438 459 475
rect 389 404 402 438
rect 436 404 459 438
rect 389 392 459 404
rect 489 580 549 592
rect 489 546 502 580
rect 536 546 549 580
rect 489 509 549 546
rect 489 475 502 509
rect 536 475 549 509
rect 489 438 549 475
rect 489 404 502 438
rect 536 404 549 438
rect 489 392 549 404
rect 579 580 726 592
rect 579 546 593 580
rect 627 546 679 580
rect 713 546 726 580
rect 579 512 726 546
rect 579 478 593 512
rect 627 478 679 512
rect 713 478 726 512
rect 579 392 726 478
rect 756 580 826 592
rect 756 546 779 580
rect 813 546 826 580
rect 756 510 826 546
rect 756 476 779 510
rect 813 476 826 510
rect 756 440 826 476
rect 756 406 779 440
rect 813 406 826 440
rect 756 392 826 406
rect 856 580 938 592
rect 856 546 879 580
rect 913 546 938 580
rect 856 508 938 546
rect 856 474 879 508
rect 913 474 938 508
rect 856 392 938 474
rect 885 368 938 392
rect 968 580 1038 592
rect 968 546 991 580
rect 1025 546 1038 580
rect 968 497 1038 546
rect 968 463 991 497
rect 1025 463 1038 497
rect 968 414 1038 463
rect 968 380 991 414
rect 1025 380 1038 414
rect 968 368 1038 380
rect 1068 580 1128 592
rect 1068 546 1081 580
rect 1115 546 1128 580
rect 1068 478 1128 546
rect 1068 444 1081 478
rect 1115 444 1128 478
rect 1068 368 1128 444
rect 1158 580 1218 592
rect 1158 546 1171 580
rect 1205 546 1218 580
rect 1158 497 1218 546
rect 1158 463 1171 497
rect 1205 463 1218 497
rect 1158 414 1218 463
rect 1158 380 1171 414
rect 1205 380 1218 414
rect 1158 368 1218 380
rect 1248 580 1317 592
rect 1248 546 1271 580
rect 1305 546 1317 580
rect 1248 497 1317 546
rect 1248 463 1271 497
rect 1305 463 1317 497
rect 1248 414 1317 463
rect 1248 380 1271 414
rect 1305 380 1317 414
rect 1248 368 1317 380
<< ndiffc >>
rect 44 201 78 235
rect 44 131 78 165
rect 130 132 164 166
rect 216 201 250 235
rect 302 132 336 166
rect 388 201 422 235
rect 388 131 422 165
rect 474 136 508 170
rect 576 90 610 124
rect 678 131 712 165
rect 764 200 798 234
rect 882 176 916 210
rect 882 86 916 120
rect 982 176 1016 210
rect 982 86 1016 120
rect 1068 108 1102 142
rect 1168 176 1202 210
rect 1168 86 1202 120
rect 1254 86 1288 120
<< pdiffc >>
rect 39 546 73 580
rect 39 475 73 509
rect 39 406 73 440
rect 129 406 163 440
rect 219 550 253 584
rect 219 482 253 516
rect 312 546 346 580
rect 312 475 346 509
rect 312 404 346 438
rect 402 546 436 580
rect 402 475 436 509
rect 402 404 436 438
rect 502 546 536 580
rect 502 475 536 509
rect 502 404 536 438
rect 593 546 627 580
rect 679 546 713 580
rect 593 478 627 512
rect 679 478 713 512
rect 779 546 813 580
rect 779 476 813 510
rect 779 406 813 440
rect 879 546 913 580
rect 879 474 913 508
rect 991 546 1025 580
rect 991 463 1025 497
rect 991 380 1025 414
rect 1081 546 1115 580
rect 1081 444 1115 478
rect 1171 546 1205 580
rect 1171 463 1205 497
rect 1171 380 1205 414
rect 1271 546 1305 580
rect 1271 463 1305 497
rect 1271 380 1305 414
<< poly >>
rect 86 592 116 618
rect 176 592 206 618
rect 266 592 296 618
rect 359 592 389 618
rect 459 592 489 618
rect 549 592 579 618
rect 726 592 756 618
rect 826 592 856 618
rect 938 592 968 618
rect 1038 592 1068 618
rect 1128 592 1158 618
rect 1218 592 1248 618
rect 86 377 116 392
rect 176 377 206 392
rect 266 377 296 392
rect 359 377 389 392
rect 459 377 489 392
rect 549 377 579 392
rect 726 377 756 392
rect 826 377 856 392
rect 83 356 119 377
rect 44 340 119 356
rect 44 306 60 340
rect 94 306 119 340
rect 44 290 119 306
rect 89 247 119 290
rect 175 356 209 377
rect 263 356 299 377
rect 175 340 299 356
rect 175 306 228 340
rect 262 306 299 340
rect 175 290 299 306
rect 356 340 392 377
rect 447 347 492 377
rect 546 360 582 377
rect 723 360 759 377
rect 356 292 386 340
rect 447 292 477 347
rect 546 344 759 360
rect 546 310 602 344
rect 636 330 759 344
rect 823 335 859 377
rect 938 353 968 368
rect 1038 353 1068 368
rect 1128 353 1158 368
rect 1218 353 1248 368
rect 636 310 667 330
rect 546 299 667 310
rect 175 247 205 290
rect 261 247 291 290
rect 347 262 386 292
rect 433 262 477 292
rect 519 269 667 299
rect 807 319 873 335
rect 807 285 823 319
rect 857 285 873 319
rect 347 247 377 262
rect 433 247 463 262
rect 519 247 549 269
rect 637 247 667 269
rect 723 247 753 273
rect 807 269 873 285
rect 935 326 971 353
rect 1035 326 1071 353
rect 1125 326 1161 353
rect 1215 326 1251 353
rect 935 310 1251 326
rect 935 276 951 310
rect 985 276 1019 310
rect 1053 276 1087 310
rect 1121 276 1251 310
rect 89 51 119 119
rect 175 93 205 119
rect 261 93 291 119
rect 347 51 377 119
rect 89 21 377 51
rect 433 51 463 119
rect 519 93 549 119
rect 637 93 667 119
rect 723 51 753 119
rect 825 51 855 269
rect 935 260 1251 276
rect 935 222 965 260
rect 1027 222 1057 260
rect 1127 222 1157 260
rect 1213 222 1243 260
rect 433 21 855 51
rect 935 48 965 74
rect 1027 48 1057 74
rect 1127 48 1157 74
rect 1213 48 1243 74
<< polycont >>
rect 60 306 94 340
rect 228 306 262 340
rect 602 310 636 344
rect 823 285 857 319
rect 951 276 985 310
rect 1019 276 1053 310
rect 1087 276 1121 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 23 580 79 649
rect 23 546 39 580
rect 73 546 79 580
rect 23 509 79 546
rect 23 475 39 509
rect 73 475 79 509
rect 203 584 269 649
rect 203 550 219 584
rect 253 550 269 584
rect 203 516 269 550
rect 203 482 219 516
rect 253 482 269 516
rect 312 580 346 596
rect 312 509 346 546
rect 23 440 79 475
rect 312 448 346 475
rect 23 406 39 440
rect 73 406 79 440
rect 23 390 79 406
rect 113 440 346 448
rect 113 406 129 440
rect 163 438 346 440
rect 163 406 312 438
rect 113 404 312 406
rect 113 390 346 404
rect 25 340 110 356
rect 25 306 60 340
rect 94 306 110 340
rect 25 290 110 306
rect 144 251 178 390
rect 212 340 278 356
rect 212 306 228 340
rect 262 306 278 340
rect 312 354 346 390
rect 386 580 452 649
rect 386 546 402 580
rect 436 546 452 580
rect 386 509 452 546
rect 386 475 402 509
rect 436 475 452 509
rect 386 438 452 475
rect 386 404 402 438
rect 436 404 452 438
rect 386 388 452 404
rect 486 580 552 596
rect 486 546 502 580
rect 536 546 552 580
rect 486 509 552 546
rect 486 475 502 509
rect 536 475 552 509
rect 486 438 552 475
rect 586 580 729 649
rect 586 546 593 580
rect 627 546 679 580
rect 713 546 729 580
rect 586 512 729 546
rect 586 478 593 512
rect 627 478 679 512
rect 713 478 729 512
rect 586 462 729 478
rect 763 580 829 596
rect 763 546 779 580
rect 813 546 829 580
rect 763 510 829 546
rect 763 476 779 510
rect 813 476 829 510
rect 486 404 502 438
rect 536 428 552 438
rect 763 440 829 476
rect 863 580 929 649
rect 863 546 879 580
rect 913 546 929 580
rect 863 508 929 546
rect 863 474 879 508
rect 913 474 929 508
rect 863 458 929 474
rect 975 580 1041 596
rect 975 546 991 580
rect 1025 546 1041 580
rect 975 497 1041 546
rect 975 463 991 497
rect 1025 463 1041 497
rect 763 428 779 440
rect 536 406 779 428
rect 813 424 829 440
rect 813 406 941 424
rect 536 404 941 406
rect 486 394 941 404
rect 486 354 552 394
rect 763 390 941 394
rect 312 320 552 354
rect 586 344 652 360
rect 212 290 278 306
rect 586 310 602 344
rect 636 310 652 344
rect 586 294 652 310
rect 796 319 873 356
rect 796 285 823 319
rect 857 285 873 319
rect 796 269 873 285
rect 907 326 941 390
rect 975 414 1041 463
rect 1081 580 1131 649
rect 1115 546 1131 580
rect 1081 478 1131 546
rect 1115 444 1131 478
rect 1081 428 1131 444
rect 1171 580 1221 596
rect 1205 546 1221 580
rect 1171 497 1221 546
rect 1205 463 1221 497
rect 975 380 991 414
rect 1025 394 1041 414
rect 1171 414 1221 463
rect 1025 380 1171 394
rect 1205 380 1221 414
rect 975 360 1221 380
rect 1255 580 1321 649
rect 1255 546 1271 580
rect 1305 546 1321 580
rect 1255 497 1321 546
rect 1255 463 1271 497
rect 1305 463 1321 497
rect 1255 414 1321 463
rect 1255 380 1271 414
rect 1305 380 1321 414
rect 1255 364 1321 380
rect 1171 330 1221 360
rect 907 310 1137 326
rect 907 276 951 310
rect 985 276 1019 310
rect 1053 276 1087 310
rect 1121 276 1137 310
rect 1171 296 1319 330
rect 907 260 1137 276
rect 28 235 78 251
rect 28 201 44 235
rect 144 235 266 251
rect 144 201 216 235
rect 250 201 266 235
rect 388 235 762 260
rect 422 234 814 235
rect 422 226 764 234
rect 28 165 78 201
rect 28 131 44 165
rect 114 166 352 167
rect 114 132 130 166
rect 164 132 302 166
rect 336 132 352 166
rect 114 131 352 132
rect 388 165 422 201
rect 728 200 764 226
rect 798 200 814 234
rect 1273 226 1319 296
rect 728 199 814 200
rect 866 210 932 226
rect 28 97 78 131
rect 388 97 422 131
rect 458 170 694 192
rect 458 136 474 170
rect 508 165 694 170
rect 866 176 882 210
rect 916 176 932 210
rect 508 158 678 165
rect 508 136 524 158
rect 458 115 524 136
rect 660 131 678 158
rect 712 131 728 165
rect 28 63 422 97
rect 560 90 576 124
rect 610 90 626 124
rect 660 115 728 131
rect 866 120 932 176
rect 560 17 626 90
rect 866 86 882 120
rect 916 86 932 120
rect 866 17 932 86
rect 966 210 1319 226
rect 966 176 982 210
rect 1016 192 1168 210
rect 966 120 1016 176
rect 1152 176 1168 192
rect 1202 192 1319 210
rect 1202 176 1218 192
rect 966 86 982 120
rect 966 70 1016 86
rect 1052 142 1118 158
rect 1052 108 1068 142
rect 1102 108 1118 142
rect 1052 17 1118 108
rect 1152 120 1218 176
rect 1152 86 1168 120
rect 1202 86 1218 120
rect 1152 70 1218 86
rect 1252 120 1304 136
rect 1252 86 1254 120
rect 1288 86 1304 120
rect 1252 17 1304 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
<< metal1 >>
rect 0 683 1344 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 0 617 1344 649
rect 0 17 1344 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
rect 0 -49 1344 -17
<< labels >>
rlabel comment s 0 0 0 0 4 and4_4
flabel pwell s 0 0 1344 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 1344 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 1344 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 1344 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 D
port 4 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 1279 242 1313 276 0 FreeSans 340 0 0 0 X
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 1344 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3371538
string GDS_START 3360608
<< end >>
