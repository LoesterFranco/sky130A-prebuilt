magic
tech sky130A
magscale 1 2
timestamp 1604502741
<< locali >>
rect 25 270 110 356
rect 212 364 329 414
rect 212 226 246 364
rect 407 270 473 356
rect 212 70 278 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 23 482 89 540
rect 130 516 196 649
rect 353 516 419 649
rect 23 448 541 482
rect 23 390 178 448
rect 144 236 178 390
rect 24 202 178 236
rect 293 260 359 326
rect 507 330 541 448
rect 575 364 655 572
rect 507 264 587 330
rect 325 230 359 260
rect 621 230 655 364
rect 24 108 90 202
rect 126 17 176 168
rect 325 196 655 230
rect 312 17 447 162
rect 481 70 547 196
rect 583 17 649 162
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel locali s 407 270 473 356 6 A
port 1 nsew signal input
rlabel locali s 25 270 110 356 6 B_N
port 2 nsew signal input
rlabel locali s 212 364 329 414 6 X
port 3 nsew signal output
rlabel locali s 212 226 246 364 6 X
port 3 nsew signal output
rlabel locali s 212 70 278 226 6 X
port 3 nsew signal output
rlabel metal1 s 0 -49 672 49 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 617 672 715 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 767442
string GDS_START 761948
<< end >>
