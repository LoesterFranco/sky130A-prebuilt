magic
tech sky130A
magscale 1 2
timestamp 1601050058
<< locali >>
rect 105 297 171 493
rect 21 215 87 265
rect 121 177 171 297
rect 105 51 171 177
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 276 561
rect 25 299 71 527
rect 205 299 247 527
rect 25 17 71 181
rect 205 17 247 181
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 276 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
<< metal1 >>
rect 0 561 276 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 276 561
rect 0 496 276 527
rect 0 17 276 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 276 17
rect 0 -48 276 -17
<< labels >>
rlabel locali s 21 215 87 265 6 A
port 1 nsew signal input
rlabel locali s 121 177 171 297 6 Y
port 2 nsew signal output
rlabel locali s 105 297 171 493 6 Y
port 2 nsew signal output
rlabel locali s 105 51 171 177 6 Y
port 2 nsew signal output
rlabel metal1 s 0 -48 276 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 276 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 276 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1608640
string GDS_START 1604892
<< end >>
