magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 25 270 359 356
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 24 390 74 649
rect 114 424 180 596
rect 220 458 254 649
rect 294 424 360 596
rect 400 458 450 649
rect 486 424 532 596
rect 114 390 427 424
rect 393 282 427 390
rect 478 390 492 424
rect 526 390 532 424
rect 566 406 632 649
rect 668 424 709 596
rect 393 236 442 282
rect 393 230 427 236
rect 109 196 427 230
rect 23 17 73 162
rect 109 70 159 196
rect 195 17 245 162
rect 285 70 335 196
rect 371 17 437 162
rect 478 70 532 390
rect 668 390 672 424
rect 706 390 709 424
rect 746 406 812 649
rect 846 424 886 596
rect 668 372 709 390
rect 846 390 849 424
rect 883 390 886 424
rect 926 406 992 649
rect 1028 424 1070 596
rect 846 372 886 390
rect 1028 390 1032 424
rect 1066 390 1070 424
rect 1106 406 1172 649
rect 1208 424 1249 596
rect 1028 372 1070 390
rect 1208 390 1212 424
rect 1246 390 1249 424
rect 1286 406 1352 649
rect 1389 424 1430 596
rect 1208 372 1249 390
rect 1389 390 1392 424
rect 1426 390 1430 424
rect 1466 406 1532 649
rect 1568 424 1610 596
rect 1389 372 1430 390
rect 1568 390 1572 424
rect 1606 390 1610 424
rect 1646 406 1712 649
rect 1750 424 1794 596
rect 1568 372 1610 390
rect 1750 390 1756 424
rect 1790 390 1794 424
rect 1830 406 1896 649
rect 1750 372 1794 390
rect 655 338 709 372
rect 834 338 886 372
rect 1005 338 1070 372
rect 1187 338 1249 372
rect 1373 338 1430 372
rect 1559 338 1610 372
rect 1745 366 1794 372
rect 567 238 621 304
rect 573 17 607 136
rect 655 70 700 338
rect 734 238 800 304
rect 834 149 868 338
rect 902 238 968 304
rect 734 17 779 145
rect 815 70 868 149
rect 902 17 967 148
rect 1005 70 1051 338
rect 1085 238 1151 304
rect 1087 17 1153 136
rect 1187 70 1237 338
rect 1273 238 1339 304
rect 1273 17 1339 136
rect 1373 70 1423 338
rect 1459 238 1525 304
rect 1459 17 1525 136
rect 1559 70 1609 338
rect 1645 238 1711 304
rect 1645 17 1711 136
rect 1745 70 1795 366
rect 1831 17 1897 149
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 492 390 526 424
rect 672 390 706 424
rect 849 390 883 424
rect 1032 390 1066 424
rect 1212 390 1246 424
rect 1392 390 1426 424
rect 1572 390 1606 424
rect 1756 390 1790 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
<< metal1 >>
rect 0 683 1920 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 0 617 1920 649
rect 478 424 1818 430
rect 478 390 492 424
rect 526 390 672 424
rect 706 390 849 424
rect 883 390 1032 424
rect 1066 390 1212 424
rect 1246 390 1392 424
rect 1426 390 1572 424
rect 1606 390 1756 424
rect 1790 390 1818 424
rect 478 384 1818 390
rect 0 17 1920 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
rect 0 -49 1920 -17
<< obsm1 >>
rect 388 236 1728 282
<< labels >>
rlabel locali s 25 270 359 356 6 A
port 1 nsew signal input
rlabel metal1 s 478 384 1818 430 6 X
port 2 nsew signal output
rlabel metal1 s 0 -49 1920 49 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1920 715 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1920 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3328040
string GDS_START 3312114
<< end >>
