magic
tech sky130A
magscale 1 2
timestamp 1599588209
<< nwell >>
rect -38 332 998 704
<< pwell >>
rect 0 0 960 49
<< scpmos >>
rect 85 392 115 592
rect 285 368 315 592
rect 375 368 405 592
rect 465 368 495 592
rect 555 368 585 592
rect 755 368 785 592
rect 845 368 875 592
<< nmoslvt >>
rect 85 74 115 202
rect 199 74 229 222
rect 288 74 318 222
rect 462 74 492 222
rect 548 74 578 222
rect 746 74 776 222
rect 842 74 872 222
<< ndiff >>
rect 149 202 199 222
rect 28 190 85 202
rect 28 156 40 190
rect 74 156 85 190
rect 28 120 85 156
rect 28 86 40 120
rect 74 86 85 120
rect 28 74 85 86
rect 115 188 199 202
rect 115 154 140 188
rect 174 154 199 188
rect 115 120 199 154
rect 115 86 140 120
rect 174 86 199 120
rect 115 74 199 86
rect 229 188 288 222
rect 229 154 240 188
rect 274 154 288 188
rect 229 120 288 154
rect 229 86 240 120
rect 274 86 288 120
rect 229 74 288 86
rect 318 120 462 222
rect 318 86 329 120
rect 363 86 417 120
rect 451 86 462 120
rect 318 74 462 86
rect 492 210 548 222
rect 492 176 503 210
rect 537 176 548 210
rect 492 120 548 176
rect 492 86 503 120
rect 537 86 548 120
rect 492 74 548 86
rect 578 138 746 222
rect 578 104 589 138
rect 623 104 701 138
rect 735 104 746 138
rect 578 74 746 104
rect 776 210 842 222
rect 776 176 787 210
rect 821 176 842 210
rect 776 120 842 176
rect 776 86 787 120
rect 821 86 842 120
rect 776 74 842 86
rect 872 210 933 222
rect 872 176 887 210
rect 921 176 933 210
rect 872 120 933 176
rect 872 86 887 120
rect 921 86 933 120
rect 872 74 933 86
<< pdiff >>
rect 27 580 85 592
rect 27 546 38 580
rect 72 546 85 580
rect 27 510 85 546
rect 27 476 38 510
rect 72 476 85 510
rect 27 440 85 476
rect 27 406 38 440
rect 72 406 85 440
rect 27 392 85 406
rect 115 580 173 592
rect 115 546 128 580
rect 162 546 173 580
rect 115 510 173 546
rect 115 476 128 510
rect 162 476 173 510
rect 115 440 173 476
rect 115 406 128 440
rect 162 406 173 440
rect 115 392 173 406
rect 227 580 285 592
rect 227 546 238 580
rect 272 546 285 580
rect 227 497 285 546
rect 227 463 238 497
rect 272 463 285 497
rect 227 414 285 463
rect 227 380 238 414
rect 272 380 285 414
rect 227 368 285 380
rect 315 531 375 592
rect 315 497 328 531
rect 362 497 375 531
rect 315 414 375 497
rect 315 380 328 414
rect 362 380 375 414
rect 315 368 375 380
rect 405 580 465 592
rect 405 546 418 580
rect 452 546 465 580
rect 405 497 465 546
rect 405 463 418 497
rect 452 463 465 497
rect 405 414 465 463
rect 405 380 418 414
rect 452 380 465 414
rect 405 368 465 380
rect 495 547 555 592
rect 495 513 508 547
rect 542 513 555 547
rect 495 424 555 513
rect 495 390 508 424
rect 542 390 555 424
rect 495 368 555 390
rect 585 576 643 592
rect 585 542 598 576
rect 632 542 643 576
rect 585 508 643 542
rect 585 474 598 508
rect 632 474 643 508
rect 585 368 643 474
rect 697 580 755 592
rect 697 546 708 580
rect 742 546 755 580
rect 697 496 755 546
rect 697 462 708 496
rect 742 462 755 496
rect 697 368 755 462
rect 785 580 845 592
rect 785 546 798 580
rect 832 546 845 580
rect 785 505 845 546
rect 785 471 798 505
rect 832 471 845 505
rect 785 424 845 471
rect 785 390 798 424
rect 832 390 845 424
rect 785 368 845 390
rect 875 580 933 592
rect 875 546 888 580
rect 922 546 933 580
rect 875 510 933 546
rect 875 476 888 510
rect 922 476 933 510
rect 875 440 933 476
rect 875 406 888 440
rect 922 406 933 440
rect 875 368 933 406
<< ndiffc >>
rect 40 156 74 190
rect 40 86 74 120
rect 140 154 174 188
rect 140 86 174 120
rect 240 154 274 188
rect 240 86 274 120
rect 329 86 363 120
rect 417 86 451 120
rect 503 176 537 210
rect 503 86 537 120
rect 589 104 623 138
rect 701 104 735 138
rect 787 176 821 210
rect 787 86 821 120
rect 887 176 921 210
rect 887 86 921 120
<< pdiffc >>
rect 38 546 72 580
rect 38 476 72 510
rect 38 406 72 440
rect 128 546 162 580
rect 128 476 162 510
rect 128 406 162 440
rect 238 546 272 580
rect 238 463 272 497
rect 238 380 272 414
rect 328 497 362 531
rect 328 380 362 414
rect 418 546 452 580
rect 418 463 452 497
rect 418 380 452 414
rect 508 513 542 547
rect 508 390 542 424
rect 598 542 632 576
rect 598 474 632 508
rect 708 546 742 580
rect 708 462 742 496
rect 798 546 832 580
rect 798 471 832 505
rect 798 390 832 424
rect 888 546 922 580
rect 888 476 922 510
rect 888 406 922 440
<< poly >>
rect 85 592 115 618
rect 285 592 315 618
rect 375 592 405 618
rect 465 592 495 618
rect 555 592 585 618
rect 755 592 785 618
rect 845 592 875 618
rect 85 377 115 392
rect 82 356 118 377
rect 82 340 151 356
rect 285 353 315 368
rect 375 353 405 368
rect 465 353 495 368
rect 555 353 585 368
rect 755 353 785 368
rect 845 353 875 368
rect 82 306 101 340
rect 135 306 151 340
rect 282 310 318 353
rect 82 290 151 306
rect 199 306 318 310
rect 372 306 408 353
rect 199 294 408 306
rect 85 202 115 290
rect 199 260 217 294
rect 251 260 408 294
rect 199 244 408 260
rect 462 336 498 353
rect 552 336 588 353
rect 752 336 788 353
rect 842 336 878 353
rect 462 320 655 336
rect 462 286 537 320
rect 571 286 605 320
rect 639 286 655 320
rect 462 270 655 286
rect 738 320 878 336
rect 738 286 754 320
rect 788 286 822 320
rect 856 286 878 320
rect 738 270 878 286
rect 199 222 229 244
rect 288 222 318 244
rect 462 222 492 270
rect 548 222 578 270
rect 746 222 776 270
rect 842 222 872 270
rect 85 48 115 74
rect 199 48 229 74
rect 288 48 318 74
rect 462 48 492 74
rect 548 48 578 74
rect 746 48 776 74
rect 842 48 872 74
<< polycont >>
rect 101 306 135 340
rect 217 260 251 294
rect 537 286 571 320
rect 605 286 639 320
rect 754 286 788 320
rect 822 286 856 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 17 580 72 596
rect 17 546 38 580
rect 17 510 72 546
rect 17 476 38 510
rect 17 440 72 476
rect 17 406 38 440
rect 17 390 72 406
rect 112 580 178 649
rect 112 546 128 580
rect 162 546 178 580
rect 112 510 178 546
rect 112 476 128 510
rect 162 476 178 510
rect 112 440 178 476
rect 112 406 128 440
rect 162 406 178 440
rect 112 390 178 406
rect 222 581 648 615
rect 222 580 288 581
rect 222 546 238 580
rect 272 546 288 580
rect 402 580 458 581
rect 222 497 288 546
rect 222 463 238 497
rect 272 463 288 497
rect 222 414 288 463
rect 17 256 51 390
rect 222 380 238 414
rect 272 380 288 414
rect 222 364 288 380
rect 328 531 362 547
rect 328 414 362 497
rect 85 340 167 356
rect 85 306 101 340
rect 135 306 167 340
rect 85 290 167 306
rect 201 294 267 310
rect 201 260 217 294
rect 251 260 267 294
rect 201 256 267 260
rect 17 222 267 256
rect 328 226 362 380
rect 402 546 418 580
rect 452 546 458 580
rect 594 576 648 581
rect 402 497 458 546
rect 402 463 418 497
rect 452 463 458 497
rect 402 414 458 463
rect 402 380 418 414
rect 452 380 458 414
rect 492 513 508 547
rect 542 513 558 547
rect 492 424 558 513
rect 594 542 598 576
rect 632 542 648 576
rect 594 508 648 542
rect 594 474 598 508
rect 632 474 648 508
rect 594 458 648 474
rect 692 580 758 649
rect 692 546 708 580
rect 742 546 758 580
rect 692 496 758 546
rect 692 462 708 496
rect 742 462 758 496
rect 692 458 758 462
rect 798 580 848 596
rect 832 546 848 580
rect 798 505 848 546
rect 832 471 848 505
rect 798 424 848 471
rect 492 390 508 424
rect 542 390 798 424
rect 832 390 848 424
rect 885 580 938 649
rect 885 546 888 580
rect 922 546 938 580
rect 885 510 938 546
rect 885 476 888 510
rect 922 476 938 510
rect 885 440 938 476
rect 885 406 888 440
rect 922 406 938 440
rect 885 390 938 406
rect 402 364 458 380
rect 521 320 655 356
rect 521 286 537 320
rect 571 286 605 320
rect 639 286 655 320
rect 521 270 655 286
rect 697 320 935 356
rect 697 286 754 320
rect 788 286 822 320
rect 856 286 935 320
rect 697 270 935 286
rect 17 190 90 222
rect 17 156 40 190
rect 74 156 90 190
rect 313 210 837 226
rect 313 188 503 210
rect 17 120 90 156
rect 17 86 40 120
rect 74 86 90 120
rect 17 70 90 86
rect 124 154 140 188
rect 174 154 190 188
rect 124 120 190 154
rect 124 86 140 120
rect 174 86 190 120
rect 124 17 190 86
rect 224 154 240 188
rect 274 176 503 188
rect 537 192 787 210
rect 537 176 539 192
rect 274 154 539 176
rect 785 176 787 192
rect 821 176 837 210
rect 224 120 279 154
rect 501 120 539 154
rect 224 86 240 120
rect 274 86 279 120
rect 224 70 279 86
rect 313 86 329 120
rect 363 86 417 120
rect 451 86 467 120
rect 313 17 467 86
rect 501 86 503 120
rect 537 86 539 120
rect 501 70 539 86
rect 573 138 751 154
rect 573 104 589 138
rect 623 104 701 138
rect 735 104 751 138
rect 573 17 751 104
rect 785 120 837 176
rect 785 86 787 120
rect 821 86 837 120
rect 785 70 837 86
rect 871 210 937 226
rect 871 176 887 210
rect 921 176 937 210
rect 871 120 937 176
rect 871 86 887 120
rect 921 86 937 120
rect 871 17 937 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
rlabel comment s 0 0 0 0 4 nor3b_2
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 319 168 353 202 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 415 168 449 202 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 C_N
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 960 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1704206
string GDS_START 1695484
<< end >>
