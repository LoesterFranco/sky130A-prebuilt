magic
tech sky130A
magscale 1 2
timestamp 1604502710
<< nwell >>
rect -38 335 3014 704
rect -38 332 710 335
rect 1194 332 3014 335
rect 1625 311 1929 332
<< pwell >>
rect 0 0 2976 49
<< scpmos >>
rect 83 464 119 592
rect 307 464 343 592
rect 391 464 427 592
rect 481 464 517 592
rect 593 464 629 592
rect 707 464 743 592
rect 911 387 947 611
rect 1001 387 1037 611
rect 1209 463 1245 547
rect 1309 463 1345 547
rect 1387 463 1423 547
rect 1515 463 1551 547
rect 1717 347 1753 547
rect 1807 347 1843 547
rect 1949 508 1985 592
rect 2033 508 2069 592
rect 2170 508 2206 592
rect 2277 508 2313 592
rect 2390 368 2426 536
rect 2480 368 2516 536
rect 2587 368 2623 592
rect 2677 368 2713 592
rect 2767 368 2803 592
rect 2857 368 2893 592
<< nmoslvt >>
rect 84 74 114 158
rect 282 81 312 165
rect 385 81 415 165
rect 525 81 555 165
rect 597 81 627 165
rect 693 81 723 165
rect 904 119 934 267
rect 1014 119 1044 267
rect 1203 138 1233 222
rect 1289 138 1319 222
rect 1367 138 1397 222
rect 1445 138 1475 222
rect 1620 74 1650 222
rect 1715 74 1745 202
rect 1925 74 1955 158
rect 2003 74 2033 158
rect 2111 74 2141 158
rect 2183 74 2213 158
rect 2396 74 2426 222
rect 2482 74 2512 222
rect 2568 74 2598 222
rect 2776 74 2806 222
rect 2862 74 2892 222
<< ndiff >>
rect 853 235 904 267
rect 27 133 84 158
rect 27 99 39 133
rect 73 99 84 133
rect 27 74 84 99
rect 114 128 171 158
rect 114 94 125 128
rect 159 94 171 128
rect 114 74 171 94
rect 225 127 282 165
rect 225 93 237 127
rect 271 93 282 127
rect 225 81 282 93
rect 312 81 385 165
rect 415 153 525 165
rect 415 119 480 153
rect 514 119 525 153
rect 415 81 525 119
rect 555 81 597 165
rect 627 130 693 165
rect 627 96 644 130
rect 678 96 693 130
rect 627 81 693 96
rect 723 134 780 165
rect 723 100 738 134
rect 772 100 780 134
rect 723 81 780 100
rect 834 150 904 235
rect 834 116 847 150
rect 881 119 904 150
rect 934 150 1014 267
rect 934 119 957 150
rect 881 116 889 119
rect 834 93 889 116
rect 949 116 957 119
rect 991 119 1014 150
rect 1044 239 1096 267
rect 1044 205 1054 239
rect 1088 205 1096 239
rect 1044 165 1096 205
rect 1044 131 1054 165
rect 1088 131 1096 165
rect 1150 197 1203 222
rect 1150 163 1158 197
rect 1192 163 1203 197
rect 1150 138 1203 163
rect 1233 191 1289 222
rect 1233 157 1244 191
rect 1278 157 1289 191
rect 1233 138 1289 157
rect 1319 138 1367 222
rect 1397 138 1445 222
rect 1475 138 1620 222
rect 1044 119 1096 131
rect 991 116 999 119
rect 949 93 999 116
rect 1490 82 1620 138
rect 1490 48 1502 82
rect 1536 74 1620 82
rect 1650 202 1700 222
rect 1650 179 1715 202
rect 1650 145 1670 179
rect 1704 145 1715 179
rect 1650 74 1715 145
rect 1745 158 1795 202
rect 2339 210 2396 222
rect 2339 176 2351 210
rect 2385 176 2396 210
rect 1745 131 1925 158
rect 1745 97 1864 131
rect 1898 97 1925 131
rect 1745 74 1925 97
rect 1955 74 2003 158
rect 2033 120 2111 158
rect 2033 86 2055 120
rect 2089 86 2111 120
rect 2033 74 2111 86
rect 2141 74 2183 158
rect 2213 127 2285 158
rect 2213 93 2231 127
rect 2265 93 2285 127
rect 2213 74 2285 93
rect 2339 120 2396 176
rect 2339 86 2351 120
rect 2385 86 2396 120
rect 2339 74 2396 86
rect 2426 204 2482 222
rect 2426 170 2437 204
rect 2471 170 2482 204
rect 2426 120 2482 170
rect 2426 86 2437 120
rect 2471 86 2482 120
rect 2426 74 2482 86
rect 2512 204 2568 222
rect 2512 170 2523 204
rect 2557 170 2568 204
rect 2512 120 2568 170
rect 2512 86 2523 120
rect 2557 86 2568 120
rect 2512 74 2568 86
rect 2598 136 2776 222
rect 2598 102 2609 136
rect 2643 102 2731 136
rect 2765 102 2776 136
rect 2598 74 2776 102
rect 2806 210 2862 222
rect 2806 176 2817 210
rect 2851 176 2862 210
rect 2806 120 2862 176
rect 2806 86 2817 120
rect 2851 86 2862 120
rect 2806 74 2862 86
rect 2892 210 2949 222
rect 2892 176 2903 210
rect 2937 176 2949 210
rect 2892 120 2949 176
rect 2892 86 2903 120
rect 2937 86 2949 120
rect 2892 74 2949 86
rect 1536 48 1548 74
rect 1490 36 1548 48
<< pdiff >>
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 510 83 546
rect 27 476 39 510
rect 73 476 83 510
rect 27 464 83 476
rect 119 580 307 592
rect 119 546 139 580
rect 173 546 263 580
rect 297 546 307 580
rect 119 510 307 546
rect 119 476 139 510
rect 173 476 263 510
rect 297 476 307 510
rect 119 464 307 476
rect 343 464 391 592
rect 427 580 481 592
rect 427 546 437 580
rect 471 546 481 580
rect 427 510 481 546
rect 427 476 437 510
rect 471 476 481 510
rect 427 464 481 476
rect 517 464 593 592
rect 629 575 707 592
rect 629 541 640 575
rect 674 541 707 575
rect 629 464 707 541
rect 743 580 800 592
rect 743 546 754 580
rect 788 546 800 580
rect 743 510 800 546
rect 743 476 754 510
rect 788 476 800 510
rect 743 464 800 476
rect 855 441 911 611
rect 855 407 867 441
rect 901 407 911 441
rect 855 387 911 407
rect 947 593 1001 611
rect 947 559 957 593
rect 991 559 1001 593
rect 947 387 1001 559
rect 1037 441 1093 611
rect 1037 407 1047 441
rect 1081 407 1093 441
rect 1037 387 1093 407
rect 1438 582 1500 594
rect 1438 548 1452 582
rect 1486 548 1500 582
rect 1438 547 1500 548
rect 1858 560 1949 592
rect 1858 547 1887 560
rect 1153 522 1209 547
rect 1153 488 1165 522
rect 1199 488 1209 522
rect 1153 463 1209 488
rect 1245 535 1309 547
rect 1245 501 1265 535
rect 1299 501 1309 535
rect 1245 463 1309 501
rect 1345 463 1387 547
rect 1423 463 1515 547
rect 1551 524 1607 547
rect 1551 490 1561 524
rect 1595 490 1607 524
rect 1551 463 1607 490
rect 1661 535 1717 547
rect 1661 501 1673 535
rect 1707 501 1717 535
rect 1661 467 1717 501
rect 1661 433 1673 467
rect 1707 433 1717 467
rect 1661 399 1717 433
rect 1661 365 1673 399
rect 1707 365 1717 399
rect 1661 347 1717 365
rect 1753 535 1807 547
rect 1753 501 1763 535
rect 1797 501 1807 535
rect 1753 464 1807 501
rect 1753 430 1763 464
rect 1797 430 1807 464
rect 1753 393 1807 430
rect 1753 359 1763 393
rect 1797 359 1807 393
rect 1753 347 1807 359
rect 1843 526 1887 547
rect 1921 526 1949 560
rect 1843 508 1949 526
rect 1985 508 2033 592
rect 2069 567 2170 592
rect 2069 533 2109 567
rect 2143 533 2170 567
rect 2069 508 2170 533
rect 2206 567 2277 592
rect 2206 533 2216 567
rect 2250 533 2277 567
rect 2206 508 2277 533
rect 2313 536 2375 592
rect 2531 580 2587 592
rect 2531 546 2543 580
rect 2577 546 2587 580
rect 2531 536 2587 546
rect 2313 524 2390 536
rect 2313 508 2346 524
rect 1843 347 1893 508
rect 2333 490 2346 508
rect 2380 490 2390 524
rect 2333 414 2390 490
rect 2333 380 2346 414
rect 2380 380 2390 414
rect 2333 368 2390 380
rect 2426 524 2480 536
rect 2426 490 2436 524
rect 2470 490 2480 524
rect 2426 414 2480 490
rect 2426 380 2436 414
rect 2470 380 2480 414
rect 2426 368 2480 380
rect 2516 497 2587 536
rect 2516 463 2543 497
rect 2577 463 2587 497
rect 2516 414 2587 463
rect 2516 380 2543 414
rect 2577 380 2587 414
rect 2516 368 2587 380
rect 2623 580 2677 592
rect 2623 546 2633 580
rect 2667 546 2677 580
rect 2623 497 2677 546
rect 2623 463 2633 497
rect 2667 463 2677 497
rect 2623 414 2677 463
rect 2623 380 2633 414
rect 2667 380 2677 414
rect 2623 368 2677 380
rect 2713 580 2767 592
rect 2713 546 2723 580
rect 2757 546 2767 580
rect 2713 472 2767 546
rect 2713 438 2723 472
rect 2757 438 2767 472
rect 2713 368 2767 438
rect 2803 580 2857 592
rect 2803 546 2813 580
rect 2847 546 2857 580
rect 2803 497 2857 546
rect 2803 463 2813 497
rect 2847 463 2857 497
rect 2803 414 2857 463
rect 2803 380 2813 414
rect 2847 380 2857 414
rect 2803 368 2857 380
rect 2893 580 2949 592
rect 2893 546 2903 580
rect 2937 546 2949 580
rect 2893 472 2949 546
rect 2893 438 2903 472
rect 2937 438 2949 472
rect 2893 368 2949 438
<< ndiffc >>
rect 39 99 73 133
rect 125 94 159 128
rect 237 93 271 127
rect 480 119 514 153
rect 644 96 678 130
rect 738 100 772 134
rect 847 116 881 150
rect 957 116 991 150
rect 1054 205 1088 239
rect 1054 131 1088 165
rect 1158 163 1192 197
rect 1244 157 1278 191
rect 1502 48 1536 82
rect 1670 145 1704 179
rect 2351 176 2385 210
rect 1864 97 1898 131
rect 2055 86 2089 120
rect 2231 93 2265 127
rect 2351 86 2385 120
rect 2437 170 2471 204
rect 2437 86 2471 120
rect 2523 170 2557 204
rect 2523 86 2557 120
rect 2609 102 2643 136
rect 2731 102 2765 136
rect 2817 176 2851 210
rect 2817 86 2851 120
rect 2903 176 2937 210
rect 2903 86 2937 120
<< pdiffc >>
rect 39 546 73 580
rect 39 476 73 510
rect 139 546 173 580
rect 263 546 297 580
rect 139 476 173 510
rect 263 476 297 510
rect 437 546 471 580
rect 437 476 471 510
rect 640 541 674 575
rect 754 546 788 580
rect 754 476 788 510
rect 867 407 901 441
rect 957 559 991 593
rect 1047 407 1081 441
rect 1452 548 1486 582
rect 1165 488 1199 522
rect 1265 501 1299 535
rect 1561 490 1595 524
rect 1673 501 1707 535
rect 1673 433 1707 467
rect 1673 365 1707 399
rect 1763 501 1797 535
rect 1763 430 1797 464
rect 1763 359 1797 393
rect 1887 526 1921 560
rect 2109 533 2143 567
rect 2216 533 2250 567
rect 2543 546 2577 580
rect 2346 490 2380 524
rect 2346 380 2380 414
rect 2436 490 2470 524
rect 2436 380 2470 414
rect 2543 463 2577 497
rect 2543 380 2577 414
rect 2633 546 2667 580
rect 2633 463 2667 497
rect 2633 380 2667 414
rect 2723 546 2757 580
rect 2723 438 2757 472
rect 2813 546 2847 580
rect 2813 463 2847 497
rect 2813 380 2847 414
rect 2903 546 2937 580
rect 2903 438 2937 472
<< poly >>
rect 83 592 119 618
rect 307 592 343 618
rect 391 592 427 618
rect 481 592 517 618
rect 593 592 629 618
rect 707 592 743 618
rect 911 611 947 637
rect 1001 611 1037 637
rect 1108 615 1843 645
rect 83 367 119 464
rect 307 367 343 464
rect 83 351 343 367
rect 83 317 137 351
rect 171 317 205 351
rect 239 317 273 351
rect 307 317 343 351
rect 83 301 343 317
rect 84 158 114 301
rect 391 253 427 464
rect 481 432 517 464
rect 593 449 629 464
rect 707 449 743 464
rect 473 416 539 432
rect 473 382 489 416
rect 523 382 539 416
rect 473 366 539 382
rect 581 406 647 449
rect 581 372 597 406
rect 631 372 647 406
rect 581 338 647 372
rect 162 237 228 253
rect 162 203 178 237
rect 212 217 228 237
rect 354 237 427 253
rect 473 302 539 318
rect 473 268 489 302
rect 523 268 539 302
rect 581 304 597 338
rect 631 304 647 338
rect 581 288 647 304
rect 693 432 743 449
rect 693 416 823 432
rect 693 382 773 416
rect 807 382 823 416
rect 693 370 823 382
rect 693 366 819 370
rect 473 252 539 268
rect 212 203 312 217
rect 162 187 312 203
rect 354 203 370 237
rect 404 203 427 237
rect 509 240 539 252
rect 509 210 555 240
rect 354 187 427 203
rect 282 165 312 187
rect 385 165 415 187
rect 525 165 555 210
rect 597 165 627 288
rect 693 165 723 366
rect 911 355 947 387
rect 1001 355 1037 387
rect 866 351 947 355
rect 862 339 947 351
rect 862 322 878 339
rect 765 306 878 322
rect 765 272 781 306
rect 815 305 878 306
rect 912 305 947 339
rect 815 282 947 305
rect 995 339 1061 355
rect 995 305 1011 339
rect 1045 319 1061 339
rect 1108 319 1138 615
rect 1209 547 1245 573
rect 1309 547 1345 615
rect 1387 547 1423 573
rect 1515 547 1551 573
rect 1717 547 1753 573
rect 1807 547 1843 615
rect 1949 592 1985 618
rect 2033 592 2069 618
rect 2170 592 2206 618
rect 2277 592 2313 618
rect 2587 592 2623 618
rect 2677 592 2713 618
rect 2767 592 2803 618
rect 2857 592 2893 618
rect 1209 383 1245 463
rect 1309 437 1345 463
rect 1387 389 1423 463
rect 1515 430 1551 463
rect 1515 414 1629 430
rect 1045 305 1138 319
rect 1180 367 1246 383
rect 1180 333 1196 367
rect 1230 347 1246 367
rect 1367 373 1471 389
rect 1230 333 1319 347
rect 1180 317 1319 333
rect 995 295 1138 305
rect 995 282 1143 295
rect 815 272 837 282
rect 765 256 837 272
rect 904 267 934 282
rect 1014 267 1044 282
rect 1109 275 1143 282
rect 904 93 934 119
rect 1111 245 1233 275
rect 1203 222 1233 245
rect 1289 222 1319 317
rect 1367 339 1421 373
rect 1455 339 1471 373
rect 1367 323 1471 339
rect 1515 380 1579 414
rect 1613 380 1629 414
rect 1515 364 1629 380
rect 1367 222 1397 323
rect 1515 267 1549 364
rect 2390 536 2426 562
rect 2480 536 2516 562
rect 1949 476 1985 508
rect 1925 460 1991 476
rect 1925 426 1941 460
rect 1975 426 1991 460
rect 1925 410 1991 426
rect 1717 319 1753 347
rect 1445 237 1549 267
rect 1597 299 1753 319
rect 1807 332 1843 347
rect 1807 302 1955 332
rect 2033 311 2069 508
rect 2170 430 2206 508
rect 1597 265 1613 299
rect 1647 289 1753 299
rect 1647 265 1663 289
rect 1597 249 1663 265
rect 1445 222 1475 237
rect 1620 222 1650 249
rect 1715 231 1883 247
rect 1014 93 1044 119
rect 1203 112 1233 138
rect 1289 112 1319 138
rect 1367 112 1397 138
rect 84 48 114 74
rect 282 55 312 81
rect 385 55 415 81
rect 525 55 555 81
rect 597 55 627 81
rect 693 51 723 81
rect 1445 51 1475 138
rect 693 21 1475 51
rect 1715 217 1833 231
rect 1715 202 1745 217
rect 1817 197 1833 217
rect 1867 197 1883 231
rect 1817 181 1883 197
rect 1925 158 1955 302
rect 2003 295 2069 311
rect 2003 261 2019 295
rect 2053 261 2069 295
rect 2003 245 2069 261
rect 2111 414 2206 430
rect 2111 380 2133 414
rect 2167 380 2206 414
rect 2111 364 2206 380
rect 2003 158 2033 245
rect 2111 158 2141 364
rect 2277 315 2313 508
rect 2390 353 2426 368
rect 2480 353 2516 368
rect 2390 323 2516 353
rect 2277 267 2307 315
rect 2396 267 2426 323
rect 2587 320 2623 368
rect 2677 320 2713 368
rect 2767 320 2803 368
rect 2857 320 2893 368
rect 2568 304 2893 320
rect 2568 275 2584 304
rect 2183 237 2426 267
rect 2183 230 2307 237
rect 2183 196 2199 230
rect 2233 196 2307 230
rect 2396 222 2426 237
rect 2482 270 2584 275
rect 2618 270 2652 304
rect 2686 270 2720 304
rect 2754 290 2893 304
rect 2754 270 2892 290
rect 2482 245 2892 270
rect 2482 222 2512 245
rect 2568 222 2598 245
rect 2776 222 2806 245
rect 2862 222 2892 245
rect 2183 180 2307 196
rect 2183 158 2213 180
rect 1620 48 1650 74
rect 1715 48 1745 74
rect 1925 48 1955 74
rect 2003 48 2033 74
rect 2111 48 2141 74
rect 2183 48 2213 74
rect 2396 48 2426 74
rect 2482 48 2512 74
rect 2568 48 2598 74
rect 2776 48 2806 74
rect 2862 48 2892 74
<< polycont >>
rect 137 317 171 351
rect 205 317 239 351
rect 273 317 307 351
rect 489 382 523 416
rect 597 372 631 406
rect 178 203 212 237
rect 489 268 523 302
rect 597 304 631 338
rect 773 382 807 416
rect 370 203 404 237
rect 781 272 815 306
rect 878 305 912 339
rect 1011 305 1045 339
rect 1196 333 1230 367
rect 1421 339 1455 373
rect 1579 380 1613 414
rect 1941 426 1975 460
rect 1613 265 1647 299
rect 1833 197 1867 231
rect 2019 261 2053 295
rect 2133 380 2167 414
rect 2199 196 2233 230
rect 2584 270 2618 304
rect 2652 270 2686 304
rect 2720 270 2754 304
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 2976 683
rect 23 580 89 596
rect 23 546 39 580
rect 73 546 89 580
rect 23 510 89 546
rect 23 476 39 510
rect 73 476 89 510
rect 23 435 89 476
rect 123 580 313 649
rect 123 546 139 580
rect 173 546 263 580
rect 297 546 313 580
rect 123 510 313 546
rect 123 476 139 510
rect 173 476 263 510
rect 297 476 313 510
rect 123 469 313 476
rect 421 580 487 596
rect 421 546 437 580
rect 471 546 487 580
rect 421 510 487 546
rect 619 575 690 649
rect 619 541 640 575
rect 674 541 690 575
rect 619 538 690 541
rect 724 580 804 611
rect 724 546 754 580
rect 788 546 804 580
rect 941 593 1007 649
rect 941 559 957 593
rect 991 559 1007 593
rect 1434 582 1504 649
rect 421 476 437 510
rect 471 503 487 510
rect 724 525 804 546
rect 1165 525 1215 545
rect 724 522 1215 525
rect 724 510 1165 522
rect 724 503 754 510
rect 471 476 754 503
rect 788 491 1165 510
rect 788 476 804 491
rect 421 469 804 476
rect 1199 488 1215 522
rect 23 416 541 435
rect 23 401 489 416
rect 23 253 57 401
rect 475 382 489 401
rect 523 382 541 416
rect 121 351 359 367
rect 475 366 541 382
rect 589 406 655 430
rect 589 372 597 406
rect 631 372 655 406
rect 121 317 137 351
rect 171 317 205 351
rect 239 317 273 351
rect 307 332 359 351
rect 589 338 655 372
rect 307 317 547 332
rect 121 302 547 317
rect 121 298 489 302
rect 481 268 489 298
rect 523 268 547 302
rect 589 304 597 338
rect 631 304 655 338
rect 589 288 655 304
rect 23 237 228 253
rect 23 203 178 237
rect 212 203 228 237
rect 23 187 228 203
rect 313 237 420 253
rect 481 252 547 268
rect 313 203 370 237
rect 404 203 420 237
rect 689 218 723 469
rect 867 441 917 457
rect 757 424 833 432
rect 757 416 799 424
rect 757 382 773 416
rect 807 382 833 390
rect 901 434 917 441
rect 1031 441 1131 455
rect 901 407 996 434
rect 867 389 996 407
rect 1031 407 1047 441
rect 1081 407 1131 441
rect 1165 451 1215 488
rect 1249 535 1377 551
rect 1249 501 1265 535
rect 1299 501 1377 535
rect 1434 548 1452 582
rect 1486 548 1504 582
rect 1434 532 1504 548
rect 1249 498 1377 501
rect 1545 524 1611 551
rect 1545 498 1561 524
rect 1249 490 1561 498
rect 1595 490 1611 524
rect 1249 485 1611 490
rect 1343 464 1611 485
rect 1673 535 1707 649
rect 1854 560 2059 576
rect 1673 467 1707 501
rect 1165 417 1309 451
rect 1031 394 1131 407
rect 757 366 833 382
rect 962 360 996 389
rect 1090 383 1131 394
rect 1090 367 1241 383
rect 867 339 928 355
rect 867 332 878 339
rect 23 133 73 187
rect 313 162 420 203
rect 513 184 723 218
rect 757 306 878 332
rect 757 272 781 306
rect 815 305 878 306
rect 912 305 928 339
rect 815 272 928 305
rect 757 252 928 272
rect 962 339 1056 360
rect 962 305 1011 339
rect 1045 305 1056 339
rect 962 289 1056 305
rect 1090 333 1196 367
rect 1230 333 1241 367
rect 1090 317 1241 333
rect 757 184 839 252
rect 962 218 1004 289
rect 1090 255 1124 317
rect 1275 283 1309 417
rect 873 184 1004 218
rect 1041 239 1124 255
rect 1041 205 1054 239
rect 1088 205 1124 239
rect 513 169 547 184
rect 464 153 547 169
rect 23 99 39 133
rect 23 70 73 99
rect 109 128 175 153
rect 109 94 125 128
rect 159 94 175 128
rect 109 17 175 94
rect 221 127 287 128
rect 221 93 237 127
rect 271 93 287 127
rect 464 119 480 153
rect 514 119 547 153
rect 873 150 907 184
rect 1041 165 1124 205
rect 628 130 694 150
rect 221 85 287 93
rect 628 96 644 130
rect 678 96 694 130
rect 628 85 694 96
rect 221 51 694 85
rect 728 134 788 150
rect 728 100 738 134
rect 772 100 788 134
rect 827 116 847 150
rect 881 116 907 150
rect 827 100 907 116
rect 941 116 957 150
rect 991 116 1007 150
rect 728 17 788 100
rect 941 17 1007 116
rect 1041 131 1054 165
rect 1088 131 1124 165
rect 1158 249 1309 283
rect 1158 197 1192 249
rect 1343 215 1377 464
rect 1158 134 1192 163
rect 1228 191 1377 215
rect 1228 157 1244 191
rect 1278 181 1377 191
rect 1411 373 1465 389
rect 1411 339 1421 373
rect 1455 339 1465 373
rect 1411 218 1465 339
rect 1499 315 1533 464
rect 1567 424 1629 430
rect 1601 414 1629 424
rect 1567 380 1579 390
rect 1613 380 1629 414
rect 1567 364 1629 380
rect 1673 399 1707 433
rect 1673 349 1707 365
rect 1747 535 1813 551
rect 1747 501 1763 535
rect 1797 501 1813 535
rect 1854 526 1887 560
rect 1921 526 2059 560
rect 1854 510 2059 526
rect 1747 464 1813 501
rect 1747 430 1763 464
rect 1797 430 1813 464
rect 1747 393 1813 430
rect 1747 359 1763 393
rect 1797 359 1813 393
rect 1747 315 1813 359
rect 1499 299 1663 315
rect 1499 265 1613 299
rect 1647 265 1663 299
rect 1499 252 1663 265
rect 1697 281 1813 315
rect 1849 460 1991 476
rect 1849 426 1941 460
rect 1975 426 1991 460
rect 1849 413 1991 426
rect 1697 218 1731 281
rect 1849 247 1883 413
rect 2025 379 2059 510
rect 2093 567 2159 649
rect 2093 533 2109 567
rect 2143 533 2159 567
rect 2093 504 2159 533
rect 2200 567 2266 596
rect 2200 533 2216 567
rect 2250 533 2266 567
rect 2200 504 2266 533
rect 1411 184 1731 218
rect 1278 157 1294 181
rect 1228 134 1294 157
rect 1654 179 1731 184
rect 1041 100 1124 131
rect 1411 116 1620 150
rect 1654 145 1670 179
rect 1704 145 1731 179
rect 1654 119 1731 145
rect 1765 231 1883 247
rect 1765 197 1833 231
rect 1867 197 1883 231
rect 1765 181 1883 197
rect 1917 345 2059 379
rect 2117 424 2183 430
rect 2117 414 2143 424
rect 2117 380 2133 414
rect 2177 390 2183 424
rect 2167 380 2183 390
rect 2117 364 2183 380
rect 1917 211 1951 345
rect 2232 311 2266 504
rect 2330 524 2380 649
rect 2527 580 2577 649
rect 2527 546 2543 580
rect 2330 490 2346 524
rect 2330 414 2380 490
rect 2330 380 2346 414
rect 2330 364 2380 380
rect 2420 524 2486 540
rect 2420 490 2436 524
rect 2470 490 2486 524
rect 2420 414 2486 490
rect 2420 380 2436 414
rect 2470 380 2486 414
rect 2420 320 2486 380
rect 2527 497 2577 546
rect 2527 463 2543 497
rect 2527 414 2577 463
rect 2527 380 2543 414
rect 2527 364 2577 380
rect 2617 580 2683 596
rect 2617 546 2633 580
rect 2667 546 2683 580
rect 2617 497 2683 546
rect 2617 463 2633 497
rect 2667 463 2683 497
rect 2617 414 2683 463
rect 2723 580 2773 649
rect 2757 546 2773 580
rect 2723 472 2773 546
rect 2757 438 2773 472
rect 2723 422 2773 438
rect 2813 580 2856 596
rect 2847 546 2856 580
rect 2813 497 2856 546
rect 2847 463 2856 497
rect 2617 380 2633 414
rect 2667 388 2683 414
rect 2813 414 2856 463
rect 2894 580 2953 649
rect 2894 546 2903 580
rect 2937 546 2953 580
rect 2894 472 2953 546
rect 2894 438 2903 472
rect 2937 438 2953 472
rect 2894 422 2953 438
rect 2667 380 2813 388
rect 2847 388 2856 414
rect 2847 380 2951 388
rect 2617 354 2951 380
rect 2003 295 2317 311
rect 2003 261 2019 295
rect 2053 277 2317 295
rect 2053 261 2069 277
rect 2003 245 2069 261
rect 2183 230 2249 243
rect 2183 211 2199 230
rect 1917 196 2199 211
rect 2233 196 2249 230
rect 1411 100 1445 116
rect 1041 66 1445 100
rect 1586 85 1620 116
rect 1765 85 1799 181
rect 1917 177 2249 196
rect 1917 147 1951 177
rect 1486 48 1502 82
rect 1536 48 1552 82
rect 1586 51 1799 85
rect 1833 131 1951 147
rect 2283 143 2317 277
rect 1833 97 1864 131
rect 1898 97 1951 131
rect 1833 81 1951 97
rect 2028 120 2116 136
rect 2028 86 2055 120
rect 2089 86 2116 120
rect 1486 17 1552 48
rect 2028 17 2116 86
rect 2208 127 2317 143
rect 2208 93 2231 127
rect 2265 93 2317 127
rect 2208 77 2317 93
rect 2351 304 2770 320
rect 2351 270 2584 304
rect 2618 270 2652 304
rect 2686 270 2720 304
rect 2754 270 2770 304
rect 2351 254 2770 270
rect 2817 260 2951 354
rect 2351 210 2385 254
rect 2817 220 2851 260
rect 2351 120 2385 176
rect 2351 70 2385 86
rect 2421 204 2473 220
rect 2421 170 2437 204
rect 2471 170 2473 204
rect 2421 120 2473 170
rect 2421 86 2437 120
rect 2471 86 2473 120
rect 2421 17 2473 86
rect 2507 210 2851 220
rect 2507 204 2817 210
rect 2507 170 2523 204
rect 2557 186 2817 204
rect 2557 170 2573 186
rect 2507 120 2573 170
rect 2507 86 2523 120
rect 2557 86 2573 120
rect 2507 70 2573 86
rect 2607 136 2781 152
rect 2607 102 2609 136
rect 2643 102 2731 136
rect 2765 102 2781 136
rect 2607 17 2781 102
rect 2817 120 2851 176
rect 2817 70 2851 86
rect 2887 210 2953 226
rect 2887 176 2903 210
rect 2937 176 2953 210
rect 2887 120 2953 176
rect 2887 86 2903 120
rect 2937 86 2953 120
rect 2887 17 2953 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 2976 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 799 416 833 424
rect 799 390 807 416
rect 807 390 833 416
rect 1567 414 1601 424
rect 1567 390 1579 414
rect 1579 390 1601 414
rect 2143 414 2177 424
rect 2143 390 2167 414
rect 2167 390 2177 414
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
<< metal1 >>
rect 0 683 2976 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 2976 683
rect 0 617 2976 649
rect 787 424 845 430
rect 787 390 799 424
rect 833 421 845 424
rect 1555 424 1613 430
rect 1555 421 1567 424
rect 833 393 1567 421
rect 833 390 845 393
rect 787 384 845 390
rect 1555 390 1567 393
rect 1601 421 1613 424
rect 2131 424 2189 430
rect 2131 421 2143 424
rect 1601 393 2143 421
rect 1601 390 1613 393
rect 1555 384 1613 390
rect 2131 390 2143 393
rect 2177 390 2189 424
rect 2131 384 2189 390
rect 0 17 2976 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 2976 17
rect 0 -49 2976 -17
<< labels >>
flabel pwell s 0 0 2976 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 0 617 2976 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel comment s 1485 630 1485 630 0 FreeSans 300 0 0 0 no_jumper_check
rlabel comment s 0 0 0 0 4 sdfrtp_4
flabel comment s 1108 36 1108 36 0 FreeSans 300 0 0 0 no_jumper_check
flabel metal1 s 2143 390 2177 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew
flabel metal1 s 0 0 2976 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel metal1 s 0 617 2976 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel corelocali s 319 168 353 202 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 SCD
port 4 nsew
flabel corelocali s 607 390 641 424 0 FreeSans 340 0 0 0 SCD
port 4 nsew
flabel corelocali s 799 242 833 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 2911 316 2945 350 0 FreeSans 340 0 0 0 Q
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 2976 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 189334
string GDS_START 168064
<< end >>
