magic
tech sky130A
magscale 1 2
timestamp 1599588238
<< locali >>
rect 121 378 209 596
rect 347 378 451 596
rect 121 344 451 378
rect 21 236 167 310
rect 203 88 269 310
rect 313 236 383 310
rect 417 202 451 344
rect 342 168 451 202
rect 342 70 408 168
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 37 364 87 649
rect 243 412 309 649
rect 64 17 130 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< metal1 >>
rect 0 683 480 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 0 617 480 649
rect 0 17 480 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
rect 0 -49 480 -17
<< labels >>
rlabel locali s 313 236 383 310 6 A
port 1 nsew signal input
rlabel locali s 203 88 269 310 6 B
port 2 nsew signal input
rlabel locali s 21 236 167 310 6 C
port 3 nsew signal input
rlabel locali s 417 202 451 344 6 Y
port 4 nsew signal output
rlabel locali s 347 378 451 596 6 Y
port 4 nsew signal output
rlabel locali s 342 168 451 202 6 Y
port 4 nsew signal output
rlabel locali s 342 70 408 168 6 Y
port 4 nsew signal output
rlabel locali s 121 378 209 596 6 Y
port 4 nsew signal output
rlabel locali s 121 344 451 378 6 Y
port 4 nsew signal output
rlabel metal1 s 0 -49 480 49 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 617 480 715 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 480 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1801126
string GDS_START 1795802
<< end >>
