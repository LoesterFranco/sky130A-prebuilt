magic
tech sky130A
magscale 1 2
timestamp 1604502701
<< nwell >>
rect -38 352 1862 704
rect -38 332 344 352
rect 1194 332 1862 352
<< pwell >>
rect 0 0 1824 49
<< scpmos >>
rect 86 392 116 592
rect 196 392 226 592
rect 442 388 472 588
rect 566 388 596 588
rect 660 388 690 588
rect 756 388 786 588
rect 866 388 896 588
rect 956 388 986 588
rect 1230 388 1260 588
rect 1331 368 1361 568
rect 1438 368 1468 592
rect 1528 368 1558 592
rect 1618 368 1648 592
rect 1708 368 1738 592
<< nmoslvt >>
rect 84 74 114 202
rect 170 74 200 202
rect 483 140 513 268
rect 569 140 599 268
rect 655 140 685 268
rect 741 140 771 268
rect 953 137 983 265
rect 1039 137 1069 265
rect 1237 94 1267 222
rect 1323 94 1353 222
rect 1423 74 1453 222
rect 1509 74 1539 222
rect 1615 74 1645 222
rect 1709 74 1739 222
<< ndiff >>
rect 412 254 483 268
rect 412 220 424 254
rect 458 220 483 254
rect 27 190 84 202
rect 27 156 39 190
rect 73 156 84 190
rect 27 120 84 156
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 184 170 202
rect 114 150 125 184
rect 159 150 170 184
rect 114 116 170 150
rect 114 82 125 116
rect 159 82 170 116
rect 114 74 170 82
rect 200 188 271 202
rect 200 154 225 188
rect 259 154 271 188
rect 200 142 271 154
rect 200 74 250 142
rect 412 140 483 220
rect 513 254 569 268
rect 513 220 524 254
rect 558 220 569 254
rect 513 140 569 220
rect 599 228 655 268
rect 599 194 610 228
rect 644 194 655 228
rect 599 140 655 194
rect 685 201 741 268
rect 685 167 696 201
rect 730 167 741 201
rect 685 140 741 167
rect 771 254 828 268
rect 771 220 782 254
rect 816 220 828 254
rect 771 140 828 220
rect 882 253 953 265
rect 882 219 894 253
rect 928 219 953 253
rect 882 137 953 219
rect 983 185 1039 265
rect 983 151 994 185
rect 1028 151 1039 185
rect 983 137 1039 151
rect 1069 256 1126 265
rect 1069 222 1080 256
rect 1114 222 1126 256
rect 1069 183 1126 222
rect 1069 149 1080 183
rect 1114 149 1126 183
rect 1069 137 1126 149
rect 1180 146 1237 222
rect 1180 112 1192 146
rect 1226 112 1237 146
rect 1180 94 1237 112
rect 1267 210 1323 222
rect 1267 176 1278 210
rect 1312 176 1323 210
rect 1267 140 1323 176
rect 1267 106 1278 140
rect 1312 106 1323 140
rect 1267 94 1323 106
rect 1353 210 1423 222
rect 1353 176 1364 210
rect 1398 176 1423 210
rect 1353 140 1423 176
rect 1353 106 1364 140
rect 1398 106 1423 140
rect 1353 94 1423 106
rect 1373 74 1423 94
rect 1453 210 1509 222
rect 1453 176 1464 210
rect 1498 176 1509 210
rect 1453 120 1509 176
rect 1453 86 1464 120
rect 1498 86 1509 120
rect 1453 74 1509 86
rect 1539 146 1615 222
rect 1539 112 1564 146
rect 1598 112 1615 146
rect 1539 74 1615 112
rect 1645 207 1709 222
rect 1645 173 1664 207
rect 1698 173 1709 207
rect 1645 74 1709 173
rect 1739 120 1797 222
rect 1739 86 1750 120
rect 1784 86 1797 120
rect 1739 74 1797 86
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 510 86 546
rect 27 476 39 510
rect 73 476 86 510
rect 27 440 86 476
rect 27 406 39 440
rect 73 406 86 440
rect 27 392 86 406
rect 116 580 196 592
rect 116 546 139 580
rect 173 546 196 580
rect 116 508 196 546
rect 116 474 139 508
rect 173 474 196 508
rect 116 392 196 474
rect 226 580 285 592
rect 226 546 239 580
rect 273 546 285 580
rect 226 508 285 546
rect 226 474 239 508
rect 273 474 285 508
rect 226 392 285 474
rect 378 567 442 588
rect 378 533 394 567
rect 428 533 442 567
rect 378 388 442 533
rect 472 576 566 588
rect 472 542 502 576
rect 536 542 566 576
rect 472 505 566 542
rect 472 471 502 505
rect 536 471 566 505
rect 472 434 566 471
rect 472 400 502 434
rect 536 400 566 434
rect 472 388 566 400
rect 596 576 660 588
rect 596 542 609 576
rect 643 542 660 576
rect 596 506 660 542
rect 596 472 609 506
rect 643 472 660 506
rect 596 437 660 472
rect 596 403 609 437
rect 643 403 660 437
rect 596 388 660 403
rect 690 576 756 588
rect 690 542 709 576
rect 743 542 756 576
rect 690 505 756 542
rect 690 471 709 505
rect 743 471 756 505
rect 690 434 756 471
rect 690 400 709 434
rect 743 400 756 434
rect 690 388 756 400
rect 786 576 866 588
rect 786 542 809 576
rect 843 542 866 576
rect 786 506 866 542
rect 786 472 809 506
rect 843 472 866 506
rect 786 437 866 472
rect 786 403 809 437
rect 843 403 866 437
rect 786 388 866 403
rect 896 576 956 588
rect 896 542 909 576
rect 943 542 956 576
rect 896 505 956 542
rect 896 471 909 505
rect 943 471 956 505
rect 896 434 956 471
rect 896 400 909 434
rect 943 400 956 434
rect 896 388 956 400
rect 986 576 1230 588
rect 986 542 1009 576
rect 1043 542 1096 576
rect 1130 542 1183 576
rect 1217 542 1230 576
rect 986 492 1230 542
rect 986 458 1009 492
rect 1043 458 1096 492
rect 1130 458 1183 492
rect 1217 458 1230 492
rect 986 388 1230 458
rect 1260 568 1313 588
rect 1379 580 1438 592
rect 1379 568 1391 580
rect 1260 556 1331 568
rect 1260 522 1283 556
rect 1317 522 1331 556
rect 1260 430 1331 522
rect 1260 396 1283 430
rect 1317 396 1331 430
rect 1260 388 1331 396
rect 1278 368 1331 388
rect 1361 546 1391 568
rect 1425 546 1438 580
rect 1361 508 1438 546
rect 1361 474 1391 508
rect 1425 474 1438 508
rect 1361 368 1438 474
rect 1468 580 1528 592
rect 1468 546 1481 580
rect 1515 546 1528 580
rect 1468 497 1528 546
rect 1468 463 1481 497
rect 1515 463 1528 497
rect 1468 414 1528 463
rect 1468 380 1481 414
rect 1515 380 1528 414
rect 1468 368 1528 380
rect 1558 584 1618 592
rect 1558 550 1571 584
rect 1605 550 1618 584
rect 1558 498 1618 550
rect 1558 464 1571 498
rect 1605 464 1618 498
rect 1558 368 1618 464
rect 1648 414 1708 592
rect 1648 380 1661 414
rect 1695 380 1708 414
rect 1648 368 1708 380
rect 1738 580 1797 592
rect 1738 546 1751 580
rect 1785 546 1797 580
rect 1738 498 1797 546
rect 1738 464 1751 498
rect 1785 464 1797 498
rect 1738 368 1797 464
<< ndiffc >>
rect 424 220 458 254
rect 39 156 73 190
rect 39 86 73 120
rect 125 150 159 184
rect 125 82 159 116
rect 225 154 259 188
rect 524 220 558 254
rect 610 194 644 228
rect 696 167 730 201
rect 782 220 816 254
rect 894 219 928 253
rect 994 151 1028 185
rect 1080 222 1114 256
rect 1080 149 1114 183
rect 1192 112 1226 146
rect 1278 176 1312 210
rect 1278 106 1312 140
rect 1364 176 1398 210
rect 1364 106 1398 140
rect 1464 176 1498 210
rect 1464 86 1498 120
rect 1564 112 1598 146
rect 1664 173 1698 207
rect 1750 86 1784 120
<< pdiffc >>
rect 39 546 73 580
rect 39 476 73 510
rect 39 406 73 440
rect 139 546 173 580
rect 139 474 173 508
rect 239 546 273 580
rect 239 474 273 508
rect 394 533 428 567
rect 502 542 536 576
rect 502 471 536 505
rect 502 400 536 434
rect 609 542 643 576
rect 609 472 643 506
rect 609 403 643 437
rect 709 542 743 576
rect 709 471 743 505
rect 709 400 743 434
rect 809 542 843 576
rect 809 472 843 506
rect 809 403 843 437
rect 909 542 943 576
rect 909 471 943 505
rect 909 400 943 434
rect 1009 542 1043 576
rect 1096 542 1130 576
rect 1183 542 1217 576
rect 1009 458 1043 492
rect 1096 458 1130 492
rect 1183 458 1217 492
rect 1283 522 1317 556
rect 1283 396 1317 430
rect 1391 546 1425 580
rect 1391 474 1425 508
rect 1481 546 1515 580
rect 1481 463 1515 497
rect 1481 380 1515 414
rect 1571 550 1605 584
rect 1571 464 1605 498
rect 1661 380 1695 414
rect 1751 546 1785 580
rect 1751 464 1785 498
<< poly >>
rect 86 592 116 618
rect 196 592 226 618
rect 442 588 472 614
rect 566 588 596 614
rect 660 588 690 614
rect 756 588 786 614
rect 866 588 896 614
rect 956 588 986 614
rect 1230 588 1260 614
rect 86 377 116 392
rect 196 377 226 392
rect 1331 568 1361 594
rect 1438 592 1468 618
rect 1528 592 1558 618
rect 1618 592 1648 618
rect 1708 592 1738 618
rect 83 356 116 377
rect 193 356 229 377
rect 442 373 472 388
rect 566 373 596 388
rect 660 373 690 388
rect 756 373 786 388
rect 866 373 896 388
rect 956 373 986 388
rect 1230 373 1260 388
rect 439 356 475 373
rect 563 356 599 373
rect 48 340 114 356
rect 48 306 64 340
rect 98 306 114 340
rect 48 290 114 306
rect 84 202 114 290
rect 170 340 267 356
rect 170 306 217 340
rect 251 306 267 340
rect 170 290 267 306
rect 386 340 599 356
rect 386 306 402 340
rect 436 306 599 340
rect 657 313 693 373
rect 753 313 789 373
rect 170 202 200 290
rect 386 284 599 306
rect 483 268 513 284
rect 569 268 599 284
rect 655 283 693 313
rect 741 283 789 313
rect 863 356 899 373
rect 953 356 989 373
rect 863 340 1127 356
rect 863 306 1009 340
rect 1043 306 1077 340
rect 1111 306 1127 340
rect 863 290 1127 306
rect 1227 336 1263 373
rect 1331 353 1361 368
rect 1438 353 1468 368
rect 1528 353 1558 368
rect 1618 353 1648 368
rect 1708 353 1738 368
rect 1328 336 1364 353
rect 1227 320 1375 336
rect 655 268 685 283
rect 741 268 771 283
rect 953 265 983 290
rect 1039 265 1069 290
rect 1227 286 1325 320
rect 1359 286 1375 320
rect 1435 330 1471 353
rect 1525 330 1561 353
rect 1615 330 1651 353
rect 1705 330 1739 353
rect 1435 314 1739 330
rect 1435 294 1459 314
rect 1227 270 1375 286
rect 1423 280 1459 294
rect 1493 280 1527 314
rect 1561 280 1595 314
rect 1629 280 1663 314
rect 1697 280 1739 314
rect 272 101 338 117
rect 483 114 513 140
rect 84 48 114 74
rect 170 48 200 74
rect 272 67 288 101
rect 322 67 338 101
rect 272 66 338 67
rect 569 66 599 140
rect 272 36 599 66
rect 655 117 685 140
rect 741 117 771 140
rect 1237 222 1267 270
rect 1323 222 1353 270
rect 1423 264 1739 280
rect 1423 222 1453 264
rect 1509 222 1539 264
rect 1615 222 1645 264
rect 1709 222 1739 264
rect 655 101 771 117
rect 953 111 983 137
rect 1039 111 1069 137
rect 655 67 671 101
rect 705 87 771 101
rect 705 67 721 87
rect 1237 68 1267 94
rect 1323 68 1353 94
rect 655 51 721 67
rect 1423 48 1453 74
rect 1509 48 1539 74
rect 1615 48 1645 74
rect 1709 48 1739 74
<< polycont >>
rect 64 306 98 340
rect 217 306 251 340
rect 402 306 436 340
rect 1009 306 1043 340
rect 1077 306 1111 340
rect 1325 286 1359 320
rect 1459 280 1493 314
rect 1527 280 1561 314
rect 1595 280 1629 314
rect 1663 280 1697 314
rect 288 67 322 101
rect 671 67 705 101
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 23 580 89 596
rect 23 546 39 580
rect 73 546 89 580
rect 23 510 89 546
rect 23 476 39 510
rect 73 476 89 510
rect 23 440 89 476
rect 123 580 189 649
rect 123 546 139 580
rect 173 546 189 580
rect 123 508 189 546
rect 123 474 139 508
rect 173 474 189 508
rect 123 458 189 474
rect 223 580 289 596
rect 223 546 239 580
rect 273 546 289 580
rect 223 508 289 546
rect 378 567 445 649
rect 378 533 394 567
rect 428 533 445 567
rect 378 526 445 533
rect 486 576 552 592
rect 486 542 502 576
rect 536 542 552 576
rect 223 474 239 508
rect 273 492 289 508
rect 486 505 552 542
rect 273 474 452 492
rect 223 458 452 474
rect 23 406 39 440
rect 73 424 89 440
rect 73 406 335 424
rect 23 390 335 406
rect 25 340 167 356
rect 25 306 64 340
rect 98 306 167 340
rect 25 290 167 306
rect 201 340 267 356
rect 201 306 217 340
rect 251 306 267 340
rect 201 290 267 306
rect 301 256 335 390
rect 386 340 452 458
rect 386 306 402 340
rect 436 306 452 340
rect 486 471 502 505
rect 536 471 552 505
rect 486 434 552 471
rect 486 400 502 434
rect 536 400 552 434
rect 486 353 552 400
rect 593 576 659 649
rect 593 542 609 576
rect 643 542 659 576
rect 593 506 659 542
rect 593 472 609 506
rect 643 472 659 506
rect 593 437 659 472
rect 593 403 609 437
rect 643 403 659 437
rect 593 387 659 403
rect 693 576 759 592
rect 693 542 709 576
rect 743 542 759 576
rect 693 505 759 542
rect 693 471 709 505
rect 743 471 759 505
rect 693 434 759 471
rect 693 400 709 434
rect 743 400 759 434
rect 693 353 759 400
rect 793 576 859 649
rect 793 542 809 576
rect 843 542 859 576
rect 793 506 859 542
rect 793 472 809 506
rect 843 472 859 506
rect 793 437 859 472
rect 793 403 809 437
rect 843 403 859 437
rect 793 387 859 403
rect 893 576 959 592
rect 893 542 909 576
rect 943 542 959 576
rect 893 505 959 542
rect 893 471 909 505
rect 943 471 959 505
rect 893 434 959 471
rect 993 576 1233 649
rect 993 542 1009 576
rect 1043 542 1096 576
rect 1130 542 1183 576
rect 1217 542 1233 576
rect 1375 580 1441 649
rect 993 492 1233 542
rect 993 458 1009 492
rect 1043 458 1096 492
rect 1130 458 1183 492
rect 1217 458 1233 492
rect 1267 556 1333 572
rect 1267 522 1283 556
rect 1317 522 1333 556
rect 893 400 909 434
rect 943 424 959 434
rect 1267 430 1333 522
rect 1375 546 1391 580
rect 1425 546 1441 580
rect 1375 508 1441 546
rect 1375 474 1391 508
rect 1425 474 1441 508
rect 1375 458 1441 474
rect 1481 580 1515 596
rect 1481 497 1515 546
rect 1555 584 1621 649
rect 1555 550 1571 584
rect 1605 550 1621 584
rect 1555 498 1621 550
rect 1555 464 1571 498
rect 1605 464 1621 498
rect 1735 580 1801 649
rect 1735 546 1751 580
rect 1785 546 1801 580
rect 1735 498 1801 546
rect 1735 464 1751 498
rect 1785 464 1801 498
rect 1267 424 1283 430
rect 943 400 1283 424
rect 893 396 1283 400
rect 1317 424 1333 430
rect 1481 430 1515 463
rect 1317 396 1447 424
rect 893 390 1447 396
rect 893 353 959 390
rect 486 319 959 353
rect 993 340 1223 356
rect 386 290 452 306
rect 508 272 552 319
rect 993 306 1009 340
rect 1043 306 1077 340
rect 1111 306 1223 340
rect 993 290 1223 306
rect 1273 320 1375 356
rect 1273 286 1325 320
rect 1359 286 1375 320
rect 23 222 374 256
rect 23 190 73 222
rect 23 156 39 190
rect 23 120 73 156
rect 23 86 39 120
rect 23 70 73 86
rect 109 184 175 188
rect 109 150 125 184
rect 159 150 175 184
rect 109 116 175 150
rect 109 82 125 116
rect 159 82 175 116
rect 109 17 175 82
rect 209 154 225 188
rect 259 154 306 188
rect 209 117 306 154
rect 340 185 374 222
rect 408 254 474 256
rect 408 220 424 254
rect 458 220 474 254
rect 408 219 474 220
rect 508 254 574 272
rect 508 220 524 254
rect 558 220 574 254
rect 508 219 574 220
rect 610 254 832 285
rect 1273 270 1375 286
rect 1413 330 1447 390
rect 1481 414 1799 430
rect 1515 380 1661 414
rect 1695 380 1799 414
rect 1481 364 1799 380
rect 1413 314 1713 330
rect 1413 280 1459 314
rect 1493 280 1527 314
rect 1561 280 1595 314
rect 1629 280 1663 314
rect 1697 280 1713 314
rect 610 251 782 254
rect 610 228 644 251
rect 440 185 474 219
rect 766 220 782 251
rect 816 220 832 254
rect 766 219 832 220
rect 878 256 944 269
rect 1413 264 1713 280
rect 878 253 1080 256
rect 878 219 894 253
rect 928 222 1080 253
rect 1114 236 1130 256
rect 1114 222 1312 236
rect 1753 230 1799 364
rect 928 219 944 222
rect 610 185 644 194
rect 340 151 406 185
rect 440 151 644 185
rect 680 201 730 217
rect 680 167 696 201
rect 1080 210 1312 222
rect 1080 202 1278 210
rect 978 185 1044 188
rect 730 167 994 185
rect 680 151 994 167
rect 1028 151 1044 185
rect 372 117 406 151
rect 978 133 1044 151
rect 1080 183 1130 202
rect 1114 149 1130 183
rect 1262 176 1278 202
rect 1080 133 1130 149
rect 1176 146 1226 168
rect 209 101 338 117
rect 209 67 288 101
rect 322 67 338 101
rect 209 51 338 67
rect 372 101 721 117
rect 372 67 671 101
rect 705 67 721 101
rect 372 51 721 67
rect 1176 112 1192 146
rect 1176 17 1226 112
rect 1262 140 1312 176
rect 1262 106 1278 140
rect 1262 90 1312 106
rect 1348 210 1414 226
rect 1348 176 1364 210
rect 1398 176 1414 210
rect 1348 140 1414 176
rect 1348 106 1364 140
rect 1398 106 1414 140
rect 1348 17 1414 106
rect 1448 210 1799 230
rect 1448 176 1464 210
rect 1498 207 1799 210
rect 1498 196 1664 207
rect 1498 176 1514 196
rect 1448 120 1514 176
rect 1648 173 1664 196
rect 1698 173 1799 207
rect 1448 86 1464 120
rect 1498 86 1514 120
rect 1448 70 1514 86
rect 1548 146 1614 162
rect 1648 154 1799 173
rect 1548 112 1564 146
rect 1598 112 1614 146
rect 1548 17 1614 112
rect 1734 86 1750 120
rect 1784 86 1801 120
rect 1734 17 1801 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
<< metal1 >>
rect 0 683 1824 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 0 617 1824 649
rect 0 17 1824 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
rect 0 -49 1824 -17
<< labels >>
rlabel comment s 0 0 0 0 4 and4bb_4
flabel comment s 575 313 575 313 0 FreeSans 200 0 0 0 no_jumper_check
flabel pwell s 0 0 1824 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 1824 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 1824 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 1824 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 B_N
port 2 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 B_N
port 2 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew
flabel corelocali s 1279 316 1313 350 0 FreeSans 340 0 0 0 D
port 4 nsew
flabel corelocali s 1087 316 1121 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 1183 316 1217 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 1759 168 1793 202 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 1759 242 1793 276 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 1759 316 1793 350 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 1759 390 1793 424 0 FreeSans 340 0 0 0 X
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 1824 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3317970
string GDS_START 3303446
<< end >>
