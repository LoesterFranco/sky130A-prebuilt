magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 207 325 275 493
rect 413 325 463 493
rect 715 325 765 425
rect 903 325 953 425
rect 207 291 953 325
rect 539 289 953 291
rect 17 215 102 257
rect 539 215 639 289
rect 673 215 995 255
rect 1029 215 1450 257
rect 539 163 585 215
rect 304 129 585 163
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 29 325 95 487
rect 139 359 173 527
rect 319 359 369 527
rect 507 359 557 527
rect 605 459 1047 493
rect 605 359 671 459
rect 809 359 859 459
rect 29 291 170 325
rect 997 325 1047 459
rect 1091 359 1141 527
rect 1185 325 1235 493
rect 1279 359 1329 527
rect 1373 325 1423 493
rect 997 291 1423 325
rect 136 257 170 291
rect 136 215 505 257
rect 136 179 189 215
rect 45 17 79 179
rect 113 58 189 179
rect 629 145 1431 181
rect 629 95 679 145
rect 236 61 679 95
rect 723 17 757 111
rect 791 51 867 145
rect 911 17 945 111
rect 979 51 1055 145
rect 1099 17 1133 111
rect 1167 51 1243 145
rect 1287 17 1321 111
rect 1355 51 1431 145
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< labels >>
rlabel locali s 1029 215 1450 257 6 A1
port 1 nsew signal input
rlabel locali s 673 215 995 255 6 A2
port 2 nsew signal input
rlabel locali s 17 215 102 257 6 B1_N
port 3 nsew signal input
rlabel locali s 903 325 953 425 6 Y
port 4 nsew signal output
rlabel locali s 715 325 765 425 6 Y
port 4 nsew signal output
rlabel locali s 539 289 953 291 6 Y
port 4 nsew signal output
rlabel locali s 539 215 639 289 6 Y
port 4 nsew signal output
rlabel locali s 539 163 585 215 6 Y
port 4 nsew signal output
rlabel locali s 413 325 463 493 6 Y
port 4 nsew signal output
rlabel locali s 304 129 585 163 6 Y
port 4 nsew signal output
rlabel locali s 207 325 275 493 6 Y
port 4 nsew signal output
rlabel locali s 207 291 953 325 6 Y
port 4 nsew signal output
rlabel metal1 s 0 -48 1472 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 1472 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1472 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1047426
string GDS_START 1036122
<< end >>
