magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1288 561
rect 103 427 169 527
rect 18 197 66 325
rect 103 17 169 93
rect 391 367 450 527
rect 750 435 818 527
rect 856 427 912 527
rect 288 191 354 265
rect 1028 375 1097 527
rect 1131 375 1185 493
rect 1151 300 1185 375
rect 1219 334 1271 527
rect 1151 285 1271 300
rect 1152 283 1271 285
rect 1153 282 1271 283
rect 1155 277 1271 282
rect 896 207 1048 265
rect 896 199 963 207
rect 1157 178 1271 277
rect 1154 173 1271 178
rect 375 17 441 89
rect 1151 153 1271 173
rect 744 17 812 106
rect 1051 17 1085 105
rect 1151 97 1185 153
rect 1119 51 1185 97
rect 1219 17 1271 119
rect 0 -17 1288 17
<< obsli1 >>
rect 35 393 69 493
rect 35 359 156 393
rect 122 323 156 359
rect 122 280 156 289
rect 203 391 248 493
rect 203 357 214 391
rect 203 337 248 357
rect 122 214 168 280
rect 122 161 156 214
rect 17 127 156 161
rect 17 69 69 127
rect 203 69 237 337
rect 287 333 357 483
rect 554 451 716 485
rect 682 417 716 451
rect 682 400 721 417
rect 683 399 721 400
rect 581 391 635 399
rect 684 397 721 399
rect 581 357 585 391
rect 619 382 635 391
rect 619 357 653 382
rect 581 356 653 357
rect 287 299 424 333
rect 390 219 424 299
rect 490 323 551 337
rect 524 289 551 323
rect 490 271 551 289
rect 586 314 653 356
rect 390 157 467 219
rect 586 208 620 314
rect 687 265 721 397
rect 960 373 994 493
rect 755 341 994 373
rect 755 307 1117 341
rect 1083 265 1117 307
rect 303 153 467 157
rect 303 123 424 153
rect 517 147 620 208
rect 654 199 844 265
rect 1083 199 1123 265
rect 303 69 341 123
rect 654 107 689 199
rect 1083 173 1117 199
rect 991 165 1117 173
rect 554 73 689 107
rect 848 139 1117 165
rect 848 131 1019 139
rect 848 51 916 131
<< obsli1c >>
rect 122 289 156 323
rect 214 357 248 391
rect 585 357 619 391
rect 490 289 524 323
<< metal1 >>
rect 0 496 1288 592
rect 0 -48 1288 48
<< obsm1 >>
rect 202 391 260 397
rect 202 357 214 391
rect 248 388 260 391
rect 573 391 631 397
rect 573 388 585 391
rect 248 360 585 388
rect 248 357 260 360
rect 202 351 260 357
rect 573 357 585 360
rect 619 357 631 391
rect 573 351 631 357
rect 110 323 168 329
rect 110 289 122 323
rect 156 320 168 323
rect 478 323 536 329
rect 478 320 490 323
rect 156 292 490 320
rect 156 289 168 292
rect 110 283 168 289
rect 478 289 490 292
rect 524 289 536 323
rect 478 283 536 289
<< labels >>
rlabel locali s 288 191 354 265 6 D
port 1 nsew signal input
rlabel locali s 1157 178 1271 277 6 Q
port 2 nsew signal output
rlabel locali s 1155 277 1271 282 6 Q
port 2 nsew signal output
rlabel locali s 1154 173 1271 178 6 Q
port 2 nsew signal output
rlabel locali s 1153 282 1271 283 6 Q
port 2 nsew signal output
rlabel locali s 1152 283 1271 285 6 Q
port 2 nsew signal output
rlabel locali s 1151 300 1185 375 6 Q
port 2 nsew signal output
rlabel locali s 1151 285 1271 300 6 Q
port 2 nsew signal output
rlabel locali s 1151 153 1271 173 6 Q
port 2 nsew signal output
rlabel locali s 1151 97 1185 153 6 Q
port 2 nsew signal output
rlabel locali s 1131 375 1185 493 6 Q
port 2 nsew signal output
rlabel locali s 1119 51 1185 97 6 Q
port 2 nsew signal output
rlabel locali s 896 207 1048 265 6 RESET_B
port 3 nsew signal input
rlabel locali s 896 199 963 207 6 RESET_B
port 3 nsew signal input
rlabel locali s 18 197 66 325 6 GATE
port 4 nsew clock input
rlabel locali s 1219 17 1271 119 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 1051 17 1085 105 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 744 17 812 106 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 375 17 441 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 103 17 169 93 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 1288 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1288 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 1219 334 1271 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 1028 375 1097 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 856 427 912 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 750 435 818 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 391 367 450 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 103 427 169 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 1288 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 1288 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1288 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2683818
string GDS_START 2672624
<< end >>
