magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 902 704
<< pwell >>
rect 0 0 864 49
<< scnmos >>
rect 97 74 127 222
rect 185 74 215 222
rect 325 74 355 222
rect 403 74 433 222
rect 517 74 547 222
rect 631 74 661 222
rect 745 74 775 222
<< pmoshvt >>
rect 86 368 116 592
rect 176 368 206 592
rect 316 368 346 568
rect 406 368 436 568
rect 548 368 578 568
rect 638 368 668 568
rect 748 368 778 568
<< ndiff >>
rect 27 210 97 222
rect 27 176 39 210
rect 73 176 97 210
rect 27 120 97 176
rect 27 86 39 120
rect 73 86 97 120
rect 27 74 97 86
rect 127 214 185 222
rect 127 180 139 214
rect 173 180 185 214
rect 127 116 185 180
rect 127 82 139 116
rect 173 82 185 116
rect 127 74 185 82
rect 215 152 325 222
rect 215 118 253 152
rect 287 118 325 152
rect 215 74 325 118
rect 355 74 403 222
rect 433 74 517 222
rect 547 210 631 222
rect 547 176 571 210
rect 605 176 631 210
rect 547 120 631 176
rect 547 86 571 120
rect 605 86 631 120
rect 547 74 631 86
rect 661 74 745 222
rect 775 210 832 222
rect 775 176 786 210
rect 820 176 832 210
rect 775 120 832 176
rect 775 86 786 120
rect 820 86 832 120
rect 775 74 832 86
<< pdiff >>
rect 27 573 86 592
rect 27 539 39 573
rect 73 539 86 573
rect 27 368 86 539
rect 116 414 176 592
rect 116 380 129 414
rect 163 380 176 414
rect 116 368 176 380
rect 206 582 298 592
rect 206 548 244 582
rect 278 568 298 582
rect 278 548 316 568
rect 206 368 316 548
rect 346 560 406 568
rect 346 526 359 560
rect 393 526 406 560
rect 346 492 406 526
rect 346 458 359 492
rect 393 458 406 492
rect 346 368 406 458
rect 436 560 548 568
rect 436 526 475 560
rect 509 526 548 560
rect 436 368 548 526
rect 578 560 638 568
rect 578 526 591 560
rect 625 526 638 560
rect 578 492 638 526
rect 578 458 591 492
rect 625 458 638 492
rect 578 368 638 458
rect 668 539 748 568
rect 668 505 691 539
rect 725 505 748 539
rect 668 430 748 505
rect 668 396 691 430
rect 725 396 748 430
rect 668 368 748 396
rect 778 556 837 568
rect 778 522 791 556
rect 825 522 837 556
rect 778 430 837 522
rect 778 396 791 430
rect 825 396 837 430
rect 778 368 837 396
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 139 180 173 214
rect 139 82 173 116
rect 253 118 287 152
rect 571 176 605 210
rect 571 86 605 120
rect 786 176 820 210
rect 786 86 820 120
<< pdiffc >>
rect 39 539 73 573
rect 129 380 163 414
rect 244 548 278 582
rect 359 526 393 560
rect 359 458 393 492
rect 475 526 509 560
rect 591 526 625 560
rect 591 458 625 492
rect 691 505 725 539
rect 691 396 725 430
rect 791 522 825 556
rect 791 396 825 430
<< poly >>
rect 86 592 116 618
rect 176 592 206 618
rect 316 568 346 594
rect 406 568 436 594
rect 548 568 578 594
rect 638 568 668 594
rect 748 568 778 594
rect 86 353 116 368
rect 176 353 206 368
rect 316 353 346 368
rect 406 353 436 368
rect 548 353 578 368
rect 638 353 668 368
rect 748 353 778 368
rect 83 330 119 353
rect 173 330 209 353
rect 313 336 349 353
rect 403 336 439 353
rect 545 336 581 353
rect 635 336 671 353
rect 45 314 209 330
rect 45 280 61 314
rect 95 294 209 314
rect 289 320 355 336
rect 95 280 215 294
rect 45 264 215 280
rect 289 286 305 320
rect 339 286 355 320
rect 289 270 355 286
rect 97 222 127 264
rect 185 222 215 264
rect 325 222 355 270
rect 403 320 469 336
rect 403 286 419 320
rect 453 286 469 320
rect 403 270 469 286
rect 517 320 583 336
rect 517 286 533 320
rect 567 286 583 320
rect 517 270 583 286
rect 631 320 697 336
rect 631 286 647 320
rect 681 286 697 320
rect 631 270 697 286
rect 745 326 781 353
rect 745 310 843 326
rect 745 276 793 310
rect 827 276 843 310
rect 403 222 433 270
rect 517 222 547 270
rect 631 222 661 270
rect 745 260 843 276
rect 745 222 775 260
rect 97 48 127 74
rect 185 48 215 74
rect 325 48 355 74
rect 403 48 433 74
rect 517 48 547 74
rect 631 48 661 74
rect 745 48 775 74
<< polycont >>
rect 61 280 95 314
rect 305 286 339 320
rect 419 286 453 320
rect 533 286 567 320
rect 647 286 681 320
rect 793 276 827 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 23 573 89 649
rect 23 539 39 573
rect 73 539 89 573
rect 23 532 89 539
rect 220 582 302 649
rect 220 548 244 582
rect 278 548 302 582
rect 220 532 302 548
rect 343 560 409 572
rect 343 526 359 560
rect 393 526 409 560
rect 453 560 529 649
rect 453 526 475 560
rect 509 526 529 560
rect 575 581 841 615
rect 575 560 641 581
rect 575 526 591 560
rect 625 526 641 560
rect 775 556 841 581
rect 45 464 255 498
rect 45 330 79 464
rect 113 414 187 430
rect 113 380 129 414
rect 163 380 187 414
rect 113 364 187 380
rect 45 314 111 330
rect 45 280 61 314
rect 95 280 111 314
rect 45 264 111 280
rect 145 230 187 364
rect 23 210 89 226
rect 23 176 39 210
rect 73 176 89 210
rect 23 120 89 176
rect 23 86 39 120
rect 73 86 89 120
rect 23 17 89 86
rect 123 214 187 230
rect 123 180 139 214
rect 173 180 187 214
rect 221 424 255 464
rect 343 492 409 526
rect 575 492 641 526
rect 343 458 359 492
rect 393 458 591 492
rect 625 458 641 492
rect 675 539 741 547
rect 675 505 691 539
rect 725 505 741 539
rect 675 430 741 505
rect 675 424 691 430
rect 221 396 691 424
rect 725 396 741 430
rect 221 390 741 396
rect 775 522 791 556
rect 825 522 841 556
rect 775 430 841 522
rect 775 396 791 430
rect 825 396 841 430
rect 775 390 841 396
rect 221 236 255 390
rect 289 320 355 356
rect 289 286 305 320
rect 339 286 355 320
rect 289 270 355 286
rect 403 320 469 356
rect 403 286 419 320
rect 453 286 469 320
rect 403 270 469 286
rect 505 320 583 356
rect 505 286 533 320
rect 567 286 583 320
rect 505 270 583 286
rect 631 320 743 356
rect 631 286 647 320
rect 681 286 743 320
rect 631 270 743 286
rect 777 310 843 356
rect 777 276 793 310
rect 827 276 843 310
rect 777 260 843 276
rect 221 210 621 236
rect 221 202 571 210
rect 123 116 187 180
rect 555 176 571 202
rect 605 176 621 210
rect 123 82 139 116
rect 173 82 187 116
rect 123 66 187 82
rect 237 152 303 168
rect 237 118 253 152
rect 287 118 303 152
rect 237 17 303 118
rect 555 120 621 176
rect 555 86 571 120
rect 605 86 621 120
rect 555 70 621 86
rect 770 210 836 226
rect 770 176 786 210
rect 820 176 836 210
rect 770 120 836 176
rect 770 86 786 120
rect 820 86 836 120
rect 770 17 836 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a32o_2
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 B2
port 5 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 B1
port 4 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 127 390 161 424 0 FreeSans 340 0 0 0 X
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 864 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3719660
string GDS_START 3712684
<< end >>
