magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 17 153 68 335
rect 208 153 297 335
rect 631 211 763 330
rect 2649 299 2731 490
rect 2670 165 2731 299
rect 2649 55 2731 165
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2852 561
rect 17 405 69 493
rect 103 439 167 527
rect 211 451 449 493
rect 211 405 245 451
rect 494 417 544 493
rect 588 428 647 527
rect 17 369 245 405
rect 279 369 369 417
rect 108 255 174 335
rect 108 221 128 255
rect 162 221 174 255
rect 108 153 174 221
rect 331 323 369 369
rect 331 289 335 323
rect 331 119 369 289
rect 413 354 544 417
rect 701 400 735 465
rect 769 455 845 527
rect 889 427 958 493
rect 701 391 859 400
rect 701 366 825 391
rect 807 357 825 366
rect 413 181 480 354
rect 514 255 590 320
rect 514 221 529 255
rect 563 221 590 255
rect 514 215 590 221
rect 413 143 544 181
rect 807 177 859 357
rect 17 17 150 119
rect 184 51 369 119
rect 405 17 458 109
rect 492 51 544 143
rect 704 143 859 177
rect 895 284 958 427
rect 993 323 1036 493
rect 1087 427 1241 493
rect 1289 455 1366 527
rect 993 318 1002 323
rect 1155 357 1173 391
rect 1121 315 1173 357
rect 895 254 968 284
rect 895 220 927 254
rect 961 220 968 254
rect 895 217 968 220
rect 588 17 670 111
rect 704 51 741 143
rect 785 17 851 109
rect 895 51 937 217
rect 1002 156 1036 289
rect 1207 279 1241 427
rect 1431 421 1484 490
rect 1542 425 1753 527
rect 1787 425 1968 492
rect 2012 447 2088 527
rect 1285 387 1484 421
rect 1934 413 1968 425
rect 2122 413 2203 490
rect 2241 447 2317 527
rect 1285 315 1319 387
rect 1577 357 1642 391
rect 1676 357 1777 391
rect 1438 323 1543 353
rect 1577 334 1777 357
rect 1438 289 1487 323
rect 1521 289 1543 323
rect 971 51 1036 156
rect 1093 255 1395 279
rect 1601 255 1683 265
rect 1093 245 1683 255
rect 1093 51 1178 245
rect 1219 161 1295 203
rect 1361 195 1683 245
rect 1717 181 1777 334
rect 1835 255 1900 381
rect 1934 379 2317 413
rect 1946 323 2199 345
rect 1946 289 1958 323
rect 1992 309 2199 323
rect 2241 321 2317 379
rect 1992 289 2007 309
rect 1946 285 2007 289
rect 2351 273 2403 493
rect 1835 221 1856 255
rect 1890 221 1900 255
rect 1835 215 1900 221
rect 1934 181 2001 251
rect 1219 127 1407 161
rect 1212 17 1319 93
rect 1357 51 1407 127
rect 1451 17 1683 161
rect 1717 144 2001 181
rect 2044 239 2403 273
rect 2044 171 2096 239
rect 2142 157 2323 203
rect 2142 109 2182 157
rect 2357 117 2403 239
rect 1853 55 2182 109
rect 2233 17 2283 109
rect 2335 51 2403 117
rect 2437 265 2505 493
rect 2553 369 2604 527
rect 2765 299 2799 527
rect 2437 199 2625 265
rect 2437 51 2489 199
rect 2523 17 2604 110
rect 2765 17 2799 177
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2852 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 128 221 162 255
rect 335 289 369 323
rect 825 357 859 391
rect 529 221 563 255
rect 1002 289 1036 323
rect 1121 357 1155 391
rect 927 220 961 254
rect 1642 357 1676 391
rect 1487 289 1521 323
rect 1958 289 1992 323
rect 1856 221 1890 255
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
<< metal1 >>
rect 0 561 2852 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2852 561
rect 0 496 2852 527
rect 1475 323 1543 329
rect 1475 289 1487 323
rect 1521 320 1543 323
rect 1946 323 2014 329
rect 1946 320 1958 323
rect 1521 292 1958 320
rect 1521 289 1543 292
rect 1475 283 1543 289
rect 1946 289 1958 292
rect 1992 289 2014 323
rect 1946 283 2014 289
rect 116 255 174 261
rect 116 221 128 255
rect 162 252 174 255
rect 517 255 575 261
rect 517 252 529 255
rect 162 224 529 252
rect 162 221 174 224
rect 116 215 174 221
rect 517 221 529 224
rect 563 221 575 255
rect 517 215 575 221
rect 0 17 2852 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2852 17
rect 0 -48 2852 -17
<< obsm1 >>
rect 813 391 881 397
rect 813 357 825 391
rect 859 388 881 391
rect 1109 391 1177 397
rect 1109 388 1121 391
rect 859 360 1121 388
rect 859 357 881 360
rect 813 351 881 357
rect 1109 357 1121 360
rect 1155 388 1177 391
rect 1630 391 1698 397
rect 1630 388 1642 391
rect 1155 360 1642 388
rect 1155 357 1177 360
rect 1109 351 1177 357
rect 1630 357 1642 360
rect 1676 357 1698 391
rect 1630 351 1698 357
rect 323 323 391 329
rect 323 289 335 323
rect 369 320 391 323
rect 990 323 1048 329
rect 990 320 1002 323
rect 369 292 1002 320
rect 369 289 391 292
rect 323 283 391 289
rect 990 289 1002 292
rect 1036 289 1048 323
rect 990 283 1048 289
rect 915 254 973 260
rect 915 220 927 254
rect 961 252 973 254
rect 1834 255 1912 261
rect 1834 252 1856 255
rect 961 224 1856 252
rect 961 220 973 224
rect 915 214 973 220
rect 1834 221 1856 224
rect 1890 221 1912 255
rect 1834 215 1912 221
<< labels >>
rlabel locali s 631 211 763 330 6 CLK
port 1 nsew signal input
rlabel locali s 208 153 297 335 6 D
port 2 nsew signal input
rlabel locali s 2670 165 2731 299 6 Q
port 3 nsew signal output
rlabel locali s 2649 299 2731 490 6 Q
port 3 nsew signal output
rlabel locali s 2649 55 2731 165 6 Q
port 3 nsew signal output
rlabel locali s 17 153 68 335 6 SCD
port 4 nsew signal input
rlabel metal1 s 517 252 575 261 6 SCE
port 5 nsew signal input
rlabel metal1 s 517 215 575 224 6 SCE
port 5 nsew signal input
rlabel metal1 s 116 252 174 261 6 SCE
port 5 nsew signal input
rlabel metal1 s 116 224 575 252 6 SCE
port 5 nsew signal input
rlabel metal1 s 116 215 174 224 6 SCE
port 5 nsew signal input
rlabel metal1 s 1946 320 2014 329 6 SET_B
port 6 nsew signal input
rlabel metal1 s 1946 283 2014 292 6 SET_B
port 6 nsew signal input
rlabel metal1 s 1475 320 1543 329 6 SET_B
port 6 nsew signal input
rlabel metal1 s 1475 292 2014 320 6 SET_B
port 6 nsew signal input
rlabel metal1 s 1475 283 1543 292 6 SET_B
port 6 nsew signal input
rlabel metal1 s 0 -48 2852 48 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 496 2852 592 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2852 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 263582
string GDS_START 243254
<< end >>
