magic
tech sky130A
magscale 1 2
timestamp 1599588201
<< nwell >>
rect -38 261 1510 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 260 47 290 119
rect 365 47 395 119
rect 487 47 517 131
rect 607 47 637 177
rect 795 47 825 131
rect 879 47 909 131
rect 1072 47 1102 131
rect 1144 47 1174 131
rect 1279 47 1309 177
rect 1363 47 1393 177
<< pmoshvt >>
rect 79 369 109 497
rect 151 369 181 497
rect 257 413 287 497
rect 353 413 383 497
rect 471 413 501 497
rect 607 297 637 497
rect 802 303 832 431
rect 912 303 942 431
rect 1100 369 1130 497
rect 1184 369 1214 497
rect 1279 297 1309 497
rect 1363 297 1393 497
<< ndiff >>
rect 27 103 79 131
rect 27 69 35 103
rect 69 69 79 103
rect 27 47 79 69
rect 109 89 163 131
rect 109 55 119 89
rect 153 55 163 89
rect 109 47 163 55
rect 193 119 245 131
rect 532 131 607 177
rect 437 119 487 131
rect 193 101 260 119
rect 193 67 203 101
rect 237 67 260 101
rect 193 47 260 67
rect 290 89 365 119
rect 290 55 310 89
rect 344 55 365 89
rect 290 47 365 55
rect 395 47 487 119
rect 517 119 607 131
rect 517 85 546 119
rect 580 85 607 119
rect 517 47 607 85
rect 637 101 689 177
rect 1229 131 1279 177
rect 637 67 647 101
rect 681 67 689 101
rect 637 47 689 67
rect 743 110 795 131
rect 743 76 751 110
rect 785 76 795 110
rect 743 47 795 76
rect 825 89 879 131
rect 825 55 835 89
rect 869 55 879 89
rect 825 47 879 55
rect 909 110 961 131
rect 909 76 919 110
rect 953 76 961 110
rect 909 47 961 76
rect 1020 109 1072 131
rect 1020 75 1028 109
rect 1062 75 1072 109
rect 1020 47 1072 75
rect 1102 47 1144 131
rect 1174 89 1279 131
rect 1174 55 1212 89
rect 1246 55 1279 89
rect 1174 47 1279 55
rect 1309 101 1363 177
rect 1309 67 1319 101
rect 1353 67 1363 101
rect 1309 47 1363 67
rect 1393 161 1445 177
rect 1393 127 1403 161
rect 1437 127 1445 161
rect 1393 93 1445 127
rect 1393 59 1403 93
rect 1437 59 1445 93
rect 1393 47 1445 59
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 369 79 383
rect 109 369 151 497
rect 181 475 257 497
rect 181 441 202 475
rect 236 441 257 475
rect 181 413 257 441
rect 287 480 353 497
rect 287 446 303 480
rect 337 446 353 480
rect 287 413 353 446
rect 383 413 471 497
rect 501 489 607 497
rect 501 455 542 489
rect 576 455 607 489
rect 501 413 607 455
rect 181 369 242 413
rect 557 297 607 413
rect 637 458 689 497
rect 637 424 647 458
rect 681 424 689 458
rect 847 485 897 497
rect 847 451 855 485
rect 889 451 897 485
rect 847 431 897 451
rect 1048 485 1100 497
rect 1048 451 1056 485
rect 1090 451 1100 485
rect 637 297 689 424
rect 750 349 802 431
rect 750 315 758 349
rect 792 315 802 349
rect 750 303 802 315
rect 832 303 912 431
rect 942 349 994 431
rect 1048 369 1100 451
rect 1130 442 1184 497
rect 1130 408 1140 442
rect 1174 408 1184 442
rect 1130 369 1184 408
rect 1214 489 1279 497
rect 1214 455 1230 489
rect 1264 455 1279 489
rect 1214 369 1279 455
rect 942 315 952 349
rect 986 315 994 349
rect 942 303 994 315
rect 1229 297 1279 369
rect 1309 448 1363 497
rect 1309 414 1319 448
rect 1353 414 1363 448
rect 1309 380 1363 414
rect 1309 346 1319 380
rect 1353 346 1363 380
rect 1309 297 1363 346
rect 1393 485 1445 497
rect 1393 451 1403 485
rect 1437 451 1445 485
rect 1393 417 1445 451
rect 1393 383 1403 417
rect 1437 383 1445 417
rect 1393 349 1445 383
rect 1393 315 1403 349
rect 1437 315 1445 349
rect 1393 297 1445 315
<< ndiffc >>
rect 35 69 69 103
rect 119 55 153 89
rect 203 67 237 101
rect 310 55 344 89
rect 546 85 580 119
rect 647 67 681 101
rect 751 76 785 110
rect 835 55 869 89
rect 919 76 953 110
rect 1028 75 1062 109
rect 1212 55 1246 89
rect 1319 67 1353 101
rect 1403 127 1437 161
rect 1403 59 1437 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 202 441 236 475
rect 303 446 337 480
rect 542 455 576 489
rect 647 424 681 458
rect 855 451 889 485
rect 1056 451 1090 485
rect 758 315 792 349
rect 1140 408 1174 442
rect 1230 455 1264 489
rect 952 315 986 349
rect 1319 414 1353 448
rect 1319 346 1353 380
rect 1403 451 1437 485
rect 1403 383 1437 417
rect 1403 315 1437 349
<< poly >>
rect 79 497 109 523
rect 151 497 181 523
rect 257 497 287 523
rect 353 497 383 523
rect 471 497 501 523
rect 607 497 637 523
rect 79 265 109 369
rect 21 249 109 265
rect 21 215 31 249
rect 65 215 109 249
rect 21 199 109 215
rect 151 265 181 369
rect 257 273 287 413
rect 353 381 383 413
rect 471 381 501 413
rect 329 365 383 381
rect 329 331 339 365
rect 373 331 383 365
rect 329 315 383 331
rect 465 365 519 381
rect 465 331 475 365
rect 509 331 519 365
rect 465 315 519 331
rect 151 249 215 265
rect 151 215 171 249
rect 205 215 215 249
rect 257 243 395 273
rect 151 199 215 215
rect 365 207 395 243
rect 79 131 109 199
rect 163 131 193 199
rect 257 191 323 201
rect 257 157 273 191
rect 307 157 323 191
rect 257 147 323 157
rect 365 191 419 207
rect 365 157 375 191
rect 409 157 419 191
rect 260 119 290 147
rect 365 141 419 157
rect 365 119 395 141
rect 487 131 517 315
rect 802 431 832 523
rect 912 431 942 523
rect 1100 497 1130 523
rect 1184 497 1214 523
rect 1279 497 1309 523
rect 1363 497 1393 523
rect 1100 331 1130 369
rect 1064 321 1130 331
rect 607 265 637 297
rect 802 265 832 303
rect 912 265 942 303
rect 1064 287 1080 321
rect 1114 287 1130 321
rect 1064 277 1130 287
rect 559 249 637 265
rect 559 215 569 249
rect 603 215 637 249
rect 559 199 637 215
rect 783 255 849 265
rect 783 221 799 255
rect 833 221 849 255
rect 783 211 849 221
rect 901 249 985 265
rect 901 215 941 249
rect 975 215 985 249
rect 607 177 637 199
rect 795 131 825 211
rect 901 176 985 215
rect 879 146 985 176
rect 879 131 909 146
rect 1072 131 1102 277
rect 1184 237 1214 369
rect 1279 265 1309 297
rect 1363 265 1393 297
rect 1144 227 1214 237
rect 1144 193 1160 227
rect 1194 193 1214 227
rect 1256 249 1393 265
rect 1256 215 1266 249
rect 1300 215 1393 249
rect 1256 199 1393 215
rect 1144 183 1214 193
rect 1144 131 1174 183
rect 1279 177 1309 199
rect 1363 177 1393 199
rect 79 21 109 47
rect 163 21 193 47
rect 260 21 290 47
rect 365 21 395 47
rect 487 21 517 47
rect 607 21 637 47
rect 795 21 825 47
rect 879 21 909 47
rect 1072 21 1102 47
rect 1144 21 1174 47
rect 1279 21 1309 47
rect 1363 21 1393 47
<< polycont >>
rect 31 215 65 249
rect 339 331 373 365
rect 475 331 509 365
rect 171 215 205 249
rect 273 157 307 191
rect 375 157 409 191
rect 1080 287 1114 321
rect 569 215 603 249
rect 799 221 833 255
rect 941 215 975 249
rect 1160 193 1194 227
rect 1266 215 1300 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 17 485 69 527
rect 17 451 35 485
rect 17 417 69 451
rect 17 383 35 417
rect 17 367 69 383
rect 103 475 252 493
rect 103 441 202 475
rect 236 441 252 475
rect 103 425 252 441
rect 286 480 441 493
rect 286 446 303 480
rect 337 446 441 480
rect 286 425 441 446
rect 17 249 68 333
rect 17 215 31 249
rect 65 215 68 249
rect 17 191 68 215
rect 103 157 137 425
rect 171 289 248 391
rect 282 365 373 391
rect 282 331 339 365
rect 282 323 373 331
rect 282 289 306 323
rect 340 289 373 323
rect 171 249 239 289
rect 282 265 373 289
rect 205 215 239 249
rect 171 191 239 215
rect 273 241 373 265
rect 407 275 441 425
rect 475 489 603 527
rect 475 455 542 489
rect 576 455 603 489
rect 475 415 603 455
rect 637 458 681 493
rect 637 424 647 458
rect 715 485 1106 527
rect 715 451 855 485
rect 889 451 1056 485
rect 1090 451 1106 485
rect 637 417 681 424
rect 1140 442 1174 493
rect 1214 489 1280 527
rect 1214 455 1230 489
rect 1264 455 1280 489
rect 1214 451 1280 455
rect 637 383 1098 417
rect 637 381 681 383
rect 475 365 681 381
rect 509 331 681 365
rect 475 327 681 331
rect 475 315 509 327
rect 407 249 603 275
rect 407 241 569 249
rect 273 191 341 241
rect 466 215 569 241
rect 307 157 341 191
rect 17 123 239 157
rect 273 141 341 157
rect 375 191 432 207
rect 409 187 432 191
rect 375 153 398 157
rect 375 141 432 153
rect 466 199 603 215
rect 17 103 69 123
rect 17 69 35 103
rect 203 101 239 123
rect 466 107 500 199
rect 17 51 69 69
rect 103 55 119 89
rect 153 55 169 89
rect 103 17 169 55
rect 237 67 239 101
rect 203 51 239 67
rect 273 89 500 107
rect 273 55 310 89
rect 344 55 500 89
rect 273 51 500 55
rect 534 119 603 165
rect 534 85 546 119
rect 580 85 603 119
rect 534 17 603 85
rect 637 101 681 327
rect 637 67 647 101
rect 637 51 681 67
rect 715 315 758 349
rect 792 315 808 349
rect 842 323 952 349
rect 715 187 749 315
rect 842 289 858 323
rect 892 315 952 323
rect 986 315 1002 349
rect 892 299 1002 315
rect 1036 321 1098 383
rect 1314 448 1368 493
rect 1174 408 1280 417
rect 1140 355 1280 408
rect 842 255 892 289
rect 1036 287 1080 321
rect 1114 287 1130 321
rect 1164 287 1280 355
rect 1314 414 1319 448
rect 1353 414 1368 448
rect 1314 380 1368 414
rect 1314 346 1319 380
rect 1353 346 1368 380
rect 1314 299 1368 346
rect 1246 265 1280 287
rect 783 221 799 255
rect 833 221 892 255
rect 715 153 766 187
rect 834 157 892 221
rect 941 253 985 265
rect 941 249 1210 253
rect 975 227 1210 249
rect 975 215 1160 227
rect 941 193 1160 215
rect 1194 193 1210 227
rect 941 191 1210 193
rect 1246 249 1300 265
rect 1246 215 1266 249
rect 1246 199 1300 215
rect 1334 263 1368 299
rect 1402 485 1455 527
rect 1402 451 1403 485
rect 1437 451 1455 485
rect 1402 417 1455 451
rect 1402 383 1403 417
rect 1437 383 1455 417
rect 1402 349 1455 383
rect 1402 315 1403 349
rect 1437 315 1455 349
rect 1402 297 1455 315
rect 1334 211 1455 263
rect 1246 157 1280 199
rect 1334 165 1368 211
rect 715 110 785 153
rect 834 123 965 157
rect 715 76 751 110
rect 919 110 965 123
rect 715 51 785 76
rect 819 55 835 89
rect 869 55 885 89
rect 819 17 885 55
rect 953 76 965 110
rect 919 51 965 76
rect 1020 123 1280 157
rect 1020 109 1062 123
rect 1020 75 1028 109
rect 1314 101 1368 165
rect 1020 51 1062 75
rect 1098 55 1212 89
rect 1246 55 1280 89
rect 1098 17 1280 55
rect 1314 67 1319 101
rect 1353 67 1368 101
rect 1314 51 1368 67
rect 1402 161 1455 177
rect 1402 127 1403 161
rect 1437 127 1455 161
rect 1402 93 1455 127
rect 1402 59 1403 93
rect 1437 59 1455 93
rect 1402 17 1455 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 306 289 340 323
rect 398 157 409 187
rect 409 157 432 187
rect 398 153 432 157
rect 858 289 892 323
rect 766 153 800 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 294 323 352 329
rect 294 289 306 323
rect 340 320 352 323
rect 846 323 904 329
rect 846 320 858 323
rect 340 292 858 320
rect 340 289 352 292
rect 294 283 352 289
rect 846 289 858 292
rect 892 289 904 323
rect 846 283 904 289
rect 386 187 444 193
rect 386 153 398 187
rect 432 184 444 187
rect 754 187 812 193
rect 754 184 766 187
rect 432 156 766 184
rect 432 153 444 156
rect 386 147 444 153
rect 754 153 766 156
rect 800 153 812 187
rect 754 147 812 153
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< labels >>
flabel corelocali s 29 289 63 323 0 FreeSans 200 0 0 0 SCE
port 3 nsew
flabel corelocali s 950 221 984 255 0 FreeSans 200 0 0 0 CLK
port 1 nsew
flabel corelocali s 1329 425 1363 459 0 FreeSans 200 0 0 0 GCLK
port 8 nsew
flabel corelocali s 1329 357 1363 391 0 FreeSans 200 0 0 0 GCLK
port 8 nsew
flabel corelocali s 214 357 248 391 0 FreeSans 200 0 0 0 GATE
port 2 nsew
flabel corelocali s 1329 85 1363 119 0 FreeSans 200 0 0 0 GCLK
port 8 nsew
flabel corelocali s 214 289 248 323 0 FreeSans 200 0 0 0 GATE
port 2 nsew
flabel corelocali s 29 221 63 255 0 FreeSans 200 0 0 0 SCE
port 3 nsew
flabel corelocali s 1421 221 1455 255 0 FreeSans 200 0 0 0 GCLK
port 8 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
rlabel comment s 0 0 0 0 4 sdlclkp_2
<< properties >>
string FIXED_BBOX 0 0 1472 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 431368
string GDS_START 419768
string path 0.000 0.000 7.360 0.000 
<< end >>
