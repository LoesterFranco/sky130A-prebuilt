magic
tech sky130A
magscale 1 2
timestamp 1601050088
<< locali >>
rect 25 236 108 310
rect 195 270 263 578
rect 309 270 375 430
rect 453 390 557 596
rect 409 270 489 356
rect 523 236 557 390
rect 156 202 557 236
rect 156 70 208 202
rect 362 70 428 202
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 51 364 117 649
rect 42 17 122 202
rect 242 17 308 168
rect 462 17 528 168
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
rlabel locali s 25 236 108 310 6 A
port 1 nsew signal input
rlabel locali s 195 270 263 578 6 B
port 2 nsew signal input
rlabel locali s 309 270 375 430 6 C
port 3 nsew signal input
rlabel locali s 409 270 489 356 6 D
port 4 nsew signal input
rlabel locali s 523 236 557 390 6 Y
port 5 nsew signal output
rlabel locali s 453 390 557 596 6 Y
port 5 nsew signal output
rlabel locali s 362 70 428 202 6 Y
port 5 nsew signal output
rlabel locali s 156 202 557 236 6 Y
port 5 nsew signal output
rlabel locali s 156 70 208 202 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -49 576 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 576 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 576 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1639498
string GDS_START 1634016
<< end >>
