magic
tech sky130A
magscale 1 2
timestamp 1604502710
<< nwell >>
rect -38 332 1670 704
<< pwell >>
rect 0 0 1632 49
<< scpmos >>
rect 82 413 118 581
rect 204 413 240 581
rect 430 392 466 560
rect 553 392 589 592
rect 631 392 667 592
rect 737 508 773 592
rect 868 508 904 592
rect 1011 368 1047 592
rect 1213 368 1249 592
rect 1314 424 1350 592
rect 1514 368 1550 592
<< nmoslvt >>
rect 85 112 115 222
rect 201 74 231 222
rect 430 82 460 230
rect 559 80 589 208
rect 637 80 667 208
rect 785 124 815 208
rect 863 124 893 208
rect 979 74 1009 222
rect 1220 78 1250 226
rect 1320 116 1350 226
rect 1518 74 1548 222
<< ndiff >>
rect 28 176 85 222
rect 28 142 40 176
rect 74 142 85 176
rect 28 112 85 142
rect 115 202 201 222
rect 115 168 142 202
rect 176 168 201 202
rect 115 121 201 168
rect 115 112 142 121
rect 130 87 142 112
rect 176 87 201 121
rect 130 74 201 87
rect 231 202 288 222
rect 231 168 242 202
rect 276 168 288 202
rect 231 121 288 168
rect 231 87 242 121
rect 276 87 288 121
rect 231 74 288 87
rect 373 218 430 230
rect 373 184 385 218
rect 419 184 430 218
rect 373 82 430 184
rect 460 208 510 230
rect 908 208 979 222
rect 460 82 559 208
rect 475 48 492 82
rect 526 80 559 82
rect 589 80 637 208
rect 667 170 785 208
rect 667 136 709 170
rect 743 136 785 170
rect 667 124 785 136
rect 815 124 863 208
rect 893 196 979 208
rect 893 162 920 196
rect 954 162 979 196
rect 893 124 979 162
rect 667 80 717 124
rect 908 120 979 124
rect 526 48 544 80
rect 475 36 544 48
rect 908 86 920 120
rect 954 86 979 120
rect 908 74 979 86
rect 1009 198 1066 222
rect 1009 164 1020 198
rect 1054 164 1066 198
rect 1009 120 1066 164
rect 1009 86 1020 120
rect 1054 86 1066 120
rect 1009 74 1066 86
rect 1164 214 1220 226
rect 1164 180 1175 214
rect 1209 180 1220 214
rect 1164 124 1220 180
rect 1164 90 1175 124
rect 1209 90 1220 124
rect 1164 78 1220 90
rect 1250 188 1320 226
rect 1250 154 1268 188
rect 1302 154 1320 188
rect 1250 116 1320 154
rect 1350 188 1407 226
rect 1350 154 1361 188
rect 1395 154 1407 188
rect 1350 116 1407 154
rect 1461 210 1518 222
rect 1461 176 1473 210
rect 1507 176 1518 210
rect 1461 120 1518 176
rect 1250 78 1300 116
rect 1461 86 1473 120
rect 1507 86 1518 120
rect 1461 74 1518 86
rect 1548 210 1605 222
rect 1548 176 1559 210
rect 1593 176 1605 210
rect 1548 120 1605 176
rect 1548 86 1559 120
rect 1593 86 1605 120
rect 1548 74 1605 86
<< pdiff >>
rect 133 627 189 639
rect 133 593 144 627
rect 178 593 189 627
rect 133 581 189 593
rect 481 606 538 618
rect 27 569 82 581
rect 27 535 38 569
rect 72 535 82 569
rect 27 462 82 535
rect 27 428 38 462
rect 72 428 82 462
rect 27 413 82 428
rect 118 413 204 581
rect 240 459 296 581
rect 481 572 492 606
rect 526 592 538 606
rect 526 572 553 592
rect 481 560 553 572
rect 240 425 250 459
rect 284 425 296 459
rect 240 413 296 425
rect 374 539 430 560
rect 374 505 386 539
rect 420 505 430 539
rect 374 392 430 505
rect 466 392 553 560
rect 589 392 631 592
rect 667 508 737 592
rect 773 508 868 592
rect 904 559 1011 592
rect 904 525 935 559
rect 969 525 1011 559
rect 904 508 1011 525
rect 667 438 722 508
rect 667 404 677 438
rect 711 404 722 438
rect 667 392 722 404
rect 961 368 1011 508
rect 1047 580 1103 592
rect 1047 546 1057 580
rect 1091 546 1103 580
rect 1047 497 1103 546
rect 1047 463 1057 497
rect 1091 463 1103 497
rect 1047 414 1103 463
rect 1047 380 1057 414
rect 1091 380 1103 414
rect 1047 368 1103 380
rect 1157 580 1213 592
rect 1157 546 1169 580
rect 1203 546 1213 580
rect 1157 497 1213 546
rect 1157 463 1169 497
rect 1203 463 1213 497
rect 1157 414 1213 463
rect 1157 380 1169 414
rect 1203 380 1213 414
rect 1157 368 1213 380
rect 1249 580 1314 592
rect 1249 546 1259 580
rect 1293 546 1314 580
rect 1249 470 1314 546
rect 1249 436 1259 470
rect 1293 436 1314 470
rect 1249 424 1314 436
rect 1350 580 1405 592
rect 1350 546 1360 580
rect 1394 546 1405 580
rect 1350 470 1405 546
rect 1350 436 1360 470
rect 1394 436 1405 470
rect 1350 424 1405 436
rect 1459 580 1514 592
rect 1459 546 1470 580
rect 1504 546 1514 580
rect 1459 497 1514 546
rect 1459 463 1470 497
rect 1504 463 1514 497
rect 1249 368 1299 424
rect 1459 414 1514 463
rect 1459 380 1470 414
rect 1504 380 1514 414
rect 1459 368 1514 380
rect 1550 580 1605 592
rect 1550 546 1560 580
rect 1594 546 1605 580
rect 1550 497 1605 546
rect 1550 463 1560 497
rect 1594 463 1605 497
rect 1550 414 1605 463
rect 1550 380 1560 414
rect 1594 380 1605 414
rect 1550 368 1605 380
<< ndiffc >>
rect 40 142 74 176
rect 142 168 176 202
rect 142 87 176 121
rect 242 168 276 202
rect 242 87 276 121
rect 385 184 419 218
rect 492 48 526 82
rect 709 136 743 170
rect 920 162 954 196
rect 920 86 954 120
rect 1020 164 1054 198
rect 1020 86 1054 120
rect 1175 180 1209 214
rect 1175 90 1209 124
rect 1268 154 1302 188
rect 1361 154 1395 188
rect 1473 176 1507 210
rect 1473 86 1507 120
rect 1559 176 1593 210
rect 1559 86 1593 120
<< pdiffc >>
rect 144 593 178 627
rect 38 535 72 569
rect 38 428 72 462
rect 492 572 526 606
rect 250 425 284 459
rect 386 505 420 539
rect 935 525 969 559
rect 677 404 711 438
rect 1057 546 1091 580
rect 1057 463 1091 497
rect 1057 380 1091 414
rect 1169 546 1203 580
rect 1169 463 1203 497
rect 1169 380 1203 414
rect 1259 546 1293 580
rect 1259 436 1293 470
rect 1360 546 1394 580
rect 1360 436 1394 470
rect 1470 546 1504 580
rect 1470 463 1504 497
rect 1470 380 1504 414
rect 1560 546 1594 580
rect 1560 463 1594 497
rect 1560 380 1594 414
<< poly >>
rect 82 581 118 607
rect 204 581 240 607
rect 430 560 466 586
rect 553 592 589 618
rect 631 592 667 618
rect 737 592 773 618
rect 868 592 904 618
rect 1011 592 1047 618
rect 1213 592 1249 618
rect 1314 592 1350 618
rect 1514 592 1550 618
rect 82 378 118 413
rect 82 362 153 378
rect 82 328 103 362
rect 137 328 153 362
rect 82 294 153 328
rect 204 310 240 413
rect 737 476 773 508
rect 737 460 820 476
rect 868 464 904 508
rect 737 426 770 460
rect 804 426 820 460
rect 737 410 820 426
rect 863 448 929 464
rect 863 414 879 448
rect 913 414 929 448
rect 430 360 466 392
rect 553 360 589 392
rect 332 344 466 360
rect 332 310 348 344
rect 382 310 416 344
rect 450 310 466 344
rect 82 260 103 294
rect 137 260 153 294
rect 82 244 153 260
rect 201 294 267 310
rect 332 294 466 310
rect 509 344 589 360
rect 509 310 525 344
rect 559 310 589 344
rect 631 368 667 392
rect 631 338 815 368
rect 509 294 589 310
rect 201 260 217 294
rect 251 260 267 294
rect 201 244 267 260
rect 85 222 115 244
rect 201 222 231 244
rect 430 230 460 294
rect 85 86 115 112
rect 559 208 589 294
rect 637 280 703 296
rect 637 246 653 280
rect 687 246 703 280
rect 637 230 703 246
rect 637 208 667 230
rect 785 208 815 338
rect 863 362 929 414
rect 863 208 893 362
rect 1011 314 1047 368
rect 1213 330 1249 368
rect 1314 330 1350 424
rect 1514 330 1550 368
rect 941 298 1047 314
rect 941 264 957 298
rect 991 284 1047 298
rect 1089 314 1350 330
rect 991 264 1009 284
rect 1089 280 1105 314
rect 1139 280 1350 314
rect 1089 264 1350 280
rect 1398 314 1550 330
rect 1398 280 1414 314
rect 1448 280 1550 314
rect 1398 264 1550 280
rect 941 248 1009 264
rect 979 222 1009 248
rect 1220 226 1250 264
rect 1320 226 1350 264
rect 201 48 231 74
rect 430 56 460 82
rect 785 102 815 124
rect 749 86 815 102
rect 863 98 893 124
rect 559 54 589 80
rect 637 54 667 80
rect 749 52 765 86
rect 799 52 815 86
rect 1518 222 1548 264
rect 1320 90 1350 116
rect 749 36 815 52
rect 979 48 1009 74
rect 1220 52 1250 78
rect 1518 48 1548 74
<< polycont >>
rect 103 328 137 362
rect 770 426 804 460
rect 879 414 913 448
rect 348 310 382 344
rect 416 310 450 344
rect 103 260 137 294
rect 525 310 559 344
rect 217 260 251 294
rect 653 246 687 280
rect 957 264 991 298
rect 1105 280 1139 314
rect 1414 280 1448 314
rect 765 52 799 86
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 128 627 194 649
rect 128 593 144 627
rect 178 593 194 627
rect 19 569 88 585
rect 128 577 194 593
rect 476 606 542 649
rect 19 535 38 569
rect 72 543 88 569
rect 476 572 492 606
rect 526 572 542 606
rect 72 535 352 543
rect 19 509 352 535
rect 19 462 88 509
rect 19 428 38 462
rect 72 428 88 462
rect 19 412 88 428
rect 234 459 284 475
rect 234 425 250 459
rect 19 210 53 412
rect 234 378 284 425
rect 318 446 352 509
rect 386 539 436 564
rect 476 556 542 572
rect 898 559 1007 649
rect 420 522 436 539
rect 898 525 935 559
rect 969 525 1007 559
rect 420 505 820 522
rect 898 509 1007 525
rect 1041 580 1107 596
rect 1041 546 1057 580
rect 1091 546 1107 580
rect 386 488 820 505
rect 386 480 436 488
rect 318 412 575 446
rect 87 362 167 378
rect 87 328 103 362
rect 137 328 167 362
rect 234 344 466 378
rect 87 294 167 328
rect 301 310 348 344
rect 382 310 416 344
rect 450 310 466 344
rect 87 260 103 294
rect 137 260 167 294
rect 87 244 167 260
rect 201 294 267 310
rect 201 260 217 294
rect 251 260 267 294
rect 201 236 267 260
rect 301 294 466 310
rect 509 344 575 412
rect 509 310 525 344
rect 559 310 575 344
rect 509 294 575 310
rect 609 296 643 488
rect 754 460 820 488
rect 1041 497 1107 546
rect 1041 464 1057 497
rect 677 438 711 454
rect 754 426 770 460
rect 804 426 820 460
rect 754 410 820 426
rect 863 463 1057 464
rect 1091 463 1107 497
rect 863 448 1107 463
rect 863 414 879 448
rect 913 414 1107 448
rect 677 364 711 404
rect 863 398 1057 414
rect 1041 380 1057 398
rect 1091 380 1107 414
rect 677 330 1007 364
rect 19 176 90 210
rect 301 202 335 294
rect 609 280 703 296
rect 609 246 653 280
rect 687 246 703 280
rect 609 238 703 246
rect 19 142 40 176
rect 74 142 90 176
rect 19 108 90 142
rect 126 168 142 202
rect 176 168 192 202
rect 126 121 192 168
rect 126 87 142 121
rect 176 87 192 121
rect 126 17 192 87
rect 226 168 242 202
rect 276 168 335 202
rect 369 218 703 238
rect 369 184 385 218
rect 419 204 703 218
rect 419 184 435 204
rect 756 170 790 330
rect 941 298 1007 330
rect 941 264 957 298
rect 991 264 1007 298
rect 941 248 1007 264
rect 1041 330 1107 380
rect 1153 580 1225 596
rect 1153 546 1169 580
rect 1203 546 1225 580
rect 1153 497 1225 546
rect 1153 463 1169 497
rect 1203 463 1225 497
rect 1153 414 1225 463
rect 1259 580 1309 649
rect 1293 546 1309 580
rect 1259 470 1309 546
rect 1293 436 1309 470
rect 1259 420 1309 436
rect 1344 580 1410 596
rect 1344 546 1360 580
rect 1394 546 1410 580
rect 1344 470 1410 546
rect 1344 436 1360 470
rect 1394 436 1410 470
rect 1153 380 1169 414
rect 1203 380 1225 414
rect 1153 364 1225 380
rect 1041 314 1155 330
rect 1041 280 1105 314
rect 1139 280 1155 314
rect 1041 264 1155 280
rect 1041 214 1075 264
rect 1191 230 1225 364
rect 1344 330 1410 436
rect 1454 580 1504 649
rect 1454 546 1470 580
rect 1454 497 1504 546
rect 1454 463 1470 497
rect 1454 414 1504 463
rect 1454 380 1470 414
rect 1454 364 1504 380
rect 1543 580 1610 596
rect 1543 546 1560 580
rect 1594 546 1610 580
rect 1543 497 1610 546
rect 1543 463 1560 497
rect 1594 463 1610 497
rect 1543 414 1610 463
rect 1543 380 1560 414
rect 1594 380 1610 414
rect 1344 314 1464 330
rect 1344 280 1414 314
rect 1448 280 1464 314
rect 1344 264 1464 280
rect 226 150 335 168
rect 226 121 616 150
rect 662 136 709 170
rect 743 136 790 170
rect 904 196 970 212
rect 904 162 920 196
rect 954 162 970 196
rect 226 87 242 121
rect 276 116 616 121
rect 276 87 335 116
rect 226 70 335 87
rect 582 102 616 116
rect 904 120 970 162
rect 582 86 815 102
rect 471 48 492 82
rect 526 48 548 82
rect 582 52 765 86
rect 799 52 815 86
rect 582 51 815 52
rect 904 86 920 120
rect 954 86 970 120
rect 471 17 548 48
rect 904 17 970 86
rect 1004 198 1075 214
rect 1004 164 1020 198
rect 1054 164 1075 198
rect 1004 120 1075 164
rect 1004 86 1020 120
rect 1054 86 1075 120
rect 1004 70 1075 86
rect 1159 214 1225 230
rect 1159 180 1175 214
rect 1209 180 1225 214
rect 1159 124 1225 180
rect 1159 90 1175 124
rect 1209 90 1225 124
rect 1159 74 1225 90
rect 1259 188 1309 230
rect 1259 154 1268 188
rect 1302 154 1309 188
rect 1259 17 1309 154
rect 1344 188 1411 264
rect 1344 154 1361 188
rect 1395 154 1411 188
rect 1344 112 1411 154
rect 1457 210 1507 226
rect 1457 176 1473 210
rect 1457 120 1507 176
rect 1457 86 1473 120
rect 1457 17 1507 86
rect 1543 210 1610 380
rect 1543 176 1559 210
rect 1593 176 1610 210
rect 1543 120 1610 176
rect 1543 86 1559 120
rect 1593 86 1610 120
rect 1543 70 1610 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
rlabel comment s 0 0 0 0 4 dlxbp_1
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 1567 94 1601 128 0 FreeSans 340 0 0 0 Q_N
port 8 nsew
flabel corelocali s 1567 168 1601 202 0 FreeSans 340 0 0 0 Q_N
port 8 nsew
flabel corelocali s 1567 242 1601 276 0 FreeSans 340 0 0 0 Q_N
port 8 nsew
flabel corelocali s 1567 316 1601 350 0 FreeSans 340 0 0 0 Q_N
port 8 nsew
flabel corelocali s 1567 390 1601 424 0 FreeSans 340 0 0 0 Q_N
port 8 nsew
flabel corelocali s 1567 464 1601 498 0 FreeSans 340 0 0 0 Q_N
port 8 nsew
flabel corelocali s 1567 538 1601 572 0 FreeSans 340 0 0 0 Q_N
port 8 nsew
flabel corelocali s 1183 94 1217 128 0 FreeSans 340 0 0 0 Q
port 7 nsew
flabel corelocali s 1183 168 1217 202 0 FreeSans 340 0 0 0 Q
port 7 nsew
flabel corelocali s 223 242 257 276 0 FreeSans 340 0 0 0 GATE
port 2 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 1632 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 2169540
string GDS_START 2156844
<< end >>
