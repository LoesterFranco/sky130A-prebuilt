magic
tech sky130A
magscale 1 2
timestamp 1599588244
<< locali >>
rect 25 290 103 356
rect 205 290 258 356
rect 1435 394 1485 596
rect 1619 394 1685 596
rect 1435 360 1799 394
rect 1177 224 1319 290
rect 1753 226 1799 360
rect 1477 176 1799 226
rect 1477 73 1529 176
rect 1663 73 1701 176
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 23 508 89 566
rect 130 542 196 649
rect 467 542 533 649
rect 569 581 797 615
rect 23 474 533 508
rect 23 390 171 474
rect 237 390 326 440
rect 360 404 448 440
rect 137 256 171 390
rect 292 356 326 390
rect 292 290 380 356
rect 23 222 171 256
rect 292 240 326 290
rect 414 256 448 404
rect 499 360 533 474
rect 569 428 603 581
rect 637 481 693 547
rect 569 394 625 428
rect 499 294 557 360
rect 591 290 625 394
rect 659 379 693 481
rect 731 413 797 581
rect 869 530 981 649
rect 1022 496 1088 540
rect 839 413 1088 496
rect 659 345 1004 379
rect 591 256 668 290
rect 23 122 89 222
rect 248 188 326 240
rect 360 222 668 256
rect 136 17 202 188
rect 248 154 601 188
rect 702 185 736 345
rect 248 84 326 154
rect 467 17 533 120
rect 567 85 601 154
rect 635 119 736 185
rect 770 245 830 311
rect 944 270 1004 345
rect 1038 358 1088 413
rect 1122 392 1188 649
rect 1222 358 1288 540
rect 1329 392 1395 649
rect 1519 428 1585 649
rect 1719 428 1785 649
rect 1038 326 1387 358
rect 1038 324 1719 326
rect 770 85 804 245
rect 567 51 804 85
rect 838 17 888 162
rect 934 90 1000 206
rect 1038 190 1072 324
rect 1353 260 1719 324
rect 1036 124 1072 190
rect 1107 154 1345 190
rect 1107 90 1157 154
rect 934 56 1157 90
rect 1193 17 1259 120
rect 1293 69 1345 154
rect 1391 17 1443 226
rect 1563 17 1629 142
rect 1735 17 1801 142
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
<< metal1 >>
rect 0 683 1824 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 0 617 1824 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 1824 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
rect 0 -49 1824 -17
<< labels >>
rlabel locali s 25 290 103 356 6 D
port 1 nsew signal input
rlabel locali s 1753 226 1799 360 6 Q
port 2 nsew signal output
rlabel locali s 1663 73 1701 176 6 Q
port 2 nsew signal output
rlabel locali s 1619 394 1685 596 6 Q
port 2 nsew signal output
rlabel locali s 1477 176 1799 226 6 Q
port 2 nsew signal output
rlabel locali s 1477 73 1529 176 6 Q
port 2 nsew signal output
rlabel locali s 1435 394 1485 596 6 Q
port 2 nsew signal output
rlabel locali s 1435 360 1799 394 6 Q
port 2 nsew signal output
rlabel locali s 1177 224 1319 290 6 RESET_B
port 3 nsew signal input
rlabel locali s 205 290 258 356 6 GATE
port 4 nsew clock input
rlabel metal1 s 0 -49 1824 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 6 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 617 1824 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1824 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 2130608
string GDS_START 2117296
<< end >>
