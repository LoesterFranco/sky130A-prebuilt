magic
tech sky130A
magscale 1 2
timestamp 1599588232
<< locali >>
rect 22 108 89 596
rect 197 581 529 615
rect 197 424 231 581
rect 463 575 529 581
rect 133 390 231 424
rect 133 180 167 390
rect 201 282 267 356
rect 133 146 335 180
rect 301 80 415 146
rect 1829 236 1895 310
rect 2564 294 2698 360
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 129 458 163 649
rect 587 593 658 649
rect 692 581 1400 615
rect 692 559 726 581
rect 265 541 335 547
rect 563 541 726 559
rect 265 525 726 541
rect 265 507 597 525
rect 265 390 335 507
rect 841 491 907 547
rect 631 473 907 491
rect 301 248 335 390
rect 226 214 335 248
rect 369 457 907 473
rect 369 439 665 457
rect 369 214 435 439
rect 699 405 800 423
rect 841 420 907 457
rect 941 546 1225 581
rect 601 371 800 405
rect 601 350 689 371
rect 941 353 975 546
rect 1266 498 1332 528
rect 500 282 566 327
rect 601 316 607 350
rect 641 316 689 350
rect 834 337 975 353
rect 500 248 621 282
rect 369 180 553 214
rect 124 17 190 112
rect 451 17 485 146
rect 519 85 553 180
rect 587 153 621 248
rect 655 237 689 316
rect 734 319 975 337
rect 1009 464 1332 498
rect 734 287 868 319
rect 1009 285 1043 464
rect 1266 458 1332 464
rect 976 253 1043 285
rect 1081 424 1127 430
rect 1366 424 1400 581
rect 1081 390 1087 424
rect 1121 390 1127 424
rect 1081 341 1127 390
rect 1211 390 1400 424
rect 1434 390 1500 585
rect 1081 275 1177 341
rect 655 187 721 237
rect 755 219 1043 253
rect 1211 241 1245 390
rect 755 153 789 219
rect 1077 207 1245 241
rect 1279 350 1319 356
rect 1313 316 1319 350
rect 1279 310 1319 316
rect 1369 350 1415 356
rect 1369 316 1375 350
rect 1409 316 1415 350
rect 1369 310 1415 316
rect 1077 187 1143 207
rect 587 119 789 153
rect 823 153 1009 185
rect 1177 153 1243 173
rect 823 151 1243 153
rect 823 85 857 151
rect 975 119 1243 151
rect 1279 134 1313 310
rect 1369 276 1413 310
rect 1347 142 1413 276
rect 1466 226 1500 390
rect 1534 353 1600 649
rect 1634 581 2348 615
rect 1634 376 1722 581
rect 1756 513 2163 547
rect 1756 424 1822 513
rect 1756 390 1768 424
rect 1802 390 1822 424
rect 1756 376 1822 390
rect 1856 424 2095 479
rect 1856 390 1977 424
rect 2011 390 2049 424
rect 2083 390 2095 424
rect 1634 242 1668 376
rect 1856 361 2095 390
rect 1702 276 1795 342
rect 1447 158 1513 226
rect 1634 192 1727 242
rect 1761 158 1795 276
rect 1929 192 1995 361
rect 2029 244 2095 310
rect 2029 158 2063 244
rect 2129 210 2163 513
rect 1447 124 2063 158
rect 519 51 857 85
rect 891 85 941 117
rect 1447 85 1513 124
rect 2097 119 2163 210
rect 2197 356 2231 547
rect 2197 350 2243 356
rect 2197 316 2203 350
rect 2237 316 2243 350
rect 2197 310 2243 316
rect 891 51 1513 85
rect 1549 17 1615 90
rect 1779 85 1877 90
rect 2197 85 2231 310
rect 2277 226 2348 581
rect 2390 466 2458 649
rect 2390 422 2444 466
rect 2504 432 2570 596
rect 2478 424 2570 432
rect 2478 390 2487 424
rect 2521 394 2570 424
rect 2610 394 2660 649
rect 2694 394 2766 596
rect 2521 390 2530 394
rect 2478 388 2530 390
rect 1779 51 2231 85
rect 2281 70 2348 226
rect 2382 344 2530 388
rect 2382 192 2416 344
rect 2450 260 2516 310
rect 2732 260 2766 394
rect 2450 226 2766 260
rect 2382 158 2561 192
rect 2383 17 2449 124
rect 2495 70 2561 158
rect 2595 17 2661 192
rect 2695 70 2766 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 607 316 641 350
rect 1087 390 1121 424
rect 1279 316 1313 350
rect 1375 316 1409 350
rect 1768 390 1802 424
rect 1977 390 2011 424
rect 2049 390 2083 424
rect 2203 316 2237 350
rect 2487 390 2521 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
<< metal1 >>
rect 0 683 2784 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 0 617 2784 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 2784 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
rect 0 -49 2784 -17
<< obsm1 >>
rect 1075 424 1133 430
rect 1075 390 1087 424
rect 1121 421 1133 424
rect 1756 424 1814 430
rect 1756 421 1768 424
rect 1121 393 1768 421
rect 1121 390 1133 393
rect 1075 384 1133 390
rect 1756 390 1768 393
rect 1802 390 1814 424
rect 1756 384 1814 390
rect 1965 424 2095 430
rect 1965 390 1977 424
rect 2011 390 2049 424
rect 2083 421 2095 424
rect 2475 424 2533 430
rect 2475 421 2487 424
rect 2083 393 2487 421
rect 2083 390 2095 393
rect 1965 384 2095 390
rect 2475 390 2487 393
rect 2521 390 2533 424
rect 2475 384 2533 390
rect 595 350 653 356
rect 595 316 607 350
rect 641 347 653 350
rect 1267 350 1325 356
rect 1267 347 1279 350
rect 641 319 1279 347
rect 641 316 653 319
rect 595 310 653 316
rect 1267 316 1279 319
rect 1313 316 1325 350
rect 1267 310 1325 316
rect 1363 350 1421 356
rect 1363 316 1375 350
rect 1409 347 1421 350
rect 2191 350 2249 356
rect 2191 347 2203 350
rect 1409 319 2203 347
rect 1409 316 1421 319
rect 1363 310 1421 316
rect 2191 316 2203 319
rect 2237 316 2249 350
rect 2191 310 2249 316
<< labels >>
rlabel locali s 2564 294 2698 360 6 A
port 1 nsew signal input
rlabel locali s 1829 236 1895 310 6 B
port 2 nsew signal input
rlabel locali s 201 282 267 356 6 CI
port 3 nsew signal input
rlabel locali s 463 575 529 581 6 COUT
port 4 nsew signal output
rlabel locali s 301 80 415 146 6 COUT
port 4 nsew signal output
rlabel locali s 197 581 529 615 6 COUT
port 4 nsew signal output
rlabel locali s 197 424 231 581 6 COUT
port 4 nsew signal output
rlabel locali s 133 390 231 424 6 COUT
port 4 nsew signal output
rlabel locali s 133 180 167 390 6 COUT
port 4 nsew signal output
rlabel locali s 133 146 335 180 6 COUT
port 4 nsew signal output
rlabel locali s 22 108 89 596 6 SUM
port 5 nsew signal output
rlabel metal1 s 0 -49 2784 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 7 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 617 2784 715 6 VPWR
port 9 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2784 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 2532620
string GDS_START 2512166
<< end >>
