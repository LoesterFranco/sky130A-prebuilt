magic
tech sky130A
magscale 1 2
timestamp 1599588218
<< nwell >>
rect -38 332 1190 704
<< pwell >>
rect 0 0 1152 49
<< scpmos >>
rect 81 368 117 592
rect 171 368 207 592
rect 261 368 297 592
rect 351 368 387 592
rect 456 392 492 592
rect 546 392 582 592
rect 745 387 781 587
rect 835 387 871 587
rect 1035 392 1071 592
<< nmoslvt >>
rect 84 74 114 222
rect 170 74 200 222
rect 270 74 300 222
rect 361 74 391 222
rect 456 74 486 202
rect 576 74 606 202
rect 676 74 706 202
rect 762 74 792 202
rect 862 74 892 202
<< ndiff >>
rect 27 186 84 222
rect 27 152 39 186
rect 73 152 84 186
rect 27 118 84 152
rect 27 84 39 118
rect 73 84 84 118
rect 27 74 84 84
rect 114 210 170 222
rect 114 176 125 210
rect 159 176 170 210
rect 114 120 170 176
rect 114 86 125 120
rect 159 86 170 120
rect 114 74 170 86
rect 200 137 270 222
rect 200 103 211 137
rect 245 103 270 137
rect 200 74 270 103
rect 300 210 361 222
rect 300 176 311 210
rect 345 176 361 210
rect 300 120 361 176
rect 300 86 311 120
rect 345 86 361 120
rect 300 74 361 86
rect 391 202 441 222
rect 391 188 456 202
rect 391 154 411 188
rect 445 154 456 188
rect 391 120 456 154
rect 391 86 411 120
rect 445 86 456 120
rect 391 74 456 86
rect 486 190 576 202
rect 486 156 511 190
rect 545 156 576 190
rect 486 120 576 156
rect 486 86 511 120
rect 545 86 576 120
rect 486 74 576 86
rect 606 188 676 202
rect 606 154 617 188
rect 651 154 676 188
rect 606 120 676 154
rect 606 86 617 120
rect 651 86 676 120
rect 606 74 676 86
rect 706 190 762 202
rect 706 156 717 190
rect 751 156 762 190
rect 706 120 762 156
rect 706 86 717 120
rect 751 86 762 120
rect 706 74 762 86
rect 792 190 862 202
rect 792 156 803 190
rect 837 156 862 190
rect 792 120 862 156
rect 792 86 803 120
rect 837 86 862 120
rect 792 74 862 86
rect 892 188 1088 202
rect 892 154 903 188
rect 937 154 972 188
rect 1006 154 1042 188
rect 1076 154 1088 188
rect 892 120 1088 154
rect 892 86 903 120
rect 937 86 972 120
rect 1006 86 1042 120
rect 1076 86 1088 120
rect 892 74 1088 86
<< pdiff >>
rect 27 580 81 592
rect 27 546 37 580
rect 71 546 81 580
rect 27 497 81 546
rect 27 463 37 497
rect 71 463 81 497
rect 27 414 81 463
rect 27 380 37 414
rect 71 380 81 414
rect 27 368 81 380
rect 117 580 171 592
rect 117 546 127 580
rect 161 546 171 580
rect 117 497 171 546
rect 117 463 127 497
rect 161 463 171 497
rect 117 414 171 463
rect 117 380 127 414
rect 161 380 171 414
rect 117 368 171 380
rect 207 580 261 592
rect 207 546 217 580
rect 251 546 261 580
rect 207 478 261 546
rect 207 444 217 478
rect 251 444 261 478
rect 207 368 261 444
rect 297 580 351 592
rect 297 546 307 580
rect 341 546 351 580
rect 297 497 351 546
rect 297 463 307 497
rect 341 463 351 497
rect 297 414 351 463
rect 297 380 307 414
rect 341 380 351 414
rect 297 368 351 380
rect 387 580 456 592
rect 387 546 397 580
rect 431 546 456 580
rect 387 509 456 546
rect 387 475 397 509
rect 431 475 456 509
rect 387 438 456 475
rect 387 404 397 438
rect 431 404 456 438
rect 387 392 456 404
rect 492 580 546 592
rect 492 546 502 580
rect 536 546 546 580
rect 492 510 546 546
rect 492 476 502 510
rect 536 476 546 510
rect 492 440 546 476
rect 492 406 502 440
rect 536 406 546 440
rect 492 392 546 406
rect 582 580 636 592
rect 582 546 592 580
rect 626 546 636 580
rect 582 508 636 546
rect 582 474 592 508
rect 626 474 636 508
rect 582 392 636 474
rect 690 575 745 587
rect 690 541 701 575
rect 735 541 745 575
rect 690 504 745 541
rect 690 470 701 504
rect 735 470 745 504
rect 690 433 745 470
rect 690 399 701 433
rect 735 399 745 433
rect 387 368 441 392
rect 690 387 745 399
rect 781 531 835 587
rect 781 497 791 531
rect 825 497 835 531
rect 781 433 835 497
rect 781 399 791 433
rect 825 399 835 433
rect 781 387 835 399
rect 871 575 926 587
rect 871 541 881 575
rect 915 541 926 575
rect 871 507 926 541
rect 871 473 881 507
rect 915 473 926 507
rect 871 439 926 473
rect 871 405 881 439
rect 915 405 926 439
rect 871 387 926 405
rect 980 580 1035 592
rect 980 546 991 580
rect 1025 546 1035 580
rect 980 511 1035 546
rect 980 477 991 511
rect 1025 477 1035 511
rect 980 442 1035 477
rect 980 408 991 442
rect 1025 408 1035 442
rect 980 392 1035 408
rect 1071 580 1125 592
rect 1071 546 1081 580
rect 1115 546 1125 580
rect 1071 509 1125 546
rect 1071 475 1081 509
rect 1115 475 1125 509
rect 1071 438 1125 475
rect 1071 404 1081 438
rect 1115 404 1125 438
rect 1071 392 1125 404
<< ndiffc >>
rect 39 152 73 186
rect 39 84 73 118
rect 125 176 159 210
rect 125 86 159 120
rect 211 103 245 137
rect 311 176 345 210
rect 311 86 345 120
rect 411 154 445 188
rect 411 86 445 120
rect 511 156 545 190
rect 511 86 545 120
rect 617 154 651 188
rect 617 86 651 120
rect 717 156 751 190
rect 717 86 751 120
rect 803 156 837 190
rect 803 86 837 120
rect 903 154 937 188
rect 972 154 1006 188
rect 1042 154 1076 188
rect 903 86 937 120
rect 972 86 1006 120
rect 1042 86 1076 120
<< pdiffc >>
rect 37 546 71 580
rect 37 463 71 497
rect 37 380 71 414
rect 127 546 161 580
rect 127 463 161 497
rect 127 380 161 414
rect 217 546 251 580
rect 217 444 251 478
rect 307 546 341 580
rect 307 463 341 497
rect 307 380 341 414
rect 397 546 431 580
rect 397 475 431 509
rect 397 404 431 438
rect 502 546 536 580
rect 502 476 536 510
rect 502 406 536 440
rect 592 546 626 580
rect 592 474 626 508
rect 701 541 735 575
rect 701 470 735 504
rect 701 399 735 433
rect 791 497 825 531
rect 791 399 825 433
rect 881 541 915 575
rect 881 473 915 507
rect 881 405 915 439
rect 991 546 1025 580
rect 991 477 1025 511
rect 991 408 1025 442
rect 1081 546 1115 580
rect 1081 475 1115 509
rect 1081 404 1115 438
<< poly >>
rect 81 592 117 618
rect 171 592 207 618
rect 261 592 297 618
rect 351 592 387 618
rect 456 592 492 618
rect 546 592 582 618
rect 745 587 781 613
rect 835 587 871 613
rect 1035 592 1071 618
rect 81 326 117 368
rect 171 326 207 368
rect 261 326 297 368
rect 351 326 387 368
rect 81 310 391 326
rect 81 296 205 310
rect 84 222 114 296
rect 170 276 205 296
rect 239 276 273 310
rect 307 276 341 310
rect 375 276 391 310
rect 170 260 391 276
rect 170 222 200 260
rect 270 222 300 260
rect 361 222 391 260
rect 456 318 492 392
rect 546 356 582 392
rect 540 340 606 356
rect 540 318 556 340
rect 456 306 556 318
rect 590 306 606 340
rect 745 319 781 387
rect 835 355 871 387
rect 1035 358 1071 392
rect 835 339 925 355
rect 835 319 875 339
rect 456 288 606 306
rect 456 202 486 288
rect 576 202 606 288
rect 676 305 875 319
rect 909 305 925 339
rect 676 289 925 305
rect 981 342 1065 358
rect 981 308 997 342
rect 1031 308 1065 342
rect 676 202 706 289
rect 762 202 792 289
rect 981 274 1065 308
rect 981 247 997 274
rect 862 240 997 247
rect 1031 240 1065 274
rect 862 217 1065 240
rect 862 202 892 217
rect 84 48 114 74
rect 170 48 200 74
rect 270 48 300 74
rect 361 48 391 74
rect 456 48 486 74
rect 576 48 606 74
rect 676 48 706 74
rect 762 48 792 74
rect 862 48 892 74
<< polycont >>
rect 205 276 239 310
rect 273 276 307 310
rect 341 276 375 310
rect 556 306 590 340
rect 875 305 909 339
rect 997 308 1031 342
rect 997 240 1031 274
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 21 580 87 649
rect 21 546 37 580
rect 71 546 87 580
rect 21 497 87 546
rect 21 463 37 497
rect 71 463 87 497
rect 21 414 87 463
rect 21 380 37 414
rect 71 380 87 414
rect 21 364 87 380
rect 121 580 161 596
rect 121 546 127 580
rect 121 497 161 546
rect 121 463 127 497
rect 121 414 161 463
rect 201 580 251 649
rect 201 546 217 580
rect 201 478 251 546
rect 201 444 217 478
rect 201 428 251 444
rect 291 580 357 596
rect 291 546 307 580
rect 341 546 357 580
rect 291 497 357 546
rect 291 463 307 497
rect 341 463 357 497
rect 121 380 127 414
rect 291 414 357 463
rect 291 394 307 414
rect 161 380 307 394
rect 341 380 357 414
rect 397 580 447 649
rect 431 546 447 580
rect 397 509 447 546
rect 431 475 447 509
rect 397 438 447 475
rect 431 404 447 438
rect 397 388 447 404
rect 486 580 552 596
rect 486 546 502 580
rect 536 546 552 580
rect 486 510 552 546
rect 486 476 502 510
rect 536 476 552 510
rect 486 440 552 476
rect 592 580 642 649
rect 626 546 642 580
rect 592 508 642 546
rect 626 474 642 508
rect 592 458 642 474
rect 685 581 931 615
rect 685 575 735 581
rect 685 541 701 575
rect 865 575 931 581
rect 685 504 735 541
rect 685 470 701 504
rect 486 406 502 440
rect 536 424 552 440
rect 685 433 735 470
rect 685 424 701 433
rect 536 406 701 424
rect 486 399 701 406
rect 486 390 735 399
rect 685 383 735 390
rect 775 531 825 547
rect 775 497 791 531
rect 775 433 825 497
rect 775 399 791 433
rect 121 360 357 380
rect 121 282 155 360
rect 505 340 647 356
rect 25 236 155 282
rect 189 310 429 326
rect 189 276 205 310
rect 239 276 273 310
rect 307 276 341 310
rect 375 276 429 310
rect 505 306 556 340
rect 590 306 647 340
rect 505 290 647 306
rect 775 290 825 399
rect 865 541 881 575
rect 915 541 931 575
rect 865 507 931 541
rect 865 473 881 507
rect 915 473 931 507
rect 865 439 931 473
rect 865 405 881 439
rect 915 405 931 439
rect 865 389 931 405
rect 975 580 1041 649
rect 975 546 991 580
rect 1025 546 1041 580
rect 975 511 1041 546
rect 975 477 991 511
rect 1025 477 1041 511
rect 975 442 1041 477
rect 975 408 991 442
rect 1025 408 1041 442
rect 975 392 1041 408
rect 1081 580 1131 596
rect 1115 546 1131 580
rect 1081 509 1131 546
rect 1115 475 1131 509
rect 1081 438 1131 475
rect 1115 404 1131 438
rect 189 260 429 276
rect 109 226 155 236
rect 395 256 429 260
rect 701 256 825 290
rect 859 339 925 355
rect 859 305 875 339
rect 909 305 925 339
rect 859 289 925 305
rect 109 210 361 226
rect 395 222 751 256
rect 23 186 73 202
rect 23 152 39 186
rect 23 118 73 152
rect 23 84 39 118
rect 23 17 73 84
rect 109 176 125 210
rect 159 192 311 210
rect 109 120 159 176
rect 295 176 311 192
rect 345 176 361 210
rect 495 190 561 222
rect 109 86 125 120
rect 109 70 159 86
rect 195 137 261 153
rect 195 103 211 137
rect 245 103 261 137
rect 195 17 261 103
rect 295 120 361 176
rect 295 86 311 120
rect 345 86 361 120
rect 295 70 361 86
rect 395 154 411 188
rect 445 154 461 188
rect 395 120 461 154
rect 395 86 411 120
rect 445 86 461 120
rect 395 17 461 86
rect 495 156 511 190
rect 545 156 561 190
rect 701 190 751 222
rect 495 120 561 156
rect 495 86 511 120
rect 545 86 561 120
rect 495 70 561 86
rect 601 154 617 188
rect 651 154 667 188
rect 601 120 667 154
rect 601 86 617 120
rect 651 86 667 120
rect 601 17 667 86
rect 701 156 717 190
rect 701 120 751 156
rect 701 86 717 120
rect 701 70 751 86
rect 787 190 853 206
rect 787 156 803 190
rect 837 156 853 190
rect 787 120 853 156
rect 787 86 803 120
rect 837 86 853 120
rect 787 17 853 86
rect 887 190 925 289
rect 981 342 1047 358
rect 981 308 997 342
rect 1031 308 1047 342
rect 981 274 1047 308
rect 981 240 997 274
rect 1031 240 1047 274
rect 981 224 1047 240
rect 1081 190 1131 404
rect 887 188 1131 190
rect 887 154 903 188
rect 937 154 972 188
rect 1006 154 1042 188
rect 1076 154 1131 188
rect 887 120 1131 154
rect 887 86 903 120
rect 937 86 972 120
rect 1006 86 1042 120
rect 1076 86 1131 120
rect 887 70 1131 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
rlabel comment s 0 0 0 0 4 or2b_4
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 991 242 1025 276 0 FreeSans 340 0 0 0 B_N
port 2 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 B_N
port 2 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 1152 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 777392
string GDS_START 767498
<< end >>
