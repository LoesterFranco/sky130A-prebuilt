magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 1075 325 1125 425
rect 1263 325 1313 425
rect 1075 291 1449 325
rect 22 215 89 257
rect 242 215 554 257
rect 657 215 940 257
rect 1381 181 1449 291
rect 201 145 1449 181
rect 201 51 277 145
rect 389 51 465 145
rect 681 51 757 145
rect 869 51 945 145
rect 1057 51 1133 145
rect 1245 51 1321 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 22 325 81 493
rect 125 359 175 527
rect 219 393 269 493
rect 313 427 363 527
rect 407 393 457 493
rect 501 427 551 527
rect 605 459 1407 493
rect 605 427 655 459
rect 793 427 843 459
rect 699 393 749 425
rect 887 393 937 425
rect 219 359 937 393
rect 981 359 1031 459
rect 1169 359 1219 459
rect 1357 359 1407 459
rect 22 291 1031 325
rect 133 181 167 291
rect 997 257 1031 291
rect 997 215 1344 257
rect 22 147 167 181
rect 22 51 89 147
rect 133 17 167 111
rect 321 17 355 111
rect 509 17 647 111
rect 801 17 835 111
rect 989 17 1023 111
rect 1177 17 1211 111
rect 1365 17 1399 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< labels >>
rlabel locali s 242 215 554 257 6 A
port 1 nsew signal input
rlabel locali s 657 215 940 257 6 B
port 2 nsew signal input
rlabel locali s 22 215 89 257 6 C_N
port 3 nsew signal input
rlabel locali s 1381 181 1449 291 6 Y
port 4 nsew signal output
rlabel locali s 1263 325 1313 425 6 Y
port 4 nsew signal output
rlabel locali s 1245 51 1321 145 6 Y
port 4 nsew signal output
rlabel locali s 1075 325 1125 425 6 Y
port 4 nsew signal output
rlabel locali s 1075 291 1449 325 6 Y
port 4 nsew signal output
rlabel locali s 1057 51 1133 145 6 Y
port 4 nsew signal output
rlabel locali s 869 51 945 145 6 Y
port 4 nsew signal output
rlabel locali s 681 51 757 145 6 Y
port 4 nsew signal output
rlabel locali s 389 51 465 145 6 Y
port 4 nsew signal output
rlabel locali s 201 145 1449 181 6 Y
port 4 nsew signal output
rlabel locali s 201 51 277 145 6 Y
port 4 nsew signal output
rlabel metal1 s 0 -48 1472 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 1472 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1472 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2474650
string GDS_START 2464006
<< end >>
