magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 644 561
rect 18 451 85 527
rect 17 153 65 415
rect 213 383 279 527
rect 459 367 525 527
rect 559 441 627 493
rect 177 72 247 265
rect 283 71 343 265
rect 379 71 435 265
rect 471 17 525 177
rect 575 161 627 441
rect 559 59 627 161
rect 0 -17 644 17
<< obsli1 >>
rect 119 333 169 493
rect 316 333 366 493
rect 99 299 537 333
rect 99 117 133 299
rect 474 265 537 299
rect 34 51 133 117
rect 474 215 540 265
<< metal1 >>
rect 0 496 644 592
rect 0 -48 644 48
<< labels >>
rlabel locali s 17 153 65 415 6 A
port 1 nsew signal input
rlabel locali s 177 72 247 265 6 B
port 2 nsew signal input
rlabel locali s 283 71 343 265 6 C
port 3 nsew signal input
rlabel locali s 379 71 435 265 6 D
port 4 nsew signal input
rlabel locali s 575 161 627 441 6 X
port 5 nsew signal output
rlabel locali s 559 441 627 493 6 X
port 5 nsew signal output
rlabel locali s 559 59 627 161 6 X
port 5 nsew signal output
rlabel locali s 471 17 525 177 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 644 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 644 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 459 367 525 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 213 383 279 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 18 451 85 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 644 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 644 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3821246
string GDS_START 3814892
<< end >>
