magic
tech sky130A
magscale 1 2
timestamp 1604502697
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 89 47 119 177
rect 183 47 213 177
rect 267 47 297 177
rect 477 47 507 177
rect 571 47 601 177
rect 665 47 695 177
rect 759 47 789 177
<< pmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 469 297 505 497
rect 563 297 599 497
rect 657 297 693 497
rect 751 297 787 497
<< ndiff >>
rect 27 165 89 177
rect 27 131 35 165
rect 69 131 89 165
rect 27 97 89 131
rect 27 63 35 97
rect 69 63 89 97
rect 27 47 89 63
rect 119 95 183 177
rect 119 61 129 95
rect 163 61 183 95
rect 119 47 183 61
rect 213 165 267 177
rect 213 131 223 165
rect 257 131 267 165
rect 213 97 267 131
rect 213 63 223 97
rect 257 63 267 97
rect 213 47 267 63
rect 297 95 477 177
rect 297 61 317 95
rect 351 61 423 95
rect 457 61 477 95
rect 297 47 477 61
rect 507 163 571 177
rect 507 129 517 163
rect 551 129 571 163
rect 507 95 571 129
rect 507 61 517 95
rect 551 61 571 95
rect 507 47 571 61
rect 601 95 665 177
rect 601 61 611 95
rect 645 61 665 95
rect 601 47 665 61
rect 695 163 759 177
rect 695 129 705 163
rect 739 129 759 163
rect 695 95 759 129
rect 695 61 705 95
rect 739 61 759 95
rect 695 47 759 61
rect 789 95 852 177
rect 789 61 799 95
rect 833 61 852 95
rect 789 47 852 61
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 297 175 497
rect 211 297 269 497
rect 305 485 469 497
rect 305 451 330 485
rect 364 451 423 485
rect 457 451 469 485
rect 305 417 469 451
rect 305 383 330 417
rect 364 383 423 417
rect 457 383 469 417
rect 305 297 469 383
rect 505 477 563 497
rect 505 443 517 477
rect 551 443 563 477
rect 505 409 563 443
rect 505 375 517 409
rect 551 375 563 409
rect 505 341 563 375
rect 505 307 517 341
rect 551 307 563 341
rect 505 297 563 307
rect 599 477 657 497
rect 599 443 611 477
rect 645 443 657 477
rect 599 409 657 443
rect 599 375 611 409
rect 645 375 657 409
rect 599 297 657 375
rect 693 477 751 497
rect 693 443 705 477
rect 739 443 751 477
rect 693 409 751 443
rect 693 375 705 409
rect 739 375 751 409
rect 693 341 751 375
rect 693 307 705 341
rect 739 307 751 341
rect 693 297 751 307
rect 787 477 861 497
rect 787 443 799 477
rect 833 443 861 477
rect 787 409 861 443
rect 787 375 799 409
rect 833 375 861 409
rect 787 297 861 375
<< ndiffc >>
rect 35 131 69 165
rect 35 63 69 97
rect 129 61 163 95
rect 223 131 257 165
rect 223 63 257 97
rect 317 61 351 95
rect 423 61 457 95
rect 517 129 551 163
rect 517 61 551 95
rect 611 61 645 95
rect 705 129 739 163
rect 705 61 739 95
rect 799 61 833 95
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 330 451 364 485
rect 423 451 457 485
rect 330 383 364 417
rect 423 383 457 417
rect 517 443 551 477
rect 517 375 551 409
rect 517 307 551 341
rect 611 443 645 477
rect 611 375 645 409
rect 705 443 739 477
rect 705 375 739 409
rect 705 307 739 341
rect 799 443 833 477
rect 799 375 833 409
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 469 497 505 523
rect 563 497 599 523
rect 657 497 693 523
rect 751 497 787 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 469 282 505 297
rect 563 282 599 297
rect 657 282 693 297
rect 751 282 787 297
rect 79 265 119 282
rect 173 265 213 282
rect 267 265 307 282
rect 467 265 507 282
rect 561 265 601 282
rect 655 265 695 282
rect 749 265 789 282
rect 25 249 119 265
rect 25 215 35 249
rect 69 215 119 249
rect 25 199 119 215
rect 161 249 225 265
rect 161 215 171 249
rect 205 215 225 249
rect 161 199 225 215
rect 267 249 335 265
rect 267 215 281 249
rect 315 215 335 249
rect 267 199 335 215
rect 410 249 789 265
rect 410 215 426 249
rect 460 215 494 249
rect 528 215 572 249
rect 606 215 650 249
rect 684 215 728 249
rect 762 215 789 249
rect 410 199 789 215
rect 89 177 119 199
rect 183 177 213 199
rect 267 177 297 199
rect 477 177 507 199
rect 571 177 601 199
rect 665 177 695 199
rect 759 177 789 199
rect 89 21 119 47
rect 183 21 213 47
rect 267 21 297 47
rect 477 21 507 47
rect 571 21 601 47
rect 665 21 695 47
rect 759 21 789 47
<< polycont >>
rect 35 215 69 249
rect 171 215 205 249
rect 281 215 315 249
rect 426 215 460 249
rect 494 215 528 249
rect 572 215 606 249
rect 650 215 684 249
rect 728 215 762 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 17 485 273 493
rect 17 451 35 485
rect 69 459 273 485
rect 69 451 85 459
rect 17 417 85 451
rect 17 383 35 417
rect 69 383 85 417
rect 17 349 85 383
rect 17 315 35 349
rect 69 315 85 349
rect 17 299 85 315
rect 119 265 166 410
rect 220 333 273 459
rect 317 485 457 527
rect 317 451 330 485
rect 364 451 423 485
rect 317 417 457 451
rect 317 383 330 417
rect 364 383 423 417
rect 317 367 457 383
rect 509 477 559 493
rect 509 443 517 477
rect 551 443 559 477
rect 509 409 559 443
rect 509 375 517 409
rect 551 375 559 409
rect 509 341 559 375
rect 603 477 653 527
rect 603 443 611 477
rect 645 443 653 477
rect 603 409 653 443
rect 603 375 611 409
rect 645 375 653 409
rect 603 359 653 375
rect 697 477 747 493
rect 697 443 705 477
rect 739 443 747 477
rect 697 409 747 443
rect 697 375 705 409
rect 739 375 747 409
rect 220 299 448 333
rect 17 249 85 265
rect 17 215 35 249
rect 69 215 85 249
rect 119 249 231 265
rect 119 215 171 249
rect 205 215 231 249
rect 265 249 370 265
rect 265 215 281 249
rect 315 215 370 249
rect 404 249 448 299
rect 509 307 517 341
rect 551 323 559 341
rect 697 341 747 375
rect 791 477 841 527
rect 791 443 799 477
rect 833 443 841 477
rect 791 409 841 443
rect 791 375 799 409
rect 833 375 841 409
rect 791 359 841 375
rect 697 323 705 341
rect 551 307 705 323
rect 739 323 747 341
rect 739 307 891 323
rect 509 289 891 307
rect 404 215 426 249
rect 460 215 494 249
rect 528 215 572 249
rect 606 215 650 249
rect 684 215 728 249
rect 762 215 789 249
rect 404 181 448 215
rect 823 181 891 289
rect 17 165 448 181
rect 17 131 35 165
rect 69 145 223 165
rect 69 131 85 145
rect 17 97 85 131
rect 197 131 223 145
rect 257 145 448 165
rect 491 163 891 181
rect 257 131 273 145
rect 17 63 35 97
rect 69 63 85 97
rect 17 51 85 63
rect 129 95 163 111
rect 129 17 163 61
rect 197 97 273 131
rect 491 129 517 163
rect 551 147 705 163
rect 551 129 567 147
rect 197 63 223 97
rect 257 63 273 97
rect 197 51 273 63
rect 317 95 457 111
rect 351 61 423 95
rect 317 17 457 61
rect 491 95 567 129
rect 679 129 705 147
rect 739 147 891 163
rect 739 129 755 147
rect 491 61 517 95
rect 551 61 567 95
rect 491 53 567 61
rect 611 95 645 111
rect 611 17 645 61
rect 679 95 755 129
rect 679 61 705 95
rect 739 61 755 95
rect 679 53 755 61
rect 799 95 833 111
rect 799 17 833 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel corelocali s 305 221 339 255 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 857 153 891 187 0 FreeSans 200 0 0 0 X
port 8 nsew
flabel corelocali s 121 357 155 391 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel corelocali s 29 221 63 255 0 FreeSans 400 0 0 0 C
port 3 nsew
flabel corelocali s 121 289 155 323 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
rlabel comment s 0 0 0 0 4 or3_4
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 472498
string GDS_START 465056
<< end >>
