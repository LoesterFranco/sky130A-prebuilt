magic
tech sky130A
magscale 1 2
timestamp 1604502741
<< locali >>
rect 21 260 223 356
rect 453 430 575 596
rect 963 430 1029 596
rect 453 390 1029 430
rect 453 370 839 390
rect 657 252 731 370
rect 889 326 1131 356
rect 769 260 1131 326
rect 325 218 731 252
rect 325 127 377 218
rect 511 127 576 218
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 87 390 212 649
rect 246 390 312 540
rect 257 336 291 390
rect 353 370 419 649
rect 609 464 929 649
rect 1063 390 1120 649
rect 257 286 615 336
rect 257 226 291 286
rect 27 192 291 226
rect 27 70 77 192
rect 113 17 179 158
rect 239 85 291 158
rect 411 85 477 184
rect 796 192 1129 226
rect 796 184 862 192
rect 610 150 862 184
rect 610 85 676 150
rect 239 51 676 85
rect 710 17 776 116
rect 810 66 862 150
rect 896 17 1029 158
rect 1063 70 1129 192
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
rlabel locali s 21 260 223 356 6 A_N
port 1 nsew signal input
rlabel locali s 889 326 1131 356 6 B
port 2 nsew signal input
rlabel locali s 769 260 1131 326 6 B
port 2 nsew signal input
rlabel locali s 963 430 1029 596 6 Y
port 3 nsew signal output
rlabel locali s 657 252 731 370 6 Y
port 3 nsew signal output
rlabel locali s 511 127 576 218 6 Y
port 3 nsew signal output
rlabel locali s 453 430 575 596 6 Y
port 3 nsew signal output
rlabel locali s 453 390 1029 430 6 Y
port 3 nsew signal output
rlabel locali s 453 370 839 390 6 Y
port 3 nsew signal output
rlabel locali s 325 218 731 252 6 Y
port 3 nsew signal output
rlabel locali s 325 127 377 218 6 Y
port 3 nsew signal output
rlabel metal1 s 0 -49 1152 49 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 617 1152 715 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1997604
string GDS_START 1988448
<< end >>
