magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 18 333 85 490
rect 18 299 155 333
rect 17 149 67 265
rect 103 165 155 299
rect 193 199 257 490
rect 291 199 349 490
rect 103 131 353 165
rect 387 131 441 333
rect 103 77 163 131
rect 319 77 353 131
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 427 367 507 527
rect 17 17 69 115
rect 207 17 273 97
rect 401 17 504 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
rlabel locali s 387 131 441 333 6 A
port 1 nsew signal input
rlabel locali s 291 199 349 490 6 B
port 2 nsew signal input
rlabel locali s 193 199 257 490 6 C
port 3 nsew signal input
rlabel locali s 17 149 67 265 6 D
port 4 nsew signal input
rlabel locali s 319 77 353 131 6 Y
port 5 nsew signal output
rlabel locali s 103 165 155 299 6 Y
port 5 nsew signal output
rlabel locali s 103 131 353 165 6 Y
port 5 nsew signal output
rlabel locali s 103 77 163 131 6 Y
port 5 nsew signal output
rlabel locali s 18 333 85 490 6 Y
port 5 nsew signal output
rlabel locali s 18 299 155 333 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -48 552 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 552 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 552 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2479588
string GDS_START 2474708
<< end >>
