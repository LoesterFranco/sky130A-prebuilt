magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 17 214 66 323
rect 112 214 188 323
rect 437 333 497 493
rect 625 333 701 493
rect 911 333 987 493
rect 1099 333 1175 493
rect 437 289 1175 333
rect 437 131 526 289
rect 699 215 809 289
rect 848 215 990 255
rect 1063 215 1259 255
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 17 396 74 488
rect 108 439 163 527
rect 197 430 335 493
rect 17 357 266 396
rect 232 180 266 357
rect 17 146 266 180
rect 17 51 69 146
rect 300 112 335 430
rect 369 299 403 527
rect 531 367 591 527
rect 745 367 877 527
rect 1031 367 1065 527
rect 1219 289 1269 527
rect 589 215 665 255
rect 625 131 987 181
rect 1031 147 1269 181
rect 103 17 163 109
rect 197 51 335 112
rect 369 97 403 117
rect 1031 97 1081 147
rect 369 51 795 97
rect 833 51 1081 97
rect 1125 17 1159 113
rect 1193 51 1269 147
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< obsm1 >>
rect 220 215 677 261
<< labels >>
rlabel locali s 112 214 188 323 6 A_N
port 1 nsew signal input
rlabel locali s 17 214 66 323 6 B_N
port 2 nsew signal input
rlabel locali s 848 215 990 255 6 C
port 3 nsew signal input
rlabel locali s 1063 215 1259 255 6 D
port 4 nsew signal input
rlabel locali s 1099 333 1175 493 6 Y
port 5 nsew signal output
rlabel locali s 911 333 987 493 6 Y
port 5 nsew signal output
rlabel locali s 699 215 809 289 6 Y
port 5 nsew signal output
rlabel locali s 625 333 701 493 6 Y
port 5 nsew signal output
rlabel locali s 437 333 497 493 6 Y
port 5 nsew signal output
rlabel locali s 437 289 1175 333 6 Y
port 5 nsew signal output
rlabel locali s 437 131 526 289 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -48 1288 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 1288 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1288 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2365382
string GDS_START 2354786
<< end >>
