magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 2484 561
rect 120 436 154 527
rect 190 215 268 255
rect 126 17 160 109
rect 302 133 348 265
rect 1052 447 1118 527
rect 1340 335 1374 357
rect 848 129 898 265
rect 1036 17 1102 161
rect 1320 185 1374 335
rect 2038 439 2072 527
rect 1320 151 1385 185
rect 1351 119 1385 151
rect 2315 357 2366 527
rect 2400 357 2467 493
rect 2104 215 2193 255
rect 2036 17 2070 113
rect 2425 165 2467 357
rect 2299 17 2365 102
rect 2399 51 2467 165
rect 0 -17 2484 17
<< obsli1 >>
rect 17 402 86 493
rect 343 477 703 493
rect 188 459 703 477
rect 188 443 394 459
rect 188 402 222 443
rect 649 422 692 459
rect 17 368 222 402
rect 256 391 290 409
rect 513 391 579 409
rect 17 300 88 368
rect 256 357 376 391
rect 513 357 514 391
rect 548 357 579 391
rect 256 334 290 357
rect 122 300 290 334
rect 17 161 51 300
rect 122 265 156 300
rect 444 270 478 357
rect 85 199 156 265
rect 122 181 156 199
rect 17 147 86 161
rect 122 147 265 181
rect 20 51 86 147
rect 199 93 265 147
rect 397 255 478 270
rect 431 221 478 255
rect 590 253 624 289
rect 560 249 624 253
rect 397 135 478 221
rect 528 219 624 249
rect 528 215 594 219
rect 658 185 692 422
rect 742 458 1013 492
rect 742 264 776 458
rect 816 391 889 424
rect 816 357 828 391
rect 862 357 889 391
rect 963 413 1013 458
rect 1165 459 1590 493
rect 1165 413 1199 459
rect 963 379 1199 413
rect 1240 391 1442 425
rect 1240 379 1306 391
rect 816 339 889 357
rect 1240 345 1274 379
rect 938 323 1034 345
rect 938 289 952 323
rect 986 289 1034 323
rect 1127 311 1274 345
rect 938 277 1034 289
rect 966 265 1034 277
rect 742 230 814 264
rect 611 181 746 185
rect 444 119 478 135
rect 524 151 746 181
rect 524 147 627 151
rect 524 131 605 147
rect 643 93 678 117
rect 199 85 420 93
rect 503 85 678 93
rect 199 51 678 85
rect 712 85 746 151
rect 780 119 814 230
rect 966 199 1126 265
rect 966 102 1000 199
rect 1160 163 1194 311
rect 848 85 914 95
rect 712 51 914 85
rect 1136 76 1194 163
rect 1228 255 1285 265
rect 1262 221 1285 255
rect 1228 148 1285 221
rect 1408 246 1442 391
rect 1476 306 1510 425
rect 1556 344 1590 459
rect 1644 459 1882 493
rect 1644 391 1678 459
rect 1712 357 1778 425
rect 1556 310 1607 344
rect 1476 272 1522 306
rect 1488 258 1522 272
rect 1408 212 1454 246
rect 1488 221 1539 258
rect 1420 185 1454 212
rect 1504 187 1539 221
rect 1573 199 1607 310
rect 1675 323 1778 357
rect 1675 289 1688 323
rect 1722 306 1778 323
rect 1848 409 1882 459
rect 1848 408 2021 409
rect 1848 407 2024 408
rect 1848 406 2026 407
rect 1848 405 2029 406
rect 2107 405 2177 493
rect 1848 375 2177 405
rect 1722 289 1734 306
rect 1420 119 1470 185
rect 1538 153 1539 187
rect 1675 185 1711 289
rect 1767 255 1814 265
rect 1767 221 1780 255
rect 1767 199 1814 221
rect 1251 85 1317 114
rect 1504 85 1539 153
rect 1251 51 1539 85
rect 1573 85 1607 148
rect 1661 119 1711 185
rect 1848 153 1882 375
rect 2011 374 2177 375
rect 2014 373 2177 374
rect 2017 372 2177 373
rect 2020 371 2177 372
rect 1745 119 1882 153
rect 1928 307 2002 341
rect 1928 165 1962 307
rect 2036 289 2177 371
rect 2215 291 2281 493
rect 2036 265 2070 289
rect 1996 199 2070 265
rect 2036 181 2070 199
rect 2231 187 2281 291
rect 2329 289 2336 323
rect 2370 289 2391 323
rect 2329 199 2391 289
rect 1928 85 1996 165
rect 2036 147 2182 181
rect 1573 51 1996 85
rect 2106 57 2182 147
rect 2231 153 2244 187
rect 2278 153 2281 187
rect 2231 136 2281 153
rect 2231 54 2265 136
<< obsli1c >>
rect 376 357 410 391
rect 514 357 548 391
rect 397 221 431 255
rect 590 289 624 323
rect 828 357 862 391
rect 952 289 986 323
rect 1228 221 1262 255
rect 1688 289 1722 323
rect 1504 153 1538 187
rect 1780 221 1814 255
rect 2336 289 2370 323
rect 2244 153 2278 187
<< metal1 >>
rect 0 496 2484 592
rect 293 184 351 193
rect 845 184 903 193
rect 293 156 903 184
rect 293 147 351 156
rect 845 147 903 156
rect 0 -48 2484 48
<< obsm1 >>
rect 364 391 422 397
rect 364 357 376 391
rect 410 388 422 391
rect 502 391 560 397
rect 502 388 514 391
rect 410 360 514 388
rect 410 357 422 360
rect 364 351 422 357
rect 502 357 514 360
rect 548 388 560 391
rect 816 391 874 397
rect 816 388 828 391
rect 548 360 828 388
rect 548 357 560 360
rect 502 351 560 357
rect 816 357 828 360
rect 862 357 874 391
rect 816 351 874 357
rect 578 323 636 329
rect 578 289 590 323
rect 624 320 636 323
rect 940 323 998 329
rect 940 320 952 323
rect 624 292 952 320
rect 624 289 636 292
rect 578 283 636 289
rect 940 289 952 292
rect 986 289 998 323
rect 940 283 998 289
rect 1676 323 1734 329
rect 1676 289 1688 323
rect 1722 320 1734 323
rect 2324 323 2382 329
rect 2324 320 2336 323
rect 1722 292 2336 320
rect 1722 289 1734 292
rect 1676 283 1734 289
rect 2324 289 2336 292
rect 2370 289 2382 323
rect 2324 283 2382 289
rect 385 255 443 261
rect 385 221 397 255
rect 431 252 443 255
rect 1216 255 1274 261
rect 1216 252 1228 255
rect 431 224 1228 252
rect 431 221 443 224
rect 385 215 443 221
rect 1216 221 1228 224
rect 1262 252 1274 255
rect 1768 255 1826 261
rect 1768 252 1780 255
rect 1262 224 1780 252
rect 1262 221 1274 224
rect 1216 215 1274 221
rect 1768 221 1780 224
rect 1814 221 1826 255
rect 1768 215 1826 221
rect 1492 187 1550 193
rect 1492 153 1504 187
rect 1538 184 1550 187
rect 2232 187 2290 193
rect 2232 184 2244 187
rect 1538 156 2244 184
rect 1538 153 1550 156
rect 1492 147 1550 153
rect 2232 153 2244 156
rect 2278 153 2290 187
rect 2232 147 2290 153
<< labels >>
rlabel locali s 190 215 268 255 6 A
port 1 nsew signal input
rlabel locali s 302 133 348 265 6 B
port 2 nsew signal input
rlabel locali s 848 129 898 265 6 B
port 2 nsew signal input
rlabel metal1 s 845 184 903 193 6 B
port 2 nsew signal input
rlabel metal1 s 845 147 903 156 6 B
port 2 nsew signal input
rlabel metal1 s 293 184 351 193 6 B
port 2 nsew signal input
rlabel metal1 s 293 156 903 184 6 B
port 2 nsew signal input
rlabel metal1 s 293 147 351 156 6 B
port 2 nsew signal input
rlabel locali s 2104 215 2193 255 6 CIN
port 3 nsew signal input
rlabel locali s 1351 119 1385 151 6 COUT
port 4 nsew signal output
rlabel locali s 1340 335 1374 357 6 COUT
port 4 nsew signal output
rlabel locali s 1320 185 1374 335 6 COUT
port 4 nsew signal output
rlabel locali s 1320 151 1385 185 6 COUT
port 4 nsew signal output
rlabel locali s 2425 165 2467 357 6 SUM
port 5 nsew signal output
rlabel locali s 2400 357 2467 493 6 SUM
port 5 nsew signal output
rlabel locali s 2399 51 2467 165 6 SUM
port 5 nsew signal output
rlabel locali s 2299 17 2365 102 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 2036 17 2070 113 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1036 17 1102 161 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 126 17 160 109 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 2484 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 2484 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 2315 357 2366 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 2038 439 2072 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1052 447 1118 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 120 436 154 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 2484 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 2484 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2484 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2087298
string GDS_START 2068014
<< end >>
