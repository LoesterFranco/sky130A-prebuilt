magic
tech sky130A
magscale 1 2
timestamp 1604502697
<< nwell >>
rect -38 261 2522 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 79 47 109 177
rect 173 47 203 177
rect 277 47 307 177
rect 361 47 391 177
rect 455 47 485 177
rect 549 47 579 177
rect 643 47 673 177
rect 737 47 767 177
rect 841 47 871 177
rect 925 47 955 177
rect 1019 47 1049 177
rect 1113 47 1143 177
rect 1207 47 1237 177
rect 1301 47 1331 177
rect 1395 47 1425 177
rect 1489 47 1519 177
rect 1583 47 1613 177
rect 1677 47 1707 177
rect 1771 47 1801 177
rect 1865 47 1895 177
rect 1959 47 1989 177
rect 2053 47 2083 177
rect 2147 47 2177 177
rect 2241 47 2271 177
rect 2345 47 2375 177
<< pmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 457 297 493 497
rect 551 297 587 497
rect 645 297 681 497
rect 739 297 775 497
rect 833 297 869 497
rect 927 297 963 497
rect 1021 297 1057 497
rect 1115 297 1151 497
rect 1209 297 1245 497
rect 1303 297 1339 497
rect 1397 297 1433 497
rect 1491 297 1527 497
rect 1585 297 1621 497
rect 1679 297 1715 497
rect 1773 297 1809 497
rect 1867 297 1903 497
rect 1961 297 1997 497
rect 2055 297 2091 497
rect 2149 297 2185 497
rect 2243 297 2279 497
rect 2337 297 2373 497
<< ndiff >>
rect 27 165 79 177
rect 27 131 35 165
rect 69 131 79 165
rect 27 97 79 131
rect 27 63 35 97
rect 69 63 79 97
rect 27 47 79 63
rect 109 97 173 177
rect 109 63 129 97
rect 163 63 173 97
rect 109 47 173 63
rect 203 165 277 177
rect 203 131 223 165
rect 257 131 277 165
rect 203 97 277 131
rect 203 63 223 97
rect 257 63 277 97
rect 203 47 277 63
rect 307 97 361 177
rect 307 63 317 97
rect 351 63 361 97
rect 307 47 361 63
rect 391 165 455 177
rect 391 131 411 165
rect 445 131 455 165
rect 391 97 455 131
rect 391 63 411 97
rect 445 63 455 97
rect 391 47 455 63
rect 485 97 549 177
rect 485 63 505 97
rect 539 63 549 97
rect 485 47 549 63
rect 579 165 643 177
rect 579 131 599 165
rect 633 131 643 165
rect 579 97 643 131
rect 579 63 599 97
rect 633 63 643 97
rect 579 47 643 63
rect 673 97 737 177
rect 673 63 693 97
rect 727 63 737 97
rect 673 47 737 63
rect 767 165 841 177
rect 767 131 787 165
rect 821 131 841 165
rect 767 97 841 131
rect 767 63 787 97
rect 821 63 841 97
rect 767 47 841 63
rect 871 97 925 177
rect 871 63 881 97
rect 915 63 925 97
rect 871 47 925 63
rect 955 165 1019 177
rect 955 131 975 165
rect 1009 131 1019 165
rect 955 97 1019 131
rect 955 63 975 97
rect 1009 63 1019 97
rect 955 47 1019 63
rect 1049 97 1113 177
rect 1049 63 1069 97
rect 1103 63 1113 97
rect 1049 47 1113 63
rect 1143 165 1207 177
rect 1143 131 1163 165
rect 1197 131 1207 165
rect 1143 97 1207 131
rect 1143 63 1163 97
rect 1197 63 1207 97
rect 1143 47 1207 63
rect 1237 97 1301 177
rect 1237 63 1257 97
rect 1291 63 1301 97
rect 1237 47 1301 63
rect 1331 165 1395 177
rect 1331 131 1351 165
rect 1385 131 1395 165
rect 1331 97 1395 131
rect 1331 63 1351 97
rect 1385 63 1395 97
rect 1331 47 1395 63
rect 1425 97 1489 177
rect 1425 63 1445 97
rect 1479 63 1489 97
rect 1425 47 1489 63
rect 1519 165 1583 177
rect 1519 131 1539 165
rect 1573 131 1583 165
rect 1519 97 1583 131
rect 1519 63 1539 97
rect 1573 63 1583 97
rect 1519 47 1583 63
rect 1613 97 1677 177
rect 1613 63 1633 97
rect 1667 63 1677 97
rect 1613 47 1677 63
rect 1707 165 1771 177
rect 1707 131 1727 165
rect 1761 131 1771 165
rect 1707 97 1771 131
rect 1707 63 1727 97
rect 1761 63 1771 97
rect 1707 47 1771 63
rect 1801 97 1865 177
rect 1801 63 1821 97
rect 1855 63 1865 97
rect 1801 47 1865 63
rect 1895 165 1959 177
rect 1895 131 1915 165
rect 1949 131 1959 165
rect 1895 97 1959 131
rect 1895 63 1915 97
rect 1949 63 1959 97
rect 1895 47 1959 63
rect 1989 97 2053 177
rect 1989 63 2009 97
rect 2043 63 2053 97
rect 1989 47 2053 63
rect 2083 165 2147 177
rect 2083 131 2103 165
rect 2137 131 2147 165
rect 2083 97 2147 131
rect 2083 63 2103 97
rect 2137 63 2147 97
rect 2083 47 2147 63
rect 2177 97 2241 177
rect 2177 63 2197 97
rect 2231 63 2241 97
rect 2177 47 2241 63
rect 2271 165 2345 177
rect 2271 131 2291 165
rect 2325 131 2345 165
rect 2271 97 2345 131
rect 2271 63 2291 97
rect 2325 63 2345 97
rect 2271 47 2345 63
rect 2375 97 2427 177
rect 2375 63 2385 97
rect 2419 63 2427 97
rect 2375 47 2427 63
<< pdiff >>
rect 27 479 81 497
rect 27 445 35 479
rect 69 445 81 479
rect 27 411 81 445
rect 27 377 35 411
rect 69 377 81 411
rect 27 343 81 377
rect 27 309 35 343
rect 69 309 81 343
rect 27 297 81 309
rect 117 485 175 497
rect 117 451 129 485
rect 163 451 175 485
rect 117 417 175 451
rect 117 383 129 417
rect 163 383 175 417
rect 117 297 175 383
rect 211 479 269 497
rect 211 445 223 479
rect 257 445 269 479
rect 211 411 269 445
rect 211 377 223 411
rect 257 377 269 411
rect 211 343 269 377
rect 211 309 223 343
rect 257 309 269 343
rect 211 297 269 309
rect 305 485 363 497
rect 305 451 317 485
rect 351 451 363 485
rect 305 417 363 451
rect 305 383 317 417
rect 351 383 363 417
rect 305 297 363 383
rect 399 479 457 497
rect 399 445 411 479
rect 445 445 457 479
rect 399 411 457 445
rect 399 377 411 411
rect 445 377 457 411
rect 399 343 457 377
rect 399 309 411 343
rect 445 309 457 343
rect 399 297 457 309
rect 493 485 551 497
rect 493 451 505 485
rect 539 451 551 485
rect 493 417 551 451
rect 493 383 505 417
rect 539 383 551 417
rect 493 297 551 383
rect 587 479 645 497
rect 587 445 599 479
rect 633 445 645 479
rect 587 411 645 445
rect 587 377 599 411
rect 633 377 645 411
rect 587 343 645 377
rect 587 309 599 343
rect 633 309 645 343
rect 587 297 645 309
rect 681 485 739 497
rect 681 451 693 485
rect 727 451 739 485
rect 681 417 739 451
rect 681 383 693 417
rect 727 383 739 417
rect 681 297 739 383
rect 775 479 833 497
rect 775 445 787 479
rect 821 445 833 479
rect 775 411 833 445
rect 775 377 787 411
rect 821 377 833 411
rect 775 343 833 377
rect 775 309 787 343
rect 821 309 833 343
rect 775 297 833 309
rect 869 485 927 497
rect 869 451 881 485
rect 915 451 927 485
rect 869 417 927 451
rect 869 383 881 417
rect 915 383 927 417
rect 869 297 927 383
rect 963 479 1021 497
rect 963 445 975 479
rect 1009 445 1021 479
rect 963 411 1021 445
rect 963 377 975 411
rect 1009 377 1021 411
rect 963 343 1021 377
rect 963 309 975 343
rect 1009 309 1021 343
rect 963 297 1021 309
rect 1057 485 1115 497
rect 1057 451 1069 485
rect 1103 451 1115 485
rect 1057 417 1115 451
rect 1057 383 1069 417
rect 1103 383 1115 417
rect 1057 297 1115 383
rect 1151 479 1209 497
rect 1151 445 1163 479
rect 1197 445 1209 479
rect 1151 411 1209 445
rect 1151 377 1163 411
rect 1197 377 1209 411
rect 1151 343 1209 377
rect 1151 309 1163 343
rect 1197 309 1209 343
rect 1151 297 1209 309
rect 1245 485 1303 497
rect 1245 451 1257 485
rect 1291 451 1303 485
rect 1245 417 1303 451
rect 1245 383 1257 417
rect 1291 383 1303 417
rect 1245 297 1303 383
rect 1339 479 1397 497
rect 1339 445 1351 479
rect 1385 445 1397 479
rect 1339 411 1397 445
rect 1339 377 1351 411
rect 1385 377 1397 411
rect 1339 343 1397 377
rect 1339 309 1351 343
rect 1385 309 1397 343
rect 1339 297 1397 309
rect 1433 485 1491 497
rect 1433 451 1445 485
rect 1479 451 1491 485
rect 1433 417 1491 451
rect 1433 383 1445 417
rect 1479 383 1491 417
rect 1433 297 1491 383
rect 1527 479 1585 497
rect 1527 445 1539 479
rect 1573 445 1585 479
rect 1527 411 1585 445
rect 1527 377 1539 411
rect 1573 377 1585 411
rect 1527 343 1585 377
rect 1527 309 1539 343
rect 1573 309 1585 343
rect 1527 297 1585 309
rect 1621 485 1679 497
rect 1621 451 1633 485
rect 1667 451 1679 485
rect 1621 417 1679 451
rect 1621 383 1633 417
rect 1667 383 1679 417
rect 1621 297 1679 383
rect 1715 479 1773 497
rect 1715 445 1727 479
rect 1761 445 1773 479
rect 1715 411 1773 445
rect 1715 377 1727 411
rect 1761 377 1773 411
rect 1715 343 1773 377
rect 1715 309 1727 343
rect 1761 309 1773 343
rect 1715 297 1773 309
rect 1809 485 1867 497
rect 1809 451 1821 485
rect 1855 451 1867 485
rect 1809 417 1867 451
rect 1809 383 1821 417
rect 1855 383 1867 417
rect 1809 297 1867 383
rect 1903 479 1961 497
rect 1903 445 1915 479
rect 1949 445 1961 479
rect 1903 411 1961 445
rect 1903 377 1915 411
rect 1949 377 1961 411
rect 1903 343 1961 377
rect 1903 309 1915 343
rect 1949 309 1961 343
rect 1903 297 1961 309
rect 1997 485 2055 497
rect 1997 451 2009 485
rect 2043 451 2055 485
rect 1997 417 2055 451
rect 1997 383 2009 417
rect 2043 383 2055 417
rect 1997 297 2055 383
rect 2091 479 2149 497
rect 2091 445 2103 479
rect 2137 445 2149 479
rect 2091 411 2149 445
rect 2091 377 2103 411
rect 2137 377 2149 411
rect 2091 343 2149 377
rect 2091 309 2103 343
rect 2137 309 2149 343
rect 2091 297 2149 309
rect 2185 485 2243 497
rect 2185 451 2197 485
rect 2231 451 2243 485
rect 2185 417 2243 451
rect 2185 383 2197 417
rect 2231 383 2243 417
rect 2185 297 2243 383
rect 2279 479 2337 497
rect 2279 445 2291 479
rect 2325 445 2337 479
rect 2279 411 2337 445
rect 2279 377 2291 411
rect 2325 377 2337 411
rect 2279 343 2337 377
rect 2279 309 2291 343
rect 2325 309 2337 343
rect 2279 297 2337 309
rect 2373 485 2427 497
rect 2373 451 2385 485
rect 2419 451 2427 485
rect 2373 417 2427 451
rect 2373 383 2385 417
rect 2419 383 2427 417
rect 2373 297 2427 383
<< ndiffc >>
rect 35 131 69 165
rect 35 63 69 97
rect 129 63 163 97
rect 223 131 257 165
rect 223 63 257 97
rect 317 63 351 97
rect 411 131 445 165
rect 411 63 445 97
rect 505 63 539 97
rect 599 131 633 165
rect 599 63 633 97
rect 693 63 727 97
rect 787 131 821 165
rect 787 63 821 97
rect 881 63 915 97
rect 975 131 1009 165
rect 975 63 1009 97
rect 1069 63 1103 97
rect 1163 131 1197 165
rect 1163 63 1197 97
rect 1257 63 1291 97
rect 1351 131 1385 165
rect 1351 63 1385 97
rect 1445 63 1479 97
rect 1539 131 1573 165
rect 1539 63 1573 97
rect 1633 63 1667 97
rect 1727 131 1761 165
rect 1727 63 1761 97
rect 1821 63 1855 97
rect 1915 131 1949 165
rect 1915 63 1949 97
rect 2009 63 2043 97
rect 2103 131 2137 165
rect 2103 63 2137 97
rect 2197 63 2231 97
rect 2291 131 2325 165
rect 2291 63 2325 97
rect 2385 63 2419 97
<< pdiffc >>
rect 35 445 69 479
rect 35 377 69 411
rect 35 309 69 343
rect 129 451 163 485
rect 129 383 163 417
rect 223 445 257 479
rect 223 377 257 411
rect 223 309 257 343
rect 317 451 351 485
rect 317 383 351 417
rect 411 445 445 479
rect 411 377 445 411
rect 411 309 445 343
rect 505 451 539 485
rect 505 383 539 417
rect 599 445 633 479
rect 599 377 633 411
rect 599 309 633 343
rect 693 451 727 485
rect 693 383 727 417
rect 787 445 821 479
rect 787 377 821 411
rect 787 309 821 343
rect 881 451 915 485
rect 881 383 915 417
rect 975 445 1009 479
rect 975 377 1009 411
rect 975 309 1009 343
rect 1069 451 1103 485
rect 1069 383 1103 417
rect 1163 445 1197 479
rect 1163 377 1197 411
rect 1163 309 1197 343
rect 1257 451 1291 485
rect 1257 383 1291 417
rect 1351 445 1385 479
rect 1351 377 1385 411
rect 1351 309 1385 343
rect 1445 451 1479 485
rect 1445 383 1479 417
rect 1539 445 1573 479
rect 1539 377 1573 411
rect 1539 309 1573 343
rect 1633 451 1667 485
rect 1633 383 1667 417
rect 1727 445 1761 479
rect 1727 377 1761 411
rect 1727 309 1761 343
rect 1821 451 1855 485
rect 1821 383 1855 417
rect 1915 445 1949 479
rect 1915 377 1949 411
rect 1915 309 1949 343
rect 2009 451 2043 485
rect 2009 383 2043 417
rect 2103 445 2137 479
rect 2103 377 2137 411
rect 2103 309 2137 343
rect 2197 451 2231 485
rect 2197 383 2231 417
rect 2291 445 2325 479
rect 2291 377 2325 411
rect 2291 309 2325 343
rect 2385 451 2419 485
rect 2385 383 2419 417
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 457 497 493 523
rect 551 497 587 523
rect 645 497 681 523
rect 739 497 775 523
rect 833 497 869 523
rect 927 497 963 523
rect 1021 497 1057 523
rect 1115 497 1151 523
rect 1209 497 1245 523
rect 1303 497 1339 523
rect 1397 497 1433 523
rect 1491 497 1527 523
rect 1585 497 1621 523
rect 1679 497 1715 523
rect 1773 497 1809 523
rect 1867 497 1903 523
rect 1961 497 1997 523
rect 2055 497 2091 523
rect 2149 497 2185 523
rect 2243 497 2279 523
rect 2337 497 2373 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 457 282 493 297
rect 551 282 587 297
rect 645 282 681 297
rect 739 282 775 297
rect 833 282 869 297
rect 927 282 963 297
rect 1021 282 1057 297
rect 1115 282 1151 297
rect 1209 282 1245 297
rect 1303 282 1339 297
rect 1397 282 1433 297
rect 1491 282 1527 297
rect 1585 282 1621 297
rect 1679 282 1715 297
rect 1773 282 1809 297
rect 1867 282 1903 297
rect 1961 282 1997 297
rect 2055 282 2091 297
rect 2149 282 2185 297
rect 2243 282 2279 297
rect 2337 282 2373 297
rect 79 259 119 282
rect 173 259 213 282
rect 267 259 307 282
rect 79 249 307 259
rect 79 215 129 249
rect 163 215 197 249
rect 231 215 307 249
rect 79 205 307 215
rect 79 177 109 205
rect 173 177 203 205
rect 277 177 307 205
rect 361 259 401 282
rect 455 259 495 282
rect 549 259 589 282
rect 643 259 683 282
rect 737 259 777 282
rect 831 259 871 282
rect 361 249 871 259
rect 361 215 385 249
rect 419 215 463 249
rect 497 215 541 249
rect 575 215 619 249
rect 653 215 697 249
rect 731 215 765 249
rect 799 215 871 249
rect 361 205 871 215
rect 361 177 391 205
rect 455 177 485 205
rect 549 177 579 205
rect 643 177 673 205
rect 737 177 767 205
rect 841 177 871 205
rect 925 259 965 282
rect 1019 259 1059 282
rect 1113 259 1153 282
rect 1207 259 1247 282
rect 1301 259 1341 282
rect 1395 259 1435 282
rect 1489 259 1529 282
rect 1583 259 1623 282
rect 1677 259 1717 282
rect 1771 259 1811 282
rect 1865 259 1905 282
rect 1959 259 1999 282
rect 2053 259 2093 282
rect 2147 259 2187 282
rect 2241 259 2281 282
rect 2335 259 2375 282
rect 925 249 2375 259
rect 925 215 945 249
rect 979 215 1023 249
rect 1057 215 1101 249
rect 1135 215 1179 249
rect 1213 215 1257 249
rect 1291 215 1325 249
rect 1359 215 1403 249
rect 1437 215 1481 249
rect 1515 215 1559 249
rect 1593 215 1637 249
rect 1671 215 1705 249
rect 1739 215 1783 249
rect 1817 215 1861 249
rect 1895 215 1939 249
rect 1973 215 2017 249
rect 2051 215 2095 249
rect 2129 215 2163 249
rect 2197 215 2241 249
rect 2275 215 2375 249
rect 925 205 2375 215
rect 925 177 955 205
rect 1019 177 1049 205
rect 1113 177 1143 205
rect 1207 177 1237 205
rect 1301 177 1331 205
rect 1395 177 1425 205
rect 1489 177 1519 205
rect 1583 177 1613 205
rect 1677 177 1707 205
rect 1771 177 1801 205
rect 1865 177 1895 205
rect 1959 177 1989 205
rect 2053 177 2083 205
rect 2147 177 2177 205
rect 2241 177 2271 205
rect 2345 177 2375 205
rect 79 21 109 47
rect 173 21 203 47
rect 277 21 307 47
rect 361 21 391 47
rect 455 21 485 47
rect 549 21 579 47
rect 643 21 673 47
rect 737 21 767 47
rect 841 21 871 47
rect 925 21 955 47
rect 1019 21 1049 47
rect 1113 21 1143 47
rect 1207 21 1237 47
rect 1301 21 1331 47
rect 1395 21 1425 47
rect 1489 21 1519 47
rect 1583 21 1613 47
rect 1677 21 1707 47
rect 1771 21 1801 47
rect 1865 21 1895 47
rect 1959 21 1989 47
rect 2053 21 2083 47
rect 2147 21 2177 47
rect 2241 21 2271 47
rect 2345 21 2375 47
<< polycont >>
rect 129 215 163 249
rect 197 215 231 249
rect 385 215 419 249
rect 463 215 497 249
rect 541 215 575 249
rect 619 215 653 249
rect 697 215 731 249
rect 765 215 799 249
rect 945 215 979 249
rect 1023 215 1057 249
rect 1101 215 1135 249
rect 1179 215 1213 249
rect 1257 215 1291 249
rect 1325 215 1359 249
rect 1403 215 1437 249
rect 1481 215 1515 249
rect 1559 215 1593 249
rect 1637 215 1671 249
rect 1705 215 1739 249
rect 1783 215 1817 249
rect 1861 215 1895 249
rect 1939 215 1973 249
rect 2017 215 2051 249
rect 2095 215 2129 249
rect 2163 215 2197 249
rect 2241 215 2275 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2484 561
rect 19 479 85 493
rect 19 445 35 479
rect 69 445 85 479
rect 19 411 85 445
rect 19 377 35 411
rect 69 377 85 411
rect 19 343 85 377
rect 129 485 163 527
rect 129 417 163 451
rect 129 357 163 383
rect 197 479 273 493
rect 197 445 223 479
rect 257 445 273 479
rect 197 411 273 445
rect 197 377 223 411
rect 257 377 273 411
rect 19 309 35 343
rect 69 323 85 343
rect 197 343 273 377
rect 317 485 351 527
rect 317 417 351 451
rect 317 357 351 383
rect 385 479 461 493
rect 385 445 411 479
rect 445 445 461 479
rect 385 411 461 445
rect 385 377 411 411
rect 445 377 461 411
rect 197 323 223 343
rect 69 309 223 323
rect 257 323 273 343
rect 385 343 461 377
rect 505 485 539 527
rect 505 417 539 451
rect 505 367 539 383
rect 573 479 649 493
rect 573 445 599 479
rect 633 445 649 479
rect 573 411 649 445
rect 573 377 599 411
rect 633 377 649 411
rect 257 309 351 323
rect 19 289 351 309
rect 385 309 411 343
rect 445 323 461 343
rect 573 343 649 377
rect 693 485 727 527
rect 693 417 727 451
rect 693 367 727 383
rect 761 479 837 493
rect 761 445 787 479
rect 821 445 837 479
rect 761 411 837 445
rect 761 377 787 411
rect 821 377 837 411
rect 573 323 599 343
rect 445 309 599 323
rect 633 323 649 343
rect 761 343 837 377
rect 881 485 915 527
rect 881 417 915 451
rect 881 367 915 383
rect 949 479 1025 493
rect 949 445 975 479
rect 1009 445 1025 479
rect 949 411 1025 445
rect 949 377 975 411
rect 1009 377 1025 411
rect 761 323 787 343
rect 633 309 787 323
rect 821 323 837 343
rect 949 343 1025 377
rect 1069 485 1103 527
rect 1069 417 1103 451
rect 1069 367 1103 383
rect 1137 479 1213 493
rect 1137 445 1163 479
rect 1197 445 1213 479
rect 1137 411 1213 445
rect 1137 377 1163 411
rect 1197 377 1213 411
rect 821 309 915 323
rect 385 289 915 309
rect 949 309 975 343
rect 1009 323 1025 343
rect 1137 343 1213 377
rect 1257 485 1291 527
rect 1257 417 1291 451
rect 1257 367 1291 383
rect 1325 479 1401 493
rect 1325 445 1351 479
rect 1385 445 1401 479
rect 1325 411 1401 445
rect 1325 377 1351 411
rect 1385 377 1401 411
rect 1137 323 1163 343
rect 1009 309 1163 323
rect 1197 323 1213 343
rect 1325 343 1401 377
rect 1445 485 1479 527
rect 1445 417 1479 451
rect 1445 367 1479 383
rect 1513 479 1589 493
rect 1513 445 1539 479
rect 1573 445 1589 479
rect 1513 411 1589 445
rect 1513 377 1539 411
rect 1573 377 1589 411
rect 1325 323 1351 343
rect 1197 309 1351 323
rect 1385 323 1401 343
rect 1513 343 1589 377
rect 1633 485 1667 527
rect 1633 417 1667 451
rect 1633 367 1667 383
rect 1701 479 1777 493
rect 1701 445 1727 479
rect 1761 445 1777 479
rect 1701 411 1777 445
rect 1701 377 1727 411
rect 1761 377 1777 411
rect 1513 323 1539 343
rect 1385 309 1539 323
rect 1573 323 1589 343
rect 1701 343 1777 377
rect 1821 485 1855 527
rect 1821 417 1855 451
rect 1821 367 1855 383
rect 1889 479 1965 493
rect 1889 445 1915 479
rect 1949 445 1965 479
rect 1889 411 1965 445
rect 1889 377 1915 411
rect 1949 377 1965 411
rect 1701 323 1727 343
rect 1573 309 1727 323
rect 1761 323 1777 343
rect 1889 343 1965 377
rect 2009 485 2043 527
rect 2009 417 2043 451
rect 2009 367 2043 383
rect 2077 479 2153 493
rect 2077 445 2103 479
rect 2137 445 2153 479
rect 2077 411 2153 445
rect 2077 377 2103 411
rect 2137 377 2153 411
rect 1889 323 1915 343
rect 1761 309 1915 323
rect 1949 323 1965 343
rect 2077 343 2153 377
rect 2197 485 2231 527
rect 2197 417 2231 451
rect 2197 367 2231 383
rect 2265 479 2341 493
rect 2265 445 2291 479
rect 2325 445 2341 479
rect 2265 411 2341 445
rect 2265 377 2291 411
rect 2325 377 2341 411
rect 2077 323 2103 343
rect 1949 309 2103 323
rect 2137 323 2153 343
rect 2265 343 2341 377
rect 2385 485 2419 527
rect 2385 417 2419 451
rect 2385 367 2419 383
rect 2265 323 2291 343
rect 2137 309 2291 323
rect 2325 323 2341 343
rect 2325 309 2441 323
rect 949 289 2441 309
rect 317 255 351 289
rect 880 255 915 289
rect 18 249 273 255
rect 18 215 129 249
rect 163 215 197 249
rect 231 215 273 249
rect 317 249 829 255
rect 317 215 385 249
rect 419 215 463 249
rect 497 215 541 249
rect 575 215 619 249
rect 653 215 697 249
rect 731 215 765 249
rect 799 215 829 249
rect 880 249 2342 255
rect 880 215 945 249
rect 979 215 1023 249
rect 1057 215 1101 249
rect 1135 215 1179 249
rect 1213 215 1257 249
rect 1291 215 1325 249
rect 1359 215 1403 249
rect 1437 215 1481 249
rect 1515 215 1559 249
rect 1593 215 1637 249
rect 1671 215 1705 249
rect 1739 215 1783 249
rect 1817 215 1861 249
rect 1895 215 1939 249
rect 1973 215 2017 249
rect 2051 215 2095 249
rect 2129 215 2163 249
rect 2197 215 2241 249
rect 2275 215 2342 249
rect 317 181 351 215
rect 880 181 915 215
rect 2386 181 2441 289
rect 19 165 351 181
rect 19 131 35 165
rect 69 147 223 165
rect 69 131 85 147
rect 19 97 85 131
rect 197 131 223 147
rect 257 147 351 165
rect 385 165 915 181
rect 257 131 273 147
rect 19 63 35 97
rect 69 63 85 97
rect 19 52 85 63
rect 129 97 163 113
rect 129 17 163 63
rect 197 97 273 131
rect 385 131 411 165
rect 445 147 599 165
rect 445 131 461 147
rect 197 63 223 97
rect 257 63 273 97
rect 197 52 273 63
rect 317 97 351 113
rect 317 17 351 63
rect 385 97 461 131
rect 573 131 599 147
rect 633 147 787 165
rect 633 131 649 147
rect 385 63 411 97
rect 445 63 461 97
rect 385 52 461 63
rect 505 97 539 113
rect 505 17 539 63
rect 573 97 649 131
rect 761 131 787 147
rect 821 147 915 165
rect 949 165 2441 181
rect 821 131 837 147
rect 573 63 599 97
rect 633 63 649 97
rect 573 52 649 63
rect 693 97 727 113
rect 693 17 727 63
rect 761 97 837 131
rect 949 131 975 165
rect 1009 147 1163 165
rect 1009 131 1025 147
rect 761 63 787 97
rect 821 63 837 97
rect 761 52 837 63
rect 881 97 915 113
rect 881 17 915 63
rect 949 97 1025 131
rect 1137 131 1163 147
rect 1197 147 1351 165
rect 1197 131 1213 147
rect 949 63 975 97
rect 1009 63 1025 97
rect 949 52 1025 63
rect 1069 97 1103 113
rect 949 51 1009 52
rect 1069 17 1103 63
rect 1137 97 1213 131
rect 1325 131 1351 147
rect 1385 147 1539 165
rect 1385 131 1401 147
rect 1137 63 1163 97
rect 1197 63 1213 97
rect 1137 52 1213 63
rect 1257 97 1291 113
rect 1163 51 1197 52
rect 1257 17 1291 63
rect 1325 97 1401 131
rect 1513 131 1539 147
rect 1573 147 1727 165
rect 1573 131 1589 147
rect 1325 63 1351 97
rect 1385 63 1401 97
rect 1325 52 1401 63
rect 1445 97 1479 113
rect 1351 51 1385 52
rect 1445 17 1479 63
rect 1513 97 1589 131
rect 1701 131 1727 147
rect 1761 147 1915 165
rect 1761 131 1777 147
rect 1513 63 1539 97
rect 1573 63 1589 97
rect 1513 52 1589 63
rect 1633 97 1667 113
rect 1633 17 1667 63
rect 1701 97 1777 131
rect 1889 131 1915 147
rect 1949 147 2103 165
rect 1949 131 1965 147
rect 1701 63 1727 97
rect 1761 63 1777 97
rect 1701 52 1777 63
rect 1821 97 1855 113
rect 1821 17 1855 63
rect 1889 97 1965 131
rect 2077 131 2103 147
rect 2137 147 2291 165
rect 2137 131 2153 147
rect 1889 63 1915 97
rect 1949 63 1965 97
rect 1889 52 1965 63
rect 2009 97 2043 113
rect 2009 17 2043 63
rect 2077 97 2153 131
rect 2265 131 2291 147
rect 2325 147 2441 165
rect 2325 131 2341 147
rect 2077 63 2103 97
rect 2137 63 2153 97
rect 2077 52 2153 63
rect 2197 97 2231 113
rect 2197 17 2231 63
rect 2265 97 2341 131
rect 2265 63 2291 97
rect 2325 63 2341 97
rect 2265 52 2341 63
rect 2385 97 2419 113
rect 2385 17 2419 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2484 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
<< metal1 >>
rect 0 561 2484 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2484 561
rect 0 496 2484 527
rect 0 17 2484 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2484 17
rect 0 -48 2484 -17
<< labels >>
flabel corelocali s 30 221 64 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 2403 238 2403 238 0 FreeSans 200 0 0 0 Y
port 6 nsew
flabel corelocali s 2403 306 2403 306 0 FreeSans 200 0 0 0 Y
port 6 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew
rlabel comment s 0 0 0 0 4 bufinv_16
<< properties >>
string FIXED_BBOX 0 0 2484 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1732416
string GDS_START 1714374
<< end >>
