magic
tech sky130A
magscale 1 2
timestamp 1599588238
<< locali >>
rect 95 196 161 398
rect 263 236 355 310
rect 2026 364 2087 594
rect 2035 70 2087 364
rect 2413 364 2485 596
rect 2451 226 2485 364
rect 2417 70 2485 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2592 683
rect 23 472 73 596
rect 113 506 179 649
rect 315 506 381 649
rect 421 581 769 615
rect 421 480 455 581
rect 23 446 359 472
rect 489 459 573 547
rect 613 459 691 547
rect 489 446 523 459
rect 23 438 523 446
rect 23 162 57 438
rect 325 412 523 438
rect 195 378 291 404
rect 195 344 455 378
rect 195 202 229 344
rect 389 260 455 344
rect 23 70 73 162
rect 109 17 159 162
rect 195 70 287 202
rect 321 17 373 202
rect 409 85 443 226
rect 489 185 523 412
rect 557 287 623 421
rect 489 119 554 185
rect 588 85 622 287
rect 657 253 691 459
rect 725 513 769 581
rect 804 547 870 649
rect 904 581 1106 615
rect 904 513 938 581
rect 725 479 938 513
rect 725 287 769 479
rect 972 459 1038 547
rect 1072 472 1106 581
rect 1140 506 1214 649
rect 1356 530 1494 596
rect 1618 530 1652 649
rect 1356 496 1584 530
rect 1692 496 1758 583
rect 1926 526 1992 649
rect 972 445 1006 459
rect 828 411 1006 445
rect 1072 438 1300 472
rect 828 371 894 411
rect 950 337 1003 377
rect 803 303 1003 337
rect 1045 350 1127 404
rect 1045 316 1087 350
rect 1121 316 1127 350
rect 803 253 837 303
rect 950 282 1003 303
rect 1266 290 1300 438
rect 1356 370 1406 496
rect 1450 404 1516 462
rect 1550 424 1758 496
rect 1803 492 1869 524
rect 1803 458 1982 492
rect 1356 336 1443 370
rect 657 219 837 253
rect 657 185 706 219
rect 871 203 916 269
rect 950 248 1183 282
rect 1117 224 1183 248
rect 1266 224 1375 290
rect 656 93 706 185
rect 409 51 622 85
rect 798 17 848 169
rect 882 70 976 203
rect 1068 17 1232 136
rect 1266 90 1300 224
rect 1409 190 1443 336
rect 1334 124 1443 190
rect 1477 90 1511 404
rect 1550 390 1914 424
rect 1545 202 1611 356
rect 1657 350 1728 356
rect 1657 316 1663 350
rect 1697 316 1728 350
rect 1657 236 1728 316
rect 1780 270 1914 390
rect 1948 236 1982 458
rect 2121 364 2172 649
rect 1821 202 1982 236
rect 1545 168 1887 202
rect 1266 56 1511 90
rect 1620 17 1769 134
rect 1821 127 1887 168
rect 1933 17 1999 168
rect 2217 326 2283 572
rect 2323 364 2373 649
rect 2519 364 2569 649
rect 2217 260 2417 326
rect 2121 17 2171 226
rect 2217 70 2283 260
rect 2317 17 2383 206
rect 2519 17 2569 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2592 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 1087 316 1121 350
rect 1663 316 1697 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
<< metal1 >>
rect 0 683 2592 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2592 683
rect 0 617 2592 649
rect 1075 350 1133 356
rect 1075 316 1087 350
rect 1121 347 1133 350
rect 1651 350 1709 356
rect 1651 347 1663 350
rect 1121 319 1663 347
rect 1121 316 1133 319
rect 1075 310 1133 316
rect 1651 316 1663 319
rect 1697 316 1709 350
rect 1651 310 1709 316
rect 0 17 2592 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2592 17
rect 0 -49 2592 -17
<< labels >>
rlabel locali s 95 196 161 398 6 D
port 1 nsew signal input
rlabel locali s 2451 226 2485 364 6 Q
port 2 nsew signal output
rlabel locali s 2417 70 2485 226 6 Q
port 2 nsew signal output
rlabel locali s 2413 364 2485 596 6 Q
port 2 nsew signal output
rlabel locali s 2035 70 2087 364 6 Q_N
port 3 nsew signal output
rlabel locali s 2026 364 2087 594 6 Q_N
port 3 nsew signal output
rlabel metal1 s 1651 347 1709 356 6 SET_B
port 4 nsew signal input
rlabel metal1 s 1651 310 1709 319 6 SET_B
port 4 nsew signal input
rlabel metal1 s 1075 347 1133 356 6 SET_B
port 4 nsew signal input
rlabel metal1 s 1075 319 1709 347 6 SET_B
port 4 nsew signal input
rlabel metal1 s 1075 310 1133 319 6 SET_B
port 4 nsew signal input
rlabel locali s 263 236 355 310 6 CLK
port 5 nsew clock input
rlabel metal1 s 0 -49 2592 49 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 617 2592 715 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2592 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2769308
string GDS_START 2749916
<< end >>
