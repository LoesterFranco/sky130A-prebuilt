magic
tech sky130A
magscale 1 2
timestamp 1599588218
<< nwell >>
rect -38 332 1286 704
<< pwell >>
rect 0 0 1248 49
<< scpmos >>
rect 88 368 124 592
rect 178 368 214 592
rect 278 368 314 592
rect 368 368 404 592
rect 468 368 504 592
rect 558 368 594 592
rect 658 368 694 592
rect 748 368 784 592
rect 848 368 884 592
rect 938 368 974 592
rect 1038 368 1074 592
rect 1128 368 1164 592
<< nmoslvt >>
rect 88 80 118 164
rect 520 80 550 164
rect 634 80 664 164
rect 720 80 750 164
rect 834 80 864 164
rect 920 80 950 164
rect 1034 80 1064 164
rect 1134 80 1164 164
<< ndiff >>
rect 27 139 88 164
rect 27 105 39 139
rect 73 105 88 139
rect 27 80 88 105
rect 118 142 520 164
rect 118 108 139 142
rect 173 108 223 142
rect 257 108 307 142
rect 341 108 391 142
rect 425 108 475 142
rect 509 108 520 142
rect 118 80 520 108
rect 550 139 634 164
rect 550 105 575 139
rect 609 105 634 139
rect 550 80 634 105
rect 664 139 720 164
rect 664 105 675 139
rect 709 105 720 139
rect 664 80 720 105
rect 750 139 834 164
rect 750 105 775 139
rect 809 105 834 139
rect 750 80 834 105
rect 864 139 920 164
rect 864 105 875 139
rect 909 105 920 139
rect 864 80 920 105
rect 950 139 1034 164
rect 950 105 975 139
rect 1009 105 1034 139
rect 950 80 1034 105
rect 1064 139 1134 164
rect 1064 105 1075 139
rect 1109 105 1134 139
rect 1064 80 1134 105
rect 1164 139 1221 164
rect 1164 105 1175 139
rect 1209 105 1221 139
rect 1164 80 1221 105
<< pdiff >>
rect 27 580 88 592
rect 27 546 41 580
rect 75 546 88 580
rect 27 508 88 546
rect 27 474 41 508
rect 75 474 88 508
rect 27 368 88 474
rect 124 580 178 592
rect 124 546 134 580
rect 168 546 178 580
rect 124 505 178 546
rect 124 471 134 505
rect 168 471 178 505
rect 124 424 178 471
rect 124 390 134 424
rect 168 390 178 424
rect 124 368 178 390
rect 214 580 278 592
rect 214 546 224 580
rect 258 546 278 580
rect 214 508 278 546
rect 214 474 224 508
rect 258 474 278 508
rect 214 368 278 474
rect 314 580 368 592
rect 314 546 324 580
rect 358 546 368 580
rect 314 505 368 546
rect 314 471 324 505
rect 358 471 368 505
rect 314 424 368 471
rect 314 390 324 424
rect 358 390 368 424
rect 314 368 368 390
rect 404 580 468 592
rect 404 546 414 580
rect 448 546 468 580
rect 404 508 468 546
rect 404 474 414 508
rect 448 474 468 508
rect 404 368 468 474
rect 504 580 558 592
rect 504 546 514 580
rect 548 546 558 580
rect 504 505 558 546
rect 504 471 514 505
rect 548 471 558 505
rect 504 424 558 471
rect 504 390 514 424
rect 548 390 558 424
rect 504 368 558 390
rect 594 580 658 592
rect 594 546 604 580
rect 638 546 658 580
rect 594 508 658 546
rect 594 474 604 508
rect 638 474 658 508
rect 594 368 658 474
rect 694 580 748 592
rect 694 546 704 580
rect 738 546 748 580
rect 694 505 748 546
rect 694 471 704 505
rect 738 471 748 505
rect 694 424 748 471
rect 694 390 704 424
rect 738 390 748 424
rect 694 368 748 390
rect 784 580 848 592
rect 784 546 794 580
rect 828 546 848 580
rect 784 508 848 546
rect 784 474 794 508
rect 828 474 848 508
rect 784 368 848 474
rect 884 580 938 592
rect 884 546 894 580
rect 928 546 938 580
rect 884 505 938 546
rect 884 471 894 505
rect 928 471 938 505
rect 884 424 938 471
rect 884 390 894 424
rect 928 390 938 424
rect 884 368 938 390
rect 974 580 1038 592
rect 974 546 984 580
rect 1018 546 1038 580
rect 974 508 1038 546
rect 974 474 984 508
rect 1018 474 1038 508
rect 974 368 1038 474
rect 1074 580 1128 592
rect 1074 546 1084 580
rect 1118 546 1128 580
rect 1074 505 1128 546
rect 1074 471 1084 505
rect 1118 471 1128 505
rect 1074 424 1128 471
rect 1074 390 1084 424
rect 1118 390 1128 424
rect 1074 368 1128 390
rect 1164 580 1220 592
rect 1164 546 1174 580
rect 1208 546 1220 580
rect 1164 508 1220 546
rect 1164 474 1174 508
rect 1208 474 1220 508
rect 1164 368 1220 474
<< ndiffc >>
rect 39 105 73 139
rect 139 108 173 142
rect 223 108 257 142
rect 307 108 341 142
rect 391 108 425 142
rect 475 108 509 142
rect 575 105 609 139
rect 675 105 709 139
rect 775 105 809 139
rect 875 105 909 139
rect 975 105 1009 139
rect 1075 105 1109 139
rect 1175 105 1209 139
<< pdiffc >>
rect 41 546 75 580
rect 41 474 75 508
rect 134 546 168 580
rect 134 471 168 505
rect 134 390 168 424
rect 224 546 258 580
rect 224 474 258 508
rect 324 546 358 580
rect 324 471 358 505
rect 324 390 358 424
rect 414 546 448 580
rect 414 474 448 508
rect 514 546 548 580
rect 514 471 548 505
rect 514 390 548 424
rect 604 546 638 580
rect 604 474 638 508
rect 704 546 738 580
rect 704 471 738 505
rect 704 390 738 424
rect 794 546 828 580
rect 794 474 828 508
rect 894 546 928 580
rect 894 471 928 505
rect 894 390 928 424
rect 984 546 1018 580
rect 984 474 1018 508
rect 1084 546 1118 580
rect 1084 471 1118 505
rect 1084 390 1118 424
rect 1174 546 1208 580
rect 1174 474 1208 508
<< poly >>
rect 88 592 124 618
rect 178 592 214 618
rect 278 592 314 618
rect 368 592 404 618
rect 468 592 504 618
rect 558 592 594 618
rect 658 592 694 618
rect 748 592 784 618
rect 848 592 884 618
rect 938 592 974 618
rect 1038 592 1074 618
rect 1128 592 1164 618
rect 88 336 124 368
rect 178 336 214 368
rect 278 336 314 368
rect 368 336 404 368
rect 468 336 504 368
rect 558 336 594 368
rect 658 336 694 368
rect 748 336 784 368
rect 848 336 884 368
rect 938 336 974 368
rect 1038 336 1074 368
rect 1128 336 1164 368
rect 88 320 1164 336
rect 88 286 141 320
rect 175 286 209 320
rect 243 286 277 320
rect 311 286 345 320
rect 379 286 413 320
rect 447 286 481 320
rect 515 286 549 320
rect 583 286 617 320
rect 651 286 685 320
rect 719 286 753 320
rect 787 286 821 320
rect 855 286 889 320
rect 923 286 957 320
rect 991 286 1025 320
rect 1059 286 1093 320
rect 1127 286 1164 320
rect 88 270 1164 286
rect 88 164 118 270
rect 520 164 550 270
rect 634 164 664 270
rect 720 164 750 270
rect 834 164 864 270
rect 920 164 950 270
rect 1034 164 1064 270
rect 1134 164 1164 270
rect 88 54 118 80
rect 520 54 550 80
rect 634 54 664 80
rect 720 54 750 80
rect 834 54 864 80
rect 920 54 950 80
rect 1034 54 1064 80
rect 1134 54 1164 80
<< polycont >>
rect 141 286 175 320
rect 209 286 243 320
rect 277 286 311 320
rect 345 286 379 320
rect 413 286 447 320
rect 481 286 515 320
rect 549 286 583 320
rect 617 286 651 320
rect 685 286 719 320
rect 753 286 787 320
rect 821 286 855 320
rect 889 286 923 320
rect 957 286 991 320
rect 1025 286 1059 320
rect 1093 286 1127 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 23 580 78 649
rect 23 546 41 580
rect 75 546 78 580
rect 23 508 78 546
rect 23 474 41 508
rect 75 474 78 508
rect 23 458 78 474
rect 118 580 184 596
rect 118 546 134 580
rect 168 546 184 580
rect 118 505 184 546
rect 118 471 134 505
rect 168 471 184 505
rect 118 424 184 471
rect 224 580 274 649
rect 258 546 274 580
rect 224 508 274 546
rect 258 474 274 508
rect 224 458 274 474
rect 308 580 374 596
rect 308 546 324 580
rect 358 546 374 580
rect 308 505 374 546
rect 308 471 324 505
rect 358 471 374 505
rect 308 424 374 471
rect 414 580 464 649
rect 448 546 464 580
rect 414 508 464 546
rect 448 474 464 508
rect 414 458 464 474
rect 498 580 564 596
rect 498 546 514 580
rect 548 546 564 580
rect 498 505 564 546
rect 498 471 514 505
rect 548 471 564 505
rect 498 424 564 471
rect 604 580 654 649
rect 638 546 654 580
rect 604 508 654 546
rect 638 474 654 508
rect 604 458 654 474
rect 688 580 754 596
rect 688 546 704 580
rect 738 546 754 580
rect 688 505 754 546
rect 688 471 704 505
rect 738 471 754 505
rect 688 424 754 471
rect 794 580 844 649
rect 828 546 844 580
rect 794 508 844 546
rect 828 474 844 508
rect 794 458 844 474
rect 878 580 944 596
rect 878 546 894 580
rect 928 546 944 580
rect 878 505 944 546
rect 878 471 894 505
rect 928 471 944 505
rect 878 424 944 471
rect 984 580 1034 649
rect 1018 546 1034 580
rect 984 508 1034 546
rect 1018 474 1034 508
rect 984 458 1034 474
rect 1068 580 1134 596
rect 1068 546 1084 580
rect 1118 546 1134 580
rect 1068 505 1134 546
rect 1068 471 1084 505
rect 1118 471 1134 505
rect 1068 424 1134 471
rect 1174 580 1224 649
rect 1208 546 1224 580
rect 1174 508 1224 546
rect 1208 474 1224 508
rect 1174 458 1224 474
rect 57 390 134 424
rect 168 390 324 424
rect 358 390 514 424
rect 548 390 704 424
rect 738 390 894 424
rect 928 390 1084 424
rect 1118 390 1223 424
rect 57 236 91 390
rect 125 320 1143 356
rect 125 286 141 320
rect 175 286 209 320
rect 243 286 277 320
rect 311 286 345 320
rect 379 286 413 320
rect 447 286 481 320
rect 515 286 549 320
rect 583 286 617 320
rect 651 286 685 320
rect 719 286 753 320
rect 787 286 821 320
rect 855 286 889 320
rect 923 286 957 320
rect 991 286 1025 320
rect 1059 286 1093 320
rect 1127 286 1143 320
rect 125 270 1143 286
rect 1177 236 1223 390
rect 57 202 1223 236
rect 23 139 89 155
rect 23 105 39 139
rect 73 105 89 139
rect 23 17 89 105
rect 123 142 525 202
rect 123 108 139 142
rect 173 108 223 142
rect 257 108 307 142
rect 341 108 391 142
rect 425 108 475 142
rect 509 108 525 142
rect 123 92 525 108
rect 559 139 625 155
rect 559 105 575 139
rect 609 105 625 139
rect 559 17 625 105
rect 659 139 725 202
rect 659 105 675 139
rect 709 105 725 139
rect 659 89 725 105
rect 759 139 825 155
rect 759 105 775 139
rect 809 105 825 139
rect 759 17 825 105
rect 859 139 925 202
rect 859 105 875 139
rect 909 105 925 139
rect 859 89 925 105
rect 959 139 1025 155
rect 959 105 975 139
rect 1009 105 1025 139
rect 959 17 1025 105
rect 1059 139 1125 202
rect 1059 105 1075 139
rect 1109 105 1125 139
rect 1059 89 1125 105
rect 1159 139 1225 155
rect 1159 105 1175 139
rect 1209 105 1225 139
rect 1159 17 1225 105
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
<< metal1 >>
rect 0 683 1248 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 0 617 1248 649
rect 0 17 1248 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
rect 0 -49 1248 -17
<< labels >>
flabel pwell s 0 0 1248 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew
flabel nwell s 0 617 1248 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew
rlabel comment s 0 0 0 0 4 clkinv_8
flabel metal1 s 0 617 1248 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew
flabel metal1 s 0 0 1248 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 1183 242 1217 276 0 FreeSans 340 0 0 0 Y
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 1248 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 2722074
string GDS_START 2712588
<< end >>
