magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 167 384 263 578
rect 25 270 119 356
rect 167 270 233 384
rect 313 336 359 578
rect 281 270 359 336
rect 395 270 461 356
rect 505 270 647 356
rect 790 282 831 596
rect 790 236 839 282
rect 790 226 837 236
rect 771 70 837 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 23 390 89 649
rect 425 424 491 596
rect 539 458 756 649
rect 425 390 747 424
rect 681 260 747 390
rect 871 364 937 649
rect 681 236 715 260
rect 23 202 525 236
rect 23 70 89 202
rect 123 17 189 168
rect 223 70 289 202
rect 323 17 425 163
rect 459 70 525 202
rect 559 202 715 236
rect 559 70 625 202
rect 671 17 737 164
rect 871 17 923 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
rlabel locali s 25 270 119 356 6 A1
port 1 nsew signal input
rlabel locali s 167 384 263 578 6 A2
port 2 nsew signal input
rlabel locali s 167 270 233 384 6 A2
port 2 nsew signal input
rlabel locali s 313 336 359 578 6 A3
port 3 nsew signal input
rlabel locali s 281 270 359 336 6 A3
port 3 nsew signal input
rlabel locali s 395 270 461 356 6 A4
port 4 nsew signal input
rlabel locali s 505 270 647 356 6 B1
port 5 nsew signal input
rlabel locali s 790 282 831 596 6 X
port 6 nsew signal output
rlabel locali s 790 236 839 282 6 X
port 6 nsew signal output
rlabel locali s 790 226 837 236 6 X
port 6 nsew signal output
rlabel locali s 771 70 837 226 6 X
port 6 nsew signal output
rlabel metal1 s 0 -49 960 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 617 960 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 725914
string GDS_START 717190
<< end >>
