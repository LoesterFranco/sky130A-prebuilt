magic
tech sky130A
magscale 1 2
timestamp 1599588209
<< nwell >>
rect -38 332 1382 704
<< pwell >>
rect 0 0 1344 49
<< scpmos >>
rect 96 368 126 592
rect 186 368 216 592
rect 296 368 326 592
rect 386 368 416 592
rect 528 391 558 559
rect 618 391 648 559
rect 731 391 761 559
rect 821 391 851 559
rect 938 391 968 591
rect 1028 391 1058 591
rect 1128 391 1158 591
rect 1218 391 1248 591
<< nmoslvt >>
rect 91 74 121 222
rect 177 74 207 222
rect 277 74 307 222
rect 363 74 393 222
rect 567 125 597 253
rect 653 125 683 253
rect 739 125 769 253
rect 839 125 869 253
rect 941 125 971 253
rect 1033 125 1063 253
rect 1130 125 1160 253
rect 1230 125 1260 253
<< ndiff >>
rect 34 131 91 222
rect 34 97 46 131
rect 80 97 91 131
rect 34 74 91 97
rect 121 210 177 222
rect 121 176 132 210
rect 166 176 177 210
rect 121 120 177 176
rect 121 86 132 120
rect 166 86 177 120
rect 121 74 177 86
rect 207 131 277 222
rect 207 97 218 131
rect 252 97 277 131
rect 207 74 277 97
rect 307 210 363 222
rect 307 176 318 210
rect 352 176 363 210
rect 307 120 363 176
rect 307 86 318 120
rect 352 86 363 120
rect 307 74 363 86
rect 393 210 450 222
rect 393 176 404 210
rect 438 176 450 210
rect 393 120 450 176
rect 393 86 404 120
rect 438 86 450 120
rect 393 74 450 86
rect 517 249 567 253
rect 510 237 567 249
rect 510 203 522 237
rect 556 203 567 237
rect 510 169 567 203
rect 510 135 522 169
rect 556 135 567 169
rect 510 125 567 135
rect 597 241 653 253
rect 597 207 608 241
rect 642 207 653 241
rect 597 171 653 207
rect 597 137 608 171
rect 642 137 653 171
rect 597 125 653 137
rect 683 238 739 253
rect 683 204 694 238
rect 728 204 739 238
rect 683 125 739 204
rect 769 171 839 253
rect 769 137 794 171
rect 828 137 839 171
rect 769 125 839 137
rect 869 241 941 253
rect 869 207 880 241
rect 914 207 941 241
rect 869 171 941 207
rect 869 137 880 171
rect 914 137 941 171
rect 869 125 941 137
rect 971 171 1033 253
rect 971 137 983 171
rect 1017 137 1033 171
rect 971 125 1033 137
rect 1063 240 1130 253
rect 1063 206 1085 240
rect 1119 206 1130 240
rect 1063 171 1130 206
rect 1063 137 1085 171
rect 1119 137 1130 171
rect 1063 125 1130 137
rect 1160 171 1230 253
rect 1160 137 1171 171
rect 1205 137 1230 171
rect 1160 125 1230 137
rect 1260 240 1317 253
rect 1260 206 1271 240
rect 1305 206 1317 240
rect 1260 171 1317 206
rect 1260 137 1271 171
rect 1305 137 1317 171
rect 1260 125 1317 137
<< pdiff >>
rect 27 580 96 592
rect 27 546 39 580
rect 73 546 96 580
rect 27 478 96 546
rect 27 444 39 478
rect 73 444 96 478
rect 27 368 96 444
rect 126 580 186 592
rect 126 546 139 580
rect 173 546 186 580
rect 126 497 186 546
rect 126 463 139 497
rect 173 463 186 497
rect 126 414 186 463
rect 126 380 139 414
rect 173 380 186 414
rect 126 368 186 380
rect 216 580 296 592
rect 216 546 239 580
rect 273 546 296 580
rect 216 478 296 546
rect 216 444 239 478
rect 273 444 296 478
rect 216 368 296 444
rect 326 580 386 592
rect 326 546 339 580
rect 373 546 386 580
rect 326 497 386 546
rect 326 463 339 497
rect 373 463 386 497
rect 326 414 386 463
rect 326 380 339 414
rect 373 380 386 414
rect 326 368 386 380
rect 416 580 485 592
rect 416 546 439 580
rect 473 559 485 580
rect 869 579 938 591
rect 869 559 881 579
rect 473 546 528 559
rect 416 498 528 546
rect 416 464 439 498
rect 473 464 528 498
rect 416 391 528 464
rect 558 547 618 559
rect 558 513 571 547
rect 605 513 618 547
rect 558 440 618 513
rect 558 406 571 440
rect 605 406 618 440
rect 558 391 618 406
rect 648 508 731 559
rect 648 474 671 508
rect 705 474 731 508
rect 648 391 731 474
rect 761 547 821 559
rect 761 513 774 547
rect 808 513 821 547
rect 761 440 821 513
rect 761 406 774 440
rect 808 406 821 440
rect 761 391 821 406
rect 851 545 881 559
rect 915 545 938 579
rect 851 499 938 545
rect 851 465 881 499
rect 915 465 938 499
rect 851 391 938 465
rect 968 579 1028 591
rect 968 545 981 579
rect 1015 545 1028 579
rect 968 499 1028 545
rect 968 465 981 499
rect 1015 465 1028 499
rect 968 391 1028 465
rect 1058 531 1128 591
rect 1058 497 1081 531
rect 1115 497 1128 531
rect 1058 440 1128 497
rect 1058 406 1081 440
rect 1115 406 1128 440
rect 1058 391 1128 406
rect 1158 579 1218 591
rect 1158 545 1171 579
rect 1205 545 1218 579
rect 1158 509 1218 545
rect 1158 475 1171 509
rect 1205 475 1218 509
rect 1158 440 1218 475
rect 1158 406 1171 440
rect 1205 406 1218 440
rect 1158 391 1218 406
rect 1248 579 1317 591
rect 1248 545 1271 579
rect 1305 545 1317 579
rect 1248 509 1317 545
rect 1248 475 1271 509
rect 1305 475 1317 509
rect 1248 440 1317 475
rect 1248 406 1271 440
rect 1305 406 1317 440
rect 1248 391 1317 406
rect 416 368 469 391
<< ndiffc >>
rect 46 97 80 131
rect 132 176 166 210
rect 132 86 166 120
rect 218 97 252 131
rect 318 176 352 210
rect 318 86 352 120
rect 404 176 438 210
rect 404 86 438 120
rect 522 203 556 237
rect 522 135 556 169
rect 608 207 642 241
rect 608 137 642 171
rect 694 204 728 238
rect 794 137 828 171
rect 880 207 914 241
rect 880 137 914 171
rect 983 137 1017 171
rect 1085 206 1119 240
rect 1085 137 1119 171
rect 1171 137 1205 171
rect 1271 206 1305 240
rect 1271 137 1305 171
<< pdiffc >>
rect 39 546 73 580
rect 39 444 73 478
rect 139 546 173 580
rect 139 463 173 497
rect 139 380 173 414
rect 239 546 273 580
rect 239 444 273 478
rect 339 546 373 580
rect 339 463 373 497
rect 339 380 373 414
rect 439 546 473 580
rect 439 464 473 498
rect 571 513 605 547
rect 571 406 605 440
rect 671 474 705 508
rect 774 513 808 547
rect 774 406 808 440
rect 881 545 915 579
rect 881 465 915 499
rect 981 545 1015 579
rect 981 465 1015 499
rect 1081 497 1115 531
rect 1081 406 1115 440
rect 1171 545 1205 579
rect 1171 475 1205 509
rect 1171 406 1205 440
rect 1271 545 1305 579
rect 1271 475 1305 509
rect 1271 406 1305 440
<< poly >>
rect 96 592 126 618
rect 186 592 216 618
rect 296 592 326 618
rect 386 592 416 618
rect 938 591 968 617
rect 1028 591 1058 617
rect 1128 591 1158 617
rect 1218 591 1248 617
rect 528 559 558 585
rect 618 559 648 585
rect 731 559 761 585
rect 821 559 851 585
rect 528 376 558 391
rect 618 376 648 391
rect 731 376 761 391
rect 821 376 851 391
rect 938 376 968 391
rect 1028 376 1058 391
rect 1128 376 1158 391
rect 1218 376 1248 391
rect 96 353 126 368
rect 186 353 216 368
rect 296 353 326 368
rect 386 353 416 368
rect 525 353 561 376
rect 93 326 129 353
rect 183 326 219 353
rect 293 326 329 353
rect 383 326 419 353
rect 93 310 419 326
rect 93 290 139 310
rect 91 276 139 290
rect 173 276 207 310
rect 241 276 275 310
rect 309 276 343 310
rect 377 276 419 310
rect 91 260 419 276
rect 465 337 567 353
rect 615 346 769 376
rect 465 303 517 337
rect 551 303 567 337
rect 465 298 567 303
rect 653 340 769 346
rect 653 306 706 340
rect 740 306 769 340
rect 465 268 597 298
rect 91 222 121 260
rect 177 222 207 260
rect 277 222 307 260
rect 363 222 393 260
rect 91 48 121 74
rect 177 48 207 74
rect 277 48 307 74
rect 363 48 393 74
rect 465 51 495 268
rect 567 253 597 268
rect 653 290 769 306
rect 653 253 683 290
rect 739 253 769 290
rect 818 298 854 376
rect 818 268 869 298
rect 935 268 971 376
rect 1025 356 1061 376
rect 1125 356 1161 376
rect 1215 356 1251 376
rect 1025 340 1167 356
rect 1025 326 1049 340
rect 839 253 869 268
rect 941 253 971 268
rect 1033 306 1049 326
rect 1083 306 1117 340
rect 1151 306 1167 340
rect 1033 290 1167 306
rect 1215 340 1281 356
rect 1215 306 1231 340
rect 1265 306 1281 340
rect 1215 290 1281 306
rect 1033 253 1063 290
rect 1130 253 1160 290
rect 1230 253 1260 290
rect 567 99 597 125
rect 653 99 683 125
rect 739 99 769 125
rect 839 51 869 125
rect 465 21 869 51
rect 941 51 971 125
rect 1033 99 1063 125
rect 1130 99 1160 125
rect 1230 51 1260 125
rect 941 21 1260 51
<< polycont >>
rect 139 276 173 310
rect 207 276 241 310
rect 275 276 309 310
rect 343 276 377 310
rect 517 303 551 337
rect 706 306 740 340
rect 1049 306 1083 340
rect 1117 306 1151 340
rect 1231 306 1265 340
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 23 580 89 649
rect 23 546 39 580
rect 73 546 89 580
rect 23 478 89 546
rect 23 444 39 478
rect 73 444 89 478
rect 23 428 89 444
rect 123 580 189 596
rect 123 546 139 580
rect 173 546 189 580
rect 123 497 189 546
rect 123 463 139 497
rect 173 463 189 497
rect 123 414 189 463
rect 223 580 289 649
rect 223 546 239 580
rect 273 546 289 580
rect 223 478 289 546
rect 223 444 239 478
rect 273 444 289 478
rect 223 428 289 444
rect 323 580 389 596
rect 323 546 339 580
rect 373 546 389 580
rect 323 497 389 546
rect 323 463 339 497
rect 373 463 389 497
rect 123 394 139 414
rect 25 380 139 394
rect 173 394 189 414
rect 323 414 389 463
rect 423 580 489 649
rect 423 546 439 580
rect 473 546 489 580
rect 423 498 489 546
rect 423 464 439 498
rect 473 464 489 498
rect 423 458 489 464
rect 555 547 621 563
rect 555 513 571 547
rect 605 513 621 547
rect 555 440 621 513
rect 655 508 721 649
rect 865 579 931 649
rect 655 474 671 508
rect 705 474 721 508
rect 655 458 721 474
rect 758 547 824 563
rect 758 513 774 547
rect 808 513 824 547
rect 555 424 571 440
rect 323 394 339 414
rect 173 380 339 394
rect 373 380 389 414
rect 25 360 389 380
rect 423 406 571 424
rect 605 424 621 440
rect 758 440 824 513
rect 865 545 881 579
rect 915 545 931 579
rect 865 499 931 545
rect 865 465 881 499
rect 915 465 931 499
rect 865 458 931 465
rect 965 581 1221 615
rect 965 579 1031 581
rect 965 545 981 579
rect 1015 545 1031 579
rect 1171 579 1221 581
rect 965 499 1031 545
rect 965 465 981 499
rect 1015 465 1031 499
rect 965 458 1031 465
rect 1065 531 1131 547
rect 1065 497 1081 531
rect 1115 497 1131 531
rect 758 424 774 440
rect 605 406 774 424
rect 808 424 824 440
rect 1065 440 1131 497
rect 1065 424 1081 440
rect 808 406 1081 424
rect 1115 406 1131 440
rect 423 390 1131 406
rect 1205 545 1221 579
rect 1171 509 1221 545
rect 1205 475 1221 509
rect 1171 440 1221 475
rect 1205 406 1221 440
rect 1171 390 1221 406
rect 1255 579 1321 649
rect 1255 545 1271 579
rect 1305 545 1321 579
rect 1255 509 1321 545
rect 1255 475 1271 509
rect 1305 475 1321 509
rect 1255 440 1321 475
rect 1255 406 1271 440
rect 1305 406 1321 440
rect 1255 390 1321 406
rect 25 226 71 360
rect 423 326 457 390
rect 123 310 457 326
rect 123 276 139 310
rect 173 276 207 310
rect 241 276 275 310
rect 309 276 343 310
rect 377 276 457 310
rect 501 337 567 356
rect 501 303 517 337
rect 551 303 567 337
rect 501 287 567 303
rect 690 340 756 356
rect 690 306 706 340
rect 740 306 756 340
rect 690 290 756 306
rect 123 260 457 276
rect 506 237 556 253
rect 25 210 352 226
rect 25 192 132 210
rect 116 176 132 192
rect 166 192 318 210
rect 30 131 80 158
rect 30 97 46 131
rect 30 17 80 97
rect 116 120 166 176
rect 302 176 318 192
rect 116 86 132 120
rect 116 70 166 86
rect 202 131 268 158
rect 202 97 218 131
rect 252 97 268 131
rect 202 17 268 97
rect 302 120 352 176
rect 302 86 318 120
rect 302 70 352 86
rect 388 210 454 226
rect 388 176 404 210
rect 438 176 454 210
rect 388 120 454 176
rect 388 86 404 120
rect 438 86 454 120
rect 388 17 454 86
rect 506 203 522 237
rect 506 169 556 203
rect 506 135 522 169
rect 506 85 556 135
rect 608 241 642 257
rect 790 256 824 390
rect 985 340 1167 356
rect 985 306 1049 340
rect 1083 306 1117 340
rect 1151 306 1167 340
rect 985 290 1167 306
rect 1215 340 1319 356
rect 1215 306 1231 340
rect 1265 306 1319 340
rect 1215 290 1319 306
rect 608 171 642 207
rect 678 238 824 256
rect 678 204 694 238
rect 728 222 824 238
rect 880 256 930 257
rect 880 241 1321 256
rect 728 204 744 222
rect 678 187 744 204
rect 914 240 1321 241
rect 914 222 1085 240
rect 914 207 930 222
rect 778 171 844 188
rect 778 153 794 171
rect 642 137 794 153
rect 828 137 844 171
rect 608 119 844 137
rect 880 171 930 207
rect 1069 206 1085 222
rect 1119 222 1271 240
rect 914 137 930 171
rect 880 85 930 137
rect 506 51 930 85
rect 966 171 1035 187
rect 966 137 983 171
rect 1017 137 1035 171
rect 966 17 1035 137
rect 1069 171 1119 206
rect 1255 206 1271 222
rect 1305 206 1321 240
rect 1069 137 1085 171
rect 1069 121 1119 137
rect 1155 171 1221 188
rect 1155 137 1171 171
rect 1205 137 1221 171
rect 1155 17 1221 137
rect 1255 171 1321 206
rect 1255 137 1271 171
rect 1305 137 1321 171
rect 1255 121 1321 137
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
<< metal1 >>
rect 0 683 1344 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 0 617 1344 649
rect 0 17 1344 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
rect 0 -49 1344 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o211a_4
flabel pwell s 0 0 1344 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nwell s 0 617 1344 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 1344 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 1344 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 1279 316 1313 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 1344 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1777828
string GDS_START 1766756
<< end >>
