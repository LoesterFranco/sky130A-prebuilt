magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 1382 704
<< pwell >>
rect 0 0 1344 49
<< scnmos >>
rect 98 74 128 222
rect 184 74 214 222
rect 284 74 314 222
rect 435 74 465 222
rect 559 74 589 222
rect 645 74 675 222
rect 929 74 959 222
rect 1029 74 1059 222
<< pmoshvt >>
rect 86 368 116 592
rect 176 368 206 592
rect 266 368 296 592
rect 356 368 386 592
rect 558 392 588 592
rect 648 392 678 592
rect 738 392 768 592
rect 832 392 862 592
rect 932 392 962 592
rect 1032 392 1062 592
rect 1122 392 1152 592
rect 1212 392 1242 592
<< ndiff >>
rect 27 210 98 222
rect 27 176 39 210
rect 73 176 98 210
rect 27 120 98 176
rect 27 86 39 120
rect 73 86 98 120
rect 27 74 98 86
rect 128 210 184 222
rect 128 176 139 210
rect 173 176 184 210
rect 128 120 184 176
rect 128 86 139 120
rect 173 86 184 120
rect 128 74 184 86
rect 214 133 284 222
rect 214 99 239 133
rect 273 99 284 133
rect 214 74 284 99
rect 314 210 435 222
rect 314 176 339 210
rect 373 176 435 210
rect 314 120 435 176
rect 314 86 339 120
rect 373 86 435 120
rect 314 74 435 86
rect 465 108 559 222
rect 465 74 495 108
rect 529 74 559 108
rect 589 192 645 222
rect 589 158 600 192
rect 634 158 645 192
rect 589 120 645 158
rect 589 86 600 120
rect 634 86 645 120
rect 589 74 645 86
rect 675 108 929 222
rect 675 74 702 108
rect 736 74 785 108
rect 819 74 868 108
rect 902 74 929 108
rect 959 210 1029 222
rect 959 176 970 210
rect 1004 176 1029 210
rect 959 120 1029 176
rect 959 86 970 120
rect 1004 86 1029 120
rect 959 74 1029 86
rect 1059 132 1109 222
rect 1059 120 1219 132
rect 1059 86 1070 120
rect 1104 86 1173 120
rect 1207 86 1219 120
rect 1059 74 1219 86
rect 480 62 544 74
rect 690 62 914 74
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 498 86 546
rect 27 464 39 498
rect 73 464 86 498
rect 27 368 86 464
rect 116 580 176 592
rect 116 546 129 580
rect 163 546 176 580
rect 116 494 176 546
rect 116 460 129 494
rect 163 460 176 494
rect 116 414 176 460
rect 116 380 129 414
rect 163 380 176 414
rect 116 368 176 380
rect 206 580 266 592
rect 206 546 219 580
rect 253 546 266 580
rect 206 498 266 546
rect 206 464 219 498
rect 253 464 266 498
rect 206 368 266 464
rect 296 580 356 592
rect 296 546 309 580
rect 343 546 356 580
rect 296 494 356 546
rect 296 460 309 494
rect 343 460 356 494
rect 296 414 356 460
rect 296 380 309 414
rect 343 380 356 414
rect 296 368 356 380
rect 386 580 445 592
rect 386 546 399 580
rect 433 546 445 580
rect 386 498 445 546
rect 386 464 399 498
rect 433 464 445 498
rect 386 368 445 464
rect 499 580 558 592
rect 499 546 511 580
rect 545 546 558 580
rect 499 506 558 546
rect 499 472 511 506
rect 545 472 558 506
rect 499 438 558 472
rect 499 404 511 438
rect 545 404 558 438
rect 499 392 558 404
rect 588 580 648 592
rect 588 546 601 580
rect 635 546 648 580
rect 588 509 648 546
rect 588 475 601 509
rect 635 475 648 509
rect 588 392 648 475
rect 678 580 738 592
rect 678 546 691 580
rect 725 546 738 580
rect 678 392 738 546
rect 768 580 832 592
rect 768 546 783 580
rect 817 546 832 580
rect 768 496 832 546
rect 768 462 783 496
rect 817 462 832 496
rect 768 392 832 462
rect 862 580 932 592
rect 862 546 885 580
rect 919 546 932 580
rect 862 509 932 546
rect 862 475 885 509
rect 919 475 932 509
rect 862 438 932 475
rect 862 404 885 438
rect 919 404 932 438
rect 862 392 932 404
rect 962 577 1032 592
rect 962 543 985 577
rect 1019 543 1032 577
rect 962 392 1032 543
rect 1062 438 1122 592
rect 1062 404 1075 438
rect 1109 404 1122 438
rect 1062 392 1122 404
rect 1152 577 1212 592
rect 1152 543 1165 577
rect 1199 543 1212 577
rect 1152 392 1212 543
rect 1242 580 1311 592
rect 1242 546 1265 580
rect 1299 546 1311 580
rect 1242 508 1311 546
rect 1242 474 1265 508
rect 1299 474 1311 508
rect 1242 392 1311 474
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 139 176 173 210
rect 139 86 173 120
rect 239 99 273 133
rect 339 176 373 210
rect 339 86 373 120
rect 495 74 529 108
rect 600 158 634 192
rect 600 86 634 120
rect 702 74 736 108
rect 785 74 819 108
rect 868 74 902 108
rect 970 176 1004 210
rect 970 86 1004 120
rect 1070 86 1104 120
rect 1173 86 1207 120
<< pdiffc >>
rect 39 546 73 580
rect 39 464 73 498
rect 129 546 163 580
rect 129 460 163 494
rect 129 380 163 414
rect 219 546 253 580
rect 219 464 253 498
rect 309 546 343 580
rect 309 460 343 494
rect 309 380 343 414
rect 399 546 433 580
rect 399 464 433 498
rect 511 546 545 580
rect 511 472 545 506
rect 511 404 545 438
rect 601 546 635 580
rect 601 475 635 509
rect 691 546 725 580
rect 783 546 817 580
rect 783 462 817 496
rect 885 546 919 580
rect 885 475 919 509
rect 885 404 919 438
rect 985 543 1019 577
rect 1075 404 1109 438
rect 1165 543 1199 577
rect 1265 546 1299 580
rect 1265 474 1299 508
<< poly >>
rect 86 592 116 618
rect 176 592 206 618
rect 266 592 296 618
rect 356 592 386 618
rect 558 592 588 618
rect 648 592 678 618
rect 738 592 768 618
rect 832 592 862 618
rect 932 592 962 618
rect 1032 592 1062 618
rect 1122 592 1152 618
rect 1212 592 1242 618
rect 558 377 588 392
rect 648 377 678 392
rect 738 377 768 392
rect 832 377 862 392
rect 932 377 962 392
rect 1032 377 1062 392
rect 1122 377 1152 392
rect 1212 377 1242 392
rect 86 353 116 368
rect 176 353 206 368
rect 266 353 296 368
rect 356 353 386 368
rect 83 314 119 353
rect 173 314 209 353
rect 263 330 299 353
rect 353 330 389 353
rect 263 314 465 330
rect 83 280 279 314
rect 313 280 347 314
rect 381 280 415 314
rect 449 280 465 314
rect 555 310 591 377
rect 645 360 681 377
rect 735 360 771 377
rect 645 344 771 360
rect 645 310 697 344
rect 731 310 771 344
rect 829 310 865 377
rect 929 354 965 377
rect 921 338 987 354
rect 83 264 465 280
rect 98 222 128 264
rect 184 222 214 264
rect 284 222 314 264
rect 435 222 465 264
rect 523 294 589 310
rect 523 260 539 294
rect 573 260 589 294
rect 523 244 589 260
rect 559 222 589 244
rect 645 294 771 310
rect 813 294 879 310
rect 645 222 675 294
rect 813 260 829 294
rect 863 260 879 294
rect 921 304 937 338
rect 971 304 987 338
rect 921 288 987 304
rect 1029 297 1065 377
rect 1119 297 1155 377
rect 1209 356 1245 377
rect 813 244 879 260
rect 929 222 959 288
rect 1029 237 1155 297
rect 1197 323 1263 356
rect 1197 289 1213 323
rect 1247 289 1263 323
rect 1197 273 1263 289
rect 1029 222 1059 237
rect 1125 185 1155 237
rect 1125 169 1323 185
rect 1125 155 1273 169
rect 1257 135 1273 155
rect 1307 135 1323 169
rect 1257 101 1323 135
rect 98 48 128 74
rect 184 48 214 74
rect 284 48 314 74
rect 435 48 465 74
rect 559 48 589 74
rect 645 48 675 74
rect 929 48 959 74
rect 1029 48 1059 74
rect 1257 67 1273 101
rect 1307 67 1323 101
rect 1257 51 1323 67
<< polycont >>
rect 279 280 313 314
rect 347 280 381 314
rect 415 280 449 314
rect 697 310 731 344
rect 539 260 573 294
rect 829 260 863 294
rect 937 304 971 338
rect 1213 289 1247 323
rect 1273 135 1307 169
rect 1273 67 1307 101
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 23 580 89 649
rect 23 546 39 580
rect 73 546 89 580
rect 23 498 89 546
rect 23 464 39 498
rect 73 464 89 498
rect 123 580 169 596
rect 123 546 129 580
rect 163 546 169 580
rect 123 494 169 546
rect 123 460 129 494
rect 163 460 169 494
rect 203 580 269 649
rect 203 546 219 580
rect 253 546 269 580
rect 203 498 269 546
rect 203 464 219 498
rect 253 464 269 498
rect 303 580 349 596
rect 303 546 309 580
rect 343 546 349 580
rect 303 494 349 546
rect 123 430 169 460
rect 303 460 309 494
rect 343 460 349 494
rect 383 580 449 649
rect 383 546 399 580
rect 433 546 449 580
rect 383 498 449 546
rect 383 464 399 498
rect 433 464 449 498
rect 495 580 551 596
rect 495 546 511 580
rect 545 546 551 580
rect 495 506 551 546
rect 495 472 511 506
rect 545 472 551 506
rect 585 580 641 596
rect 585 546 601 580
rect 635 546 641 580
rect 675 580 741 649
rect 675 546 691 580
rect 725 546 741 580
rect 779 580 835 596
rect 779 546 783 580
rect 817 546 835 580
rect 585 512 641 546
rect 779 512 835 546
rect 585 509 835 512
rect 585 475 601 509
rect 635 496 835 509
rect 635 475 783 496
rect 585 472 783 475
rect 303 430 349 460
rect 495 438 551 472
rect 765 462 783 472
rect 817 462 835 496
rect 869 580 935 596
rect 869 546 885 580
rect 919 546 935 580
rect 869 509 935 546
rect 969 577 1215 596
rect 969 543 985 577
rect 1019 543 1165 577
rect 1199 543 1215 577
rect 969 540 1215 543
rect 1249 580 1315 596
rect 1249 546 1265 580
rect 1299 546 1315 580
rect 869 475 885 509
rect 919 506 935 509
rect 1249 508 1315 546
rect 1249 506 1265 508
rect 919 475 1265 506
rect 869 474 1265 475
rect 1299 474 1315 508
rect 869 472 1315 474
rect 869 438 935 472
rect 1249 458 1315 472
rect 25 414 455 430
rect 25 380 129 414
rect 163 380 309 414
rect 343 380 455 414
rect 495 404 511 438
rect 545 428 561 438
rect 869 428 885 438
rect 545 404 885 428
rect 919 404 935 438
rect 495 394 935 404
rect 495 388 561 394
rect 869 388 935 394
rect 1059 404 1075 438
rect 1109 424 1125 438
rect 1109 404 1327 424
rect 1059 390 1327 404
rect 25 364 455 380
rect 25 260 189 364
rect 681 344 747 360
rect 985 354 1257 356
rect 263 314 465 330
rect 263 280 279 314
rect 313 280 347 314
rect 381 280 415 314
rect 449 280 465 314
rect 681 310 697 344
rect 731 310 747 344
rect 921 338 1257 354
rect 523 294 647 310
rect 681 294 747 310
rect 813 294 879 310
rect 523 282 539 294
rect 263 264 465 280
rect 123 230 189 260
rect 23 210 89 226
rect 23 176 39 210
rect 73 176 89 210
rect 23 120 89 176
rect 23 86 39 120
rect 73 86 89 120
rect 23 17 89 86
rect 123 210 389 230
rect 123 176 139 210
rect 173 196 339 210
rect 173 176 189 196
rect 123 120 189 176
rect 323 176 339 196
rect 373 176 389 210
rect 123 86 139 120
rect 173 86 189 120
rect 123 70 189 86
rect 223 133 289 162
rect 223 99 239 133
rect 273 99 289 133
rect 223 17 289 99
rect 323 120 389 176
rect 431 192 465 264
rect 505 260 539 282
rect 573 260 647 294
rect 813 260 829 294
rect 863 260 879 294
rect 921 304 937 338
rect 971 323 1257 338
rect 971 304 1213 323
rect 921 289 1213 304
rect 1247 289 1257 323
rect 921 273 1257 289
rect 505 226 879 260
rect 1293 239 1327 390
rect 954 210 1327 239
rect 954 192 970 210
rect 431 158 600 192
rect 634 176 970 192
rect 1004 205 1327 210
rect 1004 176 1020 205
rect 634 158 1020 176
rect 323 86 339 120
rect 373 86 389 120
rect 323 70 389 86
rect 476 108 548 124
rect 476 74 495 108
rect 529 74 548 108
rect 476 17 548 74
rect 584 120 650 158
rect 584 86 600 120
rect 634 86 650 120
rect 584 70 650 86
rect 686 108 918 124
rect 686 74 702 108
rect 736 74 785 108
rect 819 74 868 108
rect 902 74 918 108
rect 686 17 918 74
rect 954 120 1020 158
rect 1257 169 1323 171
rect 954 86 970 120
rect 1004 86 1020 120
rect 954 70 1020 86
rect 1054 120 1223 136
rect 1054 86 1070 120
rect 1104 86 1173 120
rect 1207 86 1223 120
rect 1054 17 1223 86
rect 1257 135 1273 169
rect 1307 135 1323 169
rect 1257 101 1323 135
rect 1257 67 1273 101
rect 1307 67 1323 101
rect 1257 51 1323 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
<< metal1 >>
rect 0 683 1344 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 0 617 1344 649
rect 0 17 1344 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
rect 0 -49 1344 -17
<< labels >>
rlabel comment s 0 0 0 0 4 or4_4
flabel pwell s 0 0 1344 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 1344 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 1344 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 1344 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 127 390 161 424 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 223 390 257 424 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 319 390 353 424 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 415 390 449 424 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 1279 94 1313 128 0 FreeSans 340 0 0 0 D
port 4 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 1087 316 1121 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 1183 316 1217 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 511 242 545 276 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 607 242 641 276 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 A
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 1344 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1100322
string GDS_START 1088782
<< end >>
