magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 368 561
rect 31 326 82 487
rect 116 360 168 527
rect 202 326 254 487
rect 288 360 339 527
rect 31 292 351 326
rect 17 213 261 258
rect 295 179 351 292
rect 205 145 351 179
rect 112 17 171 122
rect 205 56 250 145
rect 284 17 350 111
rect 0 -17 368 17
<< metal1 >>
rect 0 496 368 592
rect 0 -48 368 48
<< labels >>
rlabel locali s 17 213 261 258 6 A
port 1 nsew signal input
rlabel locali s 295 179 351 292 6 Y
port 2 nsew signal output
rlabel locali s 205 145 351 179 6 Y
port 2 nsew signal output
rlabel locali s 205 56 250 145 6 Y
port 2 nsew signal output
rlabel locali s 202 326 254 487 6 Y
port 2 nsew signal output
rlabel locali s 31 326 82 487 6 Y
port 2 nsew signal output
rlabel locali s 31 292 351 326 6 Y
port 2 nsew signal output
rlabel locali s 284 17 350 111 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 112 17 171 122 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 0 -17 368 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 368 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 288 360 339 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 116 360 168 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 0 527 368 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 496 368 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 368 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3219486
string GDS_START 3215244
<< end >>
