magic
tech sky130A
magscale 1 2
timestamp 1604502693
<< nwell >>
rect -38 261 1602 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 419 47 449 177
rect 503 47 533 177
rect 691 47 721 177
rect 775 47 805 177
rect 859 47 889 177
rect 943 47 973 177
rect 1131 47 1161 177
rect 1215 47 1245 177
rect 1299 47 1329 177
rect 1383 47 1413 177
<< pmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 519 297 549 497
rect 603 297 633 497
rect 691 297 721 497
rect 775 297 805 497
rect 859 297 889 497
rect 943 297 973 497
rect 1031 297 1061 497
rect 1215 297 1245 497
rect 1299 297 1329 497
rect 1383 297 1413 497
<< ndiff >>
rect 27 93 79 177
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 101 163 177
rect 109 67 119 101
rect 153 67 163 101
rect 109 47 163 67
rect 193 93 247 177
rect 193 59 203 93
rect 237 59 247 93
rect 193 47 247 59
rect 277 101 331 177
rect 277 67 287 101
rect 321 67 331 101
rect 277 47 331 67
rect 361 93 419 177
rect 361 59 371 93
rect 405 59 419 93
rect 361 47 419 59
rect 449 101 503 177
rect 449 67 459 101
rect 493 67 503 101
rect 449 47 503 67
rect 533 93 585 177
rect 533 59 543 93
rect 577 59 585 93
rect 533 47 585 59
rect 639 93 691 177
rect 639 59 647 93
rect 681 59 691 93
rect 639 47 691 59
rect 721 163 775 177
rect 721 129 731 163
rect 765 129 775 163
rect 721 47 775 129
rect 805 147 859 177
rect 805 113 815 147
rect 849 113 859 147
rect 805 47 859 113
rect 889 93 943 177
rect 889 59 899 93
rect 933 59 943 93
rect 889 47 943 59
rect 973 163 1025 177
rect 973 129 983 163
rect 1017 129 1025 163
rect 973 47 1025 129
rect 1079 163 1131 177
rect 1079 129 1087 163
rect 1121 129 1131 163
rect 1079 47 1131 129
rect 1161 93 1215 177
rect 1161 59 1171 93
rect 1205 59 1215 93
rect 1161 47 1215 59
rect 1245 163 1299 177
rect 1245 129 1255 163
rect 1289 129 1299 163
rect 1245 47 1299 129
rect 1329 93 1383 177
rect 1329 59 1339 93
rect 1373 59 1383 93
rect 1329 47 1383 59
rect 1413 101 1465 177
rect 1413 67 1423 101
rect 1457 67 1465 101
rect 1413 47 1465 67
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 297 79 383
rect 109 477 163 497
rect 109 443 119 477
rect 153 443 163 477
rect 109 409 163 443
rect 109 375 119 409
rect 153 375 163 409
rect 109 297 163 375
rect 193 485 247 497
rect 193 451 203 485
rect 237 451 247 485
rect 193 417 247 451
rect 193 383 203 417
rect 237 383 247 417
rect 193 297 247 383
rect 277 477 331 497
rect 277 443 287 477
rect 321 443 331 477
rect 277 409 331 443
rect 277 375 287 409
rect 321 375 331 409
rect 277 297 331 375
rect 361 485 413 497
rect 361 451 371 485
rect 405 451 413 485
rect 361 417 413 451
rect 361 383 371 417
rect 405 383 413 417
rect 361 297 413 383
rect 467 477 519 497
rect 467 443 475 477
rect 509 443 519 477
rect 467 409 519 443
rect 467 375 475 409
rect 509 375 519 409
rect 467 297 519 375
rect 549 425 603 497
rect 549 391 559 425
rect 593 391 603 425
rect 549 357 603 391
rect 549 323 559 357
rect 593 323 603 357
rect 549 297 603 323
rect 633 477 691 497
rect 633 443 647 477
rect 681 443 691 477
rect 633 409 691 443
rect 633 375 647 409
rect 681 375 691 409
rect 633 297 691 375
rect 721 485 775 497
rect 721 451 731 485
rect 765 451 775 485
rect 721 417 775 451
rect 721 383 731 417
rect 765 383 775 417
rect 721 297 775 383
rect 805 477 859 497
rect 805 443 815 477
rect 849 443 859 477
rect 805 409 859 443
rect 805 375 815 409
rect 849 375 859 409
rect 805 297 859 375
rect 889 485 943 497
rect 889 451 899 485
rect 933 451 943 485
rect 889 417 943 451
rect 889 383 899 417
rect 933 383 943 417
rect 889 297 943 383
rect 973 477 1031 497
rect 973 443 987 477
rect 1021 443 1031 477
rect 973 409 1031 443
rect 973 375 987 409
rect 1021 375 1031 409
rect 973 297 1031 375
rect 1061 485 1215 497
rect 1061 451 1085 485
rect 1119 451 1157 485
rect 1191 451 1215 485
rect 1061 417 1215 451
rect 1061 383 1085 417
rect 1119 383 1157 417
rect 1191 383 1215 417
rect 1061 297 1215 383
rect 1245 477 1299 497
rect 1245 443 1255 477
rect 1289 443 1299 477
rect 1245 409 1299 443
rect 1245 375 1255 409
rect 1289 375 1299 409
rect 1245 297 1299 375
rect 1329 485 1383 497
rect 1329 451 1339 485
rect 1373 451 1383 485
rect 1329 417 1383 451
rect 1329 383 1339 417
rect 1373 383 1383 417
rect 1329 297 1383 383
rect 1413 477 1465 497
rect 1413 443 1423 477
rect 1457 443 1465 477
rect 1413 409 1465 443
rect 1413 375 1423 409
rect 1457 375 1465 409
rect 1413 297 1465 375
<< ndiffc >>
rect 35 59 69 93
rect 119 67 153 101
rect 203 59 237 93
rect 287 67 321 101
rect 371 59 405 93
rect 459 67 493 101
rect 543 59 577 93
rect 647 59 681 93
rect 731 129 765 163
rect 815 113 849 147
rect 899 59 933 93
rect 983 129 1017 163
rect 1087 129 1121 163
rect 1171 59 1205 93
rect 1255 129 1289 163
rect 1339 59 1373 93
rect 1423 67 1457 101
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 119 443 153 477
rect 119 375 153 409
rect 203 451 237 485
rect 203 383 237 417
rect 287 443 321 477
rect 287 375 321 409
rect 371 451 405 485
rect 371 383 405 417
rect 475 443 509 477
rect 475 375 509 409
rect 559 391 593 425
rect 559 323 593 357
rect 647 443 681 477
rect 647 375 681 409
rect 731 451 765 485
rect 731 383 765 417
rect 815 443 849 477
rect 815 375 849 409
rect 899 451 933 485
rect 899 383 933 417
rect 987 443 1021 477
rect 987 375 1021 409
rect 1085 451 1119 485
rect 1157 451 1191 485
rect 1085 383 1119 417
rect 1157 383 1191 417
rect 1255 443 1289 477
rect 1255 375 1289 409
rect 1339 451 1373 485
rect 1339 383 1373 417
rect 1423 443 1457 477
rect 1423 375 1457 409
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 519 497 549 523
rect 603 497 633 523
rect 691 497 721 523
rect 775 497 805 523
rect 859 497 889 523
rect 943 497 973 523
rect 1031 497 1061 523
rect 1215 497 1245 523
rect 1299 497 1329 523
rect 1383 497 1413 523
rect 79 265 109 297
rect 163 265 193 297
rect 247 265 277 297
rect 331 265 361 297
rect 519 265 549 297
rect 603 265 633 297
rect 79 259 361 265
rect 79 249 368 259
rect 79 215 114 249
rect 148 215 182 249
rect 216 215 250 249
rect 284 215 318 249
rect 352 215 368 249
rect 79 205 368 215
rect 419 249 633 265
rect 691 265 721 297
rect 775 265 805 297
rect 691 259 805 265
rect 859 259 889 297
rect 943 259 973 297
rect 1031 259 1061 297
rect 1215 259 1245 297
rect 419 215 443 249
rect 477 215 511 249
rect 545 215 579 249
rect 613 215 633 249
rect 79 199 361 205
rect 79 177 109 199
rect 163 177 193 199
rect 247 177 277 199
rect 331 177 361 199
rect 419 199 633 215
rect 679 249 813 259
rect 679 215 695 249
rect 729 215 763 249
rect 797 215 813 249
rect 679 205 813 215
rect 855 249 989 259
rect 855 215 871 249
rect 905 215 939 249
rect 973 215 989 249
rect 855 205 989 215
rect 1031 249 1245 259
rect 1031 215 1047 249
rect 1081 215 1119 249
rect 1153 215 1187 249
rect 1221 215 1245 249
rect 1031 205 1245 215
rect 691 199 805 205
rect 419 177 449 199
rect 503 177 533 199
rect 691 177 721 199
rect 775 177 805 199
rect 859 177 889 205
rect 943 177 973 205
rect 1131 177 1161 205
rect 1215 177 1245 205
rect 1299 259 1329 297
rect 1383 259 1413 297
rect 1299 249 1501 259
rect 1299 215 1315 249
rect 1349 215 1383 249
rect 1417 215 1451 249
rect 1485 215 1501 249
rect 1299 205 1501 215
rect 1299 177 1329 205
rect 1383 177 1413 205
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 419 21 449 47
rect 503 21 533 47
rect 691 21 721 47
rect 775 21 805 47
rect 859 21 889 47
rect 943 21 973 47
rect 1131 21 1161 47
rect 1215 21 1245 47
rect 1299 21 1329 47
rect 1383 21 1413 47
<< polycont >>
rect 114 215 148 249
rect 182 215 216 249
rect 250 215 284 249
rect 318 215 352 249
rect 443 215 477 249
rect 511 215 545 249
rect 579 215 613 249
rect 695 215 729 249
rect 763 215 797 249
rect 871 215 905 249
rect 939 215 973 249
rect 1047 215 1081 249
rect 1119 215 1153 249
rect 1187 215 1221 249
rect 1315 215 1349 249
rect 1383 215 1417 249
rect 1451 215 1485 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 19 485 85 527
rect 19 451 35 485
rect 69 451 85 485
rect 19 417 85 451
rect 19 383 35 417
rect 69 383 85 417
rect 119 477 153 493
rect 119 409 153 443
rect 187 485 253 527
rect 187 451 203 485
rect 237 451 253 485
rect 187 417 253 451
rect 187 383 203 417
rect 237 383 253 417
rect 287 477 321 493
rect 287 409 321 443
rect 119 349 153 375
rect 355 485 425 527
rect 355 451 371 485
rect 405 451 425 485
rect 355 417 425 451
rect 355 383 371 417
rect 405 383 425 417
rect 475 477 681 493
rect 509 459 647 477
rect 475 409 509 443
rect 287 349 321 375
rect 543 391 559 425
rect 593 391 609 425
rect 647 409 681 443
rect 475 359 509 375
rect 30 315 321 349
rect 559 357 593 391
rect 355 323 559 325
rect 30 161 64 315
rect 355 291 593 323
rect 715 485 781 527
rect 715 451 731 485
rect 765 451 781 485
rect 715 417 781 451
rect 715 383 731 417
rect 765 383 781 417
rect 815 477 849 493
rect 815 409 849 443
rect 647 341 681 375
rect 883 485 949 527
rect 883 451 899 485
rect 933 451 949 485
rect 883 417 949 451
rect 883 383 899 417
rect 933 383 949 417
rect 987 477 1021 493
rect 987 409 1021 443
rect 815 341 849 375
rect 1069 485 1207 527
rect 1069 451 1085 485
rect 1119 451 1157 485
rect 1191 451 1207 485
rect 1069 417 1207 451
rect 1069 383 1085 417
rect 1119 383 1157 417
rect 1191 383 1207 417
rect 1255 477 1289 493
rect 1255 409 1289 443
rect 987 341 1021 375
rect 1323 485 1389 527
rect 1323 451 1339 485
rect 1373 451 1389 485
rect 1323 417 1389 451
rect 1323 383 1339 417
rect 1373 383 1389 417
rect 1423 477 1457 493
rect 1423 409 1457 443
rect 1255 341 1289 375
rect 1423 341 1457 375
rect 647 307 1474 341
rect 355 249 389 291
rect 98 215 114 249
rect 148 215 182 249
rect 216 215 250 249
rect 284 215 318 249
rect 352 215 389 249
rect 427 249 629 256
rect 427 215 443 249
rect 477 215 511 249
rect 545 215 579 249
rect 613 215 629 249
rect 679 249 813 259
rect 679 215 695 249
rect 729 215 763 249
rect 797 215 813 249
rect 855 249 995 257
rect 855 215 871 249
rect 905 215 939 249
rect 973 215 995 249
rect 1031 249 1237 259
rect 1031 215 1047 249
rect 1081 215 1119 249
rect 1153 215 1187 249
rect 1221 215 1237 249
rect 1299 249 1501 259
rect 1299 215 1315 249
rect 1349 215 1383 249
rect 1417 215 1451 249
rect 1485 215 1501 249
rect 355 163 389 215
rect 30 127 321 161
rect 355 129 731 163
rect 765 129 781 163
rect 815 147 983 163
rect 119 101 153 127
rect 19 59 35 93
rect 69 59 85 93
rect 19 17 85 59
rect 287 101 321 127
rect 119 51 153 67
rect 187 59 203 93
rect 237 59 253 93
rect 187 17 253 59
rect 459 101 493 129
rect 287 51 321 67
rect 355 59 371 93
rect 405 59 425 93
rect 355 17 425 59
rect 849 129 983 147
rect 1017 129 1033 163
rect 1071 129 1087 163
rect 1121 129 1255 163
rect 1289 129 1457 163
rect 815 93 849 113
rect 1423 101 1457 129
rect 459 51 493 67
rect 527 59 543 93
rect 577 59 593 93
rect 631 59 647 93
rect 681 59 849 93
rect 883 59 899 93
rect 933 59 1171 93
rect 1205 59 1221 93
rect 1323 59 1339 93
rect 1373 59 1389 93
rect 527 17 593 59
rect 1323 17 1389 59
rect 1423 51 1457 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
<< metal1 >>
rect 0 561 1564 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 0 496 1564 527
rect 0 17 1564 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
rect 0 -48 1564 -17
<< labels >>
flabel corelocali s 30 153 64 187 0 FreeSans 200 0 0 0 X
port 10 nsew
flabel corelocali s 1330 221 1364 255 0 FreeSans 200 0 0 0 A4
port 4 nsew
flabel corelocali s 1422 221 1456 255 0 FreeSans 200 0 0 0 A4
port 4 nsew
flabel corelocali s 1146 221 1180 255 0 FreeSans 200 0 0 0 A3
port 3 nsew
flabel corelocali s 866 221 900 255 0 FreeSans 200 0 0 0 A2
port 2 nsew
flabel corelocali s 1050 221 1084 255 0 FreeSans 200 0 0 0 A3
port 3 nsew
flabel corelocali s 682 221 716 255 0 FreeSans 200 0 0 0 A1
port 1 nsew
flabel corelocali s 958 221 992 255 0 FreeSans 200 0 0 0 A2
port 2 nsew
flabel corelocali s 494 221 528 255 0 FreeSans 200 0 0 0 B1
port 5 nsew
flabel corelocali s 774 221 808 255 0 FreeSans 200 0 0 0 A1
port 1 nsew
flabel corelocali s 586 221 620 255 0 FreeSans 200 0 0 0 B1
port 5 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 200 0 0 0 X
port 10 nsew
flabel corelocali s 30 289 64 323 0 FreeSans 200 0 0 0 X
port 10 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew
rlabel comment s 0 0 0 0 4 a41o_4
<< properties >>
string FIXED_BBOX 0 0 1564 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3703642
string GDS_START 3691176
string path 0.000 0.000 39.100 0.000 
<< end >>
