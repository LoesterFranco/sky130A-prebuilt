magic
tech sky130A
magscale 1 2
timestamp 1601050058
<< locali >>
rect 638 338 719 493
rect 17 215 107 258
rect 669 128 719 338
rect 638 51 719 128
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 17 326 86 493
rect 120 360 186 527
rect 17 292 211 326
rect 141 263 211 292
rect 276 264 346 493
rect 398 333 448 493
rect 538 367 604 527
rect 398 299 516 333
rect 482 265 516 299
rect 141 205 227 263
rect 276 214 448 264
rect 141 181 211 205
rect 17 147 211 181
rect 17 51 83 147
rect 117 17 183 113
rect 276 51 346 214
rect 482 199 635 265
rect 482 180 516 199
rect 398 146 516 180
rect 398 51 448 146
rect 538 17 604 120
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel locali s 17 215 107 258 6 A
port 1 nsew signal input
rlabel locali s 669 128 719 338 6 X
port 2 nsew signal output
rlabel locali s 638 338 719 493 6 X
port 2 nsew signal output
rlabel locali s 638 51 719 128 6 X
port 2 nsew signal output
rlabel metal1 s 0 -48 736 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 736 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3191644
string GDS_START 3185492
<< end >>
