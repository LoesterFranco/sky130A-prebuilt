magic
tech sky130A
magscale 1 2
timestamp 1604502710
<< nwell >>
rect -38 332 710 704
<< pwell >>
rect 0 0 672 49
<< scpmos >>
rect 83 368 119 592
rect 183 368 219 592
rect 305 368 341 592
rect 463 368 499 592
rect 553 368 589 592
<< nmoslvt >>
rect 89 74 119 222
rect 167 74 197 222
rect 361 74 391 222
rect 439 74 469 222
rect 553 74 583 222
<< ndiff >>
rect 27 196 89 222
rect 27 162 39 196
rect 73 162 89 196
rect 27 120 89 162
rect 27 86 39 120
rect 73 86 89 120
rect 27 74 89 86
rect 119 74 167 222
rect 197 193 361 222
rect 197 159 208 193
rect 242 159 316 193
rect 350 159 361 193
rect 197 116 361 159
rect 197 82 208 116
rect 242 82 316 116
rect 350 82 361 116
rect 197 74 361 82
rect 391 74 439 222
rect 469 74 553 222
rect 583 196 640 222
rect 583 162 594 196
rect 628 162 640 196
rect 583 120 640 162
rect 583 86 594 120
rect 628 86 640 120
rect 583 74 640 86
<< pdiff >>
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 497 83 546
rect 27 463 39 497
rect 73 463 83 497
rect 27 414 83 463
rect 27 380 39 414
rect 73 380 83 414
rect 27 368 83 380
rect 119 531 183 592
rect 119 497 139 531
rect 173 497 183 531
rect 119 414 183 497
rect 119 380 139 414
rect 173 380 183 414
rect 119 368 183 380
rect 219 580 305 592
rect 219 546 239 580
rect 273 546 305 580
rect 219 462 305 546
rect 219 428 239 462
rect 273 428 305 462
rect 219 368 305 428
rect 341 572 463 592
rect 341 538 351 572
rect 385 538 419 572
rect 453 538 463 572
rect 341 368 463 538
rect 499 580 553 592
rect 499 546 509 580
rect 543 546 553 580
rect 499 497 553 546
rect 499 463 509 497
rect 543 463 553 497
rect 499 414 553 463
rect 499 380 509 414
rect 543 380 553 414
rect 499 368 553 380
rect 589 580 645 592
rect 589 546 599 580
rect 633 546 645 580
rect 589 497 645 546
rect 589 463 599 497
rect 633 463 645 497
rect 589 414 645 463
rect 589 380 599 414
rect 633 380 645 414
rect 589 368 645 380
<< ndiffc >>
rect 39 162 73 196
rect 39 86 73 120
rect 208 159 242 193
rect 316 159 350 193
rect 208 82 242 116
rect 316 82 350 116
rect 594 162 628 196
rect 594 86 628 120
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 139 497 173 531
rect 139 380 173 414
rect 239 546 273 580
rect 239 428 273 462
rect 351 538 385 572
rect 419 538 453 572
rect 509 546 543 580
rect 509 463 543 497
rect 509 380 543 414
rect 599 546 633 580
rect 599 463 633 497
rect 599 380 633 414
<< poly >>
rect 83 592 119 618
rect 183 592 219 618
rect 305 592 341 618
rect 463 592 499 618
rect 553 592 589 618
rect 83 310 119 368
rect 183 310 219 368
rect 305 310 341 368
rect 463 310 499 368
rect 553 310 589 368
rect 23 294 119 310
rect 23 260 39 294
rect 73 260 119 294
rect 23 244 119 260
rect 89 222 119 244
rect 167 294 257 310
rect 167 260 207 294
rect 241 260 257 294
rect 167 244 257 260
rect 305 294 391 310
rect 305 260 321 294
rect 355 260 391 294
rect 305 244 391 260
rect 167 222 197 244
rect 361 222 391 244
rect 439 294 505 310
rect 439 260 455 294
rect 489 260 505 294
rect 439 244 505 260
rect 553 294 619 310
rect 553 260 569 294
rect 603 260 619 294
rect 553 244 619 260
rect 439 222 469 244
rect 553 222 583 244
rect 89 48 119 74
rect 167 48 197 74
rect 361 48 391 74
rect 439 48 469 74
rect 553 48 583 74
<< polycont >>
rect 39 260 73 294
rect 207 260 241 294
rect 321 260 355 294
rect 455 260 489 294
rect 569 260 603 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 23 581 289 615
rect 23 580 89 581
rect 23 546 39 580
rect 73 546 89 580
rect 223 580 289 581
rect 23 497 89 546
rect 23 463 39 497
rect 73 463 89 497
rect 23 414 89 463
rect 23 380 39 414
rect 73 380 89 414
rect 23 364 89 380
rect 123 531 189 547
rect 123 497 139 531
rect 173 497 189 531
rect 123 414 189 497
rect 123 380 139 414
rect 173 380 189 414
rect 223 546 239 580
rect 273 546 289 580
rect 223 498 289 546
rect 335 572 469 649
rect 335 538 351 572
rect 385 538 419 572
rect 453 538 469 572
rect 335 532 469 538
rect 503 580 559 596
rect 503 546 509 580
rect 543 546 559 580
rect 503 498 559 546
rect 223 497 559 498
rect 223 464 509 497
rect 223 462 284 464
rect 223 428 239 462
rect 273 428 284 462
rect 493 463 509 464
rect 543 463 559 497
rect 223 412 284 428
rect 123 378 189 380
rect 318 378 455 430
rect 123 344 455 378
rect 493 414 559 463
rect 493 380 509 414
rect 543 380 559 414
rect 493 364 559 380
rect 599 580 649 649
rect 633 546 649 580
rect 599 497 649 546
rect 633 463 649 497
rect 599 414 649 463
rect 633 380 649 414
rect 599 364 649 380
rect 23 294 89 310
rect 23 260 39 294
rect 73 260 89 294
rect 23 236 89 260
rect 123 202 157 344
rect 191 294 263 310
rect 191 260 207 294
rect 241 260 263 294
rect 191 236 263 260
rect 305 294 371 310
rect 305 260 321 294
rect 355 260 371 294
rect 305 236 371 260
rect 409 294 505 310
rect 409 260 455 294
rect 489 260 505 294
rect 23 196 89 202
rect 23 162 39 196
rect 73 162 89 196
rect 23 120 89 162
rect 23 86 39 120
rect 73 86 89 120
rect 23 17 89 86
rect 123 193 366 202
rect 123 159 208 193
rect 242 159 316 193
rect 350 159 366 193
rect 123 116 366 159
rect 123 82 208 116
rect 242 82 316 116
rect 350 82 366 116
rect 409 88 505 260
rect 553 294 647 310
rect 553 260 569 294
rect 603 260 647 294
rect 553 236 647 260
rect 578 196 644 202
rect 578 162 594 196
rect 628 162 644 196
rect 578 120 644 162
rect 123 70 366 82
rect 578 86 594 120
rect 628 86 644 120
rect 578 17 644 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
rlabel comment s 0 0 0 0 4 a32oi_1
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 607 242 641 276 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 B2
port 5 nsew
flabel corelocali s 223 242 257 276 0 FreeSans 340 0 0 0 B1
port 4 nsew
flabel corelocali s 415 94 449 128 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 415 168 449 202 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 415 242 449 276 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 415 390 449 424 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 319 242 353 276 0 FreeSans 340 0 0 0 A1
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 672 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3722428
string GDS_START 3716062
<< end >>
