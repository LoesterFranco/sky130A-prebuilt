magic
tech sky130A
magscale 1 2
timestamp 1604502741
<< locali >>
rect 85 322 167 390
rect 217 364 316 430
rect 85 288 409 322
rect 85 256 136 288
rect 358 252 409 288
rect 511 228 561 430
rect 663 236 743 310
rect 2713 210 2763 596
rect 2676 70 2763 210
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 17 498 72 596
rect 112 532 178 649
rect 286 532 477 582
rect 513 566 579 649
rect 443 498 681 532
rect 715 516 781 649
rect 821 579 1169 613
rect 821 516 855 579
rect 17 464 409 498
rect 17 460 72 464
rect 17 222 51 460
rect 358 366 409 464
rect 178 222 244 254
rect 17 188 244 222
rect 443 218 477 498
rect 647 482 681 498
rect 889 482 1001 545
rect 647 448 1001 482
rect 1035 453 1101 545
rect 1135 503 1169 579
rect 1245 537 1295 649
rect 1329 579 1499 613
rect 1329 503 1363 579
rect 1135 469 1363 503
rect 595 364 843 414
rect 17 70 105 188
rect 311 184 477 218
rect 595 202 629 364
rect 777 270 843 364
rect 139 17 205 154
rect 311 70 377 184
rect 475 17 541 150
rect 595 70 661 202
rect 695 17 761 202
rect 795 85 845 226
rect 889 153 923 448
rect 957 221 1001 414
rect 1035 289 1069 453
rect 1135 389 1169 469
rect 1397 435 1431 545
rect 1103 355 1169 389
rect 1203 401 1431 435
rect 1465 428 1499 579
rect 1533 462 1583 649
rect 1717 581 2086 615
rect 1623 504 1673 545
rect 1717 538 1783 581
rect 1913 504 1979 547
rect 2020 512 2086 581
rect 2126 512 2160 649
rect 1623 470 1979 504
rect 2200 478 2274 596
rect 1203 359 1269 401
rect 1465 394 1589 428
rect 1103 323 1146 355
rect 1330 321 1387 367
rect 1180 289 1387 321
rect 1429 350 1511 360
rect 1429 316 1471 350
rect 1505 316 1511 350
rect 1555 350 1589 394
rect 1623 384 1673 470
rect 1818 358 1873 436
rect 1913 392 1979 470
rect 2013 444 2274 478
rect 2308 478 2374 596
rect 2414 512 2464 649
rect 2308 444 2388 478
rect 2013 358 2047 444
rect 2240 410 2274 444
rect 1555 316 1768 350
rect 1818 324 2047 358
rect 2137 350 2206 410
rect 1429 308 1511 316
rect 1035 287 1387 289
rect 1035 255 1214 287
rect 1330 274 1387 287
rect 1734 290 1768 316
rect 1552 274 1686 282
rect 957 187 1041 221
rect 889 119 973 153
rect 1007 85 1041 187
rect 795 51 1041 85
rect 1075 77 1125 255
rect 1248 206 1296 253
rect 1330 240 1686 274
rect 1552 224 1686 240
rect 1734 224 1800 290
rect 1248 172 1401 206
rect 1839 188 1873 324
rect 2137 316 2143 350
rect 2177 316 2206 350
rect 2137 276 2206 316
rect 2240 276 2320 410
rect 1958 242 2092 262
rect 2354 242 2388 444
rect 1958 208 2388 242
rect 2506 399 2572 575
rect 2606 399 2672 649
rect 2506 310 2540 399
rect 2506 244 2679 310
rect 1958 196 2354 208
rect 2506 201 2540 244
rect 1223 17 1289 138
rect 1335 114 1401 172
rect 1491 17 1661 188
rect 1759 70 1873 188
rect 2165 17 2231 162
rect 2279 70 2354 196
rect 2474 174 2540 201
rect 2391 108 2540 174
rect 2576 17 2642 210
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 1471 316 1505 350
rect 2143 316 2177 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
<< metal1 >>
rect 0 683 2784 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 0 617 2784 649
rect 1459 350 1517 356
rect 1459 316 1471 350
rect 1505 347 1517 350
rect 2131 350 2189 356
rect 2131 347 2143 350
rect 1505 319 2143 347
rect 1505 316 1517 319
rect 1459 310 1517 316
rect 2131 316 2143 319
rect 2177 316 2189 350
rect 2131 310 2189 316
rect 0 17 2784 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
rect 0 -49 2784 -17
<< labels >>
rlabel locali s 217 364 316 430 6 D
port 1 nsew signal input
rlabel locali s 2713 210 2763 596 6 Q
port 2 nsew signal output
rlabel locali s 2676 70 2763 210 6 Q
port 2 nsew signal output
rlabel locali s 511 228 561 430 6 SCD
port 3 nsew signal input
rlabel locali s 358 252 409 288 6 SCE
port 4 nsew signal input
rlabel locali s 85 322 167 390 6 SCE
port 4 nsew signal input
rlabel locali s 85 288 409 322 6 SCE
port 4 nsew signal input
rlabel locali s 85 256 136 288 6 SCE
port 4 nsew signal input
rlabel metal1 s 2131 347 2189 356 6 SET_B
port 5 nsew signal input
rlabel metal1 s 2131 310 2189 319 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1459 347 1517 356 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1459 319 2189 347 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1459 310 1517 319 6 SET_B
port 5 nsew signal input
rlabel locali s 663 236 743 310 6 CLK
port 6 nsew clock input
rlabel metal1 s 0 -49 2784 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 617 2784 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2784 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 122894
string GDS_START 102822
<< end >>
