magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 119 367 173 527
rect 307 367 361 527
rect 495 367 549 527
rect 683 367 737 527
rect 871 367 925 527
rect 1059 297 1119 527
rect 28 215 248 255
rect 123 17 179 113
rect 301 17 361 113
rect 495 17 549 113
rect 683 17 737 113
rect 871 17 925 113
rect 1059 17 1109 177
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< obsli1 >>
rect 19 323 85 493
rect 207 323 273 493
rect 395 323 461 493
rect 583 323 649 493
rect 771 323 837 493
rect 959 323 1025 493
rect 19 289 319 323
rect 395 289 1025 323
rect 284 249 319 289
rect 284 215 809 249
rect 284 181 319 215
rect 858 181 1025 289
rect 29 147 319 181
rect 395 147 1025 181
rect 29 51 89 147
rect 213 51 267 147
rect 395 51 461 147
rect 583 51 649 147
rect 771 51 837 147
rect 959 51 1025 147
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< via1 >>
rect 699 212 751 264
rect 763 212 815 264
<< obsm1 >>
rect 693 212 699 264
rect 751 212 763 264
rect 815 261 821 264
rect 815 215 1030 261
rect 815 212 821 215
<< via2 >>
rect 689 264 745 266
rect 769 264 825 266
rect 689 212 699 264
rect 699 212 745 264
rect 769 212 815 264
rect 815 212 825 264
rect 689 210 745 212
rect 769 210 825 212
<< obsm2 >>
rect 689 266 825 275
rect 745 264 769 266
rect 751 212 763 264
rect 745 210 769 212
rect 689 201 825 210
<< obsm3 >>
rect 679 270 835 271
rect 679 206 685 270
rect 749 206 765 270
rect 829 206 835 270
rect 679 205 835 206
<< via3 >>
rect 685 266 749 270
rect 685 210 689 266
rect 689 210 745 266
rect 745 210 749 266
rect 685 206 749 210
rect 765 266 829 270
rect 765 210 769 266
rect 769 210 825 266
rect 825 210 829 266
rect 765 206 829 210
<< obsm4 >>
rect 274 136 594 372
<< via4 >>
rect 594 270 830 372
rect 594 206 685 270
rect 685 206 749 270
rect 749 206 765 270
rect 765 206 829 270
rect 829 206 830 270
rect 594 136 830 206
<< metal5 >>
rect 250 390 854 432
<< obsm5 >>
rect 250 372 854 389
rect 250 136 594 372
rect 830 136 854 372
rect 250 112 854 136
<< labels >>
rlabel locali s 28 215 248 255 6 A
port 1 nsew signal input
rlabel metal5 s 250 390 854 432 6 X
port 2 nsew signal output
rlabel viali s 1133 -17 1167 17 8 VGND
port 3 nsew ground input
rlabel viali s 1041 -17 1075 17 8 VGND
port 3 nsew ground input
rlabel viali s 949 -17 983 17 8 VGND
port 3 nsew ground input
rlabel viali s 857 -17 891 17 8 VGND
port 3 nsew ground input
rlabel viali s 765 -17 799 17 8 VGND
port 3 nsew ground input
rlabel viali s 673 -17 707 17 8 VGND
port 3 nsew ground input
rlabel viali s 581 -17 615 17 8 VGND
port 3 nsew ground input
rlabel viali s 489 -17 523 17 8 VGND
port 3 nsew ground input
rlabel viali s 397 -17 431 17 8 VGND
port 3 nsew ground input
rlabel viali s 305 -17 339 17 8 VGND
port 3 nsew ground input
rlabel viali s 213 -17 247 17 8 VGND
port 3 nsew ground input
rlabel viali s 121 -17 155 17 8 VGND
port 3 nsew ground input
rlabel viali s 29 -17 63 17 8 VGND
port 3 nsew ground input
rlabel locali s 1059 17 1109 177 6 VGND
port 3 nsew ground input
rlabel locali s 871 17 925 113 6 VGND
port 3 nsew ground input
rlabel locali s 683 17 737 113 6 VGND
port 3 nsew ground input
rlabel locali s 495 17 549 113 6 VGND
port 3 nsew ground input
rlabel locali s 301 17 361 113 6 VGND
port 3 nsew ground input
rlabel locali s 123 17 179 113 6 VGND
port 3 nsew ground input
rlabel locali s 0 -17 1196 17 8 VGND
port 3 nsew ground input
rlabel metal1 s 0 -48 1196 48 8 VGND
port 3 nsew ground input
rlabel viali s 1133 527 1167 561 6 VPWR
port 4 nsew power input
rlabel viali s 1041 527 1075 561 6 VPWR
port 4 nsew power input
rlabel viali s 949 527 983 561 6 VPWR
port 4 nsew power input
rlabel viali s 857 527 891 561 6 VPWR
port 4 nsew power input
rlabel viali s 765 527 799 561 6 VPWR
port 4 nsew power input
rlabel viali s 673 527 707 561 6 VPWR
port 4 nsew power input
rlabel viali s 581 527 615 561 6 VPWR
port 4 nsew power input
rlabel viali s 489 527 523 561 6 VPWR
port 4 nsew power input
rlabel viali s 397 527 431 561 6 VPWR
port 4 nsew power input
rlabel viali s 305 527 339 561 6 VPWR
port 4 nsew power input
rlabel viali s 213 527 247 561 6 VPWR
port 4 nsew power input
rlabel viali s 121 527 155 561 6 VPWR
port 4 nsew power input
rlabel viali s 29 527 63 561 6 VPWR
port 4 nsew power input
rlabel locali s 1059 297 1119 527 6 VPWR
port 4 nsew power input
rlabel locali s 871 367 925 527 6 VPWR
port 4 nsew power input
rlabel locali s 683 367 737 527 6 VPWR
port 4 nsew power input
rlabel locali s 495 367 549 527 6 VPWR
port 4 nsew power input
rlabel locali s 307 367 361 527 6 VPWR
port 4 nsew power input
rlabel locali s 119 367 173 527 6 VPWR
port 4 nsew power input
rlabel locali s 0 527 1196 561 6 VPWR
port 4 nsew power input
rlabel metal1 s 0 496 1196 592 6 VPWR
port 4 nsew power input
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 156830
string GDS_START 146306
<< end >>
