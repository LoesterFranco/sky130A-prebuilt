magic
tech sky130A
magscale 1 2
timestamp 1604502729
<< locali >>
rect 970 424 1004 547
rect 970 390 1127 424
rect 574 310 647 356
rect 94 244 167 310
rect 121 236 167 244
rect 217 244 418 310
rect 460 270 647 310
rect 697 270 935 356
rect 969 270 1035 356
rect 217 236 263 244
rect 1081 236 1127 390
rect 511 202 1127 236
rect 511 170 749 202
rect 699 70 749 170
rect 937 70 1127 202
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 34 364 84 649
rect 124 378 190 596
rect 230 412 264 649
rect 304 378 370 596
rect 410 412 466 649
rect 506 424 540 596
rect 580 458 646 649
rect 684 581 1110 615
rect 684 458 751 581
rect 785 424 824 547
rect 506 390 824 424
rect 864 390 930 581
rect 1044 458 1110 581
rect 506 378 540 390
rect 124 344 540 378
rect 37 202 87 210
rect 381 202 447 210
rect 37 168 447 202
rect 37 70 87 168
rect 225 154 447 168
rect 123 17 189 134
rect 225 66 259 154
rect 597 120 663 136
rect 295 70 663 120
rect 783 17 903 168
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
rlabel locali s 574 310 647 356 6 A1
port 1 nsew signal input
rlabel locali s 460 270 647 310 6 A1
port 1 nsew signal input
rlabel locali s 217 244 418 310 6 A2
port 2 nsew signal input
rlabel locali s 217 236 263 244 6 A2
port 2 nsew signal input
rlabel locali s 121 236 167 244 6 A3
port 3 nsew signal input
rlabel locali s 94 244 167 310 6 A3
port 3 nsew signal input
rlabel locali s 697 270 935 356 6 B1
port 4 nsew signal input
rlabel locali s 969 270 1035 356 6 C1
port 5 nsew signal input
rlabel locali s 1081 236 1127 390 6 Y
port 6 nsew signal output
rlabel locali s 970 424 1004 547 6 Y
port 6 nsew signal output
rlabel locali s 970 390 1127 424 6 Y
port 6 nsew signal output
rlabel locali s 937 70 1127 202 6 Y
port 6 nsew signal output
rlabel locali s 699 70 749 170 6 Y
port 6 nsew signal output
rlabel locali s 511 202 1127 236 6 Y
port 6 nsew signal output
rlabel locali s 511 170 749 202 6 Y
port 6 nsew signal output
rlabel metal1 s 0 -49 1152 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 617 1152 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3699648
string GDS_START 3689400
<< end >>
