magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3157 561
rect 3191 527 3249 561
rect 3283 527 3341 561
rect 3375 527 3433 561
rect 3467 527 3525 561
rect 3559 527 3617 561
rect 3651 527 3709 561
rect 3743 527 3801 561
rect 3835 527 3893 561
rect 3927 527 3985 561
rect 4019 527 4077 561
rect 4111 527 4169 561
rect 4203 527 4261 561
rect 4295 527 4353 561
rect 4387 527 4445 561
rect 4479 527 4537 561
rect 4571 527 4629 561
rect 4663 527 4721 561
rect 4755 527 4813 561
rect 4847 527 4905 561
rect 4939 527 4997 561
rect 5031 527 5089 561
rect 5123 527 5152 561
rect 119 421 179 527
rect 113 367 179 421
rect 19 211 183 265
rect 611 293 677 527
rect 129 17 172 109
rect 558 205 625 259
rect 663 205 730 259
rect 1109 421 1169 527
rect 1109 367 1175 421
rect 1407 421 1467 527
rect 1401 367 1467 421
rect 1105 211 1269 265
rect 1307 211 1471 265
rect 1899 293 1965 527
rect 619 17 669 132
rect 1116 17 1159 109
rect 1417 17 1460 109
rect 1846 205 1913 259
rect 1951 205 2018 259
rect 2397 421 2457 527
rect 2397 367 2463 421
rect 2695 421 2755 527
rect 2689 367 2755 421
rect 2393 211 2557 265
rect 2595 211 2759 265
rect 3187 293 3253 527
rect 1907 17 1957 132
rect 2404 17 2447 109
rect 2705 17 2748 109
rect 3134 205 3201 259
rect 3239 205 3306 259
rect 3685 421 3745 527
rect 3685 367 3751 421
rect 3983 421 4043 527
rect 3977 367 4043 421
rect 3681 211 3845 265
rect 3883 211 4047 265
rect 4475 293 4541 527
rect 3195 17 3245 132
rect 3692 17 3735 109
rect 3993 17 4036 109
rect 4422 205 4489 259
rect 4527 205 4594 259
rect 4973 421 5033 527
rect 4973 367 5039 421
rect 4969 211 5133 265
rect 4483 17 4533 132
rect 4980 17 5023 109
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3341 17
rect 3375 -17 3433 17
rect 3467 -17 3525 17
rect 3559 -17 3617 17
rect 3651 -17 3709 17
rect 3743 -17 3801 17
rect 3835 -17 3893 17
rect 3927 -17 3985 17
rect 4019 -17 4077 17
rect 4111 -17 4169 17
rect 4203 -17 4261 17
rect 4295 -17 4353 17
rect 4387 -17 4445 17
rect 4479 -17 4537 17
rect 4571 -17 4629 17
rect 4663 -17 4721 17
rect 4755 -17 4813 17
rect 4847 -17 4905 17
rect 4939 -17 4997 17
rect 5031 -17 5089 17
rect 5123 -17 5152 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 2881 527 2915 561
rect 2973 527 3007 561
rect 3065 527 3099 561
rect 3157 527 3191 561
rect 3249 527 3283 561
rect 3341 527 3375 561
rect 3433 527 3467 561
rect 3525 527 3559 561
rect 3617 527 3651 561
rect 3709 527 3743 561
rect 3801 527 3835 561
rect 3893 527 3927 561
rect 3985 527 4019 561
rect 4077 527 4111 561
rect 4169 527 4203 561
rect 4261 527 4295 561
rect 4353 527 4387 561
rect 4445 527 4479 561
rect 4537 527 4571 561
rect 4629 527 4663 561
rect 4721 527 4755 561
rect 4813 527 4847 561
rect 4905 527 4939 561
rect 4997 527 5031 561
rect 5089 527 5123 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
rect 2881 -17 2915 17
rect 2973 -17 3007 17
rect 3065 -17 3099 17
rect 3157 -17 3191 17
rect 3249 -17 3283 17
rect 3341 -17 3375 17
rect 3433 -17 3467 17
rect 3525 -17 3559 17
rect 3617 -17 3651 17
rect 3709 -17 3743 17
rect 3801 -17 3835 17
rect 3893 -17 3927 17
rect 3985 -17 4019 17
rect 4077 -17 4111 17
rect 4169 -17 4203 17
rect 4261 -17 4295 17
rect 4353 -17 4387 17
rect 4445 -17 4479 17
rect 4537 -17 4571 17
rect 4629 -17 4663 17
rect 4721 -17 4755 17
rect 4813 -17 4847 17
rect 4905 -17 4939 17
rect 4997 -17 5031 17
rect 5089 -17 5123 17
<< obsli1 >>
rect 19 442 85 493
rect 19 333 79 442
rect 223 459 456 493
rect 223 333 257 459
rect 293 391 379 425
rect 293 357 305 391
rect 339 357 379 391
rect 293 351 379 357
rect 19 299 257 333
rect 206 177 267 185
rect 317 177 351 351
rect 422 329 456 459
rect 510 327 576 493
rect 490 295 576 327
rect 420 293 576 295
rect 712 327 778 493
rect 832 459 1065 493
rect 832 329 866 459
rect 909 391 995 425
rect 909 357 949 391
rect 983 357 995 391
rect 909 351 995 357
rect 712 295 798 327
rect 712 293 868 295
rect 420 261 524 293
rect 764 261 868 293
rect 420 241 503 261
rect 29 143 267 177
rect 29 51 95 143
rect 206 85 267 143
rect 301 119 367 177
rect 401 85 435 154
rect 469 151 503 241
rect 785 241 868 261
rect 785 151 819 241
rect 937 177 971 351
rect 1031 333 1065 459
rect 1203 442 1269 493
rect 1209 333 1269 442
rect 1031 299 1269 333
rect 1307 442 1373 493
rect 1307 333 1367 442
rect 1511 459 1744 493
rect 1511 333 1545 459
rect 1581 391 1667 425
rect 1581 357 1593 391
rect 1627 357 1667 391
rect 1581 351 1667 357
rect 1307 299 1545 333
rect 1021 177 1082 185
rect 1494 177 1555 185
rect 1605 177 1639 351
rect 1710 329 1744 459
rect 1798 327 1864 493
rect 1778 295 1864 327
rect 1708 293 1864 295
rect 2000 327 2066 493
rect 2120 459 2353 493
rect 2120 329 2154 459
rect 2197 391 2283 425
rect 2197 357 2237 391
rect 2271 357 2283 391
rect 2197 351 2283 357
rect 2000 295 2086 327
rect 2000 293 2156 295
rect 1708 261 1812 293
rect 2052 261 2156 293
rect 1708 241 1791 261
rect 469 117 585 151
rect 206 51 435 85
rect 535 66 585 117
rect 703 117 819 151
rect 703 66 753 117
rect 853 85 887 154
rect 921 119 987 177
rect 1021 143 1259 177
rect 1021 85 1082 143
rect 853 51 1082 85
rect 1193 51 1259 143
rect 1317 143 1555 177
rect 1317 51 1383 143
rect 1494 85 1555 143
rect 1589 119 1655 177
rect 1689 85 1723 154
rect 1757 151 1791 241
rect 2073 241 2156 261
rect 2073 151 2107 241
rect 2225 177 2259 351
rect 2319 333 2353 459
rect 2491 442 2557 493
rect 2497 333 2557 442
rect 2319 299 2557 333
rect 2595 442 2661 493
rect 2595 333 2655 442
rect 2799 459 3032 493
rect 2799 333 2833 459
rect 2869 391 2955 425
rect 2869 357 2881 391
rect 2915 357 2955 391
rect 2869 351 2955 357
rect 2595 299 2833 333
rect 2309 177 2370 185
rect 2782 177 2843 185
rect 2893 177 2927 351
rect 2998 329 3032 459
rect 3086 327 3152 493
rect 3066 295 3152 327
rect 2996 293 3152 295
rect 3288 327 3354 493
rect 3408 459 3641 493
rect 3408 329 3442 459
rect 3485 391 3571 425
rect 3485 357 3525 391
rect 3559 357 3571 391
rect 3485 351 3571 357
rect 3288 295 3374 327
rect 3288 293 3444 295
rect 2996 261 3100 293
rect 3340 261 3444 293
rect 2996 241 3079 261
rect 1757 117 1873 151
rect 1494 51 1723 85
rect 1823 66 1873 117
rect 1991 117 2107 151
rect 1991 66 2041 117
rect 2141 85 2175 154
rect 2209 119 2275 177
rect 2309 143 2547 177
rect 2309 85 2370 143
rect 2141 51 2370 85
rect 2481 51 2547 143
rect 2605 143 2843 177
rect 2605 51 2671 143
rect 2782 85 2843 143
rect 2877 119 2943 177
rect 2977 85 3011 154
rect 3045 151 3079 241
rect 3361 241 3444 261
rect 3361 151 3395 241
rect 3513 177 3547 351
rect 3607 333 3641 459
rect 3779 442 3845 493
rect 3785 333 3845 442
rect 3607 299 3845 333
rect 3883 442 3949 493
rect 3883 333 3943 442
rect 4087 459 4320 493
rect 4087 333 4121 459
rect 4157 391 4243 425
rect 4157 357 4169 391
rect 4203 357 4243 391
rect 4157 351 4243 357
rect 3883 299 4121 333
rect 3597 177 3658 185
rect 4070 177 4131 185
rect 4181 177 4215 351
rect 4286 329 4320 459
rect 4374 327 4440 493
rect 4354 295 4440 327
rect 4284 293 4440 295
rect 4576 327 4642 493
rect 4696 459 4929 493
rect 4696 329 4730 459
rect 4773 391 4859 425
rect 4773 357 4813 391
rect 4847 357 4859 391
rect 4773 351 4859 357
rect 4576 295 4662 327
rect 4576 293 4732 295
rect 4284 261 4388 293
rect 4628 261 4732 293
rect 4284 241 4367 261
rect 3045 117 3161 151
rect 2782 51 3011 85
rect 3111 66 3161 117
rect 3279 117 3395 151
rect 3279 66 3329 117
rect 3429 85 3463 154
rect 3497 119 3563 177
rect 3597 143 3835 177
rect 3597 85 3658 143
rect 3429 51 3658 85
rect 3769 51 3835 143
rect 3893 143 4131 177
rect 3893 51 3959 143
rect 4070 85 4131 143
rect 4165 119 4231 177
rect 4265 85 4299 154
rect 4333 151 4367 241
rect 4649 241 4732 261
rect 4649 151 4683 241
rect 4801 177 4835 351
rect 4895 333 4929 459
rect 5067 442 5133 493
rect 5073 333 5133 442
rect 4895 299 5133 333
rect 4885 177 4946 185
rect 4333 117 4449 151
rect 4070 51 4299 85
rect 4399 66 4449 117
rect 4567 117 4683 151
rect 4567 66 4617 117
rect 4717 85 4751 154
rect 4785 119 4851 177
rect 4885 143 5123 177
rect 4885 85 4946 143
rect 4717 51 4946 85
rect 5057 51 5123 143
<< obsli1c >>
rect 305 357 339 391
rect 949 357 983 391
rect 1593 357 1627 391
rect 2237 357 2271 391
rect 2881 357 2915 391
rect 3525 357 3559 391
rect 4169 357 4203 391
rect 4813 357 4847 391
<< metal1 >>
rect 0 561 5152 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3157 561
rect 3191 527 3249 561
rect 3283 527 3341 561
rect 3375 527 3433 561
rect 3467 527 3525 561
rect 3559 527 3617 561
rect 3651 527 3709 561
rect 3743 527 3801 561
rect 3835 527 3893 561
rect 3927 527 3985 561
rect 4019 527 4077 561
rect 4111 527 4169 561
rect 4203 527 4261 561
rect 4295 527 4353 561
rect 4387 527 4445 561
rect 4479 527 4537 561
rect 4571 527 4629 561
rect 4663 527 4721 561
rect 4755 527 4813 561
rect 4847 527 4905 561
rect 4939 527 4997 561
rect 5031 527 5089 561
rect 5123 527 5152 561
rect 0 496 5152 527
rect 293 391 351 397
rect 293 357 305 391
rect 339 388 351 391
rect 937 391 995 397
rect 937 388 949 391
rect 339 360 949 388
rect 339 357 351 360
rect 293 351 351 357
rect 937 357 949 360
rect 983 388 995 391
rect 1581 391 1639 397
rect 1581 388 1593 391
rect 983 360 1593 388
rect 983 357 995 360
rect 937 351 995 357
rect 1581 357 1593 360
rect 1627 388 1639 391
rect 2225 391 2283 397
rect 2225 388 2237 391
rect 1627 360 2237 388
rect 1627 357 1639 360
rect 1581 351 1639 357
rect 2225 357 2237 360
rect 2271 388 2283 391
rect 2869 391 2927 397
rect 2869 388 2881 391
rect 2271 360 2881 388
rect 2271 357 2283 360
rect 2225 351 2283 357
rect 2869 357 2881 360
rect 2915 388 2927 391
rect 3513 391 3571 397
rect 3513 388 3525 391
rect 2915 360 3525 388
rect 2915 357 2927 360
rect 2869 351 2927 357
rect 3513 357 3525 360
rect 3559 388 3571 391
rect 4157 391 4215 397
rect 4157 388 4169 391
rect 3559 360 4169 388
rect 3559 357 3571 360
rect 3513 351 3571 357
rect 4157 357 4169 360
rect 4203 388 4215 391
rect 4801 391 4859 397
rect 4801 388 4813 391
rect 4203 360 4813 388
rect 4203 357 4215 360
rect 4157 351 4215 357
rect 4801 357 4813 360
rect 4847 357 4859 391
rect 4801 351 4859 357
rect 0 17 5152 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3341 17
rect 3375 -17 3433 17
rect 3467 -17 3525 17
rect 3559 -17 3617 17
rect 3651 -17 3709 17
rect 3743 -17 3801 17
rect 3835 -17 3893 17
rect 3927 -17 3985 17
rect 4019 -17 4077 17
rect 4111 -17 4169 17
rect 4203 -17 4261 17
rect 4295 -17 4353 17
rect 4387 -17 4445 17
rect 4479 -17 4537 17
rect 4571 -17 4629 17
rect 4663 -17 4721 17
rect 4755 -17 4813 17
rect 4847 -17 4905 17
rect 4939 -17 4997 17
rect 5031 -17 5089 17
rect 5123 -17 5152 17
rect 0 -48 5152 -17
<< labels >>
rlabel locali s 19 211 183 265 6 D[0]
port 1 nsew signal input
rlabel locali s 1105 211 1269 265 6 D[1]
port 2 nsew signal input
rlabel locali s 1307 211 1471 265 6 D[2]
port 3 nsew signal input
rlabel locali s 2393 211 2557 265 6 D[3]
port 4 nsew signal input
rlabel locali s 2595 211 2759 265 6 D[4]
port 5 nsew signal input
rlabel locali s 3681 211 3845 265 6 D[5]
port 6 nsew signal input
rlabel locali s 3883 211 4047 265 6 D[6]
port 7 nsew signal input
rlabel locali s 4969 211 5133 265 6 D[7]
port 8 nsew signal input
rlabel locali s 558 205 625 259 6 S[0]
port 9 nsew signal input
rlabel locali s 663 205 730 259 6 S[1]
port 10 nsew signal input
rlabel locali s 1846 205 1913 259 6 S[2]
port 11 nsew signal input
rlabel locali s 1951 205 2018 259 6 S[3]
port 12 nsew signal input
rlabel locali s 3134 205 3201 259 6 S[4]
port 13 nsew signal input
rlabel locali s 3239 205 3306 259 6 S[5]
port 14 nsew signal input
rlabel locali s 4422 205 4489 259 6 S[6]
port 15 nsew signal input
rlabel locali s 4527 205 4594 259 6 S[7]
port 16 nsew signal input
rlabel metal1 s 4801 388 4859 397 6 Z
port 17 nsew signal output
rlabel metal1 s 4801 351 4859 360 6 Z
port 17 nsew signal output
rlabel metal1 s 4157 388 4215 397 6 Z
port 17 nsew signal output
rlabel metal1 s 4157 351 4215 360 6 Z
port 17 nsew signal output
rlabel metal1 s 3513 388 3571 397 6 Z
port 17 nsew signal output
rlabel metal1 s 3513 351 3571 360 6 Z
port 17 nsew signal output
rlabel metal1 s 2869 388 2927 397 6 Z
port 17 nsew signal output
rlabel metal1 s 2869 351 2927 360 6 Z
port 17 nsew signal output
rlabel metal1 s 2225 388 2283 397 6 Z
port 17 nsew signal output
rlabel metal1 s 2225 351 2283 360 6 Z
port 17 nsew signal output
rlabel metal1 s 1581 388 1639 397 6 Z
port 17 nsew signal output
rlabel metal1 s 1581 351 1639 360 6 Z
port 17 nsew signal output
rlabel metal1 s 937 388 995 397 6 Z
port 17 nsew signal output
rlabel metal1 s 937 351 995 360 6 Z
port 17 nsew signal output
rlabel metal1 s 293 388 351 397 6 Z
port 17 nsew signal output
rlabel metal1 s 293 360 4859 388 6 Z
port 17 nsew signal output
rlabel metal1 s 293 351 351 360 6 Z
port 17 nsew signal output
rlabel viali s 5089 -17 5123 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 4997 -17 5031 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 4905 -17 4939 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 4813 -17 4847 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 4721 -17 4755 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 4629 -17 4663 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 4537 -17 4571 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 4445 -17 4479 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 4353 -17 4387 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 4261 -17 4295 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 4169 -17 4203 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 4077 -17 4111 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 3985 -17 4019 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 3893 -17 3927 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 3801 -17 3835 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 3709 -17 3743 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 3617 -17 3651 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 3525 -17 3559 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 3433 -17 3467 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 3341 -17 3375 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 3249 -17 3283 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 3157 -17 3191 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 3065 -17 3099 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 2973 -17 3007 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 2881 -17 2915 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 2789 -17 2823 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 2697 -17 2731 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 2605 -17 2639 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 2513 -17 2547 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 2421 -17 2455 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 2329 -17 2363 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 2237 -17 2271 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 2145 -17 2179 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 2053 -17 2087 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 1961 -17 1995 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 1869 -17 1903 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 1777 -17 1811 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 1685 -17 1719 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 1593 -17 1627 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 1501 -17 1535 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 1409 -17 1443 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 1317 -17 1351 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 1225 -17 1259 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 1133 -17 1167 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 1041 -17 1075 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 949 -17 983 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 857 -17 891 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 765 -17 799 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 673 -17 707 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 581 -17 615 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 489 -17 523 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 397 -17 431 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 305 -17 339 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 213 -17 247 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 121 -17 155 17 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 29 -17 63 17 8 VGND
port 18 nsew ground bidirectional
rlabel locali s 4980 17 5023 109 6 VGND
port 18 nsew ground bidirectional
rlabel locali s 4483 17 4533 132 6 VGND
port 18 nsew ground bidirectional
rlabel locali s 3993 17 4036 109 6 VGND
port 18 nsew ground bidirectional
rlabel locali s 3692 17 3735 109 6 VGND
port 18 nsew ground bidirectional
rlabel locali s 3195 17 3245 132 6 VGND
port 18 nsew ground bidirectional
rlabel locali s 2705 17 2748 109 6 VGND
port 18 nsew ground bidirectional
rlabel locali s 2404 17 2447 109 6 VGND
port 18 nsew ground bidirectional
rlabel locali s 1907 17 1957 132 6 VGND
port 18 nsew ground bidirectional
rlabel locali s 1417 17 1460 109 6 VGND
port 18 nsew ground bidirectional
rlabel locali s 1116 17 1159 109 6 VGND
port 18 nsew ground bidirectional
rlabel locali s 619 17 669 132 6 VGND
port 18 nsew ground bidirectional
rlabel locali s 129 17 172 109 6 VGND
port 18 nsew ground bidirectional
rlabel locali s 0 -17 5152 17 8 VGND
port 18 nsew ground bidirectional
rlabel metal1 s 0 -48 5152 48 8 VGND
port 18 nsew ground bidirectional
rlabel viali s 5089 527 5123 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 4997 527 5031 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 4905 527 4939 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 4813 527 4847 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 4721 527 4755 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 4629 527 4663 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 4537 527 4571 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 4445 527 4479 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 4353 527 4387 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 4261 527 4295 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 4169 527 4203 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 4077 527 4111 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 3985 527 4019 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 3893 527 3927 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 3801 527 3835 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 3709 527 3743 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 3617 527 3651 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 3525 527 3559 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 3433 527 3467 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 3341 527 3375 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 3249 527 3283 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 3157 527 3191 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 3065 527 3099 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 2973 527 3007 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 2881 527 2915 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 2789 527 2823 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 2697 527 2731 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 2605 527 2639 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 2513 527 2547 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 2421 527 2455 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 2329 527 2363 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 2237 527 2271 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 2145 527 2179 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 2053 527 2087 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 1961 527 1995 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 1869 527 1903 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 1777 527 1811 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 1685 527 1719 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 1593 527 1627 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 1501 527 1535 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 1409 527 1443 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 1317 527 1351 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 1225 527 1259 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 1133 527 1167 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 1041 527 1075 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 949 527 983 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 857 527 891 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 765 527 799 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 673 527 707 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 581 527 615 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 489 527 523 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 397 527 431 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 305 527 339 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 213 527 247 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 121 527 155 561 6 VPWR
port 19 nsew power bidirectional
rlabel viali s 29 527 63 561 6 VPWR
port 19 nsew power bidirectional
rlabel locali s 4973 421 5033 527 6 VPWR
port 19 nsew power bidirectional
rlabel locali s 4973 367 5039 421 6 VPWR
port 19 nsew power bidirectional
rlabel locali s 4475 293 4541 527 6 VPWR
port 19 nsew power bidirectional
rlabel locali s 3983 421 4043 527 6 VPWR
port 19 nsew power bidirectional
rlabel locali s 3977 367 4043 421 6 VPWR
port 19 nsew power bidirectional
rlabel locali s 3685 421 3745 527 6 VPWR
port 19 nsew power bidirectional
rlabel locali s 3685 367 3751 421 6 VPWR
port 19 nsew power bidirectional
rlabel locali s 3187 293 3253 527 6 VPWR
port 19 nsew power bidirectional
rlabel locali s 2695 421 2755 527 6 VPWR
port 19 nsew power bidirectional
rlabel locali s 2689 367 2755 421 6 VPWR
port 19 nsew power bidirectional
rlabel locali s 2397 421 2457 527 6 VPWR
port 19 nsew power bidirectional
rlabel locali s 2397 367 2463 421 6 VPWR
port 19 nsew power bidirectional
rlabel locali s 1899 293 1965 527 6 VPWR
port 19 nsew power bidirectional
rlabel locali s 1407 421 1467 527 6 VPWR
port 19 nsew power bidirectional
rlabel locali s 1401 367 1467 421 6 VPWR
port 19 nsew power bidirectional
rlabel locali s 1109 421 1169 527 6 VPWR
port 19 nsew power bidirectional
rlabel locali s 1109 367 1175 421 6 VPWR
port 19 nsew power bidirectional
rlabel locali s 611 293 677 527 6 VPWR
port 19 nsew power bidirectional
rlabel locali s 119 421 179 527 6 VPWR
port 19 nsew power bidirectional
rlabel locali s 113 367 179 421 6 VPWR
port 19 nsew power bidirectional
rlabel locali s 0 527 5152 561 6 VPWR
port 19 nsew power bidirectional
rlabel metal1 s 0 496 5152 592 6 VPWR
port 19 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 5152 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2893436
string GDS_START 2834862
<< end >>
