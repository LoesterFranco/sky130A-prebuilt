magic
tech sky130A
magscale 1 2
timestamp 1604502711
<< locali >>
rect 232 425 351 493
rect 17 199 130 345
rect 232 119 266 425
rect 300 153 351 391
rect 232 51 351 119
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 17 413 80 493
rect 114 447 198 527
rect 17 379 198 413
rect 164 165 198 379
rect 17 131 198 165
rect 17 51 72 131
rect 106 17 198 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
<< metal1 >>
rect 0 561 368 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 0 496 368 527
rect 0 17 368 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
rect 0 -48 368 -17
<< labels >>
rlabel locali s 300 153 351 391 6 A
port 1 nsew signal input
rlabel locali s 17 199 130 345 6 TE_B
port 2 nsew signal input
rlabel locali s 232 425 351 493 6 Z
port 3 nsew signal output
rlabel locali s 232 119 266 425 6 Z
port 3 nsew signal output
rlabel locali s 232 51 351 119 6 Z
port 3 nsew signal output
rlabel metal1 s 0 -48 368 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 368 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 368 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2888674
string GDS_START 2884432
<< end >>
