magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 552 561
rect 142 299 192 527
rect 226 333 292 493
rect 326 367 383 527
rect 417 333 535 493
rect 226 299 535 333
rect 85 199 155 265
rect 193 199 247 265
rect 285 199 351 265
rect 477 97 535 299
rect 142 17 208 97
rect 417 51 535 97
rect 0 -17 552 17
<< obsli1 >>
rect 17 319 102 385
rect 17 165 51 319
rect 409 165 443 265
rect 17 131 443 165
rect 17 89 102 131
<< metal1 >>
rect 0 496 552 592
rect 0 -48 552 48
<< labels >>
rlabel locali s 85 199 155 265 6 A_N
port 1 nsew signal input
rlabel locali s 285 199 351 265 6 B
port 2 nsew signal input
rlabel locali s 193 199 247 265 6 C
port 3 nsew signal input
rlabel locali s 477 97 535 299 6 Y
port 4 nsew signal output
rlabel locali s 417 333 535 493 6 Y
port 4 nsew signal output
rlabel locali s 417 51 535 97 6 Y
port 4 nsew signal output
rlabel locali s 226 333 292 493 6 Y
port 4 nsew signal output
rlabel locali s 226 299 535 333 6 Y
port 4 nsew signal output
rlabel locali s 142 17 208 97 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 552 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 552 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 326 367 383 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 142 299 192 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 552 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 552 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 552 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1817266
string GDS_START 1811732
<< end >>
