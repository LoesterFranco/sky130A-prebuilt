magic
tech sky130A
magscale 1 2
timestamp 1601050056
<< nwell >>
rect -38 332 2918 704
rect 1481 311 1694 332
<< pwell >>
rect 0 0 2880 49
<< scpmos >>
rect 83 464 119 592
rect 173 464 209 592
rect 257 464 293 592
rect 383 464 419 592
rect 467 464 503 592
rect 685 368 721 592
rect 775 368 811 592
rect 979 463 1015 547
rect 1100 478 1136 562
rect 1204 463 1240 547
rect 1341 463 1377 547
rect 1459 463 1495 547
rect 1567 347 1603 547
rect 1762 374 1798 458
rect 1870 374 1906 574
rect 2070 508 2106 592
rect 2160 508 2196 592
rect 2360 508 2396 592
rect 2461 368 2497 592
rect 2661 403 2697 571
rect 2762 368 2798 592
<< nmoslvt >>
rect 84 74 114 158
rect 198 74 228 158
rect 276 74 306 158
rect 362 74 392 158
rect 440 74 470 158
rect 651 74 681 222
rect 751 74 781 222
rect 965 74 995 158
rect 1085 74 1115 158
rect 1163 74 1193 158
rect 1381 74 1411 158
rect 1459 74 1489 158
rect 1654 74 1684 202
rect 1732 74 1762 202
rect 1846 74 1876 158
rect 1924 74 1954 158
rect 2032 74 2062 158
rect 2188 74 2218 158
rect 2400 74 2430 222
rect 2613 112 2643 222
rect 2766 74 2796 222
<< ndiff >>
rect 594 186 651 222
rect 27 133 84 158
rect 27 99 39 133
rect 73 99 84 133
rect 27 74 84 99
rect 114 130 198 158
rect 114 96 139 130
rect 173 96 198 130
rect 114 74 198 96
rect 228 74 276 158
rect 306 133 362 158
rect 306 99 317 133
rect 351 99 362 133
rect 306 74 362 99
rect 392 74 440 158
rect 470 127 527 158
rect 470 93 481 127
rect 515 93 527 127
rect 470 74 527 93
rect 594 152 606 186
rect 640 152 651 186
rect 594 118 651 152
rect 594 84 606 118
rect 640 84 651 118
rect 594 74 651 84
rect 681 186 751 222
rect 681 152 692 186
rect 726 152 751 186
rect 681 118 751 152
rect 681 84 692 118
rect 726 84 751 118
rect 681 74 751 84
rect 781 186 838 222
rect 781 152 792 186
rect 826 152 838 186
rect 781 118 838 152
rect 781 84 792 118
rect 826 84 838 118
rect 781 74 838 84
rect 892 169 950 181
rect 892 135 904 169
rect 938 158 950 169
rect 1504 158 1654 202
rect 938 135 965 158
rect 892 74 965 135
rect 995 133 1085 158
rect 995 99 1040 133
rect 1074 99 1085 133
rect 995 74 1085 99
rect 1115 74 1163 158
rect 1193 113 1270 158
rect 1193 79 1222 113
rect 1256 79 1270 113
rect 1193 74 1270 79
rect 1324 125 1381 158
rect 1324 91 1336 125
rect 1370 91 1381 125
rect 1324 74 1381 91
rect 1411 74 1459 158
rect 1489 131 1654 158
rect 1489 97 1500 131
rect 1534 97 1609 131
rect 1643 97 1654 131
rect 1489 74 1654 97
rect 1684 74 1732 202
rect 1762 188 1819 202
rect 1762 154 1773 188
rect 1807 158 1819 188
rect 2329 210 2400 222
rect 2329 176 2341 210
rect 2375 176 2400 210
rect 1807 154 1846 158
rect 1762 120 1846 154
rect 1762 86 1801 120
rect 1835 86 1846 120
rect 1762 74 1846 86
rect 1876 74 1924 158
rect 1954 74 2032 158
rect 2062 120 2188 158
rect 2062 86 2073 120
rect 2107 86 2143 120
rect 2177 86 2188 120
rect 2062 74 2188 86
rect 2218 133 2275 158
rect 2218 99 2229 133
rect 2263 99 2275 133
rect 2218 74 2275 99
rect 2329 120 2400 176
rect 2329 86 2341 120
rect 2375 86 2400 120
rect 2329 74 2400 86
rect 2430 210 2487 222
rect 2430 176 2441 210
rect 2475 176 2487 210
rect 2430 120 2487 176
rect 2430 86 2441 120
rect 2475 86 2487 120
rect 2556 184 2613 222
rect 2556 150 2568 184
rect 2602 150 2613 184
rect 2556 112 2613 150
rect 2643 194 2766 222
rect 2643 160 2707 194
rect 2741 160 2766 194
rect 2643 120 2766 160
rect 2643 112 2707 120
rect 2695 86 2707 112
rect 2741 86 2766 120
rect 2430 74 2487 86
rect 2695 74 2766 86
rect 2796 210 2853 222
rect 2796 176 2807 210
rect 2841 176 2853 210
rect 2796 120 2853 176
rect 2796 86 2807 120
rect 2841 86 2853 120
rect 2796 74 2853 86
rect 1208 67 1270 74
<< pdiff >>
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 510 83 546
rect 27 476 39 510
rect 73 476 83 510
rect 27 464 83 476
rect 119 578 173 592
rect 119 544 129 578
rect 163 544 173 578
rect 119 464 173 544
rect 209 464 257 592
rect 293 576 383 592
rect 293 542 321 576
rect 355 542 383 576
rect 293 464 383 542
rect 419 464 467 592
rect 503 582 565 592
rect 503 548 514 582
rect 548 548 565 582
rect 503 464 565 548
rect 630 414 685 592
rect 630 380 641 414
rect 675 380 685 414
rect 630 368 685 380
rect 721 573 775 592
rect 721 539 731 573
rect 765 539 775 573
rect 721 368 775 539
rect 811 570 865 592
rect 811 536 821 570
rect 855 536 865 570
rect 811 368 865 536
rect 1712 588 1766 600
rect 1030 547 1100 562
rect 925 520 979 547
rect 925 486 935 520
rect 969 486 979 520
rect 925 463 979 486
rect 1015 527 1100 547
rect 1015 493 1040 527
rect 1074 493 1100 527
rect 1015 478 1100 493
rect 1136 547 1186 562
rect 1712 554 1722 588
rect 1756 554 1766 588
rect 1136 478 1204 547
rect 1015 463 1085 478
rect 1154 463 1204 478
rect 1240 535 1341 547
rect 1240 501 1251 535
rect 1285 501 1341 535
rect 1240 463 1341 501
rect 1377 520 1459 547
rect 1377 486 1387 520
rect 1421 486 1459 520
rect 1377 463 1459 486
rect 1495 522 1567 547
rect 1495 488 1523 522
rect 1557 488 1567 522
rect 1495 463 1567 488
rect 1517 347 1567 463
rect 1603 521 1658 547
rect 1603 487 1613 521
rect 1647 487 1658 521
rect 1603 347 1658 487
rect 1712 542 1766 554
rect 1712 458 1742 542
rect 1820 458 1870 574
rect 1712 374 1762 458
rect 1798 420 1870 458
rect 1798 386 1825 420
rect 1859 386 1870 420
rect 1798 374 1870 386
rect 1906 519 1961 574
rect 1906 485 1916 519
rect 1950 485 1961 519
rect 2015 567 2070 592
rect 2015 533 2026 567
rect 2060 533 2070 567
rect 2015 508 2070 533
rect 2106 567 2160 592
rect 2106 533 2116 567
rect 2150 533 2160 567
rect 2106 508 2160 533
rect 2196 567 2251 592
rect 2196 533 2206 567
rect 2240 533 2251 567
rect 2196 508 2251 533
rect 2305 567 2360 592
rect 2305 533 2316 567
rect 2350 533 2360 567
rect 2305 508 2360 533
rect 2396 567 2461 592
rect 2396 533 2406 567
rect 2440 533 2461 567
rect 2396 508 2461 533
rect 1906 374 1961 485
rect 2411 368 2461 508
rect 2497 580 2552 592
rect 2497 546 2507 580
rect 2541 546 2552 580
rect 2712 571 2762 592
rect 2497 497 2552 546
rect 2497 463 2507 497
rect 2541 463 2552 497
rect 2497 414 2552 463
rect 2497 380 2507 414
rect 2541 380 2552 414
rect 2606 559 2661 571
rect 2606 525 2617 559
rect 2651 525 2661 559
rect 2606 449 2661 525
rect 2606 415 2617 449
rect 2651 415 2661 449
rect 2606 403 2661 415
rect 2697 559 2762 571
rect 2697 525 2707 559
rect 2741 525 2762 559
rect 2697 449 2762 525
rect 2697 415 2707 449
rect 2741 415 2762 449
rect 2697 403 2762 415
rect 2497 368 2552 380
rect 2712 368 2762 403
rect 2798 580 2853 592
rect 2798 546 2808 580
rect 2842 546 2853 580
rect 2798 497 2853 546
rect 2798 463 2808 497
rect 2842 463 2853 497
rect 2798 414 2853 463
rect 2798 380 2808 414
rect 2842 380 2853 414
rect 2798 368 2853 380
<< ndiffc >>
rect 39 99 73 133
rect 139 96 173 130
rect 317 99 351 133
rect 481 93 515 127
rect 606 152 640 186
rect 606 84 640 118
rect 692 152 726 186
rect 692 84 726 118
rect 792 152 826 186
rect 792 84 826 118
rect 904 135 938 169
rect 1040 99 1074 133
rect 1222 79 1256 113
rect 1336 91 1370 125
rect 1500 97 1534 131
rect 1609 97 1643 131
rect 1773 154 1807 188
rect 2341 176 2375 210
rect 1801 86 1835 120
rect 2073 86 2107 120
rect 2143 86 2177 120
rect 2229 99 2263 133
rect 2341 86 2375 120
rect 2441 176 2475 210
rect 2441 86 2475 120
rect 2568 150 2602 184
rect 2707 160 2741 194
rect 2707 86 2741 120
rect 2807 176 2841 210
rect 2807 86 2841 120
<< pdiffc >>
rect 39 546 73 580
rect 39 476 73 510
rect 129 544 163 578
rect 321 542 355 576
rect 514 548 548 582
rect 641 380 675 414
rect 731 539 765 573
rect 821 536 855 570
rect 935 486 969 520
rect 1040 493 1074 527
rect 1722 554 1756 588
rect 1251 501 1285 535
rect 1387 486 1421 520
rect 1523 488 1557 522
rect 1613 487 1647 521
rect 1825 386 1859 420
rect 1916 485 1950 519
rect 2026 533 2060 567
rect 2116 533 2150 567
rect 2206 533 2240 567
rect 2316 533 2350 567
rect 2406 533 2440 567
rect 2507 546 2541 580
rect 2507 463 2541 497
rect 2507 380 2541 414
rect 2617 525 2651 559
rect 2617 415 2651 449
rect 2707 525 2741 559
rect 2707 415 2741 449
rect 2808 546 2842 580
rect 2808 463 2842 497
rect 2808 380 2842 414
<< poly >>
rect 83 592 119 618
rect 173 592 209 618
rect 257 592 293 618
rect 383 592 419 618
rect 467 592 503 618
rect 685 592 721 618
rect 775 592 811 618
rect 880 615 1906 645
rect 83 370 119 464
rect 173 418 209 464
rect 257 424 293 464
rect 383 432 419 464
rect 179 370 209 418
rect 83 354 209 370
rect 251 408 317 424
rect 251 374 267 408
rect 301 374 317 408
rect 251 358 317 374
rect 359 416 425 432
rect 467 430 503 464
rect 359 382 375 416
rect 409 382 425 416
rect 359 366 425 382
rect 473 414 566 430
rect 473 380 516 414
rect 550 380 566 414
rect 83 320 117 354
rect 151 340 209 354
rect 151 320 167 340
rect 83 304 167 320
rect 84 158 114 304
rect 162 240 228 256
rect 162 206 178 240
rect 212 206 228 240
rect 162 190 228 206
rect 198 158 228 190
rect 276 158 306 358
rect 473 346 566 380
rect 685 352 721 368
rect 359 302 425 318
rect 359 268 375 302
rect 409 268 425 302
rect 359 252 425 268
rect 473 312 516 346
rect 550 312 566 346
rect 473 278 566 312
rect 679 322 721 352
rect 679 310 709 322
rect 362 158 392 252
rect 473 244 516 278
rect 550 244 566 278
rect 643 294 709 310
rect 643 260 659 294
rect 693 260 709 294
rect 775 310 811 368
rect 880 310 910 615
rect 979 547 1015 573
rect 1100 562 1136 615
rect 1204 547 1240 573
rect 1341 547 1377 573
rect 1459 547 1495 573
rect 1567 547 1603 573
rect 1870 574 1906 615
rect 2070 592 2106 618
rect 2160 592 2196 618
rect 2360 592 2396 618
rect 2461 592 2497 618
rect 979 408 1015 463
rect 1100 452 1136 478
rect 775 294 910 310
rect 775 274 793 294
rect 643 244 709 260
rect 751 260 793 274
rect 827 260 910 294
rect 952 392 1018 408
rect 952 358 968 392
rect 1002 368 1018 392
rect 1085 388 1162 404
rect 1085 368 1112 388
rect 1002 358 1112 368
rect 952 354 1112 358
rect 1146 354 1162 388
rect 1204 393 1240 463
rect 1204 377 1276 393
rect 1204 363 1226 377
rect 952 338 1162 354
rect 1210 343 1226 363
rect 1260 343 1276 377
rect 952 324 1018 338
rect 952 290 968 324
rect 1002 290 1018 324
rect 952 274 1018 290
rect 751 244 910 260
rect 473 228 566 244
rect 473 203 503 228
rect 651 222 681 244
rect 751 222 781 244
rect 880 226 910 244
rect 440 173 503 203
rect 440 158 470 173
rect 880 196 995 226
rect 965 158 995 196
rect 1085 158 1115 338
rect 1210 327 1276 343
rect 1210 246 1240 327
rect 1341 304 1377 463
rect 1459 315 1495 463
rect 1762 458 1798 484
rect 2070 463 2106 508
rect 1976 433 2106 463
rect 1762 359 1798 374
rect 1870 359 1906 374
rect 1345 288 1411 304
rect 1345 254 1361 288
rect 1395 254 1411 288
rect 1163 230 1297 246
rect 1345 238 1411 254
rect 1163 196 1179 230
rect 1213 196 1247 230
rect 1281 196 1297 230
rect 1163 180 1297 196
rect 1163 158 1193 180
rect 1381 158 1411 238
rect 1459 299 1525 315
rect 1459 265 1475 299
rect 1509 265 1525 299
rect 1459 249 1525 265
rect 1567 290 1603 347
rect 1732 320 1798 359
rect 1567 274 1684 290
rect 1459 158 1489 249
rect 1567 240 1583 274
rect 1617 240 1684 274
rect 1567 224 1684 240
rect 1654 202 1684 224
rect 1732 286 1748 320
rect 1782 286 1798 320
rect 1732 270 1798 286
rect 1846 329 1906 359
rect 1732 202 1762 270
rect 1846 158 1876 329
rect 1976 281 2006 433
rect 2160 385 2196 508
rect 2360 401 2396 508
rect 2360 394 2390 401
rect 1924 251 2006 281
rect 2110 369 2196 385
rect 2110 335 2133 369
rect 2167 355 2196 369
rect 2245 378 2390 394
rect 2167 335 2190 355
rect 2110 301 2190 335
rect 2110 267 2133 301
rect 2167 267 2190 301
rect 2110 251 2190 267
rect 2245 344 2261 378
rect 2295 344 2329 378
rect 2363 353 2390 378
rect 2661 571 2697 597
rect 2762 592 2798 618
rect 2661 388 2697 403
rect 2461 353 2497 368
rect 2613 358 2697 388
rect 2613 353 2643 358
rect 2363 344 2643 353
rect 2245 323 2643 344
rect 1924 230 1990 251
rect 1924 196 1940 230
rect 1974 196 1990 230
rect 2110 203 2140 251
rect 2245 203 2275 323
rect 2400 222 2430 323
rect 2613 222 2643 323
rect 2762 310 2798 368
rect 2691 294 2798 310
rect 2691 260 2707 294
rect 2741 260 2798 294
rect 2691 244 2798 260
rect 2766 222 2796 244
rect 1924 173 1990 196
rect 2032 173 2140 203
rect 2188 173 2275 203
rect 1924 158 1954 173
rect 2032 158 2062 173
rect 2188 158 2218 173
rect 2613 86 2643 112
rect 84 48 114 74
rect 198 48 228 74
rect 276 48 306 74
rect 362 48 392 74
rect 440 48 470 74
rect 651 48 681 74
rect 751 48 781 74
rect 965 48 995 74
rect 1085 48 1115 74
rect 1163 48 1193 74
rect 1381 48 1411 74
rect 1459 48 1489 74
rect 1654 48 1684 74
rect 1732 48 1762 74
rect 1846 48 1876 74
rect 1924 48 1954 74
rect 2032 48 2062 74
rect 2188 48 2218 74
rect 2400 48 2430 74
rect 2766 48 2796 74
<< polycont >>
rect 267 374 301 408
rect 375 382 409 416
rect 516 380 550 414
rect 117 320 151 354
rect 178 206 212 240
rect 375 268 409 302
rect 516 312 550 346
rect 516 244 550 278
rect 659 260 693 294
rect 793 260 827 294
rect 968 358 1002 392
rect 1112 354 1146 388
rect 1226 343 1260 377
rect 968 290 1002 324
rect 1361 254 1395 288
rect 1179 196 1213 230
rect 1247 196 1281 230
rect 1475 265 1509 299
rect 1583 240 1617 274
rect 1748 286 1782 320
rect 2133 335 2167 369
rect 2133 267 2167 301
rect 2261 344 2295 378
rect 2329 344 2363 378
rect 1940 196 1974 230
rect 2707 260 2741 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2880 683
rect 23 580 73 596
rect 23 546 39 580
rect 23 510 73 546
rect 113 578 179 649
rect 113 544 129 578
rect 163 544 179 578
rect 113 526 179 544
rect 287 576 389 592
rect 287 542 321 576
rect 355 560 389 576
rect 511 582 564 649
rect 355 542 477 560
rect 287 526 477 542
rect 511 548 514 582
rect 548 548 564 582
rect 511 532 564 548
rect 715 573 781 649
rect 715 539 731 573
rect 765 539 781 573
rect 715 532 781 539
rect 821 581 1162 615
rect 821 570 871 581
rect 855 536 871 570
rect 23 476 39 510
rect 443 498 477 526
rect 821 510 871 536
rect 918 520 985 547
rect 73 476 409 492
rect 23 458 409 476
rect 23 256 67 458
rect 217 408 317 424
rect 217 374 267 408
rect 301 374 317 408
rect 101 354 167 370
rect 217 358 317 374
rect 359 416 409 458
rect 359 382 375 416
rect 359 366 409 382
rect 443 476 759 498
rect 918 486 935 520
rect 969 486 985 520
rect 918 476 985 486
rect 443 464 985 476
rect 1024 527 1090 547
rect 1024 493 1040 527
rect 1074 493 1090 527
rect 1024 474 1090 493
rect 101 320 117 354
rect 151 324 167 354
rect 151 320 409 324
rect 101 302 409 320
rect 101 290 375 302
rect 359 268 375 290
rect 23 240 228 256
rect 359 252 409 268
rect 23 206 178 240
rect 212 206 228 240
rect 443 218 477 464
rect 725 442 985 464
rect 511 414 553 430
rect 511 380 516 414
rect 550 380 553 414
rect 511 346 553 380
rect 511 312 516 346
rect 550 312 553 346
rect 511 278 553 312
rect 511 244 516 278
rect 550 244 553 278
rect 511 228 553 244
rect 587 414 691 430
rect 587 380 641 414
rect 675 398 691 414
rect 675 380 843 398
rect 587 364 843 380
rect 23 190 228 206
rect 23 133 89 190
rect 301 184 477 218
rect 587 202 621 364
rect 655 294 743 310
rect 655 260 659 294
rect 693 260 743 294
rect 655 236 743 260
rect 777 294 843 364
rect 777 260 793 294
rect 827 260 843 294
rect 777 244 843 260
rect 587 186 640 202
rect 23 99 39 133
rect 73 99 89 133
rect 23 70 89 99
rect 123 130 189 156
rect 123 96 139 130
rect 173 96 189 130
rect 123 17 189 96
rect 301 133 367 184
rect 587 152 606 186
rect 301 99 317 133
rect 351 99 367 133
rect 301 70 367 99
rect 465 127 531 150
rect 465 93 481 127
rect 515 93 531 127
rect 465 17 531 93
rect 587 118 640 152
rect 587 84 606 118
rect 587 68 640 84
rect 676 186 742 202
rect 676 152 692 186
rect 726 152 742 186
rect 676 118 742 152
rect 676 84 692 118
rect 726 84 742 118
rect 676 17 742 84
rect 776 186 842 202
rect 776 152 792 186
rect 826 152 842 186
rect 776 118 842 152
rect 884 185 918 442
rect 952 392 1006 408
rect 952 358 968 392
rect 1002 358 1006 392
rect 952 324 1006 358
rect 952 290 968 324
rect 1002 290 1006 324
rect 952 274 1006 290
rect 884 169 938 185
rect 884 135 904 169
rect 884 119 938 135
rect 776 84 792 118
rect 826 85 842 118
rect 972 85 1006 274
rect 826 84 1006 85
rect 776 51 1006 84
rect 1040 304 1074 474
rect 1128 451 1162 581
rect 1235 535 1285 649
rect 1235 501 1251 535
rect 1235 485 1285 501
rect 1319 581 1489 615
rect 1319 451 1353 581
rect 1128 417 1353 451
rect 1387 520 1421 547
rect 1128 404 1162 417
rect 1108 388 1162 404
rect 1108 354 1112 388
rect 1146 354 1162 388
rect 1387 383 1421 486
rect 1455 424 1489 581
rect 1523 522 1557 649
rect 1706 588 2076 615
rect 1706 554 1722 588
rect 1756 581 2076 588
rect 1756 554 1772 581
rect 1523 459 1557 488
rect 1597 521 1663 551
rect 1706 538 1772 554
rect 2010 567 2076 581
rect 1597 487 1613 521
rect 1647 504 1663 521
rect 1916 519 1966 547
rect 1647 487 1916 504
rect 1597 485 1916 487
rect 1950 485 1966 519
rect 2010 533 2026 567
rect 2060 533 2076 567
rect 2010 504 2076 533
rect 2116 567 2150 649
rect 2116 504 2150 533
rect 2190 567 2256 596
rect 2190 533 2206 567
rect 2240 533 2256 567
rect 2190 504 2256 533
rect 1597 470 1966 485
rect 1597 458 1663 470
rect 1916 458 1966 470
rect 2222 453 2256 504
rect 1809 424 1876 436
rect 2000 424 2256 453
rect 2300 567 2350 596
rect 2300 533 2316 567
rect 2300 470 2350 533
rect 2390 567 2456 649
rect 2390 533 2406 567
rect 2440 533 2456 567
rect 2390 504 2456 533
rect 2490 580 2541 596
rect 2490 546 2507 580
rect 2490 497 2541 546
rect 2300 436 2447 470
rect 1455 390 1766 424
rect 1108 338 1162 354
rect 1210 377 1421 383
rect 1210 343 1226 377
rect 1260 343 1421 377
rect 1210 338 1421 343
rect 1459 350 1525 356
rect 1459 316 1471 350
rect 1505 316 1525 350
rect 1040 288 1422 304
rect 1040 270 1361 288
rect 1040 133 1090 270
rect 1345 254 1361 270
rect 1395 254 1422 288
rect 1345 238 1422 254
rect 1459 299 1525 316
rect 1459 265 1475 299
rect 1509 265 1525 299
rect 1732 336 1766 390
rect 1809 420 2256 424
rect 1809 386 1825 420
rect 1859 419 2256 420
rect 1859 390 2034 419
rect 2222 394 2256 419
rect 1859 386 1876 390
rect 1809 370 1876 386
rect 1732 320 1798 336
rect 1459 249 1525 265
rect 1567 274 1633 290
rect 1163 230 1297 236
rect 1163 196 1179 230
rect 1213 196 1247 230
rect 1281 196 1297 230
rect 1163 181 1297 196
rect 1388 215 1422 238
rect 1567 240 1583 274
rect 1617 240 1633 274
rect 1732 286 1748 320
rect 1782 286 1798 320
rect 1732 270 1798 286
rect 1567 215 1633 240
rect 1388 181 1633 215
rect 1842 210 1876 370
rect 2117 369 2183 385
rect 2117 356 2133 369
rect 1945 350 2133 356
rect 1945 316 1951 350
rect 1985 335 2133 350
rect 2167 335 2183 369
rect 1985 316 2183 335
rect 2222 378 2379 394
rect 2222 344 2261 378
rect 2295 344 2329 378
rect 2363 344 2379 378
rect 2222 328 2379 344
rect 1945 310 2183 316
rect 2117 301 2183 310
rect 2117 267 2133 301
rect 2167 267 2183 301
rect 2413 294 2447 436
rect 2117 251 2183 267
rect 2245 260 2447 294
rect 2490 463 2507 497
rect 2490 414 2541 463
rect 2490 380 2507 414
rect 2490 364 2541 380
rect 2601 559 2651 575
rect 2601 525 2617 559
rect 2601 449 2651 525
rect 2601 415 2617 449
rect 1757 188 1876 210
rect 1163 147 1354 181
rect 1757 154 1773 188
rect 1807 154 1876 188
rect 1924 230 1990 246
rect 1924 196 1940 230
rect 1974 214 1990 230
rect 2245 214 2279 260
rect 2490 226 2524 364
rect 2601 310 2651 415
rect 2691 559 2757 649
rect 2691 525 2707 559
rect 2741 525 2757 559
rect 2691 449 2757 525
rect 2691 415 2707 449
rect 2741 415 2757 449
rect 2691 399 2757 415
rect 2791 580 2858 596
rect 2791 546 2808 580
rect 2842 546 2858 580
rect 2791 497 2858 546
rect 2791 463 2808 497
rect 2842 463 2858 497
rect 2791 414 2858 463
rect 2791 380 2808 414
rect 2842 380 2858 414
rect 2601 294 2757 310
rect 2601 260 2707 294
rect 2741 260 2757 294
rect 2601 244 2757 260
rect 2601 226 2651 244
rect 1974 196 2279 214
rect 1924 180 2279 196
rect 1074 99 1090 133
rect 1320 125 1386 147
rect 1040 70 1090 99
rect 1204 79 1222 113
rect 1256 79 1274 113
rect 1204 17 1274 79
rect 1320 91 1336 125
rect 1370 91 1386 125
rect 1320 70 1386 91
rect 1500 131 1659 147
rect 1534 97 1609 131
rect 1643 97 1659 131
rect 1500 17 1659 97
rect 1757 120 1876 154
rect 1757 86 1801 120
rect 1835 86 1876 120
rect 1757 70 1876 86
rect 2057 120 2179 136
rect 2057 86 2073 120
rect 2107 86 2143 120
rect 2177 86 2179 120
rect 2057 17 2179 86
rect 2213 133 2279 180
rect 2213 99 2229 133
rect 2263 99 2279 133
rect 2213 70 2279 99
rect 2325 210 2391 226
rect 2325 176 2341 210
rect 2375 176 2391 210
rect 2325 120 2391 176
rect 2325 86 2341 120
rect 2375 86 2391 120
rect 2325 17 2391 86
rect 2425 210 2524 226
rect 2425 176 2441 210
rect 2475 176 2524 210
rect 2425 120 2524 176
rect 2425 86 2441 120
rect 2475 86 2524 120
rect 2568 184 2651 226
rect 2791 210 2858 380
rect 2602 150 2651 184
rect 2568 108 2651 150
rect 2691 194 2757 210
rect 2691 160 2707 194
rect 2741 160 2757 194
rect 2691 120 2757 160
rect 2425 70 2524 86
rect 2691 86 2707 120
rect 2741 86 2757 120
rect 2691 17 2757 86
rect 2791 176 2807 210
rect 2841 176 2858 210
rect 2791 120 2858 176
rect 2791 86 2807 120
rect 2841 86 2858 120
rect 2791 70 2858 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2880 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 1471 316 1505 350
rect 1951 316 1985 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
<< metal1 >>
rect 0 683 2880 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2880 683
rect 0 617 2880 649
rect 1459 350 1517 356
rect 1459 316 1471 350
rect 1505 347 1517 350
rect 1939 350 1997 356
rect 1939 347 1951 350
rect 1505 319 1951 347
rect 1505 316 1517 319
rect 1459 310 1517 316
rect 1939 316 1951 319
rect 1985 316 1997 350
rect 1939 310 1997 316
rect 0 17 2880 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2880 17
rect 0 -49 2880 -17
<< labels >>
flabel pwell s 0 0 2880 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 0 617 2880 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
rlabel comment s 0 0 0 0 4 sdfsbp_1
flabel comment s 1227 315 1227 315 0 FreeSans 200 0 0 0 no_jumper_check
flabel comment s 1084 358 1084 358 0 FreeSans 200 0 0 0 no_jumper_check
flabel metal1 s 1951 316 1985 350 0 FreeSans 340 0 0 0 SET_B
port 5 nsew
flabel metal1 s 0 617 2880 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 2880 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 2815 94 2849 128 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2815 168 2849 202 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2815 242 2849 276 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2815 316 2849 350 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2815 390 2849 424 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2815 464 2849 498 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2815 538 2849 572 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2431 94 2465 128 0 FreeSans 340 0 0 0 Q_N
port 11 nsew
flabel corelocali s 2431 168 2465 202 0 FreeSans 340 0 0 0 Q_N
port 11 nsew
flabel corelocali s 511 242 545 276 0 FreeSans 340 0 0 0 SCD
port 3 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 SCD
port 3 nsew
flabel corelocali s 511 390 545 424 0 FreeSans 340 0 0 0 SCD
port 3 nsew
flabel corelocali s 703 242 737 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 SCE
port 4 nsew
flabel corelocali s 223 390 257 424 0 FreeSans 340 0 0 0 D
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 2880 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 168006
string GDS_START 147166
<< end >>
