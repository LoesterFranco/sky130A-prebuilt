magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 2024 561
rect 106 337 172 417
rect 278 337 344 417
rect 106 331 344 337
rect 29 295 344 331
rect 1244 357 1310 527
rect 1416 361 1482 527
rect 1616 379 1682 527
rect 1806 383 1872 527
rect 29 157 64 295
rect 99 204 369 255
rect 411 204 749 255
rect 791 204 1130 255
rect 1219 204 1549 255
rect 1592 204 1998 255
rect 29 123 1524 157
rect 123 91 158 123
rect 292 91 330 123
rect 480 91 518 123
rect 652 91 702 123
rect 836 91 884 123
rect 1018 91 1055 123
rect 23 17 89 89
rect 192 17 258 89
rect 364 17 446 89
rect 552 17 618 89
rect 736 17 802 89
rect 918 17 984 89
rect 1089 17 1156 89
rect 1649 17 1715 89
rect 1821 17 1887 89
rect 0 -17 2024 17
<< obsli1 >>
rect 20 451 774 489
rect 20 367 72 451
rect 206 371 244 451
rect 378 371 416 451
rect 450 337 516 417
rect 550 371 588 451
rect 622 337 688 417
rect 722 367 774 451
rect 812 455 1210 489
rect 812 451 1036 455
rect 812 367 864 451
rect 450 331 688 337
rect 898 337 964 417
rect 998 371 1036 451
rect 1070 337 1136 417
rect 898 331 1136 337
rect 450 295 1136 331
rect 1172 323 1210 455
rect 1344 323 1382 463
rect 1516 333 1582 463
rect 1716 334 1768 458
rect 1906 334 1954 452
rect 1716 333 1954 334
rect 1516 323 1954 333
rect 1172 289 1954 323
rect 1577 123 1973 157
rect 1577 89 1615 123
rect 1196 55 1615 89
rect 1749 60 1787 123
rect 1921 58 1973 123
<< metal1 >>
rect 0 496 2024 592
rect 0 -48 2024 48
<< labels >>
rlabel locali s 1219 204 1549 255 6 A1
port 1 nsew signal input
rlabel locali s 1592 204 1998 255 6 A2
port 2 nsew signal input
rlabel locali s 791 204 1130 255 6 B1
port 3 nsew signal input
rlabel locali s 411 204 749 255 6 C1
port 4 nsew signal input
rlabel locali s 99 204 369 255 6 D1
port 5 nsew signal input
rlabel locali s 1018 91 1055 123 6 Y
port 6 nsew signal output
rlabel locali s 836 91 884 123 6 Y
port 6 nsew signal output
rlabel locali s 652 91 702 123 6 Y
port 6 nsew signal output
rlabel locali s 480 91 518 123 6 Y
port 6 nsew signal output
rlabel locali s 292 91 330 123 6 Y
port 6 nsew signal output
rlabel locali s 278 337 344 417 6 Y
port 6 nsew signal output
rlabel locali s 123 91 158 123 6 Y
port 6 nsew signal output
rlabel locali s 106 337 172 417 6 Y
port 6 nsew signal output
rlabel locali s 106 331 344 337 6 Y
port 6 nsew signal output
rlabel locali s 29 295 344 331 6 Y
port 6 nsew signal output
rlabel locali s 29 157 64 295 6 Y
port 6 nsew signal output
rlabel locali s 29 123 1524 157 6 Y
port 6 nsew signal output
rlabel locali s 1821 17 1887 89 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1649 17 1715 89 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1089 17 1156 89 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 918 17 984 89 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 736 17 802 89 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 552 17 618 89 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 364 17 446 89 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 192 17 258 89 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 23 17 89 89 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 2024 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 2024 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1806 383 1872 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1616 379 1682 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1416 361 1482 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1244 357 1310 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 2024 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 2024 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2024 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3949216
string GDS_START 3935052
<< end >>
