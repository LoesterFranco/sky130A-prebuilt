magic
tech sky130A
magscale 1 2
timestamp 1599588232
<< locali >>
rect 25 236 102 310
rect 204 364 283 414
rect 204 208 238 364
rect 545 252 647 356
rect 681 290 747 356
rect 204 168 279 208
rect 245 150 279 168
rect 245 70 313 150
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 24 482 90 540
rect 127 516 193 649
rect 307 516 373 649
rect 24 448 362 482
rect 24 364 90 448
rect 136 202 170 448
rect 54 168 170 202
rect 321 378 362 448
rect 411 412 483 596
rect 517 454 551 596
rect 591 488 641 649
rect 681 454 747 596
rect 517 420 747 454
rect 449 386 483 412
rect 681 390 747 420
rect 321 344 415 378
rect 449 352 511 386
rect 381 318 415 344
rect 272 244 347 310
rect 381 252 443 318
rect 313 218 347 244
rect 477 218 511 352
rect 313 184 562 218
rect 54 108 120 168
rect 161 17 211 134
rect 347 17 462 150
rect 496 70 562 184
rect 676 17 742 218
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel locali s 545 252 647 356 6 A1
port 1 nsew signal input
rlabel locali s 681 290 747 356 6 A2
port 2 nsew signal input
rlabel locali s 25 236 102 310 6 B1_N
port 3 nsew signal input
rlabel locali s 245 150 279 168 6 X
port 4 nsew signal output
rlabel locali s 245 70 313 150 6 X
port 4 nsew signal output
rlabel locali s 204 364 283 414 6 X
port 4 nsew signal output
rlabel locali s 204 208 238 364 6 X
port 4 nsew signal output
rlabel locali s 204 168 279 208 6 X
port 4 nsew signal output
rlabel metal1 s 0 -49 768 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 6 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 617 768 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 4039504
string GDS_START 4032776
<< end >>
