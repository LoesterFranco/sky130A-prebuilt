magic
tech sky130A
magscale 1 2
timestamp 1599588209
<< nwell >>
rect -38 332 806 704
<< pwell >>
rect 0 0 768 49
<< scpmos >>
rect 86 368 116 592
rect 218 368 248 568
rect 302 368 332 568
rect 410 368 440 568
rect 518 368 548 568
rect 637 368 667 568
<< nmoslvt >>
rect 107 74 137 222
rect 221 74 251 202
rect 307 74 337 202
rect 421 74 451 202
rect 521 74 551 202
rect 640 74 670 202
<< ndiff >>
rect 50 210 107 222
rect 50 176 62 210
rect 96 176 107 210
rect 50 120 107 176
rect 50 86 62 120
rect 96 86 107 120
rect 50 74 107 86
rect 137 202 187 222
rect 137 190 221 202
rect 137 156 162 190
rect 196 156 221 190
rect 137 120 221 156
rect 137 86 162 120
rect 196 86 221 120
rect 137 74 221 86
rect 251 190 307 202
rect 251 156 262 190
rect 296 156 307 190
rect 251 120 307 156
rect 251 86 262 120
rect 296 86 307 120
rect 251 74 307 86
rect 337 148 421 202
rect 337 114 362 148
rect 396 114 421 148
rect 337 74 421 114
rect 451 190 521 202
rect 451 156 462 190
rect 496 156 521 190
rect 451 120 521 156
rect 451 86 462 120
rect 496 86 521 120
rect 451 74 521 86
rect 551 190 640 202
rect 551 156 578 190
rect 612 156 640 190
rect 551 74 640 156
rect 670 186 737 202
rect 670 152 681 186
rect 715 152 737 186
rect 670 118 737 152
rect 670 84 681 118
rect 715 84 737 118
rect 670 74 737 84
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 497 86 546
rect 27 463 39 497
rect 73 463 86 497
rect 27 414 86 463
rect 27 380 39 414
rect 73 380 86 414
rect 27 368 86 380
rect 116 580 185 592
rect 116 546 139 580
rect 173 568 185 580
rect 173 546 218 568
rect 116 508 218 546
rect 116 474 139 508
rect 173 474 218 508
rect 116 368 218 474
rect 248 368 302 568
rect 332 368 410 568
rect 440 560 518 568
rect 440 526 462 560
rect 496 526 518 560
rect 440 492 518 526
rect 440 458 462 492
rect 496 458 518 492
rect 440 424 518 458
rect 440 390 462 424
rect 496 390 518 424
rect 440 368 518 390
rect 548 368 637 568
rect 667 556 726 568
rect 667 522 680 556
rect 714 522 726 556
rect 667 444 726 522
rect 667 410 682 444
rect 716 410 726 444
rect 667 368 726 410
<< ndiffc >>
rect 62 176 96 210
rect 62 86 96 120
rect 162 156 196 190
rect 162 86 196 120
rect 262 156 296 190
rect 262 86 296 120
rect 362 114 396 148
rect 462 156 496 190
rect 462 86 496 120
rect 578 156 612 190
rect 681 152 715 186
rect 681 84 715 118
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 139 546 173 580
rect 139 474 173 508
rect 462 526 496 560
rect 462 458 496 492
rect 462 390 496 424
rect 680 522 714 556
rect 682 410 716 444
<< poly >>
rect 86 592 116 618
rect 218 568 248 594
rect 302 568 332 594
rect 410 568 440 594
rect 518 568 548 594
rect 637 568 667 594
rect 86 353 116 368
rect 218 353 248 368
rect 302 353 332 368
rect 410 353 440 368
rect 518 353 548 368
rect 637 353 667 368
rect 83 330 119 353
rect 215 336 251 353
rect 299 336 335 353
rect 407 336 443 353
rect 515 336 551 353
rect 83 314 149 330
rect 83 280 99 314
rect 133 280 149 314
rect 83 264 149 280
rect 191 320 257 336
rect 191 286 207 320
rect 241 286 257 320
rect 191 270 257 286
rect 299 320 365 336
rect 299 286 315 320
rect 349 286 365 320
rect 299 270 365 286
rect 407 320 473 336
rect 407 286 423 320
rect 457 286 473 320
rect 407 270 473 286
rect 515 320 581 336
rect 515 286 531 320
rect 565 286 581 320
rect 515 270 581 286
rect 634 302 670 353
rect 634 286 747 302
rect 107 222 137 264
rect 221 202 251 270
rect 307 202 337 270
rect 421 202 451 270
rect 521 202 551 270
rect 634 252 697 286
rect 731 252 747 286
rect 634 236 747 252
rect 640 202 670 236
rect 107 48 137 74
rect 221 48 251 74
rect 307 48 337 74
rect 421 48 451 74
rect 521 48 551 74
rect 640 48 670 74
<< polycont >>
rect 99 280 133 314
rect 207 286 241 320
rect 315 286 349 320
rect 423 286 457 320
rect 531 286 565 320
rect 697 252 731 286
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 17 580 89 596
rect 17 546 39 580
rect 73 546 89 580
rect 17 497 89 546
rect 17 463 39 497
rect 73 463 89 497
rect 17 414 89 463
rect 123 580 189 649
rect 123 546 139 580
rect 173 546 189 580
rect 123 508 189 546
rect 123 474 139 508
rect 173 474 189 508
rect 123 458 189 474
rect 441 560 519 576
rect 441 526 462 560
rect 496 526 519 560
rect 441 492 519 526
rect 441 458 462 492
rect 496 458 519 492
rect 664 556 730 649
rect 664 522 680 556
rect 714 522 730 556
rect 664 458 730 522
rect 441 424 519 458
rect 682 444 730 458
rect 17 380 39 414
rect 73 380 89 414
rect 17 364 89 380
rect 123 390 462 424
rect 496 390 647 424
rect 716 410 730 444
rect 682 394 730 410
rect 17 226 51 364
rect 123 330 157 390
rect 85 314 157 330
rect 85 280 99 314
rect 133 280 157 314
rect 85 264 157 280
rect 191 320 263 356
rect 191 286 207 320
rect 241 286 263 320
rect 191 270 263 286
rect 299 320 365 356
rect 299 286 315 320
rect 349 286 365 320
rect 299 270 365 286
rect 407 320 473 356
rect 407 286 423 320
rect 457 286 473 320
rect 407 270 473 286
rect 507 320 579 356
rect 507 286 531 320
rect 565 286 579 320
rect 507 270 579 286
rect 613 236 647 390
rect 682 286 747 356
rect 682 252 697 286
rect 731 252 747 286
rect 682 236 747 252
rect 17 210 112 226
rect 17 176 62 210
rect 96 176 112 210
rect 17 120 112 176
rect 17 86 62 120
rect 96 86 112 120
rect 17 70 112 86
rect 146 190 212 206
rect 146 156 162 190
rect 196 156 212 190
rect 146 120 212 156
rect 146 86 162 120
rect 196 86 212 120
rect 146 17 212 86
rect 246 202 512 236
rect 246 190 312 202
rect 246 156 262 190
rect 296 156 312 190
rect 446 190 512 202
rect 246 120 312 156
rect 246 86 262 120
rect 296 86 312 120
rect 246 70 312 86
rect 346 148 412 164
rect 346 114 362 148
rect 396 114 412 148
rect 346 17 412 114
rect 446 156 462 190
rect 496 156 512 190
rect 446 120 512 156
rect 546 202 647 236
rect 546 190 645 202
rect 546 156 578 190
rect 612 156 645 190
rect 546 140 645 156
rect 681 186 731 202
rect 715 152 731 186
rect 446 86 462 120
rect 496 104 512 120
rect 681 118 731 152
rect 496 86 681 104
rect 446 84 681 86
rect 715 84 731 118
rect 446 68 731 84
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o32a_1
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 703 242 737 276 0 FreeSans 340 0 0 0 B1
port 4 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 B1
port 4 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 B2
port 5 nsew
flabel corelocali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 10 nsew
flabel corelocali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 768 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 688302
string GDS_START 681218
<< end >>
