magic
tech sky130A
magscale 1 2
timestamp 1604502705
<< nwell >>
rect -38 332 710 704
<< pwell >>
rect 0 0 672 49
<< scnmos >>
rect 87 100 117 248
rect 235 120 265 248
rect 307 120 337 248
rect 415 123 445 251
rect 533 123 563 251
<< pmoshvt >>
rect 84 368 114 592
rect 220 392 250 592
rect 310 392 340 592
rect 436 392 466 592
rect 526 392 556 592
<< ndiff >>
rect 365 248 415 251
rect 34 220 87 248
rect 34 186 42 220
rect 76 186 87 220
rect 34 146 87 186
rect 34 112 42 146
rect 76 112 87 146
rect 34 100 87 112
rect 117 196 235 248
rect 117 162 190 196
rect 224 162 235 196
rect 117 142 235 162
rect 117 108 128 142
rect 162 120 235 142
rect 265 120 307 248
rect 337 123 415 248
rect 445 208 533 251
rect 445 174 472 208
rect 506 174 533 208
rect 445 123 533 174
rect 563 196 616 251
rect 563 162 574 196
rect 608 162 616 196
rect 563 123 616 162
rect 337 120 387 123
rect 162 108 188 120
rect 117 100 188 108
<< pdiff >>
rect 29 580 84 592
rect 29 546 37 580
rect 71 546 84 580
rect 29 500 84 546
rect 29 466 37 500
rect 71 466 84 500
rect 29 420 84 466
rect 29 386 37 420
rect 71 386 84 420
rect 29 368 84 386
rect 114 580 220 592
rect 114 546 150 580
rect 184 546 220 580
rect 114 512 220 546
rect 114 478 150 512
rect 184 478 220 512
rect 114 444 220 478
rect 114 410 150 444
rect 184 410 220 444
rect 114 392 220 410
rect 250 580 310 592
rect 250 546 263 580
rect 297 546 310 580
rect 250 512 310 546
rect 250 478 263 512
rect 297 478 310 512
rect 250 444 310 478
rect 250 410 263 444
rect 297 410 310 444
rect 250 392 310 410
rect 340 580 436 592
rect 340 546 371 580
rect 405 546 436 580
rect 340 501 436 546
rect 340 467 371 501
rect 405 467 436 501
rect 340 392 436 467
rect 466 580 526 592
rect 466 546 479 580
rect 513 546 526 580
rect 466 512 526 546
rect 466 478 479 512
rect 513 478 526 512
rect 466 444 526 478
rect 466 410 479 444
rect 513 410 526 444
rect 466 392 526 410
rect 556 580 611 592
rect 556 546 569 580
rect 603 546 611 580
rect 556 509 611 546
rect 556 475 569 509
rect 603 475 611 509
rect 556 438 611 475
rect 556 404 569 438
rect 603 404 611 438
rect 556 392 611 404
rect 114 368 167 392
<< ndiffc >>
rect 42 186 76 220
rect 42 112 76 146
rect 190 162 224 196
rect 128 108 162 142
rect 472 174 506 208
rect 574 162 608 196
<< pdiffc >>
rect 37 546 71 580
rect 37 466 71 500
rect 37 386 71 420
rect 150 546 184 580
rect 150 478 184 512
rect 150 410 184 444
rect 263 546 297 580
rect 263 478 297 512
rect 263 410 297 444
rect 371 546 405 580
rect 371 467 405 501
rect 479 546 513 580
rect 479 478 513 512
rect 479 410 513 444
rect 569 546 603 580
rect 569 475 603 509
rect 569 404 603 438
<< poly >>
rect 84 592 114 618
rect 220 592 250 618
rect 310 592 340 618
rect 436 592 466 618
rect 526 592 556 618
rect 220 377 250 392
rect 310 377 340 392
rect 436 377 466 392
rect 526 377 556 392
rect 84 353 114 368
rect 217 360 253 377
rect 307 360 343 377
rect 433 360 469 377
rect 81 336 117 353
rect 199 344 265 360
rect 81 320 151 336
rect 81 286 101 320
rect 135 286 151 320
rect 199 310 215 344
rect 249 310 265 344
rect 199 294 265 310
rect 81 270 151 286
rect 87 248 117 270
rect 235 248 265 294
rect 307 344 373 360
rect 307 310 323 344
rect 357 310 373 344
rect 307 294 373 310
rect 415 344 481 360
rect 415 310 431 344
rect 465 310 481 344
rect 415 294 481 310
rect 523 317 559 377
rect 307 248 337 294
rect 415 251 445 294
rect 523 287 563 317
rect 533 251 563 287
rect 87 74 117 100
rect 235 94 265 120
rect 307 94 337 120
rect 415 97 445 123
rect 533 101 563 123
rect 497 85 563 101
rect 497 51 513 85
rect 547 51 563 85
rect 497 35 563 51
<< polycont >>
rect 101 286 135 320
rect 215 310 249 344
rect 323 310 357 344
rect 431 310 465 344
rect 513 51 547 85
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 17 580 87 596
rect 17 546 37 580
rect 71 546 87 580
rect 17 500 87 546
rect 17 466 37 500
rect 71 466 87 500
rect 17 420 87 466
rect 17 386 37 420
rect 71 386 87 420
rect 121 580 213 649
rect 121 546 150 580
rect 184 546 213 580
rect 121 512 213 546
rect 121 478 150 512
rect 184 478 213 512
rect 121 444 213 478
rect 121 410 150 444
rect 184 410 213 444
rect 121 394 213 410
rect 247 580 313 596
rect 247 546 263 580
rect 297 546 313 580
rect 247 512 313 546
rect 247 478 263 512
rect 297 478 313 512
rect 247 444 313 478
rect 347 580 429 649
rect 347 546 371 580
rect 405 546 429 580
rect 347 501 429 546
rect 347 467 371 501
rect 405 467 429 501
rect 347 462 429 467
rect 463 580 529 596
rect 463 546 479 580
rect 513 546 529 580
rect 463 512 529 546
rect 463 478 479 512
rect 513 478 529 512
rect 247 410 263 444
rect 297 428 313 444
rect 463 444 529 478
rect 463 428 479 444
rect 297 410 479 428
rect 513 410 529 444
rect 247 394 529 410
rect 569 580 619 596
rect 603 546 619 580
rect 569 509 619 546
rect 603 475 619 509
rect 569 438 619 475
rect 603 404 619 438
rect 17 370 87 386
rect 17 236 51 370
rect 199 344 265 360
rect 85 320 165 336
rect 85 286 101 320
rect 135 286 165 320
rect 199 310 215 344
rect 249 310 265 344
rect 199 298 265 310
rect 307 344 373 360
rect 307 310 323 344
rect 357 310 373 344
rect 307 298 373 310
rect 409 344 481 360
rect 409 310 431 344
rect 465 310 481 344
rect 409 298 481 310
rect 85 270 165 286
rect 124 264 165 270
rect 569 264 619 404
rect 17 220 90 236
rect 124 230 619 264
rect 17 186 42 220
rect 76 186 90 220
rect 456 208 522 230
rect 17 146 90 186
rect 17 112 42 146
rect 76 112 90 146
rect 17 96 90 112
rect 124 162 190 196
rect 224 162 240 196
rect 456 174 472 208
rect 506 174 522 208
rect 456 162 522 174
rect 558 162 574 196
rect 608 162 631 196
rect 124 142 240 162
rect 124 108 128 142
rect 162 108 240 142
rect 124 17 240 108
rect 313 85 563 128
rect 313 51 513 85
rect 547 51 563 85
rect 597 17 631 162
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a31o_1
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 319 94 353 128 0 FreeSans 340 0 0 0 B1
port 4 nsew
flabel corelocali s 415 94 449 128 0 FreeSans 340 0 0 0 B1
port 4 nsew
flabel corelocali s 511 94 545 128 0 FreeSans 340 0 0 0 B1
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 672 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3699264
string GDS_START 3692294
<< end >>
