magic
tech sky130A
magscale 1 2
timestamp 1604502710
<< nwell >>
rect -38 332 902 704
<< pwell >>
rect 0 0 864 49
<< scpmos >>
rect 83 424 119 592
rect 340 368 376 568
rect 454 368 490 568
rect 544 368 580 568
rect 652 368 688 592
rect 745 368 781 592
<< nmoslvt >>
rect 84 88 114 198
rect 346 74 376 222
rect 424 74 454 222
rect 538 74 568 222
rect 652 74 682 222
rect 738 74 768 222
<< ndiff >>
rect 289 210 346 222
rect 27 160 84 198
rect 27 126 39 160
rect 73 126 84 160
rect 27 88 84 126
rect 114 141 173 198
rect 114 107 125 141
rect 159 107 173 141
rect 114 88 173 107
rect 289 176 301 210
rect 335 176 346 210
rect 289 120 346 176
rect 289 86 301 120
rect 335 86 346 120
rect 289 74 346 86
rect 376 74 424 222
rect 454 74 538 222
rect 568 210 652 222
rect 568 176 579 210
rect 613 176 652 210
rect 568 120 652 176
rect 568 86 579 120
rect 613 86 652 120
rect 568 74 652 86
rect 682 210 738 222
rect 682 176 693 210
rect 727 176 738 210
rect 682 120 738 176
rect 682 86 693 120
rect 727 86 738 120
rect 682 74 738 86
rect 768 210 825 222
rect 768 176 779 210
rect 813 176 825 210
rect 768 120 825 176
rect 768 86 779 120
rect 813 86 825 120
rect 768 74 825 86
<< pdiff >>
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 470 83 546
rect 27 436 39 470
rect 73 436 83 470
rect 27 424 83 436
rect 119 538 177 592
rect 596 568 652 592
rect 119 504 130 538
rect 164 504 177 538
rect 119 424 177 504
rect 284 556 340 568
rect 284 522 296 556
rect 330 522 340 556
rect 284 485 340 522
rect 284 451 296 485
rect 330 451 340 485
rect 284 414 340 451
rect 284 380 296 414
rect 330 380 340 414
rect 284 368 340 380
rect 376 560 454 568
rect 376 526 396 560
rect 430 526 454 560
rect 376 492 454 526
rect 376 458 396 492
rect 430 458 454 492
rect 376 368 454 458
rect 490 560 544 568
rect 490 526 500 560
rect 534 526 544 560
rect 490 492 544 526
rect 490 458 500 492
rect 534 458 544 492
rect 490 424 544 458
rect 490 390 500 424
rect 534 390 544 424
rect 490 368 544 390
rect 580 560 652 568
rect 580 526 608 560
rect 642 526 652 560
rect 580 368 652 526
rect 688 414 745 592
rect 688 380 699 414
rect 733 380 745 414
rect 688 368 745 380
rect 781 560 837 592
rect 781 526 791 560
rect 825 526 837 560
rect 781 368 837 526
<< ndiffc >>
rect 39 126 73 160
rect 125 107 159 141
rect 301 176 335 210
rect 301 86 335 120
rect 579 176 613 210
rect 579 86 613 120
rect 693 176 727 210
rect 693 86 727 120
rect 779 176 813 210
rect 779 86 813 120
<< pdiffc >>
rect 39 546 73 580
rect 39 436 73 470
rect 130 504 164 538
rect 296 522 330 556
rect 296 451 330 485
rect 296 380 330 414
rect 396 526 430 560
rect 396 458 430 492
rect 500 526 534 560
rect 500 458 534 492
rect 500 390 534 424
rect 608 526 642 560
rect 699 380 733 414
rect 791 526 825 560
<< poly >>
rect 83 592 119 618
rect 340 568 376 594
rect 454 568 490 594
rect 544 568 580 594
rect 652 592 688 618
rect 745 592 781 618
rect 83 386 119 424
rect 44 370 114 386
rect 44 336 60 370
rect 94 336 114 370
rect 44 302 114 336
rect 44 268 60 302
rect 94 268 114 302
rect 44 252 114 268
rect 84 198 114 252
rect 180 355 246 371
rect 180 321 196 355
rect 230 322 246 355
rect 340 322 376 368
rect 230 321 376 322
rect 180 287 376 321
rect 454 310 490 368
rect 544 336 580 368
rect 180 253 196 287
rect 230 253 376 287
rect 180 237 376 253
rect 346 222 376 237
rect 424 294 490 310
rect 424 260 440 294
rect 474 260 490 294
rect 424 244 490 260
rect 538 320 604 336
rect 538 286 554 320
rect 588 286 604 320
rect 538 270 604 286
rect 652 326 688 368
rect 745 326 781 368
rect 652 310 843 326
rect 652 276 793 310
rect 827 276 843 310
rect 424 222 454 244
rect 538 222 568 270
rect 652 260 843 276
rect 652 222 682 260
rect 738 222 768 260
rect 84 62 114 88
rect 346 48 376 74
rect 424 48 454 74
rect 538 48 568 74
rect 652 48 682 74
rect 738 48 768 74
<< polycont >>
rect 60 336 94 370
rect 60 268 94 302
rect 196 321 230 355
rect 196 253 230 287
rect 440 260 474 294
rect 554 286 588 320
rect 793 276 827 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 23 580 80 596
rect 23 546 39 580
rect 73 546 80 580
rect 23 470 80 546
rect 114 538 180 649
rect 114 504 130 538
rect 164 504 180 538
rect 114 488 180 504
rect 280 556 346 572
rect 280 522 296 556
rect 330 522 346 556
rect 23 436 39 470
rect 73 454 80 470
rect 280 485 346 522
rect 73 436 214 454
rect 23 420 214 436
rect 25 370 110 386
rect 25 336 60 370
rect 94 336 110 370
rect 25 302 110 336
rect 25 268 60 302
rect 94 268 110 302
rect 25 252 110 268
rect 180 371 214 420
rect 280 451 296 485
rect 330 451 346 485
rect 380 560 446 649
rect 380 526 396 560
rect 430 526 446 560
rect 380 492 446 526
rect 380 458 396 492
rect 430 458 446 492
rect 484 560 550 572
rect 484 526 500 560
rect 534 526 550 560
rect 484 492 550 526
rect 592 560 658 649
rect 592 526 608 560
rect 642 526 658 560
rect 592 516 658 526
rect 775 560 841 649
rect 775 526 791 560
rect 825 526 841 560
rect 775 516 841 526
rect 484 458 500 492
rect 534 482 550 492
rect 534 458 843 482
rect 280 424 346 451
rect 484 448 843 458
rect 484 424 550 448
rect 280 414 500 424
rect 280 380 296 414
rect 330 390 500 414
rect 534 390 550 424
rect 330 380 351 390
rect 180 355 246 371
rect 180 321 196 355
rect 230 321 246 355
rect 180 287 246 321
rect 180 253 196 287
rect 230 253 246 287
rect 180 218 246 253
rect 23 184 246 218
rect 280 210 351 380
rect 682 380 699 414
rect 733 380 751 414
rect 682 364 751 380
rect 23 160 75 184
rect 23 126 39 160
rect 73 126 75 160
rect 280 176 301 210
rect 335 176 351 210
rect 23 84 75 126
rect 109 141 175 150
rect 109 107 125 141
rect 159 107 175 141
rect 109 17 175 107
rect 280 120 351 176
rect 280 86 301 120
rect 335 86 351 120
rect 409 294 490 356
rect 409 260 440 294
rect 474 260 490 294
rect 538 320 647 356
rect 538 286 554 320
rect 588 286 647 320
rect 538 270 647 286
rect 409 88 490 260
rect 682 226 743 364
rect 809 326 843 448
rect 777 310 843 326
rect 777 276 793 310
rect 827 276 843 310
rect 777 260 843 276
rect 563 210 629 226
rect 563 176 579 210
rect 613 176 629 210
rect 563 120 629 176
rect 280 70 351 86
rect 563 86 579 120
rect 613 86 629 120
rect 563 17 629 86
rect 677 210 743 226
rect 677 176 693 210
rect 727 176 743 210
rect 677 120 743 176
rect 677 86 693 120
rect 727 86 743 120
rect 677 70 743 86
rect 779 210 829 226
rect 813 176 829 210
rect 779 120 829 176
rect 813 86 829 120
rect 779 17 829 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
rlabel comment s 0 0 0 0 4 and3b_2
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 415 94 449 128 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 415 168 449 202 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 415 242 449 276 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 703 94 737 128 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 703 168 737 202 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 703 242 737 276 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 X
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 864 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3184732
string GDS_START 3177168
<< end >>
