magic
tech sky130A
magscale 1 2
timestamp 1604502701
<< nwell >>
rect -38 332 614 704
<< pwell >>
rect 0 0 576 49
<< scpmos >>
rect 126 368 156 592
rect 234 368 264 592
rect 324 368 354 592
rect 420 368 450 592
<< nmoslvt >>
rect 129 74 159 222
rect 201 74 231 222
rect 309 74 339 222
rect 417 74 447 222
<< ndiff >>
rect 76 210 129 222
rect 76 176 84 210
rect 118 176 129 210
rect 76 120 129 176
rect 76 86 84 120
rect 118 86 129 120
rect 76 74 129 86
rect 159 74 201 222
rect 231 210 309 222
rect 231 176 246 210
rect 280 176 309 210
rect 231 120 309 176
rect 231 86 246 120
rect 280 86 309 120
rect 231 74 309 86
rect 339 124 417 222
rect 339 90 354 124
rect 388 90 417 124
rect 339 74 417 90
rect 447 202 500 222
rect 447 168 458 202
rect 492 168 500 202
rect 447 120 500 168
rect 447 86 458 120
rect 492 86 500 120
rect 447 74 500 86
<< pdiff >>
rect 71 580 126 592
rect 71 546 79 580
rect 113 546 126 580
rect 71 508 126 546
rect 71 474 79 508
rect 113 474 126 508
rect 71 424 126 474
rect 71 390 79 424
rect 113 390 126 424
rect 71 368 126 390
rect 156 578 234 592
rect 156 544 173 578
rect 207 544 234 578
rect 156 508 234 544
rect 156 474 173 508
rect 207 474 234 508
rect 156 368 234 474
rect 264 580 324 592
rect 264 546 277 580
rect 311 546 324 580
rect 264 508 324 546
rect 264 474 277 508
rect 311 474 324 508
rect 264 424 324 474
rect 264 390 277 424
rect 311 390 324 424
rect 264 368 324 390
rect 354 368 420 592
rect 450 580 505 592
rect 450 546 463 580
rect 497 546 505 580
rect 450 497 505 546
rect 450 463 463 497
rect 497 463 505 497
rect 450 414 505 463
rect 450 380 463 414
rect 497 380 505 414
rect 450 368 505 380
<< ndiffc >>
rect 84 176 118 210
rect 84 86 118 120
rect 246 176 280 210
rect 246 86 280 120
rect 354 90 388 124
rect 458 168 492 202
rect 458 86 492 120
<< pdiffc >>
rect 79 546 113 580
rect 79 474 113 508
rect 79 390 113 424
rect 173 544 207 578
rect 173 474 207 508
rect 277 546 311 580
rect 277 474 311 508
rect 277 390 311 424
rect 463 546 497 580
rect 463 463 497 497
rect 463 380 497 414
<< poly >>
rect 126 592 156 618
rect 234 592 264 618
rect 324 592 354 618
rect 420 592 450 618
rect 126 353 156 368
rect 234 353 264 368
rect 324 353 354 368
rect 420 353 450 368
rect 123 336 159 353
rect 231 336 267 353
rect 321 336 357 353
rect 93 320 159 336
rect 93 286 109 320
rect 143 286 159 320
rect 93 270 159 286
rect 129 222 159 270
rect 201 320 267 336
rect 201 286 217 320
rect 251 286 267 320
rect 201 270 267 286
rect 309 320 375 336
rect 309 286 325 320
rect 359 286 375 320
rect 309 270 375 286
rect 417 310 453 353
rect 417 294 555 310
rect 201 222 231 270
rect 309 222 339 270
rect 417 260 505 294
rect 539 260 555 294
rect 417 244 555 260
rect 417 222 447 244
rect 129 48 159 74
rect 201 48 231 74
rect 309 48 339 74
rect 417 48 447 74
<< polycont >>
rect 109 286 143 320
rect 217 286 251 320
rect 325 286 359 320
rect 505 260 539 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 63 580 129 596
rect 63 546 79 580
rect 113 546 129 580
rect 63 508 129 546
rect 63 474 79 508
rect 113 474 129 508
rect 63 424 129 474
rect 163 578 227 649
rect 163 544 173 578
rect 207 544 227 578
rect 163 508 227 544
rect 163 474 173 508
rect 207 474 227 508
rect 163 458 227 474
rect 261 580 327 596
rect 261 546 277 580
rect 311 546 327 580
rect 261 508 327 546
rect 261 474 277 508
rect 311 474 327 508
rect 261 424 327 474
rect 63 390 79 424
rect 113 390 277 424
rect 311 390 327 424
rect 409 580 513 596
rect 409 546 463 580
rect 497 546 513 580
rect 409 497 513 546
rect 409 463 463 497
rect 497 463 513 497
rect 409 414 513 463
rect 409 380 463 414
rect 497 380 513 414
rect 409 364 513 380
rect 93 320 167 356
rect 93 286 109 320
rect 143 286 167 320
rect 93 270 167 286
rect 201 320 267 356
rect 201 286 217 320
rect 251 286 267 320
rect 201 270 267 286
rect 309 320 375 356
rect 309 286 325 320
rect 359 286 375 320
rect 309 270 375 286
rect 409 236 443 364
rect 489 294 555 310
rect 489 260 505 294
rect 539 260 555 294
rect 489 236 555 260
rect 68 210 134 226
rect 68 176 84 210
rect 118 176 134 210
rect 68 120 134 176
rect 68 86 84 120
rect 118 86 134 120
rect 68 17 134 86
rect 217 210 443 236
rect 217 176 246 210
rect 280 205 443 210
rect 280 202 455 205
rect 280 176 458 202
rect 217 168 458 176
rect 492 168 508 202
rect 217 162 508 168
rect 217 120 300 162
rect 217 86 246 120
rect 280 86 300 120
rect 217 70 300 86
rect 334 124 408 128
rect 334 90 354 124
rect 388 90 408 124
rect 334 17 408 90
rect 442 120 508 162
rect 442 86 458 120
rect 492 86 508 120
rect 442 70 508 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a211oi_1
flabel pwell s 0 0 576 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 576 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 576 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 576 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 511 242 545 276 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 223 168 257 202 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 319 168 353 202 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 415 168 449 202 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 576 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3999596
string GDS_START 3993932
<< end >>
