magic
tech sky130A
magscale 1 2
timestamp 1599588209
<< nwell >>
rect -38 332 902 704
<< pwell >>
rect 0 0 864 49
<< scpmos >>
rect 86 368 116 592
rect 179 368 209 592
rect 274 368 304 592
rect 364 368 394 592
rect 460 368 490 592
rect 568 368 598 592
rect 658 368 688 592
rect 748 368 778 592
<< nmoslvt >>
rect 277 74 307 222
rect 371 74 401 222
rect 485 74 515 222
rect 571 74 601 222
<< ndiff >>
rect 227 132 277 222
rect 125 120 277 132
rect 125 86 137 120
rect 171 86 226 120
rect 260 86 277 120
rect 125 74 277 86
rect 307 210 371 222
rect 307 176 326 210
rect 360 176 371 210
rect 307 120 371 176
rect 307 86 326 120
rect 360 86 371 120
rect 307 74 371 86
rect 401 146 485 222
rect 401 112 426 146
rect 460 112 485 146
rect 401 74 485 112
rect 515 210 571 222
rect 515 176 526 210
rect 560 176 571 210
rect 515 120 571 176
rect 515 86 526 120
rect 560 86 571 120
rect 515 74 571 86
rect 601 186 672 222
rect 601 152 612 186
rect 646 152 672 186
rect 601 118 672 152
rect 601 84 612 118
rect 646 84 672 118
rect 601 74 672 84
<< pdiff >>
rect 27 584 86 592
rect 27 550 39 584
rect 73 550 86 584
rect 27 516 86 550
rect 27 482 39 516
rect 73 482 86 516
rect 27 448 86 482
rect 27 414 39 448
rect 73 414 86 448
rect 27 368 86 414
rect 116 566 179 592
rect 116 532 130 566
rect 164 532 179 566
rect 116 368 179 532
rect 209 414 274 592
rect 209 380 224 414
rect 258 380 274 414
rect 209 368 274 380
rect 304 573 364 592
rect 304 539 317 573
rect 351 539 364 573
rect 304 368 364 539
rect 394 580 460 592
rect 394 546 407 580
rect 441 546 460 580
rect 394 497 460 546
rect 394 463 407 497
rect 441 463 460 497
rect 394 414 460 463
rect 394 380 407 414
rect 441 380 460 414
rect 394 368 460 380
rect 490 584 568 592
rect 490 550 511 584
rect 545 550 568 584
rect 490 516 568 550
rect 490 482 511 516
rect 545 482 568 516
rect 490 368 568 482
rect 598 580 658 592
rect 598 546 611 580
rect 645 546 658 580
rect 598 368 658 546
rect 688 584 748 592
rect 688 550 701 584
rect 735 550 748 584
rect 688 512 748 550
rect 688 478 701 512
rect 735 478 748 512
rect 688 368 748 478
rect 778 580 837 592
rect 778 546 791 580
rect 825 546 837 580
rect 778 444 837 546
rect 778 410 791 444
rect 825 410 837 444
rect 778 368 837 410
<< ndiffc >>
rect 137 86 171 120
rect 226 86 260 120
rect 326 176 360 210
rect 326 86 360 120
rect 426 112 460 146
rect 526 176 560 210
rect 526 86 560 120
rect 612 152 646 186
rect 612 84 646 118
<< pdiffc >>
rect 39 550 73 584
rect 39 482 73 516
rect 39 414 73 448
rect 130 532 164 566
rect 224 380 258 414
rect 317 539 351 573
rect 407 546 441 580
rect 407 463 441 497
rect 407 380 441 414
rect 511 550 545 584
rect 511 482 545 516
rect 611 546 645 580
rect 701 550 735 584
rect 701 478 735 512
rect 791 546 825 580
rect 791 410 825 444
<< poly >>
rect 86 592 116 618
rect 179 592 209 618
rect 274 592 304 618
rect 364 592 394 618
rect 460 592 490 618
rect 568 592 598 618
rect 658 592 688 618
rect 748 592 778 618
rect 86 353 116 368
rect 179 353 209 368
rect 274 353 304 368
rect 364 353 394 368
rect 460 353 490 368
rect 568 353 598 368
rect 658 353 688 368
rect 748 353 778 368
rect 83 300 119 353
rect 176 323 212 353
rect 182 304 212 323
rect 271 304 307 353
rect 361 330 397 353
rect 457 330 493 353
rect 74 284 140 300
rect 74 250 90 284
rect 124 250 140 284
rect 74 234 140 250
rect 182 237 307 304
rect 349 314 415 330
rect 349 280 365 314
rect 399 280 415 314
rect 349 264 415 280
rect 457 314 523 330
rect 457 280 473 314
rect 507 280 523 314
rect 457 264 523 280
rect 565 310 601 353
rect 655 310 691 353
rect 565 294 691 310
rect 182 177 212 237
rect 277 222 307 237
rect 371 222 401 264
rect 485 222 515 264
rect 565 260 635 294
rect 669 260 691 294
rect 565 244 691 260
rect 745 326 781 353
rect 745 310 843 326
rect 745 276 793 310
rect 827 276 843 310
rect 571 222 601 244
rect 745 242 843 276
rect 57 147 212 177
rect 57 132 87 147
rect 21 116 87 132
rect 21 82 37 116
rect 71 82 87 116
rect 21 66 87 82
rect 745 208 793 242
rect 827 208 843 242
rect 745 174 843 208
rect 745 140 793 174
rect 827 140 843 174
rect 745 106 843 140
rect 277 48 307 74
rect 371 48 401 74
rect 485 48 515 74
rect 571 48 601 74
rect 745 72 793 106
rect 827 72 843 106
rect 745 56 843 72
<< polycont >>
rect 90 250 124 284
rect 365 280 399 314
rect 473 280 507 314
rect 635 260 669 294
rect 793 276 827 310
rect 37 82 71 116
rect 793 208 827 242
rect 793 140 827 174
rect 793 72 827 106
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 23 584 73 600
rect 23 550 39 584
rect 23 516 73 550
rect 113 573 367 596
rect 113 566 317 573
rect 113 532 130 566
rect 164 539 317 566
rect 351 539 367 573
rect 164 532 367 539
rect 407 580 457 596
rect 441 546 457 580
rect 23 482 39 516
rect 407 498 457 546
rect 73 497 457 498
rect 73 482 407 497
rect 23 464 407 482
rect 23 448 89 464
rect 23 414 39 448
rect 73 414 89 448
rect 441 463 457 497
rect 495 584 561 600
rect 495 550 511 584
rect 545 550 561 584
rect 495 516 561 550
rect 595 580 661 649
rect 595 546 611 580
rect 645 546 661 580
rect 701 584 751 600
rect 735 550 751 584
rect 495 482 511 516
rect 545 512 561 516
rect 701 512 751 550
rect 545 482 701 512
rect 495 478 701 482
rect 735 478 751 512
rect 788 580 841 596
rect 788 546 791 580
rect 825 546 841 580
rect 407 444 457 463
rect 788 444 841 546
rect 23 402 89 414
rect 123 414 277 430
rect 123 380 224 414
rect 258 380 277 414
rect 123 368 277 380
rect 17 334 277 368
rect 17 200 51 334
rect 313 330 359 430
rect 407 414 791 444
rect 441 410 791 414
rect 825 410 841 444
rect 441 380 457 410
rect 407 364 457 380
rect 491 342 843 376
rect 491 330 525 342
rect 313 314 415 330
rect 313 300 365 314
rect 85 284 365 300
rect 85 250 90 284
rect 124 280 365 284
rect 399 280 415 314
rect 124 264 415 280
rect 457 314 525 330
rect 457 280 473 314
rect 507 280 525 314
rect 777 310 843 342
rect 457 264 525 280
rect 619 294 743 308
rect 124 250 140 264
rect 85 234 140 250
rect 619 260 635 294
rect 669 260 743 294
rect 619 236 743 260
rect 777 276 793 310
rect 827 276 843 310
rect 777 242 843 276
rect 310 210 576 230
rect 310 200 326 210
rect 17 176 326 200
rect 360 196 526 210
rect 360 176 376 196
rect 17 166 376 176
rect 21 116 87 132
rect 310 120 376 166
rect 510 176 526 196
rect 560 176 576 210
rect 777 208 793 242
rect 827 208 843 242
rect 21 82 37 116
rect 71 82 87 116
rect 21 66 87 82
rect 121 86 137 120
rect 171 86 226 120
rect 260 86 276 120
rect 121 17 276 86
rect 310 86 326 120
rect 360 86 376 120
rect 310 70 376 86
rect 410 146 476 162
rect 410 112 426 146
rect 460 112 476 146
rect 410 17 476 112
rect 510 120 576 176
rect 510 86 526 120
rect 560 86 576 120
rect 510 70 576 86
rect 610 186 676 202
rect 610 152 612 186
rect 646 152 676 186
rect 610 118 676 152
rect 610 84 612 118
rect 646 84 676 118
rect 610 17 676 84
rect 777 174 843 208
rect 777 140 793 174
rect 827 140 843 174
rect 777 106 843 140
rect 777 72 793 106
rect 827 72 843 106
rect 777 56 843 72
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel comment s 0 0 0 0 4 nor4_2
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 319 390 353 424 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 703 242 737 276 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 799 94 833 128 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 799 168 833 202 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 799 242 833 276 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 31 94 65 128 0 FreeSans 340 0 0 0 D
port 4 nsew
flabel corelocali s 127 390 161 424 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 223 390 257 424 0 FreeSans 340 0 0 0 Y
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 864 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1677912
string GDS_START 1669792
<< end >>
