magic
tech sky130A
magscale 1 2
timestamp 1599588218
<< nwell >>
rect -38 335 3014 704
rect -38 332 772 335
rect 1177 332 3014 335
rect 1594 319 2508 332
rect 1594 311 1894 319
<< pwell >>
rect 0 0 2976 49
<< scpmos >>
rect 83 464 119 592
rect 274 464 310 592
rect 358 464 394 592
rect 505 483 541 611
rect 589 483 625 611
rect 699 483 735 611
rect 911 387 947 611
rect 1001 387 1037 611
rect 1202 457 1238 541
rect 1292 457 1328 541
rect 1370 457 1406 541
rect 1487 457 1523 541
rect 1682 347 1718 547
rect 1772 347 1808 547
rect 1922 471 1958 555
rect 2006 471 2042 555
rect 2183 471 2219 555
rect 2273 471 2309 555
rect 2380 368 2416 592
rect 2470 368 2506 592
rect 2571 392 2607 592
rect 2769 368 2805 592
rect 2859 368 2895 592
<< nmoslvt >>
rect 84 79 114 163
rect 280 79 310 163
rect 358 79 388 163
rect 517 79 547 163
rect 595 79 625 163
rect 699 79 729 163
rect 909 119 939 267
rect 995 119 1025 267
rect 1193 119 1223 203
rect 1293 119 1323 203
rect 1371 119 1401 203
rect 1449 119 1479 203
rect 1674 74 1704 202
rect 1760 74 1790 202
rect 1970 74 2000 158
rect 2042 74 2072 158
rect 2128 74 2158 158
rect 2200 74 2230 158
rect 2402 74 2432 222
rect 2488 74 2518 222
rect 2583 74 2613 202
rect 2779 74 2809 222
rect 2865 74 2895 222
<< ndiff >>
rect 859 180 909 267
rect 852 167 909 180
rect 27 138 84 163
rect 27 104 39 138
rect 73 104 84 138
rect 27 79 84 104
rect 114 138 169 163
rect 114 104 125 138
rect 159 104 169 138
rect 114 79 169 104
rect 223 138 280 163
rect 223 104 235 138
rect 269 104 280 138
rect 223 79 280 104
rect 310 79 358 163
rect 388 153 517 163
rect 388 119 470 153
rect 504 119 517 153
rect 388 79 517 119
rect 547 79 595 163
rect 625 138 699 163
rect 625 104 636 138
rect 670 104 699 138
rect 625 79 699 104
rect 729 138 790 163
rect 729 104 744 138
rect 778 104 790 138
rect 852 133 864 167
rect 898 133 909 167
rect 852 119 909 133
rect 939 239 995 267
rect 939 205 950 239
rect 984 205 995 239
rect 939 165 995 205
rect 939 131 950 165
rect 984 131 995 165
rect 939 119 995 131
rect 1025 239 1082 267
rect 1025 205 1036 239
rect 1070 205 1082 239
rect 1025 165 1082 205
rect 1025 131 1036 165
rect 1070 131 1082 165
rect 1025 119 1082 131
rect 1136 164 1193 203
rect 1136 130 1148 164
rect 1182 130 1193 164
rect 1136 119 1193 130
rect 1223 177 1293 203
rect 1223 143 1248 177
rect 1282 143 1293 177
rect 1223 119 1293 143
rect 1323 119 1371 203
rect 1401 119 1449 203
rect 1479 202 1611 203
rect 1479 119 1674 202
rect 729 79 790 104
rect 1494 82 1674 119
rect 1494 48 1526 82
rect 1560 74 1674 82
rect 1704 179 1760 202
rect 1704 145 1715 179
rect 1749 145 1760 179
rect 1704 74 1760 145
rect 1790 158 1840 202
rect 1790 131 1970 158
rect 1790 97 1914 131
rect 1948 97 1970 131
rect 1790 74 1970 97
rect 2000 74 2042 158
rect 2072 133 2128 158
rect 2072 99 2083 133
rect 2117 99 2128 133
rect 2072 74 2128 99
rect 2158 74 2200 158
rect 2230 133 2283 158
rect 2230 99 2241 133
rect 2275 99 2283 133
rect 2230 74 2283 99
rect 2337 91 2402 222
rect 1560 48 1593 74
rect 2337 57 2345 91
rect 2379 74 2402 91
rect 2432 190 2488 222
rect 2432 156 2443 190
rect 2477 156 2488 190
rect 2432 120 2488 156
rect 2432 86 2443 120
rect 2477 86 2488 120
rect 2432 74 2488 86
rect 2518 202 2568 222
rect 2720 210 2779 222
rect 2518 194 2583 202
rect 2518 160 2529 194
rect 2563 160 2583 194
rect 2518 126 2583 160
rect 2518 92 2529 126
rect 2563 92 2583 126
rect 2518 74 2583 92
rect 2613 188 2666 202
rect 2613 154 2624 188
rect 2658 154 2666 188
rect 2613 120 2666 154
rect 2613 86 2624 120
rect 2658 86 2666 120
rect 2613 74 2666 86
rect 2720 176 2734 210
rect 2768 176 2779 210
rect 2720 120 2779 176
rect 2720 86 2734 120
rect 2768 86 2779 120
rect 2720 74 2779 86
rect 2809 210 2865 222
rect 2809 176 2820 210
rect 2854 176 2865 210
rect 2809 120 2865 176
rect 2809 86 2820 120
rect 2854 86 2865 120
rect 2809 74 2865 86
rect 2895 210 2949 222
rect 2895 176 2906 210
rect 2940 176 2949 210
rect 2895 120 2949 176
rect 2895 86 2906 120
rect 2940 86 2949 120
rect 2895 74 2949 86
rect 2379 57 2387 74
rect 1494 36 1593 48
rect 2337 45 2387 57
<< pdiff >>
rect 409 592 505 611
rect 27 547 83 592
rect 27 513 39 547
rect 73 513 83 547
rect 27 464 83 513
rect 119 580 274 592
rect 119 546 139 580
rect 173 546 230 580
rect 264 546 274 580
rect 119 464 274 546
rect 310 464 358 592
rect 394 566 505 592
rect 394 532 432 566
rect 466 532 505 566
rect 394 483 505 532
rect 541 483 589 611
rect 625 573 699 611
rect 625 539 639 573
rect 673 539 699 573
rect 625 483 699 539
rect 735 593 795 611
rect 735 559 749 593
rect 783 559 795 593
rect 735 483 795 559
rect 394 464 490 483
rect 855 439 911 611
rect 855 405 867 439
rect 901 405 911 439
rect 855 387 911 405
rect 947 593 1001 611
rect 947 559 957 593
rect 991 559 1001 593
rect 947 387 1001 559
rect 1037 439 1089 611
rect 1037 405 1047 439
rect 1081 405 1089 439
rect 1037 387 1089 405
rect 1421 586 1472 598
rect 1421 552 1430 586
rect 1464 552 1472 586
rect 1421 541 1472 552
rect 2057 582 2168 594
rect 2057 555 2095 582
rect 1872 547 1922 555
rect 1149 522 1202 541
rect 1149 488 1158 522
rect 1192 488 1202 522
rect 1149 457 1202 488
rect 1238 523 1292 541
rect 1238 489 1248 523
rect 1282 489 1292 523
rect 1238 457 1292 489
rect 1328 457 1370 541
rect 1406 457 1487 541
rect 1523 521 1576 541
rect 1523 487 1533 521
rect 1567 487 1576 521
rect 1523 457 1576 487
rect 1630 535 1682 547
rect 1630 501 1638 535
rect 1672 501 1682 535
rect 1630 467 1682 501
rect 1630 433 1638 467
rect 1672 433 1682 467
rect 1630 399 1682 433
rect 1630 365 1638 399
rect 1672 365 1682 399
rect 1630 347 1682 365
rect 1718 535 1772 547
rect 1718 501 1728 535
rect 1762 501 1772 535
rect 1718 467 1772 501
rect 1718 433 1728 467
rect 1762 433 1772 467
rect 1718 399 1772 433
rect 1718 365 1728 399
rect 1762 365 1772 399
rect 1718 347 1772 365
rect 1808 523 1922 547
rect 1808 489 1857 523
rect 1891 489 1922 523
rect 1808 471 1922 489
rect 1958 471 2006 555
rect 2042 548 2095 555
rect 2129 555 2168 582
rect 2328 580 2380 592
rect 2328 555 2336 580
rect 2129 548 2183 555
rect 2042 471 2183 548
rect 2219 530 2273 555
rect 2219 496 2229 530
rect 2263 496 2273 530
rect 2219 471 2273 496
rect 2309 546 2336 555
rect 2370 546 2380 580
rect 2309 495 2380 546
rect 2309 471 2336 495
rect 1808 347 1858 471
rect 2328 461 2336 471
rect 2370 461 2380 495
rect 2328 414 2380 461
rect 2328 380 2336 414
rect 2370 380 2380 414
rect 2328 368 2380 380
rect 2416 580 2470 592
rect 2416 546 2426 580
rect 2460 546 2470 580
rect 2416 498 2470 546
rect 2416 464 2426 498
rect 2460 464 2470 498
rect 2416 414 2470 464
rect 2416 380 2426 414
rect 2460 380 2470 414
rect 2416 368 2470 380
rect 2506 580 2571 592
rect 2506 546 2516 580
rect 2550 546 2571 580
rect 2506 507 2571 546
rect 2506 473 2516 507
rect 2550 473 2571 507
rect 2506 434 2571 473
rect 2506 400 2516 434
rect 2550 400 2571 434
rect 2506 392 2571 400
rect 2607 580 2659 592
rect 2607 546 2617 580
rect 2651 546 2659 580
rect 2607 508 2659 546
rect 2607 474 2617 508
rect 2651 474 2659 508
rect 2607 438 2659 474
rect 2607 404 2617 438
rect 2651 404 2659 438
rect 2607 392 2659 404
rect 2713 580 2769 592
rect 2713 546 2725 580
rect 2759 546 2769 580
rect 2713 497 2769 546
rect 2713 463 2725 497
rect 2759 463 2769 497
rect 2713 414 2769 463
rect 2506 368 2556 392
rect 2713 380 2725 414
rect 2759 380 2769 414
rect 2713 368 2769 380
rect 2805 580 2859 592
rect 2805 546 2815 580
rect 2849 546 2859 580
rect 2805 497 2859 546
rect 2805 463 2815 497
rect 2849 463 2859 497
rect 2805 414 2859 463
rect 2805 380 2815 414
rect 2849 380 2859 414
rect 2805 368 2859 380
rect 2895 580 2949 592
rect 2895 546 2905 580
rect 2939 546 2949 580
rect 2895 497 2949 546
rect 2895 463 2905 497
rect 2939 463 2949 497
rect 2895 414 2949 463
rect 2895 380 2905 414
rect 2939 380 2949 414
rect 2895 368 2949 380
<< ndiffc >>
rect 39 104 73 138
rect 125 104 159 138
rect 235 104 269 138
rect 470 119 504 153
rect 636 104 670 138
rect 744 104 778 138
rect 864 133 898 167
rect 950 205 984 239
rect 950 131 984 165
rect 1036 205 1070 239
rect 1036 131 1070 165
rect 1148 130 1182 164
rect 1248 143 1282 177
rect 1526 48 1560 82
rect 1715 145 1749 179
rect 1914 97 1948 131
rect 2083 99 2117 133
rect 2241 99 2275 133
rect 2345 57 2379 91
rect 2443 156 2477 190
rect 2443 86 2477 120
rect 2529 160 2563 194
rect 2529 92 2563 126
rect 2624 154 2658 188
rect 2624 86 2658 120
rect 2734 176 2768 210
rect 2734 86 2768 120
rect 2820 176 2854 210
rect 2820 86 2854 120
rect 2906 176 2940 210
rect 2906 86 2940 120
<< pdiffc >>
rect 39 513 73 547
rect 139 546 173 580
rect 230 546 264 580
rect 432 532 466 566
rect 639 539 673 573
rect 749 559 783 593
rect 867 405 901 439
rect 957 559 991 593
rect 1047 405 1081 439
rect 1430 552 1464 586
rect 1158 488 1192 522
rect 1248 489 1282 523
rect 1533 487 1567 521
rect 1638 501 1672 535
rect 1638 433 1672 467
rect 1638 365 1672 399
rect 1728 501 1762 535
rect 1728 433 1762 467
rect 1728 365 1762 399
rect 1857 489 1891 523
rect 2095 548 2129 582
rect 2229 496 2263 530
rect 2336 546 2370 580
rect 2336 461 2370 495
rect 2336 380 2370 414
rect 2426 546 2460 580
rect 2426 464 2460 498
rect 2426 380 2460 414
rect 2516 546 2550 580
rect 2516 473 2550 507
rect 2516 400 2550 434
rect 2617 546 2651 580
rect 2617 474 2651 508
rect 2617 404 2651 438
rect 2725 546 2759 580
rect 2725 463 2759 497
rect 2725 380 2759 414
rect 2815 546 2849 580
rect 2815 463 2849 497
rect 2815 380 2849 414
rect 2905 546 2939 580
rect 2905 463 2939 497
rect 2905 380 2939 414
<< poly >>
rect 83 592 119 618
rect 274 592 310 618
rect 358 592 394 618
rect 505 611 541 637
rect 589 611 625 637
rect 699 611 735 637
rect 911 611 947 637
rect 1001 611 1037 637
rect 1104 615 1808 645
rect 83 430 119 464
rect 274 430 310 464
rect 83 414 310 430
rect 83 394 124 414
rect 67 380 124 394
rect 158 380 192 414
rect 226 380 260 414
rect 294 380 310 414
rect 67 364 310 380
rect 67 208 97 364
rect 145 300 310 316
rect 145 266 161 300
rect 195 266 229 300
rect 263 266 310 300
rect 145 250 310 266
rect 358 251 394 464
rect 505 432 541 483
rect 455 416 541 432
rect 455 382 471 416
rect 505 382 541 416
rect 455 366 541 382
rect 589 422 625 483
rect 699 430 735 483
rect 589 406 655 422
rect 589 372 605 406
rect 639 372 655 406
rect 589 338 655 372
rect 481 308 547 324
rect 481 274 497 308
rect 531 274 547 308
rect 589 304 605 338
rect 639 304 655 338
rect 589 288 655 304
rect 699 414 823 430
rect 699 380 773 414
rect 807 380 823 414
rect 699 364 823 380
rect 481 258 547 274
rect 67 178 114 208
rect 84 163 114 178
rect 280 163 310 250
rect 352 235 418 251
rect 352 201 368 235
rect 402 201 418 235
rect 352 185 418 201
rect 358 163 388 185
rect 517 163 547 258
rect 595 163 625 288
rect 699 163 729 364
rect 911 355 947 387
rect 1001 355 1037 387
rect 865 322 947 355
rect 771 306 947 322
rect 771 272 787 306
rect 821 289 947 306
rect 995 339 1061 355
rect 995 305 1011 339
rect 1045 319 1061 339
rect 1104 319 1134 615
rect 1202 541 1238 567
rect 1292 541 1328 615
rect 1370 541 1406 567
rect 1487 541 1523 567
rect 1682 547 1718 573
rect 1772 547 1808 615
rect 2380 592 2416 618
rect 2470 592 2506 618
rect 2571 592 2607 618
rect 2769 592 2805 618
rect 2859 592 2895 618
rect 1922 555 1958 581
rect 2006 555 2042 581
rect 1202 366 1238 457
rect 1292 431 1328 457
rect 1045 305 1134 319
rect 995 289 1134 305
rect 1176 350 1242 366
rect 1176 316 1192 350
rect 1226 330 1242 350
rect 1370 356 1406 457
rect 1487 433 1523 457
rect 1487 409 1598 433
rect 1487 403 1548 409
rect 1532 375 1548 403
rect 1582 375 1598 409
rect 1532 359 1598 375
rect 1370 340 1454 356
rect 1226 316 1323 330
rect 1176 300 1323 316
rect 821 272 837 289
rect 771 238 837 272
rect 909 267 939 289
rect 995 267 1025 289
rect 771 204 787 238
rect 821 204 837 238
rect 771 188 837 204
rect 1104 252 1134 289
rect 1104 222 1223 252
rect 1193 203 1223 222
rect 1293 203 1323 300
rect 1370 306 1404 340
rect 1438 306 1454 340
rect 1370 290 1454 306
rect 1371 203 1401 290
rect 1532 248 1562 359
rect 2183 555 2219 581
rect 2273 555 2309 581
rect 1922 439 1958 471
rect 1890 423 1958 439
rect 1890 389 1906 423
rect 1940 389 1958 423
rect 1890 373 1958 389
rect 2006 439 2042 471
rect 2006 423 2114 439
rect 2183 430 2219 471
rect 2006 389 2064 423
rect 2098 389 2114 423
rect 2006 373 2114 389
rect 2156 414 2222 430
rect 2156 380 2172 414
rect 2206 380 2222 414
rect 1682 315 1718 347
rect 1652 299 1718 315
rect 1652 265 1668 299
rect 1702 265 1718 299
rect 1772 325 1808 347
rect 1772 295 2000 325
rect 1652 249 1718 265
rect 1449 218 1562 248
rect 1449 203 1479 218
rect 1674 202 1704 249
rect 1760 231 1928 247
rect 1760 217 1878 231
rect 1760 202 1790 217
rect 909 93 939 119
rect 995 93 1025 119
rect 1193 93 1223 119
rect 1293 93 1323 119
rect 1371 93 1401 119
rect 84 53 114 79
rect 280 53 310 79
rect 358 53 388 79
rect 517 53 547 79
rect 595 53 625 79
rect 699 51 729 79
rect 1449 51 1479 119
rect 699 21 1479 51
rect 1862 197 1878 217
rect 1912 197 1928 231
rect 1862 181 1928 197
rect 1970 158 2000 295
rect 2042 158 2072 373
rect 2156 364 2222 380
rect 2156 325 2186 364
rect 2128 295 2186 325
rect 2273 318 2309 471
rect 2380 318 2416 368
rect 2273 317 2416 318
rect 2470 317 2506 368
rect 2571 317 2607 392
rect 2769 326 2805 368
rect 2859 326 2895 368
rect 2128 158 2158 295
rect 2273 268 2613 317
rect 2238 252 2613 268
rect 2659 310 2895 326
rect 2659 276 2675 310
rect 2709 276 2743 310
rect 2777 276 2895 310
rect 2659 260 2895 276
rect 2238 232 2254 252
rect 2200 218 2254 232
rect 2288 251 2613 252
rect 2288 218 2309 251
rect 2402 222 2432 251
rect 2488 222 2518 251
rect 2200 202 2309 218
rect 2200 158 2230 202
rect 1674 48 1704 74
rect 1760 48 1790 74
rect 1970 48 2000 74
rect 2042 48 2072 74
rect 2128 48 2158 74
rect 2200 48 2230 74
rect 2583 202 2613 251
rect 2779 222 2809 260
rect 2865 222 2895 260
rect 2402 48 2432 74
rect 2488 48 2518 74
rect 2583 48 2613 74
rect 2779 48 2809 74
rect 2865 48 2895 74
<< polycont >>
rect 124 380 158 414
rect 192 380 226 414
rect 260 380 294 414
rect 161 266 195 300
rect 229 266 263 300
rect 471 382 505 416
rect 605 372 639 406
rect 497 274 531 308
rect 605 304 639 338
rect 773 380 807 414
rect 368 201 402 235
rect 787 272 821 306
rect 1011 305 1045 339
rect 1192 316 1226 350
rect 1548 375 1582 409
rect 787 204 821 238
rect 1404 306 1438 340
rect 1906 389 1940 423
rect 2064 389 2098 423
rect 2172 380 2206 414
rect 1668 265 1702 299
rect 1878 197 1912 231
rect 2675 276 2709 310
rect 2743 276 2777 310
rect 2254 218 2288 252
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 2976 683
rect 23 547 89 596
rect 23 513 39 547
rect 73 513 89 547
rect 123 580 280 649
rect 123 546 139 580
rect 173 546 230 580
rect 264 546 280 580
rect 388 566 589 582
rect 388 532 432 566
rect 466 532 589 566
rect 623 573 689 649
rect 623 539 639 573
rect 673 539 689 573
rect 623 538 689 539
rect 723 593 799 611
rect 723 559 749 593
rect 783 559 799 593
rect 941 593 1007 649
rect 941 559 957 593
rect 991 559 1007 593
rect 1414 586 1464 649
rect 23 498 89 513
rect 555 504 589 532
rect 723 525 799 559
rect 1414 552 1430 586
rect 1142 525 1197 545
rect 723 522 1197 525
rect 723 504 1158 522
rect 23 464 521 498
rect 555 489 1158 504
rect 555 464 799 489
rect 1151 488 1158 489
rect 1192 488 1197 522
rect 23 316 57 464
rect 108 414 359 430
rect 108 380 124 414
rect 158 380 192 414
rect 226 380 260 414
rect 294 380 359 414
rect 108 364 359 380
rect 455 416 521 464
rect 455 382 471 416
rect 505 382 521 416
rect 455 366 521 382
rect 589 406 655 430
rect 589 372 605 406
rect 639 372 655 406
rect 325 324 359 364
rect 589 338 655 372
rect 23 300 279 316
rect 23 266 161 300
rect 195 266 229 300
rect 263 266 279 300
rect 325 308 547 324
rect 325 274 497 308
rect 531 274 547 308
rect 589 304 605 338
rect 639 304 655 338
rect 589 288 655 304
rect 325 272 547 274
rect 23 250 279 266
rect 23 138 73 250
rect 313 235 418 238
rect 689 235 723 464
rect 867 439 917 455
rect 757 424 833 430
rect 757 414 799 424
rect 757 380 773 414
rect 807 380 833 390
rect 757 364 833 380
rect 901 405 917 439
rect 867 398 917 405
rect 1031 439 1117 455
rect 1031 405 1047 439
rect 1081 405 1117 439
rect 867 364 997 398
rect 1031 389 1117 405
rect 1151 434 1197 488
rect 1232 523 1332 545
rect 1414 536 1464 552
rect 1232 489 1248 523
rect 1282 502 1332 523
rect 1510 521 1583 545
rect 1510 502 1533 521
rect 1282 489 1533 502
rect 1232 487 1533 489
rect 1567 487 1583 521
rect 1232 468 1583 487
rect 1151 400 1298 434
rect 881 355 997 364
rect 1081 366 1117 389
rect 881 339 1047 355
rect 313 201 368 235
rect 402 201 418 235
rect 23 104 39 138
rect 23 75 73 104
rect 109 138 175 167
rect 109 104 125 138
rect 159 104 175 138
rect 109 17 175 104
rect 219 138 269 167
rect 313 162 418 201
rect 452 201 723 235
rect 771 306 847 310
rect 771 272 787 306
rect 821 272 847 306
rect 771 238 847 272
rect 771 204 787 238
rect 821 204 847 238
rect 771 201 847 204
rect 881 305 1011 339
rect 1045 305 1047 339
rect 881 289 1047 305
rect 1081 350 1230 366
rect 1081 316 1192 350
rect 1226 316 1230 350
rect 1081 300 1230 316
rect 219 104 235 138
rect 452 153 522 201
rect 881 167 915 289
rect 1081 255 1129 300
rect 1264 258 1298 400
rect 452 119 470 153
rect 504 119 522 153
rect 620 138 686 167
rect 219 85 269 104
rect 620 104 636 138
rect 670 104 686 138
rect 620 85 686 104
rect 219 51 686 85
rect 728 138 794 167
rect 728 104 744 138
rect 778 104 794 138
rect 848 133 864 167
rect 898 133 915 167
rect 848 117 915 133
rect 950 239 984 255
rect 950 165 984 205
rect 728 17 794 104
rect 950 17 984 131
rect 1020 239 1129 255
rect 1020 205 1036 239
rect 1070 205 1129 239
rect 1020 198 1129 205
rect 1164 224 1298 258
rect 1020 165 1086 198
rect 1020 131 1036 165
rect 1070 131 1086 165
rect 1164 164 1198 224
rect 1332 190 1366 468
rect 1476 464 1583 468
rect 1638 535 1688 649
rect 2053 582 2172 649
rect 1672 501 1688 535
rect 1638 467 1688 501
rect 1020 96 1086 131
rect 1132 130 1148 164
rect 1182 130 1198 164
rect 1232 177 1366 190
rect 1400 340 1442 356
rect 1400 306 1404 340
rect 1438 306 1442 340
rect 1400 218 1442 306
rect 1476 315 1510 464
rect 1672 433 1688 467
rect 1544 424 1604 430
rect 1544 409 1567 424
rect 1544 375 1548 409
rect 1601 390 1604 424
rect 1582 375 1604 390
rect 1544 359 1604 375
rect 1638 399 1688 433
rect 1672 365 1688 399
rect 1638 349 1688 365
rect 1728 535 1786 551
rect 2053 548 2095 582
rect 2129 548 2172 582
rect 2320 580 2370 649
rect 1762 501 1786 535
rect 1728 467 1786 501
rect 1820 523 2019 539
rect 2053 532 2172 548
rect 1820 489 1857 523
rect 1891 489 2019 523
rect 2213 530 2279 559
rect 2213 498 2229 530
rect 1820 473 2019 489
rect 1762 433 1786 467
rect 1728 399 1786 433
rect 1762 365 1786 399
rect 1728 349 1786 365
rect 1476 299 1718 315
rect 1476 265 1668 299
rect 1702 265 1718 299
rect 1476 252 1718 265
rect 1752 218 1786 349
rect 1862 423 1951 439
rect 1862 389 1906 423
rect 1940 389 1951 423
rect 1862 373 1951 389
rect 1862 247 1928 373
rect 1400 184 1786 218
rect 1232 143 1248 177
rect 1282 143 1366 177
rect 1699 179 1786 184
rect 1232 130 1366 143
rect 1400 116 1665 150
rect 1699 145 1715 179
rect 1749 145 1786 179
rect 1699 119 1786 145
rect 1820 231 1928 247
rect 1820 197 1878 231
rect 1912 197 1928 231
rect 1820 181 1928 197
rect 1985 262 2019 473
rect 2053 496 2229 498
rect 2263 496 2279 530
rect 2053 464 2279 496
rect 2320 546 2336 580
rect 2320 495 2370 546
rect 2053 423 2109 464
rect 2320 461 2336 495
rect 2053 389 2064 423
rect 2098 389 2109 423
rect 2053 330 2109 389
rect 2143 424 2279 430
rect 2177 414 2279 424
rect 2143 380 2172 390
rect 2206 380 2279 414
rect 2143 364 2279 380
rect 2320 414 2370 461
rect 2320 380 2336 414
rect 2320 364 2370 380
rect 2406 580 2472 596
rect 2406 546 2426 580
rect 2460 546 2472 580
rect 2406 498 2472 546
rect 2406 464 2426 498
rect 2460 464 2472 498
rect 2406 414 2472 464
rect 2406 380 2426 414
rect 2460 380 2472 414
rect 2508 580 2566 649
rect 2508 546 2516 580
rect 2550 546 2566 580
rect 2508 507 2566 546
rect 2508 473 2516 507
rect 2550 473 2566 507
rect 2508 434 2566 473
rect 2508 400 2516 434
rect 2550 400 2566 434
rect 2508 384 2566 400
rect 2613 580 2665 596
rect 2613 546 2617 580
rect 2651 546 2665 580
rect 2613 508 2665 546
rect 2613 474 2617 508
rect 2651 474 2665 508
rect 2613 438 2665 474
rect 2613 404 2617 438
rect 2651 404 2665 438
rect 2053 296 2372 330
rect 1985 252 2304 262
rect 1985 218 2254 252
rect 2288 218 2304 252
rect 1985 209 2304 218
rect 1400 96 1434 116
rect 1020 62 1434 96
rect 1631 85 1665 116
rect 1820 85 1854 181
rect 1985 147 2019 209
rect 2338 175 2372 296
rect 2406 217 2472 380
rect 2613 326 2665 404
rect 2709 580 2775 649
rect 2709 546 2725 580
rect 2759 546 2775 580
rect 2709 497 2775 546
rect 2709 463 2725 497
rect 2759 463 2775 497
rect 2709 414 2775 463
rect 2709 380 2725 414
rect 2759 380 2775 414
rect 2709 364 2775 380
rect 2811 580 2865 596
rect 2811 546 2815 580
rect 2849 546 2865 580
rect 2811 497 2865 546
rect 2811 463 2815 497
rect 2849 463 2865 497
rect 2811 414 2865 463
rect 2811 380 2815 414
rect 2849 380 2865 414
rect 2613 310 2777 326
rect 2613 276 2675 310
rect 2709 276 2743 310
rect 2613 260 2777 276
rect 2406 190 2493 217
rect 2406 183 2443 190
rect 1490 48 1526 82
rect 1560 48 1597 82
rect 1631 51 1854 85
rect 1888 131 2019 147
rect 1888 97 1914 131
rect 1948 97 2019 131
rect 1888 81 2019 97
rect 2067 133 2133 162
rect 2067 99 2083 133
rect 2117 99 2133 133
rect 1490 17 1597 48
rect 2067 17 2133 99
rect 2225 141 2372 175
rect 2427 156 2443 183
rect 2477 156 2493 190
rect 2225 133 2291 141
rect 2225 99 2241 133
rect 2275 99 2291 133
rect 2427 120 2493 156
rect 2225 70 2291 99
rect 2329 91 2379 107
rect 2329 57 2345 91
rect 2427 86 2443 120
rect 2477 86 2493 120
rect 2427 70 2493 86
rect 2527 194 2579 210
rect 2527 160 2529 194
rect 2563 160 2579 194
rect 2527 126 2579 160
rect 2527 92 2529 126
rect 2563 92 2579 126
rect 2329 17 2379 57
rect 2527 17 2579 92
rect 2613 188 2665 260
rect 2613 154 2624 188
rect 2658 154 2665 188
rect 2613 120 2665 154
rect 2613 86 2624 120
rect 2658 86 2665 120
rect 2613 70 2665 86
rect 2734 210 2768 226
rect 2734 120 2768 176
rect 2734 17 2768 86
rect 2811 210 2865 380
rect 2899 580 2955 649
rect 2899 546 2905 580
rect 2939 546 2955 580
rect 2899 497 2955 546
rect 2899 463 2905 497
rect 2939 463 2955 497
rect 2899 414 2955 463
rect 2899 380 2905 414
rect 2939 380 2955 414
rect 2899 364 2955 380
rect 2811 176 2820 210
rect 2854 176 2865 210
rect 2811 120 2865 176
rect 2811 86 2820 120
rect 2854 86 2865 120
rect 2811 70 2865 86
rect 2899 210 2956 226
rect 2899 176 2906 210
rect 2940 176 2956 210
rect 2899 120 2956 176
rect 2899 86 2906 120
rect 2940 86 2956 120
rect 2899 17 2956 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 2976 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 799 414 833 424
rect 799 390 807 414
rect 807 390 833 414
rect 1567 409 1601 424
rect 1567 390 1582 409
rect 1582 390 1601 409
rect 2143 414 2177 424
rect 2143 390 2172 414
rect 2172 390 2177 414
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
<< metal1 >>
rect 0 683 2976 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 2976 683
rect 0 617 2976 649
rect 787 424 845 430
rect 787 390 799 424
rect 833 421 845 424
rect 1555 424 1613 430
rect 1555 421 1567 424
rect 833 393 1567 421
rect 833 390 845 393
rect 787 384 845 390
rect 1555 390 1567 393
rect 1601 421 1613 424
rect 2131 424 2189 430
rect 2131 421 2143 424
rect 1601 393 2143 421
rect 1601 390 1613 393
rect 1555 384 1613 390
rect 2131 390 2143 393
rect 2177 390 2189 424
rect 2131 384 2189 390
rect 0 17 2976 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 2976 17
rect 0 -49 2976 -17
<< labels >>
flabel pwell s 0 0 2976 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nwell s 0 617 2976 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
rlabel comment s 0 0 0 0 4 sdfrbp_2
flabel comment s 1397 630 1397 630 0 FreeSans 300 0 0 0 no_jumper_check
flabel comment s 1086 36 1086 36 0 FreeSans 300 0 0 0 no_jumper_check
flabel metal1 s 2143 390 2177 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew
flabel metal1 s 0 617 2976 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 2976 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 319 168 353 202 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 799 242 833 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 127 390 161 424 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 223 390 257 424 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 319 390 353 424 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 SCD
port 4 nsew
flabel corelocali s 607 390 641 424 0 FreeSans 340 0 0 0 SCD
port 4 nsew
flabel corelocali s 2815 390 2849 424 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2431 168 2465 202 0 FreeSans 340 0 0 0 Q_N
port 11 nsew
flabel corelocali s 2431 242 2465 276 0 FreeSans 340 0 0 0 Q_N
port 11 nsew
flabel corelocali s 2431 316 2465 350 0 FreeSans 340 0 0 0 Q_N
port 11 nsew
<< properties >>
string FIXED_BBOX 0 0 2976 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 21850
string GDS_START 132
<< end >>
