magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 113 299 179 493
rect 295 299 367 493
rect 490 459 959 493
rect 118 265 170 299
rect 295 265 349 299
rect 490 265 530 459
rect 118 213 349 265
rect 118 51 170 213
rect 295 51 349 213
rect 475 199 530 265
rect 632 323 891 357
rect 632 162 666 323
rect 734 51 799 283
rect 833 51 891 323
rect 925 326 959 459
rect 925 288 1075 326
rect 1037 211 1075 288
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 27 299 79 527
rect 213 299 261 527
rect 401 299 456 527
rect 35 17 84 131
rect 211 17 261 131
rect 383 165 417 265
rect 564 391 853 425
rect 564 165 598 391
rect 383 131 598 165
rect 563 124 598 131
rect 383 17 455 97
rect 563 51 700 124
rect 993 367 1039 527
rect 1073 367 1153 493
rect 941 173 975 237
rect 1119 173 1153 367
rect 941 139 1153 173
rect 926 17 1029 105
rect 1083 51 1132 139
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
rlabel locali s 734 51 799 283 6 A0
port 1 nsew signal input
rlabel locali s 833 51 891 323 6 A1
port 2 nsew signal input
rlabel locali s 632 323 891 357 6 A1
port 2 nsew signal input
rlabel locali s 632 162 666 323 6 A1
port 2 nsew signal input
rlabel locali s 1037 211 1075 288 6 S
port 3 nsew signal input
rlabel locali s 925 326 959 459 6 S
port 3 nsew signal input
rlabel locali s 925 288 1075 326 6 S
port 3 nsew signal input
rlabel locali s 490 459 959 493 6 S
port 3 nsew signal input
rlabel locali s 490 265 530 459 6 S
port 3 nsew signal input
rlabel locali s 475 199 530 265 6 S
port 3 nsew signal input
rlabel locali s 295 299 367 493 6 X
port 4 nsew signal output
rlabel locali s 295 265 349 299 6 X
port 4 nsew signal output
rlabel locali s 295 51 349 213 6 X
port 4 nsew signal output
rlabel locali s 118 265 170 299 6 X
port 4 nsew signal output
rlabel locali s 118 213 349 265 6 X
port 4 nsew signal output
rlabel locali s 118 51 170 213 6 X
port 4 nsew signal output
rlabel locali s 113 299 179 493 6 X
port 4 nsew signal output
rlabel metal1 s 0 -48 1196 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 1196 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3293112
string GDS_START 3284120
<< end >>
