magic
tech sky130A
magscale 1 2
timestamp 1604502697
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 79 47 109 131
rect 194 47 224 131
rect 484 47 514 177
rect 568 47 598 177
rect 685 47 715 177
rect 789 47 819 177
<< pmoshvt >>
rect 81 369 117 497
rect 196 369 232 497
rect 394 309 430 497
rect 488 309 524 497
rect 687 297 723 497
rect 781 297 817 497
<< ndiff >>
rect 27 106 79 131
rect 27 72 35 106
rect 69 72 79 106
rect 27 47 79 72
rect 109 89 194 131
rect 109 55 129 89
rect 163 55 194 89
rect 109 47 194 55
rect 224 106 286 131
rect 224 72 244 106
rect 278 72 286 106
rect 224 47 286 72
rect 412 129 484 177
rect 412 95 420 129
rect 454 95 484 129
rect 412 47 484 95
rect 514 89 568 177
rect 514 55 524 89
rect 558 55 568 89
rect 514 47 568 55
rect 598 129 685 177
rect 598 95 629 129
rect 663 95 685 129
rect 598 47 685 95
rect 715 169 789 177
rect 715 135 735 169
rect 769 135 789 169
rect 715 47 789 135
rect 819 93 871 177
rect 819 59 829 93
rect 863 59 871 93
rect 819 47 871 59
<< pdiff >>
rect 27 461 81 497
rect 27 427 35 461
rect 69 427 81 461
rect 27 369 81 427
rect 117 489 196 497
rect 117 455 140 489
rect 174 455 196 489
rect 117 421 196 455
rect 117 387 140 421
rect 174 387 196 421
rect 117 369 196 387
rect 232 461 286 497
rect 232 427 244 461
rect 278 427 286 461
rect 232 369 286 427
rect 340 477 394 497
rect 340 443 348 477
rect 382 443 394 477
rect 340 309 394 443
rect 430 489 488 497
rect 430 455 442 489
rect 476 455 488 489
rect 430 309 488 455
rect 524 477 687 497
rect 524 443 548 477
rect 582 443 626 477
rect 660 443 687 477
rect 524 309 687 443
rect 541 297 687 309
rect 723 416 781 497
rect 723 382 735 416
rect 769 382 781 416
rect 723 348 781 382
rect 723 314 735 348
rect 769 314 781 348
rect 723 297 781 314
rect 817 477 875 497
rect 817 443 833 477
rect 867 443 875 477
rect 817 409 875 443
rect 817 375 833 409
rect 867 375 875 409
rect 817 297 875 375
<< ndiffc >>
rect 35 72 69 106
rect 129 55 163 89
rect 244 72 278 106
rect 420 95 454 129
rect 524 55 558 89
rect 629 95 663 129
rect 735 135 769 169
rect 829 59 863 93
<< pdiffc >>
rect 35 427 69 461
rect 140 455 174 489
rect 140 387 174 421
rect 244 427 278 461
rect 348 443 382 477
rect 442 455 476 489
rect 548 443 582 477
rect 626 443 660 477
rect 735 382 769 416
rect 735 314 769 348
rect 833 443 867 477
rect 833 375 867 409
<< poly >>
rect 81 497 117 523
rect 196 497 232 523
rect 394 497 430 523
rect 488 497 524 523
rect 687 497 723 523
rect 781 497 817 523
rect 81 354 117 369
rect 196 354 232 369
rect 79 265 119 354
rect 194 294 234 354
rect 394 294 430 309
rect 488 294 524 309
rect 79 249 147 265
rect 79 215 103 249
rect 137 215 147 249
rect 79 199 147 215
rect 194 264 526 294
rect 687 282 723 297
rect 781 282 817 297
rect 194 249 260 264
rect 194 215 210 249
rect 244 215 260 249
rect 568 249 627 265
rect 568 222 583 249
rect 194 203 260 215
rect 484 215 583 222
rect 617 215 627 249
rect 79 131 109 199
rect 194 131 224 203
rect 484 192 627 215
rect 685 259 725 282
rect 779 259 819 282
rect 685 249 819 259
rect 685 215 735 249
rect 769 215 819 249
rect 685 205 819 215
rect 484 177 514 192
rect 568 177 598 192
rect 685 177 715 205
rect 789 177 819 205
rect 79 21 109 47
rect 194 21 224 47
rect 484 21 514 47
rect 568 21 598 47
rect 685 21 715 47
rect 789 21 819 47
<< polycont >>
rect 103 215 137 249
rect 210 215 244 249
rect 583 215 617 249
rect 735 215 769 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 17 461 69 493
rect 17 427 35 461
rect 17 246 69 427
rect 103 489 200 527
rect 103 455 140 489
rect 174 455 200 489
rect 103 421 200 455
rect 103 387 140 421
rect 174 387 200 421
rect 103 369 200 387
rect 244 461 302 493
rect 278 427 302 461
rect 244 353 302 427
rect 340 477 382 493
rect 340 443 348 477
rect 416 489 492 527
rect 416 455 442 489
rect 476 455 492 489
rect 536 477 885 493
rect 340 421 382 443
rect 536 443 548 477
rect 582 443 626 477
rect 660 459 833 477
rect 660 443 675 459
rect 536 421 675 443
rect 867 443 885 477
rect 340 387 675 421
rect 719 416 799 425
rect 719 382 735 416
rect 769 382 799 416
rect 719 353 799 382
rect 833 409 885 443
rect 867 375 885 409
rect 833 359 885 375
rect 17 212 30 246
rect 64 212 69 246
rect 17 106 69 212
rect 103 249 155 335
rect 244 289 363 353
rect 397 348 799 353
rect 397 314 735 348
rect 769 325 799 348
rect 769 314 892 325
rect 397 289 892 314
rect 310 255 363 289
rect 137 215 155 249
rect 103 153 155 215
rect 189 249 260 255
rect 189 215 210 249
rect 244 215 260 249
rect 189 153 260 215
rect 310 249 643 255
rect 310 215 583 249
rect 617 215 643 249
rect 310 205 643 215
rect 699 249 791 255
rect 699 215 735 249
rect 769 246 791 249
rect 699 212 736 215
rect 770 212 791 246
rect 699 205 791 212
rect 310 119 366 205
rect 846 171 892 289
rect 17 72 35 106
rect 17 56 69 72
rect 103 89 180 119
rect 103 55 129 89
rect 163 55 180 89
rect 103 17 180 55
rect 214 106 366 119
rect 214 72 244 106
rect 278 72 366 106
rect 214 51 366 72
rect 400 131 675 171
rect 400 129 464 131
rect 400 95 420 129
rect 454 95 464 129
rect 618 129 675 131
rect 400 51 464 95
rect 498 89 574 97
rect 498 55 524 89
rect 558 55 574 89
rect 618 95 629 129
rect 663 95 675 129
rect 709 169 892 171
rect 709 135 735 169
rect 769 135 892 169
rect 709 127 892 135
rect 618 93 675 95
rect 618 59 829 93
rect 863 59 880 93
rect 618 55 880 59
rect 498 17 574 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 30 212 64 246
rect 736 215 769 246
rect 769 215 770 246
rect 736 212 770 215
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 17 246 782 252
rect 17 212 30 246
rect 64 224 736 246
rect 64 212 76 224
rect 17 206 76 212
rect 714 212 736 224
rect 770 212 782 246
rect 714 206 782 212
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel corelocali s 849 221 883 255 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 849 289 883 323 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 121 153 155 187 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 736 357 770 391 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 121 289 155 323 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 210 170 210 170 0 FreeSans 200 0 0 0 TE_B
port 2 nsew
flabel corelocali s 601 306 601 306 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 509 306 509 306 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 419 306 419 306 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 849 153 883 187 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew
rlabel comment s 0 0 0 0 4 ebufn_2
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1980844
string GDS_START 1973424
<< end >>
