magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 828 561
rect 195 435 261 527
rect 507 367 572 527
rect 85 299 614 333
rect 657 299 723 493
rect 757 299 811 527
rect 85 199 155 299
rect 483 283 614 299
rect 201 199 339 265
rect 373 199 431 265
rect 689 181 723 299
rect 195 17 261 97
rect 527 17 593 97
rect 657 51 723 181
rect 757 17 811 181
rect 0 -17 828 17
<< obsli1 >>
rect 17 401 123 493
rect 351 401 417 493
rect 17 367 417 401
rect 17 165 51 367
rect 585 215 655 249
rect 585 165 621 215
rect 17 131 621 165
rect 17 56 105 131
rect 351 51 417 131
<< metal1 >>
rect 0 496 828 592
rect 0 -48 828 48
<< labels >>
rlabel locali s 201 199 339 265 6 A
port 1 nsew signal input
rlabel locali s 373 199 431 265 6 B
port 2 nsew signal input
rlabel locali s 483 283 614 299 6 C
port 3 nsew signal input
rlabel locali s 85 299 614 333 6 C
port 3 nsew signal input
rlabel locali s 85 199 155 299 6 C
port 3 nsew signal input
rlabel locali s 689 181 723 299 6 X
port 4 nsew signal output
rlabel locali s 657 299 723 493 6 X
port 4 nsew signal output
rlabel locali s 657 51 723 181 6 X
port 4 nsew signal output
rlabel locali s 757 17 811 181 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 527 17 593 97 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 195 17 261 97 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 828 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 828 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 757 299 811 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 507 367 572 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 195 435 261 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 828 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 828 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1628674
string GDS_START 1622226
<< end >>
