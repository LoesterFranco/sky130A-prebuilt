magic
tech sky130A
magscale 1 2
timestamp 1604502710
<< nwell >>
rect -38 332 1286 704
<< pwell >>
rect 0 0 1248 49
<< scpmos >>
rect 83 368 119 592
rect 173 368 209 592
rect 263 368 299 592
rect 353 368 389 592
rect 555 368 591 592
rect 645 368 681 592
rect 735 368 771 592
rect 825 368 861 592
rect 1037 368 1073 592
rect 1128 368 1164 592
<< nmoslvt >>
rect 84 74 114 222
rect 170 74 200 222
rect 270 74 300 222
rect 370 74 400 222
rect 470 74 500 222
rect 636 74 666 222
rect 735 74 765 222
rect 831 74 861 222
rect 922 74 952 222
rect 1134 74 1164 222
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 172 170 222
rect 114 138 125 172
rect 159 138 170 172
rect 114 74 170 138
rect 200 149 270 222
rect 200 115 225 149
rect 259 115 270 149
rect 200 74 270 115
rect 300 172 370 222
rect 300 138 325 172
rect 359 138 370 172
rect 300 74 370 138
rect 400 136 470 222
rect 400 102 425 136
rect 459 102 470 136
rect 400 74 470 102
rect 500 84 636 222
rect 500 74 551 84
rect 515 50 551 74
rect 585 74 636 84
rect 666 210 735 222
rect 666 176 677 210
rect 711 176 735 210
rect 666 120 735 176
rect 666 86 677 120
rect 711 86 735 120
rect 666 74 735 86
rect 765 144 831 222
rect 765 110 777 144
rect 811 110 831 144
rect 765 74 831 110
rect 861 210 922 222
rect 861 176 877 210
rect 911 176 922 210
rect 861 120 922 176
rect 861 86 877 120
rect 911 86 922 120
rect 861 74 922 86
rect 952 145 1134 222
rect 952 111 963 145
rect 997 111 1089 145
rect 1123 111 1134 145
rect 952 74 1134 111
rect 1164 210 1221 222
rect 1164 176 1175 210
rect 1209 176 1221 210
rect 1164 120 1221 176
rect 1164 86 1175 120
rect 1209 86 1221 120
rect 1164 74 1221 86
rect 585 50 621 74
rect 515 38 621 50
<< pdiff >>
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 510 83 546
rect 27 476 39 510
rect 73 476 83 510
rect 27 440 83 476
rect 27 406 39 440
rect 73 406 83 440
rect 27 368 83 406
rect 119 531 173 592
rect 119 497 129 531
rect 163 497 173 531
rect 119 440 173 497
rect 119 406 129 440
rect 163 406 173 440
rect 119 368 173 406
rect 209 580 263 592
rect 209 546 219 580
rect 253 546 263 580
rect 209 508 263 546
rect 209 474 219 508
rect 253 474 263 508
rect 209 368 263 474
rect 299 578 353 592
rect 299 544 309 578
rect 343 544 353 578
rect 299 368 353 544
rect 389 580 445 592
rect 389 546 399 580
rect 433 546 445 580
rect 389 508 445 546
rect 389 474 399 508
rect 433 474 445 508
rect 389 368 445 474
rect 499 580 555 592
rect 499 546 511 580
rect 545 546 555 580
rect 499 508 555 546
rect 499 474 511 508
rect 545 474 555 508
rect 499 368 555 474
rect 591 531 645 592
rect 591 497 601 531
rect 635 497 645 531
rect 591 414 645 497
rect 591 380 601 414
rect 635 380 645 414
rect 591 368 645 380
rect 681 580 735 592
rect 681 546 691 580
rect 725 546 735 580
rect 681 510 735 546
rect 681 476 691 510
rect 725 476 735 510
rect 681 440 735 476
rect 681 406 691 440
rect 725 406 735 440
rect 681 368 735 406
rect 771 531 825 592
rect 771 497 781 531
rect 815 497 825 531
rect 771 440 825 497
rect 771 406 781 440
rect 815 406 825 440
rect 771 368 825 406
rect 861 580 917 592
rect 861 546 871 580
rect 905 546 917 580
rect 861 508 917 546
rect 861 474 871 508
rect 905 474 917 508
rect 861 368 917 474
rect 971 580 1037 592
rect 971 546 983 580
rect 1017 546 1037 580
rect 971 508 1037 546
rect 971 474 983 508
rect 1017 474 1037 508
rect 971 368 1037 474
rect 1073 580 1128 592
rect 1073 546 1083 580
rect 1117 546 1128 580
rect 1073 499 1128 546
rect 1073 465 1083 499
rect 1117 465 1128 499
rect 1073 424 1128 465
rect 1073 390 1083 424
rect 1117 390 1128 424
rect 1073 368 1128 390
rect 1164 580 1220 592
rect 1164 546 1174 580
rect 1208 546 1220 580
rect 1164 510 1220 546
rect 1164 476 1174 510
rect 1208 476 1220 510
rect 1164 440 1220 476
rect 1164 406 1174 440
rect 1208 406 1220 440
rect 1164 368 1220 406
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 125 138 159 172
rect 225 115 259 149
rect 325 138 359 172
rect 425 102 459 136
rect 551 50 585 84
rect 677 176 711 210
rect 677 86 711 120
rect 777 110 811 144
rect 877 176 911 210
rect 877 86 911 120
rect 963 111 997 145
rect 1089 111 1123 145
rect 1175 176 1209 210
rect 1175 86 1209 120
<< pdiffc >>
rect 39 546 73 580
rect 39 476 73 510
rect 39 406 73 440
rect 129 497 163 531
rect 129 406 163 440
rect 219 546 253 580
rect 219 474 253 508
rect 309 544 343 578
rect 399 546 433 580
rect 399 474 433 508
rect 511 546 545 580
rect 511 474 545 508
rect 601 497 635 531
rect 601 380 635 414
rect 691 546 725 580
rect 691 476 725 510
rect 691 406 725 440
rect 781 497 815 531
rect 781 406 815 440
rect 871 546 905 580
rect 871 474 905 508
rect 983 546 1017 580
rect 983 474 1017 508
rect 1083 546 1117 580
rect 1083 465 1117 499
rect 1083 390 1117 424
rect 1174 546 1208 580
rect 1174 476 1208 510
rect 1174 406 1208 440
<< poly >>
rect 83 592 119 618
rect 173 592 209 618
rect 263 592 299 618
rect 353 592 389 618
rect 555 592 591 618
rect 645 592 681 618
rect 735 592 771 618
rect 825 592 861 618
rect 1037 592 1073 618
rect 1128 592 1164 618
rect 83 336 119 368
rect 173 336 209 368
rect 66 320 209 336
rect 66 286 82 320
rect 116 286 150 320
rect 184 286 209 320
rect 66 270 209 286
rect 263 336 299 368
rect 353 336 389 368
rect 555 336 591 368
rect 645 336 681 368
rect 263 320 389 336
rect 263 286 313 320
rect 347 300 389 320
rect 470 320 681 336
rect 347 286 400 300
rect 263 270 400 286
rect 84 222 114 270
rect 170 222 200 270
rect 270 222 300 270
rect 370 222 400 270
rect 470 286 486 320
rect 520 306 681 320
rect 735 336 771 368
rect 825 336 861 368
rect 1037 336 1073 368
rect 1128 336 1164 368
rect 735 320 861 336
rect 520 286 666 306
rect 470 270 666 286
rect 470 222 500 270
rect 636 222 666 270
rect 735 286 751 320
rect 785 286 861 320
rect 735 270 861 286
rect 735 222 765 270
rect 831 222 861 270
rect 922 320 1164 336
rect 922 286 938 320
rect 972 286 1006 320
rect 1040 286 1074 320
rect 1108 286 1164 320
rect 922 270 1164 286
rect 922 222 952 270
rect 1134 222 1164 270
rect 84 48 114 74
rect 170 48 200 74
rect 270 48 300 74
rect 370 48 400 74
rect 470 48 500 74
rect 636 48 666 74
rect 735 48 765 74
rect 831 48 861 74
rect 922 48 952 74
rect 1134 48 1164 74
<< polycont >>
rect 82 286 116 320
rect 150 286 184 320
rect 313 286 347 320
rect 486 286 520 320
rect 751 286 785 320
rect 938 286 972 320
rect 1006 286 1040 320
rect 1074 286 1108 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 23 581 253 615
rect 23 580 73 581
rect 23 546 39 580
rect 219 580 253 581
rect 23 510 73 546
rect 23 476 39 510
rect 23 440 73 476
rect 23 406 39 440
rect 23 390 73 406
rect 113 531 179 547
rect 113 497 129 531
rect 163 497 179 531
rect 113 440 179 497
rect 219 508 253 546
rect 293 578 343 649
rect 293 544 309 578
rect 293 526 343 544
rect 383 580 449 596
rect 383 546 399 580
rect 433 546 449 580
rect 383 508 449 546
rect 383 492 399 508
rect 253 474 399 492
rect 433 474 449 508
rect 219 458 449 474
rect 495 581 921 615
rect 495 580 545 581
rect 495 546 511 580
rect 691 580 725 581
rect 495 508 545 546
rect 495 474 511 508
rect 495 458 545 474
rect 585 531 651 547
rect 585 497 601 531
rect 635 497 651 531
rect 113 406 129 440
rect 163 424 179 440
rect 585 424 651 497
rect 163 414 651 424
rect 163 406 601 414
rect 113 390 601 406
rect 585 380 601 390
rect 635 380 651 414
rect 855 580 921 581
rect 691 510 725 546
rect 691 440 725 476
rect 691 390 725 406
rect 765 531 815 547
rect 765 497 781 531
rect 765 440 815 497
rect 855 546 871 580
rect 905 546 921 580
rect 855 508 921 546
rect 855 474 871 508
rect 905 474 921 508
rect 855 458 921 474
rect 967 580 1033 649
rect 967 546 983 580
rect 1017 546 1033 580
rect 967 508 1033 546
rect 967 474 983 508
rect 1017 474 1033 508
rect 967 458 1033 474
rect 1067 580 1134 596
rect 1067 546 1083 580
rect 1117 546 1134 580
rect 1067 499 1134 546
rect 1067 465 1083 499
rect 1117 465 1134 499
rect 765 406 781 440
rect 1067 424 1134 465
rect 815 406 1083 424
rect 765 390 1083 406
rect 1117 390 1134 424
rect 1174 580 1224 649
rect 1208 546 1224 580
rect 1174 510 1224 546
rect 1208 476 1224 510
rect 1174 440 1224 476
rect 1208 406 1224 440
rect 1174 390 1224 406
rect 585 364 651 380
rect 25 320 263 356
rect 25 286 82 320
rect 116 286 150 320
rect 184 286 263 320
rect 25 270 263 286
rect 297 320 363 356
rect 297 286 313 320
rect 347 286 363 320
rect 297 270 363 286
rect 409 320 551 356
rect 409 286 486 320
rect 520 286 551 320
rect 409 270 551 286
rect 585 236 619 364
rect 697 320 839 356
rect 697 286 751 320
rect 785 286 839 320
rect 697 270 839 286
rect 889 320 1223 356
rect 889 286 938 320
rect 972 286 1006 320
rect 1040 286 1074 320
rect 1108 286 1223 320
rect 889 270 1223 286
rect 23 210 73 226
rect 23 176 39 210
rect 23 120 73 176
rect 109 202 619 236
rect 661 210 1225 236
rect 109 172 175 202
rect 109 138 125 172
rect 159 138 175 172
rect 309 172 375 202
rect 109 122 175 138
rect 209 149 275 165
rect 23 86 39 120
rect 23 85 73 86
rect 209 115 225 149
rect 259 115 275 149
rect 309 138 325 172
rect 359 138 375 172
rect 661 176 677 210
rect 711 202 877 210
rect 711 176 727 202
rect 661 168 727 176
rect 309 122 375 138
rect 409 136 727 168
rect 861 176 877 202
rect 911 202 1175 210
rect 911 176 927 202
rect 209 85 275 115
rect 409 102 425 136
rect 459 134 727 136
rect 459 102 475 134
rect 409 85 475 102
rect 661 120 727 134
rect 23 51 475 85
rect 511 84 625 100
rect 511 50 551 84
rect 585 50 625 84
rect 661 86 677 120
rect 711 86 727 120
rect 661 70 727 86
rect 761 144 827 160
rect 761 110 777 144
rect 811 110 827 144
rect 511 17 625 50
rect 761 17 827 110
rect 861 120 927 176
rect 1159 176 1175 202
rect 1209 176 1225 210
rect 861 86 877 120
rect 911 86 927 120
rect 861 70 927 86
rect 961 145 1125 161
rect 961 111 963 145
rect 997 111 1089 145
rect 1123 111 1125 145
rect 961 17 1125 111
rect 1159 120 1225 176
rect 1159 86 1175 120
rect 1209 86 1225 120
rect 1159 70 1225 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
<< metal1 >>
rect 0 683 1248 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 0 617 1248 649
rect 0 17 1248 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
rect 0 -49 1248 -17
<< labels >>
flabel pwell s 0 0 1248 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 0 617 1248 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
rlabel comment s 0 0 0 0 4 o32ai_2
flabel metal1 s 0 617 1248 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 1248 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 B2
port 5 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 B2
port 5 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 B2
port 5 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 B1
port 4 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 1183 316 1217 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 607 390 641 424 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 607 464 641 498 0 FreeSans 340 0 0 0 Y
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 1248 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 638324
string GDS_START 627714
<< end >>
