magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 1050 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 89 47 119 131
rect 184 47 214 177
rect 278 47 308 177
rect 372 47 402 177
rect 466 47 496 177
rect 594 47 624 177
rect 688 47 718 177
rect 784 47 814 177
rect 890 47 920 177
<< pmoshvt >>
rect 81 413 117 497
rect 186 297 222 497
rect 280 297 316 497
rect 374 297 410 497
rect 468 297 504 497
rect 586 297 622 497
rect 680 297 716 497
rect 786 297 822 497
rect 892 297 928 497
<< ndiff >>
rect 134 131 184 177
rect 27 101 89 131
rect 27 67 35 101
rect 69 67 89 101
rect 27 47 89 67
rect 119 93 184 131
rect 119 59 129 93
rect 163 59 184 93
rect 119 47 184 59
rect 214 101 278 177
rect 214 67 234 101
rect 268 67 278 101
rect 214 47 278 67
rect 308 94 372 177
rect 308 60 328 94
rect 362 60 372 94
rect 308 47 372 60
rect 402 101 466 177
rect 402 67 422 101
rect 456 67 466 101
rect 402 47 466 67
rect 496 89 594 177
rect 496 55 523 89
rect 557 55 594 89
rect 496 47 594 55
rect 624 47 688 177
rect 718 47 784 177
rect 814 47 890 177
rect 920 162 972 177
rect 920 128 930 162
rect 964 128 972 162
rect 920 47 972 128
<< pdiff >>
rect 27 477 81 497
rect 27 443 35 477
rect 69 443 81 477
rect 27 413 81 443
rect 117 485 186 497
rect 117 451 129 485
rect 163 451 186 485
rect 117 413 186 451
rect 134 297 186 413
rect 222 343 280 497
rect 222 309 234 343
rect 268 309 280 343
rect 222 297 280 309
rect 316 485 374 497
rect 316 451 328 485
rect 362 451 374 485
rect 316 297 374 451
rect 410 343 468 497
rect 410 309 422 343
rect 456 309 468 343
rect 410 297 468 309
rect 504 485 586 497
rect 504 451 516 485
rect 550 451 586 485
rect 504 297 586 451
rect 622 343 680 497
rect 622 309 634 343
rect 668 309 680 343
rect 622 297 680 309
rect 716 485 786 497
rect 716 451 728 485
rect 762 451 786 485
rect 716 297 786 451
rect 822 343 892 497
rect 822 309 839 343
rect 873 309 892 343
rect 822 297 892 309
rect 928 485 982 497
rect 928 451 940 485
rect 974 451 982 485
rect 928 297 982 451
<< ndiffc >>
rect 35 67 69 101
rect 129 59 163 93
rect 234 67 268 101
rect 328 60 362 94
rect 422 67 456 101
rect 523 55 557 89
rect 930 128 964 162
<< pdiffc >>
rect 35 443 69 477
rect 129 451 163 485
rect 234 309 268 343
rect 328 451 362 485
rect 422 309 456 343
rect 516 451 550 485
rect 634 309 668 343
rect 728 451 762 485
rect 839 309 873 343
rect 940 451 974 485
<< poly >>
rect 81 497 117 523
rect 186 497 222 523
rect 280 497 316 523
rect 374 497 410 523
rect 468 497 504 523
rect 586 497 622 523
rect 680 497 716 523
rect 786 497 822 523
rect 892 497 928 523
rect 81 398 117 413
rect 79 265 119 398
rect 186 282 222 297
rect 280 282 316 297
rect 374 282 410 297
rect 468 282 504 297
rect 586 282 622 297
rect 680 282 716 297
rect 786 282 822 297
rect 892 282 928 297
rect 184 265 224 282
rect 278 265 318 282
rect 372 265 412 282
rect 466 265 504 282
rect 584 265 624 282
rect 678 265 718 282
rect 784 265 824 282
rect 890 265 930 282
rect 78 249 142 265
rect 78 215 88 249
rect 122 215 142 249
rect 78 199 142 215
rect 184 249 502 265
rect 184 215 306 249
rect 340 215 384 249
rect 418 215 452 249
rect 486 215 502 249
rect 184 199 502 215
rect 560 249 624 265
rect 560 215 574 249
rect 608 215 624 249
rect 560 199 624 215
rect 666 249 730 265
rect 666 215 676 249
rect 710 215 730 249
rect 666 199 730 215
rect 784 249 848 265
rect 784 215 794 249
rect 828 215 848 249
rect 784 199 848 215
rect 890 249 987 265
rect 890 215 943 249
rect 977 215 987 249
rect 890 199 987 215
rect 89 131 119 199
rect 184 177 214 199
rect 278 177 308 199
rect 372 177 402 199
rect 466 177 496 199
rect 594 177 624 199
rect 688 177 718 199
rect 784 177 814 199
rect 890 177 920 199
rect 89 21 119 47
rect 184 21 214 47
rect 278 21 308 47
rect 372 21 402 47
rect 466 21 496 47
rect 594 21 624 47
rect 688 21 718 47
rect 784 21 814 47
rect 890 21 920 47
<< polycont >>
rect 88 215 122 249
rect 306 215 340 249
rect 384 215 418 249
rect 452 215 486 249
rect 574 215 608 249
rect 676 215 710 249
rect 794 215 828 249
rect 943 215 977 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 17 477 69 493
rect 17 443 35 477
rect 103 485 179 527
rect 103 451 129 485
rect 163 451 179 485
rect 302 485 378 527
rect 302 451 328 485
rect 362 451 378 485
rect 490 485 566 527
rect 490 451 516 485
rect 550 451 566 485
rect 702 485 778 527
rect 702 451 728 485
rect 762 451 778 485
rect 914 485 990 527
rect 914 451 940 485
rect 974 451 990 485
rect 17 417 69 443
rect 17 383 977 417
rect 17 117 52 383
rect 88 249 168 327
rect 122 215 168 249
rect 88 153 168 215
rect 206 309 234 343
rect 268 309 422 343
rect 456 309 472 343
rect 506 309 634 343
rect 668 309 839 343
rect 873 309 906 343
rect 206 164 272 309
rect 506 265 540 309
rect 306 249 540 265
rect 340 215 384 249
rect 418 215 452 249
rect 486 215 540 249
rect 306 199 540 215
rect 574 249 624 265
rect 608 215 624 249
rect 574 199 624 215
rect 666 249 728 265
rect 666 215 676 249
rect 710 215 728 249
rect 206 130 456 164
rect 666 151 728 215
rect 762 249 838 265
rect 762 215 794 249
rect 828 215 838 249
rect 762 147 838 215
rect 872 162 906 309
rect 943 249 977 383
rect 943 199 977 215
rect 17 101 69 117
rect 17 67 35 101
rect 17 51 69 67
rect 113 93 163 109
rect 113 59 129 93
rect 113 17 163 59
rect 206 101 268 130
rect 206 67 234 101
rect 422 101 456 130
rect 872 128 930 162
rect 964 128 980 162
rect 206 51 268 67
rect 302 60 328 94
rect 362 60 378 94
rect 302 17 378 60
rect 422 51 456 67
rect 507 55 523 89
rect 557 55 573 89
rect 507 17 573 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
flabel corelocali s 231 306 231 306 0 FreeSans 200 0 0 0 X
port 9 nsew
flabel corelocali s 579 221 613 255 0 FreeSans 200 0 0 0 D
port 4 nsew
flabel corelocali s 681 153 715 187 0 FreeSans 200 0 0 0 C
port 3 nsew
flabel corelocali s 681 221 715 255 0 FreeSans 200 0 0 0 C
port 3 nsew
flabel corelocali s 765 221 799 255 0 FreeSans 200 0 0 0 B
port 2 nsew
flabel corelocali s 132 153 166 187 0 FreeSans 200 0 0 0 A_N
port 1 nsew
flabel corelocali s 132 289 166 323 0 FreeSans 200 0 0 0 A_N
port 1 nsew
flabel corelocali s 231 170 231 170 0 FreeSans 200 0 0 0 X
port 9 nsew
flabel corelocali s 132 221 166 255 0 FreeSans 200 0 0 0 A_N
port 1 nsew
flabel corelocali s 231 238 231 238 0 FreeSans 200 0 0 0 X
port 9 nsew
flabel corelocali s 765 153 799 187 0 FreeSans 200 0 0 0 B
port 2 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
rlabel comment s 0 0 0 0 4 and4b_4
<< properties >>
string FIXED_BBOX 0 0 1012 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1597714
string GDS_START 1589860
<< end >>
