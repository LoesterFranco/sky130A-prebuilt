magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 1766 704
<< pwell >>
rect 0 0 1728 49
<< scnmos >>
rect 84 94 114 222
rect 199 74 229 222
rect 285 74 315 222
rect 403 74 433 222
rect 564 74 594 222
rect 666 94 696 222
rect 932 74 962 222
rect 1251 74 1281 222
rect 1380 74 1410 222
rect 1503 74 1533 222
<< pmoshvt >>
rect 86 368 116 568
rect 196 368 226 592
rect 286 368 316 592
rect 395 368 425 592
rect 541 368 571 592
rect 648 368 678 568
rect 850 392 880 592
rect 940 392 970 592
rect 1030 392 1060 592
rect 1130 392 1160 592
rect 1332 392 1362 592
rect 1422 392 1452 592
rect 1512 392 1542 592
rect 1612 392 1642 592
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 140 84 176
rect 27 106 39 140
rect 73 106 84 140
rect 27 94 84 106
rect 114 210 199 222
rect 114 176 139 210
rect 173 176 199 210
rect 114 140 199 176
rect 114 106 139 140
rect 173 106 199 140
rect 114 94 199 106
rect 149 74 199 94
rect 229 210 285 222
rect 229 176 240 210
rect 274 176 285 210
rect 229 120 285 176
rect 229 86 240 120
rect 274 86 285 120
rect 229 74 285 86
rect 315 82 403 222
rect 315 74 342 82
rect 330 48 342 74
rect 376 74 403 82
rect 433 134 564 222
rect 433 100 444 134
rect 478 100 519 134
rect 553 100 564 134
rect 433 74 564 100
rect 594 127 666 222
rect 594 93 605 127
rect 639 94 666 127
rect 696 162 746 222
rect 696 145 753 162
rect 696 111 707 145
rect 741 111 753 145
rect 696 94 753 111
rect 882 94 932 222
rect 639 93 651 94
rect 594 74 651 93
rect 376 48 388 74
rect 807 82 932 94
rect 807 48 845 82
rect 879 74 932 82
rect 962 202 1251 222
rect 962 168 973 202
rect 1007 168 1050 202
rect 1084 168 1129 202
rect 1163 168 1206 202
rect 1240 168 1251 202
rect 962 120 1251 168
rect 962 86 973 120
rect 1007 86 1050 120
rect 1084 86 1129 120
rect 1163 86 1206 120
rect 1240 86 1251 120
rect 962 74 1251 86
rect 1281 184 1380 222
rect 1281 150 1306 184
rect 1340 150 1380 184
rect 1281 116 1380 150
rect 1281 82 1306 116
rect 1340 82 1380 116
rect 1281 74 1380 82
rect 1410 210 1503 222
rect 1410 176 1421 210
rect 1455 176 1503 210
rect 1410 120 1503 176
rect 1410 86 1421 120
rect 1455 86 1503 120
rect 1410 74 1503 86
rect 1533 197 1658 222
rect 1533 163 1544 197
rect 1578 163 1612 197
rect 1646 163 1658 197
rect 1533 120 1658 163
rect 1533 86 1544 120
rect 1578 86 1612 120
rect 1646 86 1658 120
rect 1533 74 1658 86
rect 879 48 917 74
rect 330 36 388 48
rect 807 36 917 48
<< pdiff >>
rect 134 580 196 592
rect 134 568 147 580
rect 27 556 86 568
rect 27 522 39 556
rect 73 522 86 556
rect 27 440 86 522
rect 27 406 39 440
rect 73 406 86 440
rect 27 368 86 406
rect 116 546 147 568
rect 181 546 196 580
rect 116 368 196 546
rect 226 421 286 592
rect 226 387 239 421
rect 273 387 286 421
rect 226 368 286 387
rect 316 580 395 592
rect 316 546 338 580
rect 372 546 395 580
rect 316 368 395 546
rect 425 444 541 592
rect 425 410 446 444
rect 480 410 541 444
rect 425 368 541 410
rect 571 580 630 592
rect 571 546 584 580
rect 618 568 630 580
rect 791 578 850 592
rect 618 546 648 568
rect 571 368 648 546
rect 678 424 737 568
rect 678 390 691 424
rect 725 390 737 424
rect 791 544 803 578
rect 837 544 850 578
rect 791 392 850 544
rect 880 457 940 592
rect 880 423 893 457
rect 927 423 940 457
rect 880 392 940 423
rect 970 578 1030 592
rect 970 544 983 578
rect 1017 544 1030 578
rect 970 392 1030 544
rect 1060 547 1130 592
rect 1060 513 1083 547
rect 1117 513 1130 547
rect 1060 454 1130 513
rect 1060 420 1083 454
rect 1117 420 1130 454
rect 1060 392 1130 420
rect 1160 538 1219 592
rect 1160 504 1173 538
rect 1207 504 1219 538
rect 1160 392 1219 504
rect 1273 538 1332 592
rect 1273 504 1285 538
rect 1319 504 1332 538
rect 1273 392 1332 504
rect 1362 531 1422 592
rect 1362 497 1375 531
rect 1409 497 1422 531
rect 1362 440 1422 497
rect 1362 406 1375 440
rect 1409 406 1422 440
rect 1362 392 1422 406
rect 1452 580 1512 592
rect 1452 546 1465 580
rect 1499 546 1512 580
rect 1452 510 1512 546
rect 1452 476 1465 510
rect 1499 476 1512 510
rect 1452 440 1512 476
rect 1452 406 1465 440
rect 1499 406 1512 440
rect 1452 392 1512 406
rect 1542 584 1612 592
rect 1542 550 1565 584
rect 1599 550 1612 584
rect 1542 516 1612 550
rect 1542 482 1565 516
rect 1599 482 1612 516
rect 1542 392 1612 482
rect 1642 582 1701 592
rect 1642 548 1655 582
rect 1689 548 1701 582
rect 1642 508 1701 548
rect 1642 474 1655 508
rect 1689 474 1701 508
rect 1642 438 1701 474
rect 1642 404 1655 438
rect 1689 404 1701 438
rect 1642 392 1701 404
rect 678 368 737 390
<< ndiffc >>
rect 39 176 73 210
rect 39 106 73 140
rect 139 176 173 210
rect 139 106 173 140
rect 240 176 274 210
rect 240 86 274 120
rect 342 48 376 82
rect 444 100 478 134
rect 519 100 553 134
rect 605 93 639 127
rect 707 111 741 145
rect 845 48 879 82
rect 973 168 1007 202
rect 1050 168 1084 202
rect 1129 168 1163 202
rect 1206 168 1240 202
rect 973 86 1007 120
rect 1050 86 1084 120
rect 1129 86 1163 120
rect 1206 86 1240 120
rect 1306 150 1340 184
rect 1306 82 1340 116
rect 1421 176 1455 210
rect 1421 86 1455 120
rect 1544 163 1578 197
rect 1612 163 1646 197
rect 1544 86 1578 120
rect 1612 86 1646 120
<< pdiffc >>
rect 39 522 73 556
rect 39 406 73 440
rect 147 546 181 580
rect 239 387 273 421
rect 338 546 372 580
rect 446 410 480 444
rect 584 546 618 580
rect 691 390 725 424
rect 803 544 837 578
rect 893 423 927 457
rect 983 544 1017 578
rect 1083 513 1117 547
rect 1083 420 1117 454
rect 1173 504 1207 538
rect 1285 504 1319 538
rect 1375 497 1409 531
rect 1375 406 1409 440
rect 1465 546 1499 580
rect 1465 476 1499 510
rect 1465 406 1499 440
rect 1565 550 1599 584
rect 1565 482 1599 516
rect 1655 548 1689 582
rect 1655 474 1689 508
rect 1655 404 1689 438
<< poly >>
rect 86 568 116 594
rect 196 592 226 618
rect 286 592 316 618
rect 395 592 425 618
rect 541 592 571 618
rect 648 568 678 594
rect 850 592 880 618
rect 940 592 970 618
rect 1030 592 1060 618
rect 1130 592 1160 618
rect 1332 592 1362 618
rect 1422 592 1452 618
rect 1512 592 1542 618
rect 1612 592 1642 618
rect 850 377 880 392
rect 940 377 970 392
rect 1030 377 1060 392
rect 1130 377 1160 392
rect 1332 377 1362 392
rect 1422 377 1452 392
rect 1512 377 1542 392
rect 1612 377 1642 392
rect 86 353 116 368
rect 196 353 226 368
rect 286 353 316 368
rect 395 353 425 368
rect 541 353 571 368
rect 648 353 678 368
rect 83 336 119 353
rect 83 320 151 336
rect 83 286 101 320
rect 135 286 151 320
rect 83 270 151 286
rect 193 313 229 353
rect 283 313 319 353
rect 392 313 428 353
rect 538 313 574 353
rect 645 336 681 353
rect 645 320 741 336
rect 193 297 594 313
rect 193 277 408 297
rect 84 222 114 270
rect 199 263 408 277
rect 442 263 476 297
rect 510 263 544 297
rect 578 263 594 297
rect 645 286 691 320
rect 725 286 741 320
rect 847 294 883 377
rect 937 294 973 377
rect 645 270 741 286
rect 199 247 594 263
rect 199 222 229 247
rect 285 222 315 247
rect 403 222 433 247
rect 564 222 594 247
rect 666 222 696 270
rect 789 237 973 294
rect 1027 318 1063 377
rect 1127 318 1163 377
rect 1027 302 1163 318
rect 1027 268 1043 302
rect 1077 268 1111 302
rect 1145 282 1163 302
rect 1329 356 1365 377
rect 1419 356 1455 377
rect 1329 340 1455 356
rect 1329 306 1345 340
rect 1379 306 1455 340
rect 1509 310 1545 377
rect 1609 310 1645 377
rect 1329 290 1455 306
rect 1503 294 1707 310
rect 1145 268 1281 282
rect 1027 252 1281 268
rect 789 234 855 237
rect 84 68 114 94
rect 199 48 229 74
rect 285 48 315 74
rect 789 200 805 234
rect 839 200 855 234
rect 932 222 962 237
rect 1251 222 1281 252
rect 1380 222 1410 290
rect 1503 260 1521 294
rect 1555 260 1589 294
rect 1623 260 1657 294
rect 1691 260 1707 294
rect 1503 244 1707 260
rect 1503 222 1533 244
rect 789 184 855 200
rect 403 48 433 74
rect 564 48 594 74
rect 666 68 696 94
rect 932 48 962 74
rect 1251 48 1281 74
rect 1380 48 1410 74
rect 1503 48 1533 74
<< polycont >>
rect 101 286 135 320
rect 408 263 442 297
rect 476 263 510 297
rect 544 263 578 297
rect 691 286 725 320
rect 1043 268 1077 302
rect 1111 268 1145 302
rect 1345 306 1379 340
rect 805 200 839 234
rect 1521 260 1555 294
rect 1589 260 1623 294
rect 1657 260 1691 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 130 580 199 649
rect 17 556 89 572
rect 17 522 39 556
rect 73 522 89 556
rect 130 546 147 580
rect 181 546 199 580
rect 313 580 398 649
rect 313 546 338 580
rect 372 546 398 580
rect 568 580 634 649
rect 967 596 1223 615
rect 568 546 584 580
rect 618 546 634 580
rect 787 581 1223 596
rect 787 578 1033 581
rect 787 544 803 578
rect 837 544 983 578
rect 1017 544 1033 578
rect 787 526 1033 544
rect 17 512 89 522
rect 1067 513 1083 547
rect 1117 513 1133 547
rect 17 478 573 512
rect 17 440 89 478
rect 17 406 39 440
rect 73 406 89 440
rect 17 390 89 406
rect 217 421 446 444
rect 17 226 51 390
rect 217 387 239 421
rect 273 410 446 421
rect 480 410 505 444
rect 273 387 290 410
rect 85 320 167 356
rect 85 286 101 320
rect 135 286 167 320
rect 85 270 167 286
rect 217 236 290 387
rect 539 376 573 478
rect 17 210 89 226
rect 17 176 39 210
rect 73 176 89 210
rect 17 140 89 176
rect 17 106 39 140
rect 73 106 89 140
rect 17 90 89 106
rect 123 210 183 226
rect 123 176 139 210
rect 173 176 183 210
rect 123 140 183 176
rect 123 106 139 140
rect 173 106 183 140
rect 123 17 183 106
rect 224 210 290 236
rect 224 176 240 210
rect 274 176 290 210
rect 324 342 573 376
rect 607 458 943 492
rect 324 218 358 342
rect 607 308 641 458
rect 877 457 943 458
rect 675 390 691 424
rect 725 390 811 424
rect 392 297 641 308
rect 392 263 408 297
rect 442 263 476 297
rect 510 263 544 297
rect 578 263 641 297
rect 675 320 743 356
rect 675 286 691 320
rect 725 286 743 320
rect 675 270 743 286
rect 777 318 811 390
rect 877 423 893 457
rect 927 423 943 457
rect 877 386 943 423
rect 1067 454 1133 513
rect 1173 538 1223 581
rect 1207 504 1223 538
rect 1173 488 1223 504
rect 1269 581 1515 615
rect 1269 538 1335 581
rect 1449 580 1515 581
rect 1269 504 1285 538
rect 1319 504 1335 538
rect 1269 488 1335 504
rect 1375 531 1409 547
rect 1375 454 1409 497
rect 1067 420 1083 454
rect 1117 440 1409 454
rect 1117 420 1375 440
rect 1315 406 1375 420
rect 1315 390 1409 406
rect 1449 546 1465 580
rect 1499 546 1515 580
rect 1449 510 1515 546
rect 1449 476 1465 510
rect 1499 476 1515 510
rect 1549 584 1615 649
rect 1549 550 1565 584
rect 1599 550 1615 584
rect 1549 516 1615 550
rect 1549 482 1565 516
rect 1599 482 1615 516
rect 1650 582 1705 598
rect 1650 548 1655 582
rect 1689 548 1705 582
rect 1650 508 1705 548
rect 1449 448 1515 476
rect 1650 474 1655 508
rect 1689 474 1705 508
rect 1650 448 1705 474
rect 1449 440 1705 448
rect 1449 406 1465 440
rect 1499 438 1705 440
rect 1499 406 1655 438
rect 1449 404 1655 406
rect 1689 404 1705 438
rect 1449 390 1705 404
rect 1639 388 1705 390
rect 877 352 1229 386
rect 777 302 1161 318
rect 777 284 1043 302
rect 392 252 641 263
rect 889 268 1043 284
rect 1077 268 1111 302
rect 1145 268 1161 302
rect 889 252 1161 268
rect 1195 252 1229 352
rect 1273 340 1415 356
rect 1273 306 1345 340
rect 1379 306 1415 340
rect 1273 290 1415 306
rect 1505 294 1707 310
rect 1505 260 1521 294
rect 1555 260 1589 294
rect 1623 260 1657 294
rect 1691 260 1707 294
rect 789 234 855 250
rect 789 218 805 234
rect 324 200 805 218
rect 839 200 855 234
rect 324 184 855 200
rect 224 150 290 176
rect 889 150 923 252
rect 1195 218 1471 252
rect 1505 236 1707 260
rect 224 134 555 150
rect 224 120 444 134
rect 224 86 240 120
rect 274 116 444 120
rect 274 86 290 116
rect 224 70 290 86
rect 428 100 444 116
rect 478 100 519 134
rect 553 100 555 134
rect 428 84 555 100
rect 589 127 655 150
rect 589 93 605 127
rect 639 93 655 127
rect 326 48 342 82
rect 376 48 392 82
rect 326 17 392 48
rect 589 17 655 93
rect 691 145 923 150
rect 691 111 707 145
rect 741 116 923 145
rect 957 202 1256 218
rect 957 168 973 202
rect 1007 168 1050 202
rect 1084 168 1129 202
rect 1163 168 1206 202
rect 1240 168 1256 202
rect 1405 210 1471 218
rect 957 120 1256 168
rect 741 111 757 116
rect 691 90 757 111
rect 957 86 973 120
rect 1007 86 1050 120
rect 1084 86 1129 120
rect 1163 86 1206 120
rect 1240 86 1256 120
rect 803 48 845 82
rect 879 48 921 82
rect 957 70 1256 86
rect 1290 150 1306 184
rect 1340 150 1356 184
rect 1290 116 1356 150
rect 1290 82 1306 116
rect 1340 82 1356 116
rect 803 17 921 48
rect 1290 17 1356 82
rect 1405 176 1421 210
rect 1455 176 1471 210
rect 1405 120 1471 176
rect 1405 86 1421 120
rect 1455 86 1471 120
rect 1405 70 1471 86
rect 1528 163 1544 197
rect 1578 163 1612 197
rect 1646 163 1662 197
rect 1528 120 1662 163
rect 1528 86 1544 120
rect 1578 86 1612 120
rect 1646 86 1662 120
rect 1528 17 1662 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
<< metal1 >>
rect 0 683 1728 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 0 617 1728 649
rect 0 17 1728 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
rect 0 -49 1728 -17
<< labels >>
rlabel comment s 0 0 0 0 4 or4bb_4
flabel pwell s 0 0 1728 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nwell s 0 617 1728 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 1728 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 1728 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 D_N
port 4 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 C_N
port 3 nsew
flabel corelocali s 1567 242 1601 276 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 1663 242 1697 276 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 223 242 257 276 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 223 390 257 424 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 1279 316 1313 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 1375 316 1409 350 0 FreeSans 340 0 0 0 B
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 1728 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1149582
string GDS_START 1136766
<< end >>
