magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 17 51 69 493
rect 103 447 179 527
rect 189 199 265 323
rect 299 199 346 275
rect 631 435 683 527
rect 579 208 631 331
rect 673 153 725 331
rect 103 17 199 106
rect 334 17 478 97
rect 698 17 788 119
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< obsli1 >>
rect 426 474 477 493
rect 231 440 477 474
rect 521 451 589 485
rect 231 395 275 440
rect 103 361 275 395
rect 426 413 477 440
rect 103 199 137 361
rect 338 343 372 381
rect 426 379 520 413
rect 338 309 442 343
rect 408 165 442 309
rect 253 131 442 165
rect 476 174 520 379
rect 555 401 589 451
rect 727 401 763 493
rect 555 367 763 401
rect 476 140 571 174
rect 253 51 287 131
rect 537 51 571 140
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
rlabel locali s 189 199 265 323 6 A1_N
port 1 nsew signal input
rlabel locali s 299 199 346 275 6 A2_N
port 2 nsew signal input
rlabel locali s 673 153 725 331 6 B1
port 3 nsew signal input
rlabel locali s 579 208 631 331 6 B2
port 4 nsew signal input
rlabel locali s 17 51 69 493 6 X
port 5 nsew signal output
rlabel metal1 s 0 -48 828 48 8 VGND
port 6 nsew ground bidirectional
rlabel locali s 698 17 788 119 6 VGND
port 6 nsew ground bidirectional
rlabel locali s 334 17 478 97 6 VGND
port 6 nsew ground bidirectional
rlabel locali s 103 17 199 106 6 VGND
port 6 nsew ground bidirectional
rlabel locali s 0 -17 828 17 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 828 592 6 VPWR
port 7 nsew power bidirectional
rlabel locali s 631 435 683 527 6 VPWR
port 7 nsew power bidirectional
rlabel locali s 103 447 179 527 6 VPWR
port 7 nsew power bidirectional
rlabel locali s 0 527 828 561 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1311918
string GDS_START 1304590
<< end >>
