magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 25 222 121 356
rect 383 238 455 578
rect 650 364 751 596
rect 503 260 569 356
rect 717 226 751 364
rect 679 70 751 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 23 420 89 649
rect 123 420 189 596
rect 155 376 189 420
rect 155 242 241 376
rect 155 188 189 242
rect 275 204 341 595
rect 550 390 616 649
rect 611 260 683 326
rect 611 204 645 260
rect 23 17 89 188
rect 123 70 189 188
rect 235 170 645 204
rect 235 70 301 170
rect 335 17 401 136
rect 435 70 501 170
rect 535 17 645 136
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel locali s 503 260 569 356 6 A
port 1 nsew signal input
rlabel locali s 383 238 455 578 6 B
port 2 nsew signal input
rlabel locali s 25 222 121 356 6 C_N
port 3 nsew signal input
rlabel locali s 717 226 751 364 6 X
port 4 nsew signal output
rlabel locali s 679 70 751 226 6 X
port 4 nsew signal output
rlabel locali s 650 364 751 596 6 X
port 4 nsew signal output
rlabel metal1 s 0 -49 768 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 617 768 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 820256
string GDS_START 813042
<< end >>
