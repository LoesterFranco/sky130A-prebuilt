magic
tech sky130A
magscale 1 2
timestamp 1604502741
<< locali >>
rect 109 398 180 547
rect 304 398 370 547
rect 484 398 550 547
rect 674 398 740 547
rect 109 364 740 398
rect 109 230 167 364
rect 109 196 752 230
rect 109 119 175 196
rect 286 119 352 196
rect 486 119 552 196
rect 686 119 752 196
rect 1653 236 1895 310
rect 1929 236 1995 310
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 24 581 840 615
rect 24 364 74 581
rect 217 432 270 581
rect 410 432 444 581
rect 584 432 638 581
rect 774 512 840 581
rect 874 546 940 649
rect 974 512 1040 596
rect 1074 546 1140 649
rect 1174 512 1240 596
rect 1274 546 1340 649
rect 1374 546 1440 596
rect 1481 580 1547 649
rect 1588 546 1654 596
rect 1374 512 1654 546
rect 1833 512 1899 649
rect 774 478 1440 512
rect 1933 478 1989 596
rect 1517 444 1989 478
rect 774 410 1551 444
rect 774 330 808 410
rect 207 296 808 330
rect 1585 360 1809 410
rect 1933 378 1989 444
rect 2023 412 2089 649
rect 207 264 731 296
rect 944 262 1510 294
rect 788 260 1510 262
rect 23 85 73 226
rect 211 85 245 162
rect 386 85 452 162
rect 586 85 652 162
rect 788 228 1010 260
rect 788 85 822 228
rect 23 51 822 85
rect 858 17 924 194
rect 960 70 1010 228
rect 1046 17 1080 226
rect 1116 70 1166 260
rect 1202 17 1252 226
rect 1288 70 1338 260
rect 1374 17 1424 226
rect 1460 70 1510 260
rect 1585 202 1619 360
rect 1933 344 2063 378
rect 2029 202 2063 344
rect 1585 134 1830 202
rect 1544 68 1830 134
rect 1866 17 1900 202
rect 1936 168 2063 202
rect 1936 68 1986 168
rect 2022 17 2089 120
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
<< metal1 >>
rect 0 683 2112 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 0 617 2112 649
rect 0 17 2112 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
rect 0 -49 2112 -17
<< labels >>
rlabel locali s 1929 236 1995 310 6 A
port 1 nsew signal input
rlabel locali s 1653 236 1895 310 6 TE_B
port 2 nsew signal input
rlabel locali s 686 119 752 196 6 Z
port 3 nsew signal output
rlabel locali s 674 398 740 547 6 Z
port 3 nsew signal output
rlabel locali s 486 119 552 196 6 Z
port 3 nsew signal output
rlabel locali s 484 398 550 547 6 Z
port 3 nsew signal output
rlabel locali s 304 398 370 547 6 Z
port 3 nsew signal output
rlabel locali s 286 119 352 196 6 Z
port 3 nsew signal output
rlabel locali s 109 398 180 547 6 Z
port 3 nsew signal output
rlabel locali s 109 364 740 398 6 Z
port 3 nsew signal output
rlabel locali s 109 230 167 364 6 Z
port 3 nsew signal output
rlabel locali s 109 196 752 230 6 Z
port 3 nsew signal output
rlabel locali s 109 119 175 196 6 Z
port 3 nsew signal output
rlabel metal1 s 0 -49 2112 49 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 617 2112 715 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2112 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 2344920
string GDS_START 2330498
<< end >>
