magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 2852 561
rect 26 299 107 527
rect 17 215 123 264
rect 687 367 737 527
rect 839 367 905 527
rect 1031 299 1097 493
rect 49 17 107 181
rect 1203 299 1269 493
rect 1375 299 1441 493
rect 1475 347 1520 492
rect 1554 381 1606 493
rect 1640 347 1692 492
rect 1726 381 1778 493
rect 1812 347 1864 492
rect 1898 381 1950 493
rect 1984 347 2036 492
rect 2070 381 2119 493
rect 2153 347 2205 492
rect 2242 381 2291 493
rect 2325 347 2377 492
rect 2414 381 2463 493
rect 2497 347 2549 492
rect 2586 381 2637 493
rect 1475 344 2549 347
rect 2671 344 2729 492
rect 2763 378 2817 493
rect 1475 299 2817 344
rect 652 215 940 255
rect 243 17 301 181
rect 435 17 469 111
rect 603 17 637 111
rect 771 17 805 111
rect 939 113 995 181
rect 939 17 1090 113
rect 1210 17 1262 122
rect 2584 181 2817 299
rect 1468 147 2817 181
rect 1382 17 1434 129
rect 1468 56 1520 147
rect 1554 17 1606 113
rect 1640 56 1692 147
rect 1726 17 1778 113
rect 1812 56 1864 147
rect 1898 17 1947 113
rect 1981 56 2036 147
rect 2070 17 2119 113
rect 2153 56 2205 147
rect 2241 17 2291 113
rect 2325 56 2377 147
rect 2413 17 2463 113
rect 2497 56 2549 147
rect 2585 17 2637 113
rect 2671 56 2723 147
rect 2757 17 2817 113
rect 0 -17 2852 17
<< obsli1 >>
rect 141 315 207 493
rect 241 459 653 493
rect 241 315 317 459
rect 351 349 385 425
rect 419 387 485 459
rect 519 349 553 425
rect 157 255 207 315
rect 351 289 553 349
rect 587 333 653 459
rect 771 333 805 493
rect 939 333 995 493
rect 587 291 995 333
rect 157 215 453 255
rect 157 163 207 215
rect 487 193 553 289
rect 1131 265 1169 493
rect 1303 265 1341 492
rect 487 187 619 193
rect 487 181 505 187
rect 141 51 207 163
rect 335 153 505 181
rect 539 153 577 187
rect 611 181 619 187
rect 1029 187 1092 265
rect 611 153 905 181
rect 335 145 905 153
rect 335 51 401 145
rect 503 51 569 145
rect 671 51 737 145
rect 839 51 905 145
rect 1029 153 1042 187
rect 1076 153 1092 187
rect 1029 147 1092 153
rect 1131 215 2550 265
rect 1131 53 1176 215
rect 1298 53 1348 215
<< obsli1c >>
rect 505 153 539 187
rect 577 153 611 187
rect 1042 153 1076 187
<< metal1 >>
rect 0 496 2852 592
rect 14 428 2838 468
rect 1035 416 1093 428
rect 1207 416 1265 428
rect 1378 416 1436 428
rect 1548 416 1606 428
rect 1724 416 1782 428
rect 1896 416 1954 428
rect 2067 416 2125 428
rect 2239 416 2297 428
rect 2410 416 2468 428
rect 2580 416 2638 428
rect 2756 416 2814 428
rect 0 -48 2852 48
<< obsm1 >>
rect 493 187 623 193
rect 493 153 505 187
rect 539 153 577 187
rect 611 184 623 187
rect 1030 187 1088 193
rect 1030 184 1042 187
rect 611 156 1042 184
rect 611 153 623 156
rect 493 147 623 153
rect 1030 153 1042 156
rect 1076 153 1088 187
rect 1030 147 1088 153
<< labels >>
rlabel locali s 17 215 123 264 6 A
port 1 nsew signal input
rlabel locali s 652 215 940 255 6 SLEEP
port 2 nsew signal input
rlabel locali s 2671 344 2729 492 6 X
port 3 nsew signal output
rlabel locali s 2671 56 2723 147 6 X
port 3 nsew signal output
rlabel locali s 2584 181 2817 299 6 X
port 3 nsew signal output
rlabel locali s 2497 347 2549 492 6 X
port 3 nsew signal output
rlabel locali s 2497 56 2549 147 6 X
port 3 nsew signal output
rlabel locali s 2325 347 2377 492 6 X
port 3 nsew signal output
rlabel locali s 2325 56 2377 147 6 X
port 3 nsew signal output
rlabel locali s 2153 347 2205 492 6 X
port 3 nsew signal output
rlabel locali s 2153 56 2205 147 6 X
port 3 nsew signal output
rlabel locali s 1984 347 2036 492 6 X
port 3 nsew signal output
rlabel locali s 1981 56 2036 147 6 X
port 3 nsew signal output
rlabel locali s 1812 347 1864 492 6 X
port 3 nsew signal output
rlabel locali s 1812 56 1864 147 6 X
port 3 nsew signal output
rlabel locali s 1640 347 1692 492 6 X
port 3 nsew signal output
rlabel locali s 1640 56 1692 147 6 X
port 3 nsew signal output
rlabel locali s 1475 347 1520 492 6 X
port 3 nsew signal output
rlabel locali s 1475 344 2549 347 6 X
port 3 nsew signal output
rlabel locali s 1475 299 2817 344 6 X
port 3 nsew signal output
rlabel locali s 1468 147 2817 181 6 X
port 3 nsew signal output
rlabel locali s 1468 56 1520 147 6 X
port 3 nsew signal output
rlabel locali s 2070 381 2119 493 6 KAPWR
port 4 nsew power bidirectional abutment
rlabel locali s 2242 381 2291 493 6 KAPWR
port 4 nsew power bidirectional abutment
rlabel locali s 2414 381 2463 493 6 KAPWR
port 4 nsew power bidirectional abutment
rlabel locali s 2586 381 2637 493 6 KAPWR
port 4 nsew power bidirectional abutment
rlabel locali s 2763 378 2817 493 6 KAPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1031 299 1097 493 6 KAPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1203 299 1269 493 6 KAPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1375 299 1441 493 6 KAPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1554 381 1606 493 6 KAPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1726 381 1778 493 6 KAPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1898 381 1950 493 6 KAPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 2756 416 2814 428 6 KAPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 2580 416 2638 428 6 KAPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 2410 416 2468 428 6 KAPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 2239 416 2297 428 6 KAPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 2067 416 2125 428 6 KAPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 1896 416 1954 428 6 KAPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 1724 416 1782 428 6 KAPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 1548 416 1606 428 6 KAPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 1378 416 1436 428 6 KAPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 1207 416 1265 428 6 KAPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 1035 416 1093 428 6 KAPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 14 428 2838 468 6 KAPWR
port 4 nsew power bidirectional abutment
rlabel locali s 2757 17 2817 113 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 2585 17 2637 113 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 2413 17 2463 113 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 2241 17 2291 113 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 2070 17 2119 113 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 1898 17 1947 113 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 1726 17 1778 113 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 1554 17 1606 113 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 1382 17 1434 129 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 1210 17 1262 122 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 939 113 995 181 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 939 17 1090 113 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 771 17 805 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 603 17 637 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 435 17 469 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 243 17 301 181 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 49 17 107 181 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 2852 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 2852 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 839 367 905 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 687 367 737 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 26 299 107 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 2852 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 2852 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2852 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2399020
string GDS_START 2377104
<< end >>
