magic
tech sky130A
magscale 1 2
timestamp 1601050088
<< locali >>
rect 85 236 167 354
rect 201 233 267 578
rect 309 270 375 578
rect 572 394 638 596
rect 572 360 743 394
rect 409 270 491 356
rect 697 226 743 360
rect 593 192 743 226
rect 593 70 643 192
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 81 422 147 596
rect 17 388 147 422
rect 17 199 51 388
rect 472 390 538 649
rect 672 428 738 649
rect 525 260 608 326
rect 525 236 559 260
rect 372 202 559 236
rect 372 199 438 202
rect 17 165 438 199
rect 23 17 102 131
rect 138 70 204 165
rect 240 17 336 131
rect 372 70 438 165
rect 472 17 559 165
rect 679 17 745 155
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel locali s 409 270 491 356 6 A
port 1 nsew signal input
rlabel locali s 309 270 375 578 6 B
port 2 nsew signal input
rlabel locali s 201 233 267 578 6 C
port 3 nsew signal input
rlabel locali s 85 236 167 354 6 D
port 4 nsew signal input
rlabel locali s 697 226 743 360 6 X
port 5 nsew signal output
rlabel locali s 593 192 743 226 6 X
port 5 nsew signal output
rlabel locali s 593 70 643 192 6 X
port 5 nsew signal output
rlabel locali s 572 394 638 596 6 X
port 5 nsew signal output
rlabel locali s 572 360 743 394 6 X
port 5 nsew signal output
rlabel metal1 s 0 -49 768 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 768 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 808034
string GDS_START 800782
<< end >>
