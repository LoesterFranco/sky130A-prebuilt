magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 149 409 183 493
rect 337 409 371 493
rect 149 291 371 409
rect 149 288 314 291
rect 241 185 314 288
rect 129 132 351 185
rect 129 70 163 132
rect 317 70 351 132
rect 626 199 763 265
rect 1651 289 1728 323
rect 1651 199 1695 289
rect 1835 215 1927 265
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 55 427 89 527
rect 227 443 293 527
rect 415 443 481 527
rect 515 447 843 481
rect 896 447 977 481
rect 1011 447 1077 527
rect 1164 455 1823 489
rect 1923 455 1989 527
rect 515 409 559 447
rect 943 413 977 447
rect 1164 413 1198 455
rect 415 375 559 409
rect 628 379 909 413
rect 943 379 1198 413
rect 415 265 449 375
rect 514 307 831 341
rect 404 193 449 265
rect 415 173 449 193
rect 415 139 513 173
rect 35 17 69 109
rect 197 17 273 93
rect 411 17 445 105
rect 479 85 513 139
rect 558 119 592 307
rect 797 265 831 307
rect 875 339 909 379
rect 875 305 981 339
rect 924 275 981 305
rect 797 199 881 265
rect 648 131 890 165
rect 732 85 812 91
rect 479 51 812 85
rect 846 85 890 131
rect 924 119 958 275
rect 1015 241 1049 379
rect 1095 289 1198 343
rect 992 210 1049 241
rect 992 209 1048 210
rect 992 208 1046 209
rect 992 207 1043 208
rect 992 85 1026 207
rect 846 51 1026 85
rect 1060 17 1094 177
rect 1140 83 1198 289
rect 1233 119 1267 421
rect 1305 178 1339 455
rect 2033 421 2085 493
rect 1383 323 1466 409
rect 1583 387 2085 421
rect 1383 289 1549 323
rect 1386 199 1471 254
rect 1305 165 1355 178
rect 1305 144 1394 165
rect 1311 131 1394 144
rect 1233 97 1277 119
rect 1233 53 1316 97
rect 1360 64 1394 131
rect 1428 126 1471 199
rect 1515 85 1549 289
rect 1583 119 1617 387
rect 1978 375 2085 387
rect 1821 299 1995 341
rect 1961 265 1995 299
rect 1729 189 1791 255
rect 1961 199 2007 265
rect 1729 146 1770 189
rect 1961 181 1995 199
rect 1837 150 1995 181
rect 1829 147 1995 150
rect 1651 85 1754 93
rect 1515 51 1754 85
rect 1829 59 1887 147
rect 2051 117 2085 375
rect 1939 17 1973 113
rect 2033 51 2085 117
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
<< metal1 >>
rect 0 561 2116 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 0 496 2116 527
rect 0 17 2116 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
rect 0 -48 2116 -17
<< obsm1 >>
rect 935 320 993 329
rect 1425 320 1483 329
rect 935 292 1483 320
rect 935 283 993 292
rect 1425 283 1483 292
rect 1129 184 1197 193
rect 1425 184 1483 193
rect 1721 184 1779 193
rect 1129 156 1779 184
rect 1129 147 1197 156
rect 1425 147 1483 156
rect 1721 147 1779 156
rect 1231 116 1289 125
rect 1823 116 1881 125
rect 1231 88 1881 116
rect 1231 79 1289 88
rect 1823 79 1881 88
<< labels >>
rlabel locali s 1835 215 1927 265 6 A
port 1 nsew signal input
rlabel locali s 1651 289 1728 323 6 B
port 2 nsew signal input
rlabel locali s 1651 199 1695 289 6 B
port 2 nsew signal input
rlabel locali s 626 199 763 265 6 C
port 3 nsew signal input
rlabel locali s 337 409 371 493 6 X
port 4 nsew signal output
rlabel locali s 317 70 351 132 6 X
port 4 nsew signal output
rlabel locali s 241 185 314 288 6 X
port 4 nsew signal output
rlabel locali s 149 409 183 493 6 X
port 4 nsew signal output
rlabel locali s 149 291 371 409 6 X
port 4 nsew signal output
rlabel locali s 149 288 314 291 6 X
port 4 nsew signal output
rlabel locali s 129 132 351 185 6 X
port 4 nsew signal output
rlabel locali s 129 70 163 132 6 X
port 4 nsew signal output
rlabel metal1 s 0 -48 2116 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 2116 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2116 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 820024
string GDS_START 806038
<< end >>
