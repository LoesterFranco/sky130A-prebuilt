magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 920 561
rect 17 327 87 527
rect 17 17 87 177
rect 121 51 179 478
rect 213 299 263 527
rect 392 265 451 471
rect 213 89 265 173
rect 377 199 451 265
rect 485 199 547 471
rect 718 451 784 527
rect 581 199 639 348
rect 673 191 755 348
rect 789 199 903 348
rect 701 165 755 191
rect 213 17 402 89
rect 518 17 584 89
rect 701 58 799 165
rect 833 17 903 161
rect 0 -17 920 17
<< obsli1 >>
rect 299 299 357 493
rect 299 265 341 299
rect 213 215 341 265
rect 299 157 341 215
rect 614 417 680 493
rect 818 417 903 493
rect 614 383 903 417
rect 299 123 667 157
rect 436 51 484 123
rect 618 51 667 123
<< metal1 >>
rect 0 496 920 592
rect 0 -48 920 48
<< labels >>
rlabel locali s 701 165 755 191 6 A1
port 1 nsew signal input
rlabel locali s 701 58 799 165 6 A1
port 1 nsew signal input
rlabel locali s 673 191 755 348 6 A1
port 1 nsew signal input
rlabel locali s 789 199 903 348 6 A2
port 2 nsew signal input
rlabel locali s 581 199 639 348 6 B1
port 3 nsew signal input
rlabel locali s 485 199 547 471 6 C1
port 4 nsew signal input
rlabel locali s 392 265 451 471 6 D1
port 5 nsew signal input
rlabel locali s 377 199 451 265 6 D1
port 5 nsew signal input
rlabel locali s 121 51 179 478 6 X
port 6 nsew signal output
rlabel locali s 833 17 903 161 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 518 17 584 89 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 213 89 265 173 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 213 17 402 89 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 17 17 87 177 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 920 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 920 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 718 451 784 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 213 299 263 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 17 327 87 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 920 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 920 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 920 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3876812
string GDS_START 3867752
<< end >>
