magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 0 1071 29 1105
rect 63 1071 121 1105
rect 155 1071 213 1105
rect 247 1071 305 1105
rect 339 1071 397 1105
rect 431 1071 489 1105
rect 523 1071 581 1105
rect 615 1071 673 1105
rect 707 1071 765 1105
rect 799 1071 857 1105
rect 891 1071 949 1105
rect 983 1071 1041 1105
rect 1075 1071 1133 1105
rect 1167 1071 1225 1105
rect 1259 1071 1317 1105
rect 1351 1071 1409 1105
rect 1443 1071 1501 1105
rect 1535 1071 1593 1105
rect 1627 1071 1685 1105
rect 1719 1071 1777 1105
rect 1811 1071 1869 1105
rect 1903 1071 1961 1105
rect 1995 1071 2053 1105
rect 2087 1071 2145 1105
rect 2179 1071 2237 1105
rect 2271 1071 2329 1105
rect 2363 1071 2421 1105
rect 2455 1071 2513 1105
rect 2547 1071 2605 1105
rect 2639 1071 2697 1105
rect 2731 1071 2789 1105
rect 2823 1071 2881 1105
rect 2915 1071 2973 1105
rect 3007 1071 3065 1105
rect 3099 1071 3157 1105
rect 3191 1071 3249 1105
rect 3283 1071 3341 1105
rect 3375 1071 3433 1105
rect 3467 1071 3525 1105
rect 3559 1071 3617 1105
rect 3651 1071 3709 1105
rect 3743 1071 3801 1105
rect 3835 1071 3893 1105
rect 3927 1071 3985 1105
rect 4019 1071 4077 1105
rect 4111 1071 4169 1105
rect 4203 1071 4261 1105
rect 4295 1071 4353 1105
rect 4387 1071 4445 1105
rect 4479 1071 4537 1105
rect 4571 1071 4629 1105
rect 4663 1071 4721 1105
rect 4755 1071 4813 1105
rect 4847 1071 4905 1105
rect 4939 1071 4997 1105
rect 5031 1071 5089 1105
rect 5123 1071 5181 1105
rect 5215 1071 5273 1105
rect 5307 1071 5365 1105
rect 5399 1071 5457 1105
rect 5491 1071 5549 1105
rect 5583 1071 5641 1105
rect 5675 1071 5733 1105
rect 5767 1071 5825 1105
rect 5859 1071 5917 1105
rect 5951 1071 6009 1105
rect 6043 1071 6101 1105
rect 6135 1071 6193 1105
rect 6227 1071 6285 1105
rect 6319 1071 6377 1105
rect 6411 1071 6469 1105
rect 6503 1071 6561 1105
rect 6595 1071 6653 1105
rect 6687 1071 6745 1105
rect 6779 1071 6837 1105
rect 6871 1071 6929 1105
rect 6963 1071 7021 1105
rect 7055 1071 7113 1105
rect 7147 1071 7205 1105
rect 7239 1071 7297 1105
rect 7331 1071 7389 1105
rect 7423 1071 7481 1105
rect 7515 1071 7573 1105
rect 7607 1071 7665 1105
rect 7699 1071 7757 1105
rect 7791 1071 7849 1105
rect 7883 1071 7941 1105
rect 7975 1071 8033 1105
rect 8067 1071 8125 1105
rect 8159 1071 8217 1105
rect 8251 1071 8309 1105
rect 8343 1071 8401 1105
rect 8435 1071 8493 1105
rect 8527 1071 8585 1105
rect 8619 1071 8677 1105
rect 8711 1071 8769 1105
rect 8803 1071 8861 1105
rect 8895 1071 8953 1105
rect 8987 1071 9045 1105
rect 9079 1071 9137 1105
rect 9171 1071 9229 1105
rect 9263 1071 9321 1105
rect 9355 1071 9413 1105
rect 9447 1071 9505 1105
rect 9539 1071 9597 1105
rect 9631 1071 9689 1105
rect 9723 1071 9781 1105
rect 9815 1071 9873 1105
rect 9907 1071 9965 1105
rect 9999 1071 10057 1105
rect 10091 1071 10149 1105
rect 10183 1071 10241 1105
rect 10275 1071 10333 1105
rect 10367 1071 10396 1105
rect 29 911 79 1071
rect 213 979 267 1071
rect 401 979 451 1071
rect 573 911 639 969
rect 79 823 357 877
rect 593 875 639 911
rect 741 875 807 969
rect 992 966 1050 1071
rect 1176 966 1234 1071
rect 1342 966 1400 1071
rect 1526 966 1584 1071
rect 593 815 847 875
rect 25 561 79 789
rect 213 561 267 721
rect 401 561 455 721
rect 593 731 659 815
rect 593 697 609 731
rect 643 697 659 731
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 559 561
rect 25 299 79 527
rect 213 367 267 527
rect 401 367 455 527
rect 593 391 659 697
rect 781 731 847 815
rect 1152 823 1271 889
rect 1305 823 1424 889
rect 2125 979 2175 1071
rect 2309 979 2363 1071
rect 2497 911 2547 1071
rect 2605 911 2655 1071
rect 2789 979 2843 1071
rect 2977 979 3027 1071
rect 781 697 797 731
rect 831 697 847 731
rect 593 357 609 391
rect 643 357 659 391
rect 593 273 659 357
rect 781 391 847 697
rect 2219 823 2497 877
rect 2655 823 2933 877
rect 3568 966 3626 1071
rect 3752 966 3810 1071
rect 3918 966 3976 1071
rect 4102 966 4160 1071
rect 781 357 797 391
rect 831 357 847 391
rect 781 273 847 357
rect 79 211 357 265
rect 593 213 847 273
rect 593 177 639 213
rect 29 17 79 177
rect 213 17 267 109
rect 401 17 451 109
rect 573 119 639 177
rect 741 119 807 213
rect 1152 199 1271 265
rect 1305 199 1424 265
rect 2121 561 2175 721
rect 2309 561 2363 721
rect 2497 561 2551 789
rect 2601 561 2655 789
rect 2789 561 2843 721
rect 2977 561 3031 721
rect 2017 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3135 561
rect 2121 367 2175 527
rect 2309 367 2363 527
rect 2497 299 2551 527
rect 2601 299 2655 527
rect 2789 367 2843 527
rect 2977 367 3031 527
rect 3728 823 3847 889
rect 3881 823 4000 889
rect 4701 979 4751 1071
rect 4885 979 4939 1071
rect 5073 911 5123 1071
rect 5169 926 5227 1035
rect 5273 911 5323 1071
rect 5457 979 5511 1071
rect 5645 979 5695 1071
rect 4795 823 5073 877
rect 5323 823 5601 877
rect 6236 966 6294 1071
rect 6420 966 6478 1071
rect 6586 966 6644 1071
rect 6770 966 6828 1071
rect 992 17 1050 122
rect 1176 17 1234 122
rect 1342 17 1400 122
rect 1526 17 1584 122
rect 2219 211 2497 265
rect 2655 211 2933 265
rect 2125 17 2175 109
rect 2309 17 2363 109
rect 2497 17 2547 177
rect 2605 17 2655 177
rect 2789 17 2843 109
rect 2977 17 3027 109
rect 3728 199 3847 265
rect 3881 199 4000 265
rect 4697 561 4751 721
rect 4885 561 4939 721
rect 5073 561 5127 789
rect 5169 597 5227 794
rect 5269 561 5323 789
rect 5457 561 5511 721
rect 5645 561 5699 721
rect 4593 527 4629 561
rect 4663 527 4721 561
rect 4755 527 4813 561
rect 4847 527 4905 561
rect 4939 527 4997 561
rect 5031 527 5089 561
rect 5123 527 5181 561
rect 5215 527 5273 561
rect 5307 527 5365 561
rect 5399 527 5457 561
rect 5491 527 5549 561
rect 5583 527 5641 561
rect 5675 527 5733 561
rect 5767 527 5803 561
rect 4697 367 4751 527
rect 4885 367 4939 527
rect 5073 299 5127 527
rect 5169 294 5227 491
rect 5269 299 5323 527
rect 5457 367 5511 527
rect 5645 367 5699 527
rect 6396 823 6515 889
rect 6549 823 6668 889
rect 7369 979 7419 1071
rect 7553 979 7607 1071
rect 7741 911 7791 1071
rect 7849 911 7899 1071
rect 8033 979 8087 1071
rect 8221 979 8271 1071
rect 7463 823 7741 877
rect 7899 823 8177 877
rect 8812 966 8870 1071
rect 8996 966 9054 1071
rect 9162 966 9220 1071
rect 9346 966 9404 1071
rect 3568 17 3626 122
rect 3752 17 3810 122
rect 3918 17 3976 122
rect 4102 17 4160 122
rect 4795 211 5073 265
rect 5323 211 5601 265
rect 4701 17 4751 109
rect 4885 17 4939 109
rect 5073 17 5123 177
rect 5169 53 5227 162
rect 5273 17 5323 177
rect 5457 17 5511 109
rect 5645 17 5695 109
rect 6396 199 6515 265
rect 6549 199 6668 265
rect 7365 561 7419 721
rect 7553 561 7607 721
rect 7741 561 7795 789
rect 7845 561 7899 789
rect 8033 561 8087 721
rect 8221 561 8275 721
rect 7261 527 7297 561
rect 7331 527 7389 561
rect 7423 527 7481 561
rect 7515 527 7573 561
rect 7607 527 7665 561
rect 7699 527 7757 561
rect 7791 527 7849 561
rect 7883 527 7941 561
rect 7975 527 8033 561
rect 8067 527 8125 561
rect 8159 527 8217 561
rect 8251 527 8309 561
rect 8343 527 8379 561
rect 7365 367 7419 527
rect 7553 367 7607 527
rect 7741 299 7795 527
rect 7845 299 7899 527
rect 8033 367 8087 527
rect 8221 367 8275 527
rect 8972 823 9091 889
rect 9125 823 9244 889
rect 9945 979 9995 1071
rect 10129 979 10183 1071
rect 10317 911 10367 1071
rect 10039 823 10317 877
rect 6236 17 6294 122
rect 6420 17 6478 122
rect 6586 17 6644 122
rect 6770 17 6828 122
rect 7463 211 7741 265
rect 7899 211 8177 265
rect 7369 17 7419 109
rect 7553 17 7607 109
rect 7741 17 7791 177
rect 7849 17 7899 177
rect 8033 17 8087 109
rect 8221 17 8271 109
rect 8972 199 9091 265
rect 9125 199 9244 265
rect 9941 561 9995 721
rect 10129 561 10183 721
rect 10317 561 10371 789
rect 9837 527 9873 561
rect 9907 527 9965 561
rect 9999 527 10057 561
rect 10091 527 10149 561
rect 10183 527 10241 561
rect 10275 527 10333 561
rect 10367 527 10396 561
rect 9941 367 9995 527
rect 10129 367 10183 527
rect 10317 299 10371 527
rect 8812 17 8870 122
rect 8996 17 9054 122
rect 9162 17 9220 122
rect 9346 17 9404 122
rect 10039 211 10317 265
rect 9945 17 9995 109
rect 10129 17 10183 109
rect 10317 17 10367 177
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3341 17
rect 3375 -17 3433 17
rect 3467 -17 3525 17
rect 3559 -17 3617 17
rect 3651 -17 3709 17
rect 3743 -17 3801 17
rect 3835 -17 3893 17
rect 3927 -17 3985 17
rect 4019 -17 4077 17
rect 4111 -17 4169 17
rect 4203 -17 4261 17
rect 4295 -17 4353 17
rect 4387 -17 4445 17
rect 4479 -17 4537 17
rect 4571 -17 4629 17
rect 4663 -17 4721 17
rect 4755 -17 4813 17
rect 4847 -17 4905 17
rect 4939 -17 4997 17
rect 5031 -17 5089 17
rect 5123 -17 5181 17
rect 5215 -17 5273 17
rect 5307 -17 5365 17
rect 5399 -17 5457 17
rect 5491 -17 5549 17
rect 5583 -17 5641 17
rect 5675 -17 5733 17
rect 5767 -17 5825 17
rect 5859 -17 5917 17
rect 5951 -17 6009 17
rect 6043 -17 6101 17
rect 6135 -17 6193 17
rect 6227 -17 6285 17
rect 6319 -17 6377 17
rect 6411 -17 6469 17
rect 6503 -17 6561 17
rect 6595 -17 6653 17
rect 6687 -17 6745 17
rect 6779 -17 6837 17
rect 6871 -17 6929 17
rect 6963 -17 7021 17
rect 7055 -17 7113 17
rect 7147 -17 7205 17
rect 7239 -17 7297 17
rect 7331 -17 7389 17
rect 7423 -17 7481 17
rect 7515 -17 7573 17
rect 7607 -17 7665 17
rect 7699 -17 7757 17
rect 7791 -17 7849 17
rect 7883 -17 7941 17
rect 7975 -17 8033 17
rect 8067 -17 8125 17
rect 8159 -17 8217 17
rect 8251 -17 8309 17
rect 8343 -17 8401 17
rect 8435 -17 8493 17
rect 8527 -17 8585 17
rect 8619 -17 8677 17
rect 8711 -17 8769 17
rect 8803 -17 8861 17
rect 8895 -17 8953 17
rect 8987 -17 9045 17
rect 9079 -17 9137 17
rect 9171 -17 9229 17
rect 9263 -17 9321 17
rect 9355 -17 9413 17
rect 9447 -17 9505 17
rect 9539 -17 9597 17
rect 9631 -17 9689 17
rect 9723 -17 9781 17
rect 9815 -17 9873 17
rect 9907 -17 9965 17
rect 9999 -17 10057 17
rect 10091 -17 10149 17
rect 10183 -17 10241 17
rect 10275 -17 10333 17
rect 10367 -17 10396 17
<< viali >>
rect 29 1071 63 1105
rect 121 1071 155 1105
rect 213 1071 247 1105
rect 305 1071 339 1105
rect 397 1071 431 1105
rect 489 1071 523 1105
rect 581 1071 615 1105
rect 673 1071 707 1105
rect 765 1071 799 1105
rect 857 1071 891 1105
rect 949 1071 983 1105
rect 1041 1071 1075 1105
rect 1133 1071 1167 1105
rect 1225 1071 1259 1105
rect 1317 1071 1351 1105
rect 1409 1071 1443 1105
rect 1501 1071 1535 1105
rect 1593 1071 1627 1105
rect 1685 1071 1719 1105
rect 1777 1071 1811 1105
rect 1869 1071 1903 1105
rect 1961 1071 1995 1105
rect 2053 1071 2087 1105
rect 2145 1071 2179 1105
rect 2237 1071 2271 1105
rect 2329 1071 2363 1105
rect 2421 1071 2455 1105
rect 2513 1071 2547 1105
rect 2605 1071 2639 1105
rect 2697 1071 2731 1105
rect 2789 1071 2823 1105
rect 2881 1071 2915 1105
rect 2973 1071 3007 1105
rect 3065 1071 3099 1105
rect 3157 1071 3191 1105
rect 3249 1071 3283 1105
rect 3341 1071 3375 1105
rect 3433 1071 3467 1105
rect 3525 1071 3559 1105
rect 3617 1071 3651 1105
rect 3709 1071 3743 1105
rect 3801 1071 3835 1105
rect 3893 1071 3927 1105
rect 3985 1071 4019 1105
rect 4077 1071 4111 1105
rect 4169 1071 4203 1105
rect 4261 1071 4295 1105
rect 4353 1071 4387 1105
rect 4445 1071 4479 1105
rect 4537 1071 4571 1105
rect 4629 1071 4663 1105
rect 4721 1071 4755 1105
rect 4813 1071 4847 1105
rect 4905 1071 4939 1105
rect 4997 1071 5031 1105
rect 5089 1071 5123 1105
rect 5181 1071 5215 1105
rect 5273 1071 5307 1105
rect 5365 1071 5399 1105
rect 5457 1071 5491 1105
rect 5549 1071 5583 1105
rect 5641 1071 5675 1105
rect 5733 1071 5767 1105
rect 5825 1071 5859 1105
rect 5917 1071 5951 1105
rect 6009 1071 6043 1105
rect 6101 1071 6135 1105
rect 6193 1071 6227 1105
rect 6285 1071 6319 1105
rect 6377 1071 6411 1105
rect 6469 1071 6503 1105
rect 6561 1071 6595 1105
rect 6653 1071 6687 1105
rect 6745 1071 6779 1105
rect 6837 1071 6871 1105
rect 6929 1071 6963 1105
rect 7021 1071 7055 1105
rect 7113 1071 7147 1105
rect 7205 1071 7239 1105
rect 7297 1071 7331 1105
rect 7389 1071 7423 1105
rect 7481 1071 7515 1105
rect 7573 1071 7607 1105
rect 7665 1071 7699 1105
rect 7757 1071 7791 1105
rect 7849 1071 7883 1105
rect 7941 1071 7975 1105
rect 8033 1071 8067 1105
rect 8125 1071 8159 1105
rect 8217 1071 8251 1105
rect 8309 1071 8343 1105
rect 8401 1071 8435 1105
rect 8493 1071 8527 1105
rect 8585 1071 8619 1105
rect 8677 1071 8711 1105
rect 8769 1071 8803 1105
rect 8861 1071 8895 1105
rect 8953 1071 8987 1105
rect 9045 1071 9079 1105
rect 9137 1071 9171 1105
rect 9229 1071 9263 1105
rect 9321 1071 9355 1105
rect 9413 1071 9447 1105
rect 9505 1071 9539 1105
rect 9597 1071 9631 1105
rect 9689 1071 9723 1105
rect 9781 1071 9815 1105
rect 9873 1071 9907 1105
rect 9965 1071 9999 1105
rect 10057 1071 10091 1105
rect 10149 1071 10183 1105
rect 10241 1071 10275 1105
rect 10333 1071 10367 1105
rect 609 697 643 731
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 797 697 831 731
rect 609 357 643 391
rect 797 357 831 391
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 2881 527 2915 561
rect 2973 527 3007 561
rect 3065 527 3099 561
rect 4629 527 4663 561
rect 4721 527 4755 561
rect 4813 527 4847 561
rect 4905 527 4939 561
rect 4997 527 5031 561
rect 5089 527 5123 561
rect 5181 527 5215 561
rect 5273 527 5307 561
rect 5365 527 5399 561
rect 5457 527 5491 561
rect 5549 527 5583 561
rect 5641 527 5675 561
rect 5733 527 5767 561
rect 7297 527 7331 561
rect 7389 527 7423 561
rect 7481 527 7515 561
rect 7573 527 7607 561
rect 7665 527 7699 561
rect 7757 527 7791 561
rect 7849 527 7883 561
rect 7941 527 7975 561
rect 8033 527 8067 561
rect 8125 527 8159 561
rect 8217 527 8251 561
rect 8309 527 8343 561
rect 9873 527 9907 561
rect 9965 527 9999 561
rect 10057 527 10091 561
rect 10149 527 10183 561
rect 10241 527 10275 561
rect 10333 527 10367 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
rect 2881 -17 2915 17
rect 2973 -17 3007 17
rect 3065 -17 3099 17
rect 3157 -17 3191 17
rect 3249 -17 3283 17
rect 3341 -17 3375 17
rect 3433 -17 3467 17
rect 3525 -17 3559 17
rect 3617 -17 3651 17
rect 3709 -17 3743 17
rect 3801 -17 3835 17
rect 3893 -17 3927 17
rect 3985 -17 4019 17
rect 4077 -17 4111 17
rect 4169 -17 4203 17
rect 4261 -17 4295 17
rect 4353 -17 4387 17
rect 4445 -17 4479 17
rect 4537 -17 4571 17
rect 4629 -17 4663 17
rect 4721 -17 4755 17
rect 4813 -17 4847 17
rect 4905 -17 4939 17
rect 4997 -17 5031 17
rect 5089 -17 5123 17
rect 5181 -17 5215 17
rect 5273 -17 5307 17
rect 5365 -17 5399 17
rect 5457 -17 5491 17
rect 5549 -17 5583 17
rect 5641 -17 5675 17
rect 5733 -17 5767 17
rect 5825 -17 5859 17
rect 5917 -17 5951 17
rect 6009 -17 6043 17
rect 6101 -17 6135 17
rect 6193 -17 6227 17
rect 6285 -17 6319 17
rect 6377 -17 6411 17
rect 6469 -17 6503 17
rect 6561 -17 6595 17
rect 6653 -17 6687 17
rect 6745 -17 6779 17
rect 6837 -17 6871 17
rect 6929 -17 6963 17
rect 7021 -17 7055 17
rect 7113 -17 7147 17
rect 7205 -17 7239 17
rect 7297 -17 7331 17
rect 7389 -17 7423 17
rect 7481 -17 7515 17
rect 7573 -17 7607 17
rect 7665 -17 7699 17
rect 7757 -17 7791 17
rect 7849 -17 7883 17
rect 7941 -17 7975 17
rect 8033 -17 8067 17
rect 8125 -17 8159 17
rect 8217 -17 8251 17
rect 8309 -17 8343 17
rect 8401 -17 8435 17
rect 8493 -17 8527 17
rect 8585 -17 8619 17
rect 8677 -17 8711 17
rect 8769 -17 8803 17
rect 8861 -17 8895 17
rect 8953 -17 8987 17
rect 9045 -17 9079 17
rect 9137 -17 9171 17
rect 9229 -17 9263 17
rect 9321 -17 9355 17
rect 9413 -17 9447 17
rect 9505 -17 9539 17
rect 9597 -17 9631 17
rect 9689 -17 9723 17
rect 9781 -17 9815 17
rect 9873 -17 9907 17
rect 9965 -17 9999 17
rect 10057 -17 10091 17
rect 10149 -17 10183 17
rect 10241 -17 10275 17
rect 10333 -17 10367 17
<< obsli1 >>
rect 113 945 179 1037
rect 301 945 367 1037
rect 485 1003 891 1037
rect 485 945 539 1003
rect 113 911 539 945
rect 673 934 707 1003
rect 841 934 891 1003
rect 1084 923 1134 1032
rect 1442 923 1492 1032
rect 1685 1003 2091 1037
rect 1685 934 1735 1003
rect 1084 875 1118 923
rect 113 755 559 789
rect 113 595 179 755
rect 301 595 367 755
rect 499 595 559 755
rect 113 333 179 493
rect 301 333 367 493
rect 499 333 559 493
rect 113 299 559 333
rect 693 595 747 781
rect 881 809 1118 875
rect 1458 875 1492 923
rect 1769 875 1835 969
rect 1869 934 1903 1003
rect 1937 911 2003 969
rect 2037 945 2091 1003
rect 2209 945 2275 1037
rect 2397 945 2463 1037
rect 2037 911 2463 945
rect 2689 945 2755 1037
rect 2877 945 2943 1037
rect 3061 1003 3467 1037
rect 3061 945 3115 1003
rect 2689 911 3115 945
rect 3149 911 3215 969
rect 3249 934 3283 1003
rect 1937 875 1983 911
rect 693 307 747 493
rect 881 595 941 775
rect 1084 767 1118 809
rect 1458 809 1695 875
rect 1729 815 1983 875
rect 3169 875 3215 911
rect 3317 875 3383 969
rect 3417 934 3467 1003
rect 3660 923 3710 1032
rect 4018 923 4068 1032
rect 4261 1003 4667 1037
rect 4261 934 4311 1003
rect 3660 875 3694 923
rect 1458 767 1492 809
rect 990 561 1045 767
rect 1084 595 1150 767
rect 1184 561 1244 767
rect 1332 561 1392 767
rect 1426 595 1492 767
rect 1531 561 1586 767
rect 1635 595 1695 775
rect 1729 731 1795 815
rect 1729 697 1745 731
rect 1779 697 1795 731
rect 881 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1695 561
rect 881 313 941 493
rect 990 321 1045 527
rect 1084 321 1150 493
rect 1184 321 1244 527
rect 1332 321 1392 527
rect 1426 321 1492 493
rect 1531 321 1586 527
rect 1084 279 1118 321
rect 881 213 1118 279
rect 1458 279 1492 321
rect 1635 313 1695 493
rect 1729 391 1795 697
rect 1829 595 1883 781
rect 1917 731 1983 815
rect 3169 815 3423 875
rect 1917 697 1933 731
rect 1967 697 1983 731
rect 1729 357 1745 391
rect 1779 357 1795 391
rect 113 143 539 177
rect 113 51 179 143
rect 301 51 367 143
rect 485 85 539 143
rect 673 85 707 154
rect 1084 165 1118 213
rect 1458 213 1695 279
rect 1729 273 1795 357
rect 1829 307 1883 493
rect 1917 391 1983 697
rect 2017 755 2463 789
rect 2017 595 2077 755
rect 2209 595 2275 755
rect 2397 595 2463 755
rect 2689 755 3135 789
rect 2689 595 2755 755
rect 2877 595 2943 755
rect 3075 595 3135 755
rect 3169 731 3235 815
rect 3169 697 3185 731
rect 3219 697 3235 731
rect 1917 357 1933 391
rect 1967 357 1983 391
rect 1917 273 1983 357
rect 2017 333 2077 493
rect 2209 333 2275 493
rect 2397 333 2463 493
rect 2017 299 2463 333
rect 2689 333 2755 493
rect 2877 333 2943 493
rect 3075 333 3135 493
rect 2689 299 3135 333
rect 3169 391 3235 697
rect 3269 595 3323 781
rect 3357 731 3423 815
rect 3457 809 3694 875
rect 4034 875 4068 923
rect 4345 875 4411 969
rect 4445 934 4479 1003
rect 4513 911 4579 969
rect 4613 945 4667 1003
rect 4785 945 4851 1037
rect 4973 945 5039 1037
rect 4613 911 5039 945
rect 5357 945 5423 1037
rect 5545 945 5611 1037
rect 5729 1003 6135 1037
rect 5729 945 5783 1003
rect 5357 911 5783 945
rect 5817 911 5883 969
rect 5917 934 5951 1003
rect 4513 875 4559 911
rect 3357 697 3373 731
rect 3407 697 3423 731
rect 3169 357 3185 391
rect 3219 357 3235 391
rect 1729 213 1983 273
rect 3169 273 3235 357
rect 3269 307 3323 493
rect 3357 391 3423 697
rect 3457 595 3517 775
rect 3660 767 3694 809
rect 4034 809 4271 875
rect 4305 815 4559 875
rect 5837 875 5883 911
rect 5985 875 6051 969
rect 6085 934 6135 1003
rect 6328 923 6378 1032
rect 6686 923 6736 1032
rect 6929 1003 7335 1037
rect 6929 934 6979 1003
rect 6328 875 6362 923
rect 4034 767 4068 809
rect 3566 561 3621 767
rect 3660 595 3726 767
rect 3760 561 3820 767
rect 3908 561 3968 767
rect 4002 595 4068 767
rect 4107 561 4162 767
rect 4211 595 4271 775
rect 4305 731 4371 815
rect 4305 697 4321 731
rect 4355 697 4371 731
rect 3457 527 3525 561
rect 3559 527 3617 561
rect 3651 527 3709 561
rect 3743 527 3801 561
rect 3835 527 3893 561
rect 3927 527 3985 561
rect 4019 527 4077 561
rect 4111 527 4169 561
rect 4203 527 4271 561
rect 3357 357 3373 391
rect 3407 357 3423 391
rect 3357 273 3423 357
rect 3457 313 3517 493
rect 3566 321 3621 527
rect 3660 321 3726 493
rect 3760 321 3820 527
rect 3908 321 3968 527
rect 4002 321 4068 493
rect 4107 321 4162 527
rect 3660 279 3694 321
rect 1458 165 1492 213
rect 841 85 891 154
rect 485 51 891 85
rect 1084 56 1134 165
rect 1442 56 1492 165
rect 1685 85 1735 154
rect 1769 119 1835 213
rect 1937 177 1983 213
rect 3169 213 3423 273
rect 3457 213 3694 279
rect 4034 279 4068 321
rect 4211 313 4271 493
rect 4305 391 4371 697
rect 4405 595 4459 781
rect 4493 731 4559 815
rect 5837 815 6091 875
rect 4493 697 4509 731
rect 4543 697 4559 731
rect 4305 357 4321 391
rect 4355 357 4371 391
rect 3169 177 3215 213
rect 1869 85 1903 154
rect 1937 119 2003 177
rect 2037 143 2463 177
rect 2037 85 2091 143
rect 1685 51 2091 85
rect 2209 51 2275 143
rect 2397 51 2463 143
rect 2689 143 3115 177
rect 2689 51 2755 143
rect 2877 51 2943 143
rect 3061 85 3115 143
rect 3149 119 3215 177
rect 3249 85 3283 154
rect 3317 119 3383 213
rect 3660 165 3694 213
rect 4034 213 4271 279
rect 4305 273 4371 357
rect 4405 307 4459 493
rect 4493 391 4559 697
rect 4593 755 5039 789
rect 4593 595 4653 755
rect 4785 595 4851 755
rect 4973 595 5039 755
rect 5357 755 5803 789
rect 5357 595 5423 755
rect 5545 595 5611 755
rect 5743 595 5803 755
rect 5837 731 5903 815
rect 5837 697 5853 731
rect 5887 697 5903 731
rect 4493 357 4509 391
rect 4543 357 4559 391
rect 4493 273 4559 357
rect 4593 333 4653 493
rect 4785 333 4851 493
rect 4973 333 5039 493
rect 4593 299 5039 333
rect 5357 333 5423 493
rect 5545 333 5611 493
rect 5743 333 5803 493
rect 5357 299 5803 333
rect 5837 391 5903 697
rect 5937 595 5991 781
rect 6025 731 6091 815
rect 6125 809 6362 875
rect 6702 875 6736 923
rect 7013 875 7079 969
rect 7113 934 7147 1003
rect 7181 911 7247 969
rect 7281 945 7335 1003
rect 7453 945 7519 1037
rect 7641 945 7707 1037
rect 7281 911 7707 945
rect 7933 945 7999 1037
rect 8121 945 8187 1037
rect 8305 1003 8711 1037
rect 8305 945 8359 1003
rect 7933 911 8359 945
rect 8393 911 8459 969
rect 8493 934 8527 1003
rect 7181 875 7227 911
rect 6025 697 6041 731
rect 6075 697 6091 731
rect 5837 357 5853 391
rect 5887 357 5903 391
rect 4305 213 4559 273
rect 5837 273 5903 357
rect 5937 307 5991 493
rect 6025 391 6091 697
rect 6125 595 6185 775
rect 6328 767 6362 809
rect 6702 809 6939 875
rect 6973 815 7227 875
rect 8413 875 8459 911
rect 8561 875 8627 969
rect 8661 934 8711 1003
rect 8904 923 8954 1032
rect 9262 923 9312 1032
rect 9505 1003 9911 1037
rect 9505 934 9555 1003
rect 8904 875 8938 923
rect 6702 767 6736 809
rect 6234 561 6289 767
rect 6328 595 6394 767
rect 6428 561 6488 767
rect 6576 561 6636 767
rect 6670 595 6736 767
rect 6775 561 6830 767
rect 6879 595 6939 775
rect 6973 731 7039 815
rect 6973 697 6989 731
rect 7023 697 7039 731
rect 6125 527 6193 561
rect 6227 527 6285 561
rect 6319 527 6377 561
rect 6411 527 6469 561
rect 6503 527 6561 561
rect 6595 527 6653 561
rect 6687 527 6745 561
rect 6779 527 6837 561
rect 6871 527 6939 561
rect 6025 357 6041 391
rect 6075 357 6091 391
rect 6025 273 6091 357
rect 6125 313 6185 493
rect 6234 321 6289 527
rect 6328 321 6394 493
rect 6428 321 6488 527
rect 6576 321 6636 527
rect 6670 321 6736 493
rect 6775 321 6830 527
rect 6328 279 6362 321
rect 4034 165 4068 213
rect 3417 85 3467 154
rect 3061 51 3467 85
rect 3660 56 3710 165
rect 4018 56 4068 165
rect 4261 85 4311 154
rect 4345 119 4411 213
rect 4513 177 4559 213
rect 5837 213 6091 273
rect 6125 213 6362 279
rect 6702 279 6736 321
rect 6879 313 6939 493
rect 6973 391 7039 697
rect 7073 595 7127 781
rect 7161 731 7227 815
rect 8413 815 8667 875
rect 7161 697 7177 731
rect 7211 697 7227 731
rect 6973 357 6989 391
rect 7023 357 7039 391
rect 5837 177 5883 213
rect 4445 85 4479 154
rect 4513 119 4579 177
rect 4613 143 5039 177
rect 4613 85 4667 143
rect 4261 51 4667 85
rect 4785 51 4851 143
rect 4973 51 5039 143
rect 5357 143 5783 177
rect 5357 51 5423 143
rect 5545 51 5611 143
rect 5729 85 5783 143
rect 5817 119 5883 177
rect 5917 85 5951 154
rect 5985 119 6051 213
rect 6328 165 6362 213
rect 6702 213 6939 279
rect 6973 273 7039 357
rect 7073 307 7127 493
rect 7161 391 7227 697
rect 7261 755 7707 789
rect 7261 595 7321 755
rect 7453 595 7519 755
rect 7641 595 7707 755
rect 7933 755 8379 789
rect 7933 595 7999 755
rect 8121 595 8187 755
rect 8319 595 8379 755
rect 8413 731 8479 815
rect 8413 697 8429 731
rect 8463 697 8479 731
rect 7161 357 7177 391
rect 7211 357 7227 391
rect 7161 273 7227 357
rect 7261 333 7321 493
rect 7453 333 7519 493
rect 7641 333 7707 493
rect 7261 299 7707 333
rect 7933 333 7999 493
rect 8121 333 8187 493
rect 8319 333 8379 493
rect 7933 299 8379 333
rect 8413 391 8479 697
rect 8513 595 8567 781
rect 8601 731 8667 815
rect 8701 809 8938 875
rect 9278 875 9312 923
rect 9589 875 9655 969
rect 9689 934 9723 1003
rect 9757 911 9823 969
rect 9857 945 9911 1003
rect 10029 945 10095 1037
rect 10217 945 10283 1037
rect 9857 911 10283 945
rect 9757 875 9803 911
rect 8601 697 8617 731
rect 8651 697 8667 731
rect 8413 357 8429 391
rect 8463 357 8479 391
rect 6973 213 7227 273
rect 8413 273 8479 357
rect 8513 307 8567 493
rect 8601 391 8667 697
rect 8701 595 8761 775
rect 8904 767 8938 809
rect 9278 809 9515 875
rect 9549 815 9803 875
rect 9278 767 9312 809
rect 8810 561 8865 767
rect 8904 595 8970 767
rect 9004 561 9064 767
rect 9152 561 9212 767
rect 9246 595 9312 767
rect 9351 561 9406 767
rect 9455 595 9515 775
rect 9549 731 9615 815
rect 9549 697 9565 731
rect 9599 697 9615 731
rect 8701 527 8769 561
rect 8803 527 8861 561
rect 8895 527 8953 561
rect 8987 527 9045 561
rect 9079 527 9137 561
rect 9171 527 9229 561
rect 9263 527 9321 561
rect 9355 527 9413 561
rect 9447 527 9515 561
rect 8601 357 8617 391
rect 8651 357 8667 391
rect 8601 273 8667 357
rect 8701 313 8761 493
rect 8810 321 8865 527
rect 8904 321 8970 493
rect 9004 321 9064 527
rect 9152 321 9212 527
rect 9246 321 9312 493
rect 9351 321 9406 527
rect 8904 279 8938 321
rect 6702 165 6736 213
rect 6085 85 6135 154
rect 5729 51 6135 85
rect 6328 56 6378 165
rect 6686 56 6736 165
rect 6929 85 6979 154
rect 7013 119 7079 213
rect 7181 177 7227 213
rect 8413 213 8667 273
rect 8701 213 8938 279
rect 9278 279 9312 321
rect 9455 313 9515 493
rect 9549 391 9615 697
rect 9649 595 9703 781
rect 9737 731 9803 815
rect 9737 697 9753 731
rect 9787 697 9803 731
rect 9549 357 9565 391
rect 9599 357 9615 391
rect 8413 177 8459 213
rect 7113 85 7147 154
rect 7181 119 7247 177
rect 7281 143 7707 177
rect 7281 85 7335 143
rect 6929 51 7335 85
rect 7453 51 7519 143
rect 7641 51 7707 143
rect 7933 143 8359 177
rect 7933 51 7999 143
rect 8121 51 8187 143
rect 8305 85 8359 143
rect 8393 119 8459 177
rect 8493 85 8527 154
rect 8561 119 8627 213
rect 8904 165 8938 213
rect 9278 213 9515 279
rect 9549 273 9615 357
rect 9649 307 9703 493
rect 9737 391 9803 697
rect 9837 755 10283 789
rect 9837 595 9897 755
rect 10029 595 10095 755
rect 10217 595 10283 755
rect 9737 357 9753 391
rect 9787 357 9803 391
rect 9737 273 9803 357
rect 9837 333 9897 493
rect 10029 333 10095 493
rect 10217 333 10283 493
rect 9837 299 10283 333
rect 9549 213 9803 273
rect 9278 165 9312 213
rect 8661 85 8711 154
rect 8305 51 8711 85
rect 8904 56 8954 165
rect 9262 56 9312 165
rect 9505 85 9555 154
rect 9589 119 9655 213
rect 9757 177 9803 213
rect 9689 85 9723 154
rect 9757 119 9823 177
rect 9857 143 10283 177
rect 9857 85 9911 143
rect 9505 51 9911 85
rect 10029 51 10095 143
rect 10217 51 10283 143
<< obsli1c >>
rect 1745 697 1779 731
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1933 697 1967 731
rect 1745 357 1779 391
rect 3185 697 3219 731
rect 1933 357 1967 391
rect 3373 697 3407 731
rect 3185 357 3219 391
rect 4321 697 4355 731
rect 3525 527 3559 561
rect 3617 527 3651 561
rect 3709 527 3743 561
rect 3801 527 3835 561
rect 3893 527 3927 561
rect 3985 527 4019 561
rect 4077 527 4111 561
rect 4169 527 4203 561
rect 3373 357 3407 391
rect 4509 697 4543 731
rect 4321 357 4355 391
rect 5853 697 5887 731
rect 4509 357 4543 391
rect 6041 697 6075 731
rect 5853 357 5887 391
rect 6989 697 7023 731
rect 6193 527 6227 561
rect 6285 527 6319 561
rect 6377 527 6411 561
rect 6469 527 6503 561
rect 6561 527 6595 561
rect 6653 527 6687 561
rect 6745 527 6779 561
rect 6837 527 6871 561
rect 6041 357 6075 391
rect 7177 697 7211 731
rect 6989 357 7023 391
rect 8429 697 8463 731
rect 7177 357 7211 391
rect 8617 697 8651 731
rect 8429 357 8463 391
rect 9565 697 9599 731
rect 8769 527 8803 561
rect 8861 527 8895 561
rect 8953 527 8987 561
rect 9045 527 9079 561
rect 9137 527 9171 561
rect 9229 527 9263 561
rect 9321 527 9355 561
rect 9413 527 9447 561
rect 8617 357 8651 391
rect 9753 697 9787 731
rect 9565 357 9599 391
rect 9753 357 9787 391
<< metal1 >>
rect 0 1105 10396 1136
rect 0 1071 29 1105
rect 63 1071 121 1105
rect 155 1071 213 1105
rect 247 1071 305 1105
rect 339 1071 397 1105
rect 431 1071 489 1105
rect 523 1071 581 1105
rect 615 1071 673 1105
rect 707 1071 765 1105
rect 799 1071 857 1105
rect 891 1071 949 1105
rect 983 1071 1041 1105
rect 1075 1071 1133 1105
rect 1167 1071 1225 1105
rect 1259 1071 1317 1105
rect 1351 1071 1409 1105
rect 1443 1071 1501 1105
rect 1535 1071 1593 1105
rect 1627 1071 1685 1105
rect 1719 1071 1777 1105
rect 1811 1071 1869 1105
rect 1903 1071 1961 1105
rect 1995 1071 2053 1105
rect 2087 1071 2145 1105
rect 2179 1071 2237 1105
rect 2271 1071 2329 1105
rect 2363 1071 2421 1105
rect 2455 1071 2513 1105
rect 2547 1071 2605 1105
rect 2639 1071 2697 1105
rect 2731 1071 2789 1105
rect 2823 1071 2881 1105
rect 2915 1071 2973 1105
rect 3007 1071 3065 1105
rect 3099 1071 3157 1105
rect 3191 1071 3249 1105
rect 3283 1071 3341 1105
rect 3375 1071 3433 1105
rect 3467 1071 3525 1105
rect 3559 1071 3617 1105
rect 3651 1071 3709 1105
rect 3743 1071 3801 1105
rect 3835 1071 3893 1105
rect 3927 1071 3985 1105
rect 4019 1071 4077 1105
rect 4111 1071 4169 1105
rect 4203 1071 4261 1105
rect 4295 1071 4353 1105
rect 4387 1071 4445 1105
rect 4479 1071 4537 1105
rect 4571 1071 4629 1105
rect 4663 1071 4721 1105
rect 4755 1071 4813 1105
rect 4847 1071 4905 1105
rect 4939 1071 4997 1105
rect 5031 1071 5089 1105
rect 5123 1071 5181 1105
rect 5215 1071 5273 1105
rect 5307 1071 5365 1105
rect 5399 1071 5457 1105
rect 5491 1071 5549 1105
rect 5583 1071 5641 1105
rect 5675 1071 5733 1105
rect 5767 1071 5825 1105
rect 5859 1071 5917 1105
rect 5951 1071 6009 1105
rect 6043 1071 6101 1105
rect 6135 1071 6193 1105
rect 6227 1071 6285 1105
rect 6319 1071 6377 1105
rect 6411 1071 6469 1105
rect 6503 1071 6561 1105
rect 6595 1071 6653 1105
rect 6687 1071 6745 1105
rect 6779 1071 6837 1105
rect 6871 1071 6929 1105
rect 6963 1071 7021 1105
rect 7055 1071 7113 1105
rect 7147 1071 7205 1105
rect 7239 1071 7297 1105
rect 7331 1071 7389 1105
rect 7423 1071 7481 1105
rect 7515 1071 7573 1105
rect 7607 1071 7665 1105
rect 7699 1071 7757 1105
rect 7791 1071 7849 1105
rect 7883 1071 7941 1105
rect 7975 1071 8033 1105
rect 8067 1071 8125 1105
rect 8159 1071 8217 1105
rect 8251 1071 8309 1105
rect 8343 1071 8401 1105
rect 8435 1071 8493 1105
rect 8527 1071 8585 1105
rect 8619 1071 8677 1105
rect 8711 1071 8769 1105
rect 8803 1071 8861 1105
rect 8895 1071 8953 1105
rect 8987 1071 9045 1105
rect 9079 1071 9137 1105
rect 9171 1071 9229 1105
rect 9263 1071 9321 1105
rect 9355 1071 9413 1105
rect 9447 1071 9505 1105
rect 9539 1071 9597 1105
rect 9631 1071 9689 1105
rect 9723 1071 9781 1105
rect 9815 1071 9873 1105
rect 9907 1071 9965 1105
rect 9999 1071 10057 1105
rect 10091 1071 10149 1105
rect 10183 1071 10241 1105
rect 10275 1071 10333 1105
rect 10367 1071 10396 1105
rect 0 1040 10396 1071
rect 597 731 655 737
rect 597 697 609 731
rect 643 728 655 731
rect 785 731 843 737
rect 785 728 797 731
rect 643 700 797 728
rect 643 697 655 700
rect 597 691 655 697
rect 785 697 797 700
rect 831 728 843 731
rect 1733 731 1791 737
rect 1733 728 1745 731
rect 831 700 1745 728
rect 831 697 843 700
rect 785 691 843 697
rect 1733 697 1745 700
rect 1779 728 1791 731
rect 1921 731 1979 737
rect 1921 728 1933 731
rect 1779 700 1933 728
rect 1779 697 1791 700
rect 1733 691 1791 697
rect 1921 697 1933 700
rect 1967 728 1979 731
rect 3173 731 3231 737
rect 3173 728 3185 731
rect 1967 700 3185 728
rect 1967 697 1979 700
rect 1921 691 1979 697
rect 3173 697 3185 700
rect 3219 728 3231 731
rect 3361 731 3419 737
rect 3361 728 3373 731
rect 3219 700 3373 728
rect 3219 697 3231 700
rect 3173 691 3231 697
rect 3361 697 3373 700
rect 3407 728 3419 731
rect 4309 731 4367 737
rect 4309 728 4321 731
rect 3407 700 4321 728
rect 3407 697 3419 700
rect 3361 691 3419 697
rect 4309 697 4321 700
rect 4355 728 4367 731
rect 4497 731 4555 737
rect 4497 728 4509 731
rect 4355 700 4509 728
rect 4355 697 4367 700
rect 4309 691 4367 697
rect 4497 697 4509 700
rect 4543 728 4555 731
rect 5841 731 5899 737
rect 5841 728 5853 731
rect 4543 700 5853 728
rect 4543 697 4555 700
rect 4497 691 4555 697
rect 5841 697 5853 700
rect 5887 728 5899 731
rect 6029 731 6087 737
rect 6029 728 6041 731
rect 5887 700 6041 728
rect 5887 697 5899 700
rect 5841 691 5899 697
rect 6029 697 6041 700
rect 6075 728 6087 731
rect 6977 731 7035 737
rect 6977 728 6989 731
rect 6075 700 6989 728
rect 6075 697 6087 700
rect 6029 691 6087 697
rect 6977 697 6989 700
rect 7023 728 7035 731
rect 7165 731 7223 737
rect 7165 728 7177 731
rect 7023 700 7177 728
rect 7023 697 7035 700
rect 6977 691 7035 697
rect 7165 697 7177 700
rect 7211 728 7223 731
rect 8417 731 8475 737
rect 8417 728 8429 731
rect 7211 700 8429 728
rect 7211 697 7223 700
rect 7165 691 7223 697
rect 8417 697 8429 700
rect 8463 728 8475 731
rect 8605 731 8663 737
rect 8605 728 8617 731
rect 8463 700 8617 728
rect 8463 697 8475 700
rect 8417 691 8475 697
rect 8605 697 8617 700
rect 8651 728 8663 731
rect 9553 731 9611 737
rect 9553 728 9565 731
rect 8651 700 9565 728
rect 8651 697 8663 700
rect 8605 691 8663 697
rect 9553 697 9565 700
rect 9599 728 9611 731
rect 9741 731 9799 737
rect 9741 728 9753 731
rect 9599 700 9753 728
rect 9599 697 9611 700
rect 9553 691 9611 697
rect 9741 697 9753 700
rect 9787 697 9799 731
rect 9741 691 9799 697
rect 0 561 10396 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3525 561
rect 3559 527 3617 561
rect 3651 527 3709 561
rect 3743 527 3801 561
rect 3835 527 3893 561
rect 3927 527 3985 561
rect 4019 527 4077 561
rect 4111 527 4169 561
rect 4203 527 4629 561
rect 4663 527 4721 561
rect 4755 527 4813 561
rect 4847 527 4905 561
rect 4939 527 4997 561
rect 5031 527 5089 561
rect 5123 527 5181 561
rect 5215 527 5273 561
rect 5307 527 5365 561
rect 5399 527 5457 561
rect 5491 527 5549 561
rect 5583 527 5641 561
rect 5675 527 5733 561
rect 5767 527 6193 561
rect 6227 527 6285 561
rect 6319 527 6377 561
rect 6411 527 6469 561
rect 6503 527 6561 561
rect 6595 527 6653 561
rect 6687 527 6745 561
rect 6779 527 6837 561
rect 6871 527 7297 561
rect 7331 527 7389 561
rect 7423 527 7481 561
rect 7515 527 7573 561
rect 7607 527 7665 561
rect 7699 527 7757 561
rect 7791 527 7849 561
rect 7883 527 7941 561
rect 7975 527 8033 561
rect 8067 527 8125 561
rect 8159 527 8217 561
rect 8251 527 8309 561
rect 8343 527 8769 561
rect 8803 527 8861 561
rect 8895 527 8953 561
rect 8987 527 9045 561
rect 9079 527 9137 561
rect 9171 527 9229 561
rect 9263 527 9321 561
rect 9355 527 9413 561
rect 9447 527 9873 561
rect 9907 527 9965 561
rect 9999 527 10057 561
rect 10091 527 10149 561
rect 10183 527 10241 561
rect 10275 527 10333 561
rect 10367 527 10396 561
rect 0 496 10396 527
rect 597 391 655 397
rect 597 357 609 391
rect 643 388 655 391
rect 785 391 843 397
rect 785 388 797 391
rect 643 360 797 388
rect 643 357 655 360
rect 597 351 655 357
rect 785 357 797 360
rect 831 388 843 391
rect 1733 391 1791 397
rect 1733 388 1745 391
rect 831 360 1745 388
rect 831 357 843 360
rect 785 351 843 357
rect 1733 357 1745 360
rect 1779 388 1791 391
rect 1921 391 1979 397
rect 1921 388 1933 391
rect 1779 360 1933 388
rect 1779 357 1791 360
rect 1733 351 1791 357
rect 1921 357 1933 360
rect 1967 388 1979 391
rect 3173 391 3231 397
rect 3173 388 3185 391
rect 1967 360 3185 388
rect 1967 357 1979 360
rect 1921 351 1979 357
rect 3173 357 3185 360
rect 3219 388 3231 391
rect 3361 391 3419 397
rect 3361 388 3373 391
rect 3219 360 3373 388
rect 3219 357 3231 360
rect 3173 351 3231 357
rect 3361 357 3373 360
rect 3407 388 3419 391
rect 4309 391 4367 397
rect 4309 388 4321 391
rect 3407 360 4321 388
rect 3407 357 3419 360
rect 3361 351 3419 357
rect 4309 357 4321 360
rect 4355 388 4367 391
rect 4497 391 4555 397
rect 4497 388 4509 391
rect 4355 360 4509 388
rect 4355 357 4367 360
rect 4309 351 4367 357
rect 4497 357 4509 360
rect 4543 388 4555 391
rect 5841 391 5899 397
rect 5841 388 5853 391
rect 4543 360 5853 388
rect 4543 357 4555 360
rect 4497 351 4555 357
rect 5841 357 5853 360
rect 5887 388 5899 391
rect 6029 391 6087 397
rect 6029 388 6041 391
rect 5887 360 6041 388
rect 5887 357 5899 360
rect 5841 351 5899 357
rect 6029 357 6041 360
rect 6075 388 6087 391
rect 6977 391 7035 397
rect 6977 388 6989 391
rect 6075 360 6989 388
rect 6075 357 6087 360
rect 6029 351 6087 357
rect 6977 357 6989 360
rect 7023 388 7035 391
rect 7165 391 7223 397
rect 7165 388 7177 391
rect 7023 360 7177 388
rect 7023 357 7035 360
rect 6977 351 7035 357
rect 7165 357 7177 360
rect 7211 388 7223 391
rect 8417 391 8475 397
rect 8417 388 8429 391
rect 7211 360 8429 388
rect 7211 357 7223 360
rect 7165 351 7223 357
rect 8417 357 8429 360
rect 8463 388 8475 391
rect 8605 391 8663 397
rect 8605 388 8617 391
rect 8463 360 8617 388
rect 8463 357 8475 360
rect 8417 351 8475 357
rect 8605 357 8617 360
rect 8651 388 8663 391
rect 9553 391 9611 397
rect 9553 388 9565 391
rect 8651 360 9565 388
rect 8651 357 8663 360
rect 8605 351 8663 357
rect 9553 357 9565 360
rect 9599 388 9611 391
rect 9741 391 9799 397
rect 9741 388 9753 391
rect 9599 360 9753 388
rect 9599 357 9611 360
rect 9553 351 9611 357
rect 9741 357 9753 360
rect 9787 357 9799 391
rect 9741 351 9799 357
rect 0 17 10396 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3341 17
rect 3375 -17 3433 17
rect 3467 -17 3525 17
rect 3559 -17 3617 17
rect 3651 -17 3709 17
rect 3743 -17 3801 17
rect 3835 -17 3893 17
rect 3927 -17 3985 17
rect 4019 -17 4077 17
rect 4111 -17 4169 17
rect 4203 -17 4261 17
rect 4295 -17 4353 17
rect 4387 -17 4445 17
rect 4479 -17 4537 17
rect 4571 -17 4629 17
rect 4663 -17 4721 17
rect 4755 -17 4813 17
rect 4847 -17 4905 17
rect 4939 -17 4997 17
rect 5031 -17 5089 17
rect 5123 -17 5181 17
rect 5215 -17 5273 17
rect 5307 -17 5365 17
rect 5399 -17 5457 17
rect 5491 -17 5549 17
rect 5583 -17 5641 17
rect 5675 -17 5733 17
rect 5767 -17 5825 17
rect 5859 -17 5917 17
rect 5951 -17 6009 17
rect 6043 -17 6101 17
rect 6135 -17 6193 17
rect 6227 -17 6285 17
rect 6319 -17 6377 17
rect 6411 -17 6469 17
rect 6503 -17 6561 17
rect 6595 -17 6653 17
rect 6687 -17 6745 17
rect 6779 -17 6837 17
rect 6871 -17 6929 17
rect 6963 -17 7021 17
rect 7055 -17 7113 17
rect 7147 -17 7205 17
rect 7239 -17 7297 17
rect 7331 -17 7389 17
rect 7423 -17 7481 17
rect 7515 -17 7573 17
rect 7607 -17 7665 17
rect 7699 -17 7757 17
rect 7791 -17 7849 17
rect 7883 -17 7941 17
rect 7975 -17 8033 17
rect 8067 -17 8125 17
rect 8159 -17 8217 17
rect 8251 -17 8309 17
rect 8343 -17 8401 17
rect 8435 -17 8493 17
rect 8527 -17 8585 17
rect 8619 -17 8677 17
rect 8711 -17 8769 17
rect 8803 -17 8861 17
rect 8895 -17 8953 17
rect 8987 -17 9045 17
rect 9079 -17 9137 17
rect 9171 -17 9229 17
rect 9263 -17 9321 17
rect 9355 -17 9413 17
rect 9447 -17 9505 17
rect 9539 -17 9597 17
rect 9631 -17 9689 17
rect 9723 -17 9781 17
rect 9815 -17 9873 17
rect 9907 -17 9965 17
rect 9999 -17 10057 17
rect 10091 -17 10149 17
rect 10183 -17 10241 17
rect 10275 -17 10333 17
rect 10367 -17 10396 17
rect 0 -48 10396 -17
<< obsm1 >>
rect 117 657 175 666
rect 305 657 363 666
rect 501 657 559 666
rect 691 657 749 666
rect 881 657 939 666
rect 117 629 939 657
rect 117 620 175 629
rect 305 620 363 629
rect 501 620 559 629
rect 691 620 749 629
rect 881 620 939 629
rect 1637 657 1695 666
rect 1827 657 1885 666
rect 2017 657 2075 666
rect 2213 657 2271 666
rect 2401 657 2459 666
rect 1637 629 2459 657
rect 1637 620 1695 629
rect 1827 620 1885 629
rect 2017 620 2075 629
rect 2213 620 2271 629
rect 2401 620 2459 629
rect 2693 657 2751 666
rect 2881 657 2939 666
rect 3077 657 3135 666
rect 3267 657 3325 666
rect 3457 657 3515 666
rect 2693 629 3515 657
rect 2693 620 2751 629
rect 2881 620 2939 629
rect 3077 620 3135 629
rect 3267 620 3325 629
rect 3457 620 3515 629
rect 4213 657 4271 666
rect 4403 657 4461 666
rect 4593 657 4651 666
rect 4789 657 4847 666
rect 4977 657 5035 666
rect 4213 629 5035 657
rect 4213 620 4271 629
rect 4403 620 4461 629
rect 4593 620 4651 629
rect 4789 620 4847 629
rect 4977 620 5035 629
rect 5361 657 5419 666
rect 5549 657 5607 666
rect 5745 657 5803 666
rect 5935 657 5993 666
rect 6125 657 6183 666
rect 5361 629 6183 657
rect 5361 620 5419 629
rect 5549 620 5607 629
rect 5745 620 5803 629
rect 5935 620 5993 629
rect 6125 620 6183 629
rect 6881 657 6939 666
rect 7071 657 7129 666
rect 7261 657 7319 666
rect 7457 657 7515 666
rect 7645 657 7703 666
rect 6881 629 7703 657
rect 6881 620 6939 629
rect 7071 620 7129 629
rect 7261 620 7319 629
rect 7457 620 7515 629
rect 7645 620 7703 629
rect 7937 657 7995 666
rect 8125 657 8183 666
rect 8321 657 8379 666
rect 8511 657 8569 666
rect 8701 657 8759 666
rect 7937 629 8759 657
rect 7937 620 7995 629
rect 8125 620 8183 629
rect 8321 620 8379 629
rect 8511 620 8569 629
rect 8701 620 8759 629
rect 9457 657 9515 666
rect 9647 657 9705 666
rect 9837 657 9895 666
rect 10033 657 10091 666
rect 10221 657 10279 666
rect 9457 629 10279 657
rect 9457 620 9515 629
rect 9647 620 9705 629
rect 9837 620 9895 629
rect 10033 620 10091 629
rect 10221 620 10279 629
rect 117 459 175 468
rect 305 459 363 468
rect 501 459 559 468
rect 691 459 749 468
rect 881 459 939 468
rect 117 431 939 459
rect 117 422 175 431
rect 305 422 363 431
rect 501 422 559 431
rect 691 422 749 431
rect 881 422 939 431
rect 1637 459 1695 468
rect 1827 459 1885 468
rect 2017 459 2075 468
rect 2213 459 2271 468
rect 2401 459 2459 468
rect 1637 431 2459 459
rect 1637 422 1695 431
rect 1827 422 1885 431
rect 2017 422 2075 431
rect 2213 422 2271 431
rect 2401 422 2459 431
rect 2693 459 2751 468
rect 2881 459 2939 468
rect 3077 459 3135 468
rect 3267 459 3325 468
rect 3457 459 3515 468
rect 2693 431 3515 459
rect 2693 422 2751 431
rect 2881 422 2939 431
rect 3077 422 3135 431
rect 3267 422 3325 431
rect 3457 422 3515 431
rect 4213 459 4271 468
rect 4403 459 4461 468
rect 4593 459 4651 468
rect 4789 459 4847 468
rect 4977 459 5035 468
rect 4213 431 5035 459
rect 4213 422 4271 431
rect 4403 422 4461 431
rect 4593 422 4651 431
rect 4789 422 4847 431
rect 4977 422 5035 431
rect 5361 459 5419 468
rect 5549 459 5607 468
rect 5745 459 5803 468
rect 5935 459 5993 468
rect 6125 459 6183 468
rect 5361 431 6183 459
rect 5361 422 5419 431
rect 5549 422 5607 431
rect 5745 422 5803 431
rect 5935 422 5993 431
rect 6125 422 6183 431
rect 6881 459 6939 468
rect 7071 459 7129 468
rect 7261 459 7319 468
rect 7457 459 7515 468
rect 7645 459 7703 468
rect 6881 431 7703 459
rect 6881 422 6939 431
rect 7071 422 7129 431
rect 7261 422 7319 431
rect 7457 422 7515 431
rect 7645 422 7703 431
rect 7937 459 7995 468
rect 8125 459 8183 468
rect 8321 459 8379 468
rect 8511 459 8569 468
rect 8701 459 8759 468
rect 7937 431 8759 459
rect 7937 422 7995 431
rect 8125 422 8183 431
rect 8321 422 8379 431
rect 8511 422 8569 431
rect 8701 422 8759 431
rect 9457 459 9515 468
rect 9647 459 9705 468
rect 9837 459 9895 468
rect 10033 459 10091 468
rect 10221 459 10279 468
rect 9457 431 10279 459
rect 9457 422 9515 431
rect 9647 422 9705 431
rect 9837 422 9895 431
rect 10033 422 10091 431
rect 10221 422 10279 431
<< labels >>
rlabel locali s 79 211 357 265 6 D[0]
port 1 nsew signal input
rlabel locali s 2219 211 2497 265 6 D[1]
port 2 nsew signal input
rlabel locali s 2655 211 2933 265 6 D[2]
port 3 nsew signal input
rlabel locali s 4795 211 5073 265 6 D[3]
port 4 nsew signal input
rlabel locali s 5323 211 5601 265 6 D[4]
port 5 nsew signal input
rlabel locali s 7463 211 7741 265 6 D[5]
port 6 nsew signal input
rlabel locali s 7899 211 8177 265 6 D[6]
port 7 nsew signal input
rlabel locali s 10039 211 10317 265 6 D[7]
port 8 nsew signal input
rlabel locali s 79 823 357 877 6 D[8]
port 9 nsew signal input
rlabel locali s 2219 823 2497 877 6 D[9]
port 10 nsew signal input
rlabel locali s 2655 823 2933 877 6 D[10]
port 11 nsew signal input
rlabel locali s 4795 823 5073 877 6 D[11]
port 12 nsew signal input
rlabel locali s 5323 823 5601 877 6 D[12]
port 13 nsew signal input
rlabel locali s 7463 823 7741 877 6 D[13]
port 14 nsew signal input
rlabel locali s 7899 823 8177 877 6 D[14]
port 15 nsew signal input
rlabel locali s 10039 823 10317 877 6 D[15]
port 16 nsew signal input
rlabel locali s 1152 199 1271 265 6 S[0]
port 17 nsew signal input
rlabel locali s 1305 199 1424 265 6 S[1]
port 18 nsew signal input
rlabel locali s 3728 199 3847 265 6 S[2]
port 19 nsew signal input
rlabel locali s 3881 199 4000 265 6 S[3]
port 20 nsew signal input
rlabel locali s 6396 199 6515 265 6 S[4]
port 21 nsew signal input
rlabel locali s 6549 199 6668 265 6 S[5]
port 22 nsew signal input
rlabel locali s 8972 199 9091 265 6 S[6]
port 23 nsew signal input
rlabel locali s 9125 199 9244 265 6 S[7]
port 24 nsew signal input
rlabel locali s 1152 823 1271 889 6 S[8]
port 25 nsew signal input
rlabel locali s 1305 823 1424 889 6 S[9]
port 26 nsew signal input
rlabel locali s 3728 823 3847 889 6 S[10]
port 27 nsew signal input
rlabel locali s 3881 823 4000 889 6 S[11]
port 28 nsew signal input
rlabel locali s 6396 823 6515 889 6 S[12]
port 29 nsew signal input
rlabel locali s 6549 823 6668 889 6 S[13]
port 30 nsew signal input
rlabel locali s 8972 823 9091 889 6 S[14]
port 31 nsew signal input
rlabel locali s 9125 823 9244 889 6 S[15]
port 32 nsew signal input
rlabel locali s 5169 53 5227 162 6 VNB
port 33 nsew
rlabel locali s 5169 926 5227 1035 6 VNB
port 33 nsew
rlabel locali s 5169 597 5227 794 6 VPB
port 34 nsew
rlabel locali s 5169 294 5227 491 6 VPB
port 34 nsew
rlabel viali s 797 697 831 731 6 Z
port 35 nsew signal output
rlabel viali s 797 357 831 391 6 Z
port 35 nsew signal output
rlabel viali s 609 697 643 731 6 Z
port 35 nsew signal output
rlabel viali s 609 357 643 391 6 Z
port 35 nsew signal output
rlabel locali s 781 273 847 815 6 Z
port 35 nsew signal output
rlabel locali s 741 875 807 969 6 Z
port 35 nsew signal output
rlabel locali s 741 119 807 213 6 Z
port 35 nsew signal output
rlabel locali s 593 875 639 911 6 Z
port 35 nsew signal output
rlabel locali s 593 815 847 875 6 Z
port 35 nsew signal output
rlabel locali s 593 273 659 815 6 Z
port 35 nsew signal output
rlabel locali s 593 213 847 273 6 Z
port 35 nsew signal output
rlabel locali s 593 177 639 213 6 Z
port 35 nsew signal output
rlabel locali s 573 911 639 969 6 Z
port 35 nsew signal output
rlabel locali s 573 119 639 177 6 Z
port 35 nsew signal output
rlabel metal1 s 9741 728 9799 737 6 Z
port 35 nsew signal output
rlabel metal1 s 9741 691 9799 700 6 Z
port 35 nsew signal output
rlabel metal1 s 9741 388 9799 397 6 Z
port 35 nsew signal output
rlabel metal1 s 9741 351 9799 360 6 Z
port 35 nsew signal output
rlabel metal1 s 9553 728 9611 737 6 Z
port 35 nsew signal output
rlabel metal1 s 9553 691 9611 700 6 Z
port 35 nsew signal output
rlabel metal1 s 9553 388 9611 397 6 Z
port 35 nsew signal output
rlabel metal1 s 9553 351 9611 360 6 Z
port 35 nsew signal output
rlabel metal1 s 8605 728 8663 737 6 Z
port 35 nsew signal output
rlabel metal1 s 8605 691 8663 700 6 Z
port 35 nsew signal output
rlabel metal1 s 8605 388 8663 397 6 Z
port 35 nsew signal output
rlabel metal1 s 8605 351 8663 360 6 Z
port 35 nsew signal output
rlabel metal1 s 8417 728 8475 737 6 Z
port 35 nsew signal output
rlabel metal1 s 8417 691 8475 700 6 Z
port 35 nsew signal output
rlabel metal1 s 8417 388 8475 397 6 Z
port 35 nsew signal output
rlabel metal1 s 8417 351 8475 360 6 Z
port 35 nsew signal output
rlabel metal1 s 7165 728 7223 737 6 Z
port 35 nsew signal output
rlabel metal1 s 7165 691 7223 700 6 Z
port 35 nsew signal output
rlabel metal1 s 7165 388 7223 397 6 Z
port 35 nsew signal output
rlabel metal1 s 7165 351 7223 360 6 Z
port 35 nsew signal output
rlabel metal1 s 6977 728 7035 737 6 Z
port 35 nsew signal output
rlabel metal1 s 6977 691 7035 700 6 Z
port 35 nsew signal output
rlabel metal1 s 6977 388 7035 397 6 Z
port 35 nsew signal output
rlabel metal1 s 6977 351 7035 360 6 Z
port 35 nsew signal output
rlabel metal1 s 6029 728 6087 737 6 Z
port 35 nsew signal output
rlabel metal1 s 6029 691 6087 700 6 Z
port 35 nsew signal output
rlabel metal1 s 6029 388 6087 397 6 Z
port 35 nsew signal output
rlabel metal1 s 6029 351 6087 360 6 Z
port 35 nsew signal output
rlabel metal1 s 5841 728 5899 737 6 Z
port 35 nsew signal output
rlabel metal1 s 5841 691 5899 700 6 Z
port 35 nsew signal output
rlabel metal1 s 5841 388 5899 397 6 Z
port 35 nsew signal output
rlabel metal1 s 5841 351 5899 360 6 Z
port 35 nsew signal output
rlabel metal1 s 4497 728 4555 737 6 Z
port 35 nsew signal output
rlabel metal1 s 4497 691 4555 700 6 Z
port 35 nsew signal output
rlabel metal1 s 4497 388 4555 397 6 Z
port 35 nsew signal output
rlabel metal1 s 4497 351 4555 360 6 Z
port 35 nsew signal output
rlabel metal1 s 4309 728 4367 737 6 Z
port 35 nsew signal output
rlabel metal1 s 4309 691 4367 700 6 Z
port 35 nsew signal output
rlabel metal1 s 4309 388 4367 397 6 Z
port 35 nsew signal output
rlabel metal1 s 4309 351 4367 360 6 Z
port 35 nsew signal output
rlabel metal1 s 3361 728 3419 737 6 Z
port 35 nsew signal output
rlabel metal1 s 3361 691 3419 700 6 Z
port 35 nsew signal output
rlabel metal1 s 3361 388 3419 397 6 Z
port 35 nsew signal output
rlabel metal1 s 3361 351 3419 360 6 Z
port 35 nsew signal output
rlabel metal1 s 3173 728 3231 737 6 Z
port 35 nsew signal output
rlabel metal1 s 3173 691 3231 700 6 Z
port 35 nsew signal output
rlabel metal1 s 3173 388 3231 397 6 Z
port 35 nsew signal output
rlabel metal1 s 3173 351 3231 360 6 Z
port 35 nsew signal output
rlabel metal1 s 1921 728 1979 737 6 Z
port 35 nsew signal output
rlabel metal1 s 1921 691 1979 700 6 Z
port 35 nsew signal output
rlabel metal1 s 1921 388 1979 397 6 Z
port 35 nsew signal output
rlabel metal1 s 1921 351 1979 360 6 Z
port 35 nsew signal output
rlabel metal1 s 1733 728 1791 737 6 Z
port 35 nsew signal output
rlabel metal1 s 1733 691 1791 700 6 Z
port 35 nsew signal output
rlabel metal1 s 1733 388 1791 397 6 Z
port 35 nsew signal output
rlabel metal1 s 1733 351 1791 360 6 Z
port 35 nsew signal output
rlabel metal1 s 785 728 843 737 6 Z
port 35 nsew signal output
rlabel metal1 s 785 691 843 700 6 Z
port 35 nsew signal output
rlabel metal1 s 785 388 843 397 6 Z
port 35 nsew signal output
rlabel metal1 s 785 351 843 360 6 Z
port 35 nsew signal output
rlabel metal1 s 597 728 655 737 6 Z
port 35 nsew signal output
rlabel metal1 s 597 700 9799 728 6 Z
port 35 nsew signal output
rlabel metal1 s 597 691 655 700 6 Z
port 35 nsew signal output
rlabel metal1 s 597 388 655 397 6 Z
port 35 nsew signal output
rlabel metal1 s 597 360 9799 388 6 Z
port 35 nsew signal output
rlabel metal1 s 597 351 655 360 6 Z
port 35 nsew signal output
rlabel viali s 10333 -17 10367 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 10241 -17 10275 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 10149 -17 10183 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 10057 -17 10091 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 9965 -17 9999 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 9873 -17 9907 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 9781 -17 9815 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 9689 -17 9723 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 9597 -17 9631 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 9505 -17 9539 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 9413 -17 9447 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 9321 -17 9355 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 9229 -17 9263 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 9137 -17 9171 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 9045 -17 9079 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 8953 -17 8987 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 8861 -17 8895 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 8769 -17 8803 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 8677 -17 8711 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 8585 -17 8619 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 8493 -17 8527 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 8401 -17 8435 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 8309 -17 8343 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 8217 -17 8251 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 8125 -17 8159 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 8033 -17 8067 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 7941 -17 7975 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 7849 -17 7883 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 7757 -17 7791 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 7665 -17 7699 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 7573 -17 7607 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 7481 -17 7515 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 7389 -17 7423 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 7297 -17 7331 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 7205 -17 7239 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 7113 -17 7147 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 7021 -17 7055 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 6929 -17 6963 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 6837 -17 6871 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 6745 -17 6779 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 6653 -17 6687 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 6561 -17 6595 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 6469 -17 6503 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 6377 -17 6411 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 6285 -17 6319 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 6193 -17 6227 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 6101 -17 6135 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 6009 -17 6043 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 5917 -17 5951 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 5825 -17 5859 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 5733 -17 5767 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 5641 -17 5675 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 5549 -17 5583 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 5457 -17 5491 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 5365 -17 5399 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 5273 -17 5307 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 5181 -17 5215 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 5089 -17 5123 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 4997 -17 5031 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 4905 -17 4939 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 4813 -17 4847 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 4721 -17 4755 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 4629 -17 4663 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 4537 -17 4571 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 4445 -17 4479 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 4353 -17 4387 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 4261 -17 4295 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 4169 -17 4203 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 4077 -17 4111 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 3985 -17 4019 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 3893 -17 3927 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 3801 -17 3835 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 3709 -17 3743 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 3617 -17 3651 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 3525 -17 3559 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 3433 -17 3467 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 3341 -17 3375 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 3249 -17 3283 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 3157 -17 3191 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 3065 -17 3099 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 2973 -17 3007 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 2881 -17 2915 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 2789 -17 2823 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 2697 -17 2731 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 2605 -17 2639 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 2513 -17 2547 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 2421 -17 2455 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 2329 -17 2363 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 2237 -17 2271 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 2145 -17 2179 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 2053 -17 2087 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 1961 -17 1995 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 1869 -17 1903 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 1777 -17 1811 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 1685 -17 1719 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 1593 -17 1627 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 1501 -17 1535 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 1409 -17 1443 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 1317 -17 1351 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 1225 -17 1259 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 1133 -17 1167 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 1041 -17 1075 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 949 -17 983 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 857 -17 891 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 765 -17 799 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 673 -17 707 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 581 -17 615 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 489 -17 523 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 397 -17 431 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 305 -17 339 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 213 -17 247 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 121 -17 155 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 29 -17 63 17 8 VGND
port 36 nsew ground bidirectional
rlabel locali s 10317 17 10367 177 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 10129 17 10183 109 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 9945 17 9995 109 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 9346 17 9404 122 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 9162 17 9220 122 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 8996 17 9054 122 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 8812 17 8870 122 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 8221 17 8271 109 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 8033 17 8087 109 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 7849 17 7899 177 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 7741 17 7791 177 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 7553 17 7607 109 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 7369 17 7419 109 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 6770 17 6828 122 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 6586 17 6644 122 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 6420 17 6478 122 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 6236 17 6294 122 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 5645 17 5695 109 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 5457 17 5511 109 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 5273 17 5323 177 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 5073 17 5123 177 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 4885 17 4939 109 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 4701 17 4751 109 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 4102 17 4160 122 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 3918 17 3976 122 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 3752 17 3810 122 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 3568 17 3626 122 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 2977 17 3027 109 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 2789 17 2843 109 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 2605 17 2655 177 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 2497 17 2547 177 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 2309 17 2363 109 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 2125 17 2175 109 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 1526 17 1584 122 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 1342 17 1400 122 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 1176 17 1234 122 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 992 17 1050 122 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 401 17 451 109 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 213 17 267 109 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 29 17 79 177 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 0 -17 10396 17 8 VGND
port 36 nsew ground bidirectional
rlabel viali s 10333 1071 10367 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 10241 1071 10275 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 10149 1071 10183 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 10057 1071 10091 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 9965 1071 9999 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 9873 1071 9907 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 9781 1071 9815 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 9689 1071 9723 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 9597 1071 9631 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 9505 1071 9539 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 9413 1071 9447 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 9321 1071 9355 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 9229 1071 9263 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 9137 1071 9171 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 9045 1071 9079 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 8953 1071 8987 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 8861 1071 8895 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 8769 1071 8803 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 8677 1071 8711 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 8585 1071 8619 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 8493 1071 8527 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 8401 1071 8435 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 8309 1071 8343 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 8217 1071 8251 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 8125 1071 8159 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 8033 1071 8067 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 7941 1071 7975 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 7849 1071 7883 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 7757 1071 7791 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 7665 1071 7699 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 7573 1071 7607 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 7481 1071 7515 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 7389 1071 7423 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 7297 1071 7331 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 7205 1071 7239 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 7113 1071 7147 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 7021 1071 7055 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 6929 1071 6963 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 6837 1071 6871 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 6745 1071 6779 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 6653 1071 6687 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 6561 1071 6595 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 6469 1071 6503 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 6377 1071 6411 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 6285 1071 6319 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 6193 1071 6227 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 6101 1071 6135 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 6009 1071 6043 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 5917 1071 5951 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 5825 1071 5859 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 5733 1071 5767 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 5641 1071 5675 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 5549 1071 5583 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 5457 1071 5491 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 5365 1071 5399 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 5273 1071 5307 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 5181 1071 5215 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 5089 1071 5123 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 4997 1071 5031 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 4905 1071 4939 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 4813 1071 4847 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 4721 1071 4755 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 4629 1071 4663 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 4537 1071 4571 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 4445 1071 4479 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 4353 1071 4387 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 4261 1071 4295 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 4169 1071 4203 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 4077 1071 4111 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 3985 1071 4019 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 3893 1071 3927 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 3801 1071 3835 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 3709 1071 3743 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 3617 1071 3651 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 3525 1071 3559 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 3433 1071 3467 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 3341 1071 3375 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 3249 1071 3283 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 3157 1071 3191 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 3065 1071 3099 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 2973 1071 3007 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 2881 1071 2915 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 2789 1071 2823 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 2697 1071 2731 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 2605 1071 2639 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 2513 1071 2547 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 2421 1071 2455 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 2329 1071 2363 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 2237 1071 2271 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 2145 1071 2179 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 2053 1071 2087 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 1961 1071 1995 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 1869 1071 1903 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 1777 1071 1811 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 1685 1071 1719 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 1593 1071 1627 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 1501 1071 1535 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 1409 1071 1443 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 1317 1071 1351 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 1225 1071 1259 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 1133 1071 1167 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 1041 1071 1075 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 949 1071 983 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 857 1071 891 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 765 1071 799 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 673 1071 707 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 581 1071 615 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 489 1071 523 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 397 1071 431 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 305 1071 339 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 213 1071 247 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 121 1071 155 1105 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 29 1071 63 1105 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 10317 911 10367 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 10129 979 10183 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 9945 979 9995 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 9346 966 9404 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 9162 966 9220 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 8996 966 9054 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 8812 966 8870 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 8221 979 8271 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 8033 979 8087 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 7849 911 7899 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 7741 911 7791 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 7553 979 7607 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 7369 979 7419 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 6770 966 6828 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 6586 966 6644 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 6420 966 6478 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 6236 966 6294 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 5645 979 5695 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 5457 979 5511 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 5273 911 5323 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 5073 911 5123 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 4885 979 4939 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 4701 979 4751 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 4102 966 4160 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 3918 966 3976 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 3752 966 3810 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 3568 966 3626 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 2977 979 3027 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 2789 979 2843 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 2605 911 2655 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 2497 911 2547 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 2309 979 2363 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 2125 979 2175 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 1526 966 1584 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 1342 966 1400 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 1176 966 1234 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 992 966 1050 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 401 979 451 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 213 979 267 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 29 911 79 1071 6 VGND
port 36 nsew ground bidirectional
rlabel locali s 0 1071 10396 1105 6 VGND
port 36 nsew ground bidirectional
rlabel metal1 s 0 -48 10396 48 8 VGND
port 36 nsew ground bidirectional
rlabel metal1 s 0 1040 10396 1136 6 VGND
port 36 nsew ground bidirectional
rlabel viali s 489 527 523 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 397 527 431 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 305 527 339 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 213 527 247 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 121 527 155 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 29 527 63 561 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 401 561 455 721 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 401 367 455 527 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 213 561 267 721 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 213 367 267 527 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 25 561 79 789 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 25 299 79 527 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 0 527 559 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 3065 527 3099 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 2973 527 3007 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 2881 527 2915 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 2789 527 2823 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 2697 527 2731 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 2605 527 2639 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 2513 527 2547 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 2421 527 2455 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 2329 527 2363 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 2237 527 2271 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 2145 527 2179 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 2053 527 2087 561 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 2977 561 3031 721 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 2977 367 3031 527 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 2789 561 2843 721 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 2789 367 2843 527 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 2601 561 2655 789 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 2601 299 2655 527 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 2497 561 2551 789 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 2497 299 2551 527 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 2309 561 2363 721 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 2309 367 2363 527 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 2121 561 2175 721 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 2121 367 2175 527 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 2017 527 3135 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 5733 527 5767 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 5641 527 5675 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 5549 527 5583 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 5457 527 5491 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 5365 527 5399 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 5273 527 5307 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 5181 527 5215 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 5089 527 5123 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 4997 527 5031 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 4905 527 4939 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 4813 527 4847 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 4721 527 4755 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 4629 527 4663 561 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 5645 561 5699 721 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 5645 367 5699 527 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 5457 561 5511 721 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 5457 367 5511 527 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 5269 561 5323 789 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 5269 299 5323 527 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 5073 561 5127 789 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 5073 299 5127 527 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 4885 561 4939 721 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 4885 367 4939 527 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 4697 561 4751 721 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 4697 367 4751 527 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 4593 527 5803 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 8309 527 8343 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 8217 527 8251 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 8125 527 8159 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 8033 527 8067 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 7941 527 7975 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 7849 527 7883 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 7757 527 7791 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 7665 527 7699 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 7573 527 7607 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 7481 527 7515 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 7389 527 7423 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 7297 527 7331 561 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 8221 561 8275 721 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 8221 367 8275 527 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 8033 561 8087 721 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 8033 367 8087 527 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 7845 561 7899 789 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 7845 299 7899 527 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 7741 561 7795 789 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 7741 299 7795 527 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 7553 561 7607 721 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 7553 367 7607 527 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 7365 561 7419 721 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 7365 367 7419 527 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 7261 527 8379 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 10333 527 10367 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 10241 527 10275 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 10149 527 10183 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 10057 527 10091 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 9965 527 9999 561 6 VPWR
port 37 nsew power bidirectional
rlabel viali s 9873 527 9907 561 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 10317 561 10371 789 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 10317 299 10371 527 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 10129 561 10183 721 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 10129 367 10183 527 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 9941 561 9995 721 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 9941 367 9995 527 6 VPWR
port 37 nsew power bidirectional
rlabel locali s 9837 527 10396 561 6 VPWR
port 37 nsew power bidirectional
rlabel metal1 s 0 496 10396 592 6 VPWR
port 37 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 10396 1088
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3268980
string GDS_START 3118284
<< end >>
