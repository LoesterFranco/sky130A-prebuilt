magic
tech sky130A
magscale 1 2
timestamp 1601050056
<< nwell >>
rect -38 332 806 704
<< pwell >>
rect 0 0 768 49
<< scpmos >>
rect 83 368 119 536
rect 192 368 228 592
rect 282 368 318 592
rect 459 368 495 568
rect 549 368 585 568
rect 651 368 687 568
<< nmoslvt >>
rect 82 74 112 184
rect 177 74 207 222
rect 263 74 293 222
rect 457 74 487 222
rect 543 74 573 222
rect 657 74 687 222
<< ndiff >>
rect 127 184 177 222
rect 27 146 82 184
rect 27 112 37 146
rect 71 112 82 146
rect 27 74 82 112
rect 112 139 177 184
rect 112 105 123 139
rect 157 105 177 139
rect 112 74 177 105
rect 207 210 263 222
rect 207 176 218 210
rect 252 176 263 210
rect 207 120 263 176
rect 207 86 218 120
rect 252 86 263 120
rect 207 74 263 86
rect 293 145 348 222
rect 293 111 304 145
rect 338 111 348 145
rect 293 74 348 111
rect 402 210 457 222
rect 402 176 412 210
rect 446 176 457 210
rect 402 120 457 176
rect 402 86 412 120
rect 446 86 457 120
rect 402 74 457 86
rect 487 136 543 222
rect 487 102 498 136
rect 532 102 543 136
rect 487 74 543 102
rect 573 84 657 222
rect 573 74 598 84
rect 588 50 598 74
rect 632 74 657 84
rect 687 202 741 222
rect 687 168 698 202
rect 732 168 741 202
rect 687 120 741 168
rect 687 86 698 120
rect 732 86 741 120
rect 687 74 741 86
rect 632 50 642 74
rect 588 38 642 50
<< pdiff >>
rect 134 566 192 592
rect 134 536 146 566
rect 27 524 83 536
rect 27 490 39 524
rect 73 490 83 524
rect 27 440 83 490
rect 27 406 39 440
rect 73 406 83 440
rect 27 368 83 406
rect 119 532 146 536
rect 180 532 192 566
rect 119 368 192 532
rect 228 414 282 592
rect 228 380 238 414
rect 272 380 282 414
rect 228 368 282 380
rect 318 568 438 592
rect 318 560 459 568
rect 318 526 329 560
rect 363 526 397 560
rect 431 526 459 560
rect 318 368 459 526
rect 495 556 549 568
rect 495 522 505 556
rect 539 522 549 556
rect 495 485 549 522
rect 495 451 505 485
rect 539 451 549 485
rect 495 414 549 451
rect 495 380 505 414
rect 539 380 549 414
rect 495 368 549 380
rect 585 368 651 568
rect 687 556 741 568
rect 687 522 697 556
rect 731 522 741 556
rect 687 485 741 522
rect 687 451 697 485
rect 731 451 741 485
rect 687 414 741 451
rect 687 380 697 414
rect 731 380 741 414
rect 687 368 741 380
<< ndiffc >>
rect 37 112 71 146
rect 123 105 157 139
rect 218 176 252 210
rect 218 86 252 120
rect 304 111 338 145
rect 412 176 446 210
rect 412 86 446 120
rect 498 102 532 136
rect 598 50 632 84
rect 698 168 732 202
rect 698 86 732 120
<< pdiffc >>
rect 39 490 73 524
rect 39 406 73 440
rect 146 532 180 566
rect 238 380 272 414
rect 329 526 363 560
rect 397 526 431 560
rect 505 522 539 556
rect 505 451 539 485
rect 505 380 539 414
rect 697 522 731 556
rect 697 451 731 485
rect 697 380 731 414
<< poly >>
rect 192 592 228 618
rect 282 592 318 618
rect 83 536 119 562
rect 459 568 495 594
rect 549 568 585 594
rect 651 568 687 594
rect 83 326 119 368
rect 25 310 119 326
rect 192 320 228 368
rect 282 326 318 368
rect 459 336 495 368
rect 270 320 336 326
rect 25 276 41 310
rect 75 276 119 310
rect 25 260 119 276
rect 177 310 336 320
rect 177 276 286 310
rect 320 276 336 310
rect 177 269 336 276
rect 378 320 495 336
rect 378 286 394 320
rect 428 286 495 320
rect 549 310 585 368
rect 651 310 687 368
rect 378 270 495 286
rect 543 294 609 310
rect 82 184 112 260
rect 177 222 207 269
rect 263 260 336 269
rect 263 222 293 260
rect 457 222 487 270
rect 543 260 559 294
rect 593 260 609 294
rect 543 244 609 260
rect 657 294 747 310
rect 657 260 697 294
rect 731 260 747 294
rect 657 244 747 260
rect 543 222 573 244
rect 657 222 687 244
rect 82 48 112 74
rect 177 48 207 74
rect 263 48 293 74
rect 457 48 487 74
rect 543 48 573 74
rect 657 48 687 74
<< polycont >>
rect 41 276 75 310
rect 286 276 320 310
rect 394 286 428 320
rect 559 260 593 294
rect 697 260 731 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 130 566 196 649
rect 23 524 89 540
rect 23 490 39 524
rect 73 490 89 524
rect 130 532 146 566
rect 180 532 196 566
rect 130 516 196 532
rect 313 560 447 649
rect 313 526 329 560
rect 363 526 397 560
rect 431 526 447 560
rect 313 516 447 526
rect 489 556 555 572
rect 489 522 505 556
rect 539 522 555 556
rect 23 482 89 490
rect 489 485 555 522
rect 489 482 505 485
rect 23 448 442 482
rect 23 440 159 448
rect 23 406 39 440
rect 73 406 159 440
rect 23 390 159 406
rect 25 310 91 356
rect 25 276 41 310
rect 75 276 91 310
rect 25 260 91 276
rect 125 226 159 390
rect 21 192 159 226
rect 202 380 238 414
rect 272 380 288 414
rect 202 364 288 380
rect 202 226 236 364
rect 270 310 336 326
rect 270 276 286 310
rect 320 276 336 310
rect 270 260 336 276
rect 378 320 442 448
rect 378 286 394 320
rect 428 286 442 320
rect 378 270 442 286
rect 476 451 505 482
rect 539 451 555 485
rect 476 414 555 451
rect 476 380 505 414
rect 539 380 555 414
rect 476 364 555 380
rect 681 556 747 649
rect 681 522 697 556
rect 731 522 747 556
rect 681 485 747 522
rect 681 451 697 485
rect 731 451 747 485
rect 681 414 747 451
rect 681 380 697 414
rect 731 380 747 414
rect 681 364 747 380
rect 302 236 336 260
rect 476 236 510 364
rect 544 294 647 310
rect 544 260 559 294
rect 593 260 647 294
rect 544 236 647 260
rect 681 294 747 310
rect 681 260 697 294
rect 731 260 747 294
rect 681 236 747 260
rect 202 210 268 226
rect 21 146 71 192
rect 202 176 218 210
rect 252 176 268 210
rect 302 210 510 236
rect 302 202 412 210
rect 21 112 37 146
rect 21 91 71 112
rect 107 139 157 158
rect 107 105 123 139
rect 107 17 157 105
rect 202 120 268 176
rect 396 176 412 202
rect 446 202 510 210
rect 202 86 218 120
rect 252 86 268 120
rect 202 70 268 86
rect 304 145 354 164
rect 338 111 354 145
rect 304 17 354 111
rect 396 120 446 176
rect 682 168 698 202
rect 732 168 748 202
rect 396 86 412 120
rect 396 70 446 86
rect 482 136 748 168
rect 482 102 498 136
rect 532 134 748 136
rect 532 102 548 134
rect 482 70 548 102
rect 682 120 748 134
rect 582 84 648 100
rect 582 50 598 84
rect 632 50 648 84
rect 682 86 698 120
rect 732 86 748 120
rect 682 70 748 86
rect 582 17 648 50
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
rlabel comment s 0 0 0 0 4 o21ba_2
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 703 242 737 276 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 223 94 257 128 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 223 168 257 202 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 607 242 641 276 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 B1_N
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 768 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1017820
string GDS_START 1011190
<< end >>
