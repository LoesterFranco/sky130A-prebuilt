magic
tech sky130A
magscale 1 2
timestamp 1601050082
<< locali >>
rect 505 446 593 598
rect 727 446 773 598
rect 907 446 963 596
rect 505 412 963 446
rect 88 290 167 356
rect 897 404 963 412
rect 1103 404 1137 596
rect 897 398 1137 404
rect 1267 424 1333 596
rect 1467 424 1533 596
rect 1657 424 1723 596
rect 1837 424 1903 596
rect 1267 398 1903 424
rect 897 390 1903 398
rect 293 310 359 376
rect 897 370 1333 390
rect 1103 364 1333 370
rect 1467 364 1533 390
rect 1103 252 1137 364
rect 1369 330 1415 356
rect 1237 264 1522 330
rect 1653 260 1991 356
rect 667 218 1137 252
rect 667 208 701 218
rect 464 174 701 208
rect 464 119 530 174
rect 667 119 701 174
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 23 458 89 649
rect 129 424 163 596
rect 203 478 269 649
rect 303 444 359 596
rect 401 478 467 649
rect 627 480 693 649
rect 807 480 873 649
rect 20 390 163 424
rect 225 410 427 444
rect 997 438 1063 649
rect 20 256 54 390
rect 225 266 259 410
rect 393 378 427 410
rect 1177 432 1227 649
rect 1367 458 1433 649
rect 1573 458 1623 649
rect 1763 458 1797 649
rect 1943 390 1993 649
rect 393 344 863 378
rect 829 336 863 344
rect 431 276 633 310
rect 829 286 1069 336
rect 20 166 89 256
rect 225 200 284 266
rect 318 242 633 276
rect 318 166 352 242
rect 1225 226 1619 230
rect 20 132 352 166
rect 20 110 89 132
rect 125 17 191 98
rect 386 85 420 208
rect 1225 196 1993 226
rect 564 85 630 140
rect 737 150 1179 184
rect 737 85 787 150
rect 1113 119 1179 150
rect 1225 119 1275 196
rect 386 51 787 85
rect 823 85 1077 116
rect 1311 85 1377 162
rect 1413 119 1447 196
rect 1585 192 1993 196
rect 1483 85 1549 162
rect 823 51 1549 85
rect 1585 70 1619 192
rect 1655 17 1721 158
rect 1757 70 1791 192
rect 1827 17 1893 158
rect 1927 70 1993 192
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
rlabel locali s 88 290 167 356 6 A_N
port 1 nsew signal input
rlabel locali s 293 310 359 376 6 B_N
port 2 nsew signal input
rlabel locali s 1369 330 1415 356 6 C
port 3 nsew signal input
rlabel locali s 1237 264 1522 330 6 C
port 3 nsew signal input
rlabel locali s 1653 260 1991 356 6 D
port 4 nsew signal input
rlabel locali s 1837 424 1903 596 6 Y
port 5 nsew signal output
rlabel locali s 1657 424 1723 596 6 Y
port 5 nsew signal output
rlabel locali s 1467 424 1533 596 6 Y
port 5 nsew signal output
rlabel locali s 1467 364 1533 390 6 Y
port 5 nsew signal output
rlabel locali s 1267 424 1333 596 6 Y
port 5 nsew signal output
rlabel locali s 1267 398 1903 424 6 Y
port 5 nsew signal output
rlabel locali s 1103 404 1137 596 6 Y
port 5 nsew signal output
rlabel locali s 1103 364 1333 370 6 Y
port 5 nsew signal output
rlabel locali s 1103 252 1137 364 6 Y
port 5 nsew signal output
rlabel locali s 907 446 963 596 6 Y
port 5 nsew signal output
rlabel locali s 897 404 963 412 6 Y
port 5 nsew signal output
rlabel locali s 897 398 1137 404 6 Y
port 5 nsew signal output
rlabel locali s 897 390 1903 398 6 Y
port 5 nsew signal output
rlabel locali s 897 370 1333 390 6 Y
port 5 nsew signal output
rlabel locali s 727 446 773 598 6 Y
port 5 nsew signal output
rlabel locali s 667 218 1137 252 6 Y
port 5 nsew signal output
rlabel locali s 667 208 701 218 6 Y
port 5 nsew signal output
rlabel locali s 667 119 701 174 6 Y
port 5 nsew signal output
rlabel locali s 505 446 593 598 6 Y
port 5 nsew signal output
rlabel locali s 505 412 963 446 6 Y
port 5 nsew signal output
rlabel locali s 464 174 701 208 6 Y
port 5 nsew signal output
rlabel locali s 464 119 530 174 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -49 2016 49 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 617 2016 715 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2016 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1856124
string GDS_START 1840250
<< end >>
