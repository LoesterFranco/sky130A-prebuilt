magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1380 561
rect 103 427 169 527
rect 18 197 66 325
rect 103 17 169 93
rect 396 367 459 527
rect 756 435 790 527
rect 289 191 357 265
rect 944 366 994 527
rect 1028 334 1096 493
rect 1062 149 1096 334
rect 375 17 446 89
rect 753 17 819 122
rect 928 17 994 99
rect 1028 83 1096 149
rect 1218 367 1277 527
rect 1311 301 1363 493
rect 1325 165 1363 301
rect 1218 17 1277 109
rect 1311 51 1363 165
rect 0 -17 1380 17
<< obsli1 >>
rect 35 393 69 493
rect 35 359 156 393
rect 122 323 156 359
rect 122 280 156 289
rect 203 391 248 493
rect 203 357 214 391
rect 203 337 248 357
rect 122 214 168 280
rect 122 161 156 214
rect 35 127 156 161
rect 35 69 69 127
rect 203 69 237 337
rect 296 333 362 483
rect 584 426 722 455
rect 584 423 723 426
rect 584 421 724 423
rect 672 418 725 421
rect 672 415 726 418
rect 675 412 726 415
rect 684 406 726 412
rect 686 403 726 406
rect 499 391 556 401
rect 533 357 556 391
rect 296 299 433 333
rect 399 247 433 299
rect 499 271 556 357
rect 590 323 658 382
rect 590 289 591 323
rect 625 289 658 323
rect 590 283 658 289
rect 399 181 473 247
rect 590 207 624 283
rect 692 265 726 403
rect 860 373 910 487
rect 760 324 910 373
rect 760 307 916 324
rect 879 265 916 307
rect 692 233 845 265
rect 399 157 433 181
rect 307 123 433 157
rect 513 141 624 207
rect 671 199 845 233
rect 879 199 1028 265
rect 307 69 341 123
rect 671 107 705 199
rect 879 168 916 199
rect 860 132 916 168
rect 558 73 705 107
rect 860 83 894 132
rect 1132 265 1182 493
rect 1132 199 1291 265
rect 1132 51 1182 199
<< obsli1c >>
rect 122 289 156 323
rect 214 357 248 391
rect 499 357 533 391
rect 591 289 625 323
<< metal1 >>
rect 0 496 1380 592
rect 0 -48 1380 48
<< obsm1 >>
rect 202 391 260 397
rect 202 357 214 391
rect 248 388 260 391
rect 487 391 545 397
rect 487 388 499 391
rect 248 360 499 388
rect 248 357 260 360
rect 202 351 260 357
rect 487 357 499 360
rect 533 357 545 391
rect 487 351 545 357
rect 110 323 168 329
rect 110 289 122 323
rect 156 320 168 323
rect 579 323 637 329
rect 579 320 591 323
rect 156 292 591 320
rect 156 289 168 292
rect 110 283 168 289
rect 579 289 591 292
rect 625 289 637 323
rect 579 283 637 289
<< labels >>
rlabel locali s 289 191 357 265 6 D
port 1 nsew signal input
rlabel locali s 1062 149 1096 334 6 Q
port 2 nsew signal output
rlabel locali s 1028 334 1096 493 6 Q
port 2 nsew signal output
rlabel locali s 1028 83 1096 149 6 Q
port 2 nsew signal output
rlabel locali s 1325 165 1363 301 6 Q_N
port 3 nsew signal output
rlabel locali s 1311 301 1363 493 6 Q_N
port 3 nsew signal output
rlabel locali s 1311 51 1363 165 6 Q_N
port 3 nsew signal output
rlabel locali s 18 197 66 325 6 GATE_N
port 4 nsew clock input
rlabel locali s 1218 17 1277 109 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 928 17 994 99 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 753 17 819 122 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 375 17 446 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 103 17 169 93 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 1380 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1380 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 1218 367 1277 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 944 366 994 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 756 435 790 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 396 367 459 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 103 427 169 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 1380 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 1380 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1380 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2737950
string GDS_START 2724948
<< end >>
