magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1564 561
rect 17 367 69 527
rect 103 333 169 493
rect 203 367 237 527
rect 271 333 337 493
rect 17 293 337 333
rect 371 293 405 527
rect 543 367 593 527
rect 17 181 69 293
rect 1331 357 1397 527
rect 567 215 633 255
rect 682 215 808 255
rect 866 215 992 255
rect 1030 215 1272 255
rect 1330 215 1547 255
rect 17 143 337 181
rect 17 17 69 109
rect 103 51 169 143
rect 203 17 237 109
rect 271 51 337 143
rect 371 17 421 177
rect 731 17 775 109
rect 889 17 943 109
rect 1061 17 1183 109
rect 1337 17 1391 109
rect 0 -17 1564 17
<< obsli1 >>
rect 439 323 509 493
rect 627 459 865 493
rect 627 367 681 459
rect 715 323 765 425
rect 439 289 765 323
rect 799 323 865 459
rect 899 459 1229 493
rect 899 357 933 459
rect 967 323 1033 423
rect 799 289 1033 323
rect 1079 323 1129 423
rect 1163 357 1229 459
rect 1263 323 1297 491
rect 1453 323 1519 493
rect 1079 289 1519 323
rect 439 259 509 289
rect 103 249 509 259
rect 103 215 533 249
rect 459 181 533 215
rect 459 127 609 181
rect 647 147 1519 181
rect 647 93 697 147
rect 459 51 697 93
rect 815 51 849 147
rect 983 51 1017 147
rect 1248 51 1282 147
rect 1453 51 1519 147
<< metal1 >>
rect 0 496 1564 592
rect 0 -48 1564 48
<< labels >>
rlabel locali s 1330 215 1547 255 6 A1
port 1 nsew signal input
rlabel locali s 1030 215 1272 255 6 A2
port 2 nsew signal input
rlabel locali s 866 215 992 255 6 A3
port 3 nsew signal input
rlabel locali s 682 215 808 255 6 A4
port 4 nsew signal input
rlabel locali s 567 215 633 255 6 B1
port 5 nsew signal input
rlabel locali s 271 333 337 493 6 X
port 6 nsew signal output
rlabel locali s 271 51 337 143 6 X
port 6 nsew signal output
rlabel locali s 103 333 169 493 6 X
port 6 nsew signal output
rlabel locali s 103 51 169 143 6 X
port 6 nsew signal output
rlabel locali s 17 293 337 333 6 X
port 6 nsew signal output
rlabel locali s 17 181 69 293 6 X
port 6 nsew signal output
rlabel locali s 17 143 337 181 6 X
port 6 nsew signal output
rlabel locali s 1337 17 1391 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1061 17 1183 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 889 17 943 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 731 17 775 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 371 17 421 177 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 203 17 237 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 17 17 69 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 1564 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1564 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1331 357 1397 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 543 367 593 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 371 293 405 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 203 367 237 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 17 367 69 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 1564 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 1564 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1564 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 862506
string GDS_START 849402
<< end >>
