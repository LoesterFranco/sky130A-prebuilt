magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 276 561
rect 19 333 85 490
rect 19 299 155 333
rect 191 299 257 527
rect 17 215 87 265
rect 121 179 155 299
rect 189 215 259 265
rect 21 17 69 179
rect 103 51 169 179
rect 203 17 257 179
rect 0 -17 276 17
<< metal1 >>
rect 0 496 276 592
rect 0 -48 276 48
<< labels >>
rlabel locali s 189 215 259 265 6 A
port 1 nsew signal input
rlabel locali s 17 215 87 265 6 B
port 2 nsew signal input
rlabel locali s 121 179 155 299 6 Y
port 3 nsew signal output
rlabel locali s 103 51 169 179 6 Y
port 3 nsew signal output
rlabel locali s 19 333 85 490 6 Y
port 3 nsew signal output
rlabel locali s 19 299 155 333 6 Y
port 3 nsew signal output
rlabel locali s 203 17 257 179 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 21 17 69 179 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 276 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 276 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 191 299 257 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 276 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 276 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 276 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1930962
string GDS_START 1927356
<< end >>
