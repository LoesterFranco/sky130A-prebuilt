magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 37 289 71 527
rect 105 305 166 493
rect 200 447 276 527
rect 37 17 71 186
rect 105 162 149 305
rect 289 199 363 323
rect 397 199 467 275
rect 105 51 166 162
rect 735 435 785 527
rect 660 210 752 331
rect 816 153 891 331
rect 200 17 296 106
rect 431 17 578 97
rect 781 17 871 119
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< obsli1 >>
rect 540 474 574 493
rect 328 440 574 474
rect 625 451 691 485
rect 328 395 372 440
rect 200 361 372 395
rect 528 413 574 440
rect 200 265 244 361
rect 435 343 469 381
rect 528 379 620 413
rect 183 199 244 265
rect 435 309 542 343
rect 508 165 542 309
rect 353 131 542 165
rect 576 174 620 379
rect 657 401 691 451
rect 829 401 863 493
rect 657 367 863 401
rect 576 140 656 174
rect 353 51 387 131
rect 622 51 656 140
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
rlabel locali s 289 199 363 323 6 A1_N
port 1 nsew signal input
rlabel locali s 397 199 467 275 6 A2_N
port 2 nsew signal input
rlabel locali s 816 153 891 331 6 B1
port 3 nsew signal input
rlabel locali s 660 210 752 331 6 B2
port 4 nsew signal input
rlabel locali s 105 305 166 493 6 X
port 5 nsew signal output
rlabel locali s 105 162 149 305 6 X
port 5 nsew signal output
rlabel locali s 105 51 166 162 6 X
port 5 nsew signal output
rlabel metal1 s 0 -48 920 48 8 VGND
port 6 nsew ground bidirectional
rlabel locali s 781 17 871 119 6 VGND
port 6 nsew ground bidirectional
rlabel locali s 431 17 578 97 6 VGND
port 6 nsew ground bidirectional
rlabel locali s 200 17 296 106 6 VGND
port 6 nsew ground bidirectional
rlabel locali s 37 17 71 186 6 VGND
port 6 nsew ground bidirectional
rlabel locali s 0 -17 920 17 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 920 592 6 VPWR
port 7 nsew power bidirectional
rlabel locali s 735 435 785 527 6 VPWR
port 7 nsew power bidirectional
rlabel locali s 200 447 276 527 6 VPWR
port 7 nsew power bidirectional
rlabel locali s 37 289 71 527 6 VPWR
port 7 nsew power bidirectional
rlabel locali s 0 527 920 561 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 920 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1320010
string GDS_START 1311978
<< end >>
