magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1564 561
rect 103 383 169 527
rect 271 383 337 527
rect 439 383 505 527
rect 607 383 673 527
rect 779 383 845 527
rect 947 451 1013 527
rect 1215 383 1449 417
rect 24 199 347 265
rect 387 199 710 265
rect 765 199 1084 265
rect 1134 199 1371 326
rect 1409 161 1449 383
rect 795 127 1517 161
rect 103 17 169 93
rect 271 17 337 93
rect 1215 17 1281 93
rect 1315 51 1349 127
rect 1383 17 1449 93
rect 1483 51 1517 127
rect 0 -17 1564 17
<< obsli1 >>
rect 35 333 69 493
rect 203 333 237 493
rect 371 333 405 493
rect 539 333 573 493
rect 707 333 741 493
rect 879 333 913 493
rect 1047 485 1081 493
rect 1047 451 1533 485
rect 1047 333 1081 451
rect 35 299 1081 333
rect 1483 299 1533 451
rect 35 127 757 161
rect 35 51 69 127
rect 203 51 237 127
rect 371 51 405 127
rect 439 59 1113 93
<< metal1 >>
rect 0 496 1564 592
rect 0 -48 1564 48
<< labels >>
rlabel locali s 765 199 1084 265 6 A1
port 1 nsew signal input
rlabel locali s 387 199 710 265 6 A2
port 2 nsew signal input
rlabel locali s 24 199 347 265 6 A3
port 3 nsew signal input
rlabel locali s 1134 199 1371 326 6 B1
port 4 nsew signal input
rlabel locali s 1483 51 1517 127 6 Y
port 5 nsew signal output
rlabel locali s 1409 161 1449 383 6 Y
port 5 nsew signal output
rlabel locali s 1315 51 1349 127 6 Y
port 5 nsew signal output
rlabel locali s 1215 383 1449 417 6 Y
port 5 nsew signal output
rlabel locali s 795 127 1517 161 6 Y
port 5 nsew signal output
rlabel locali s 1383 17 1449 93 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1215 17 1281 93 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 271 17 337 93 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 103 17 169 93 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 1564 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1564 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 947 451 1013 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 779 383 845 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 607 383 673 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 439 383 505 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 271 383 337 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 103 383 169 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 1564 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 1564 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1564 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3531936
string GDS_START 3519070
<< end >>
