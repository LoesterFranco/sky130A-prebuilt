magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 93 47 123 177
rect 177 47 207 177
rect 281 47 311 177
rect 365 47 395 177
rect 573 47 603 177
rect 657 47 687 177
rect 761 47 791 177
rect 845 47 875 177
rect 949 47 979 177
rect 1033 47 1063 177
<< pmoshvt >>
rect 85 297 121 497
rect 179 297 215 497
rect 273 297 309 497
rect 367 297 403 497
rect 565 297 601 497
rect 659 297 695 497
rect 753 297 789 497
rect 847 297 883 497
rect 941 297 977 497
rect 1035 297 1071 497
<< ndiff >>
rect 27 163 93 177
rect 27 129 39 163
rect 73 129 93 163
rect 27 95 93 129
rect 27 61 39 95
rect 73 61 93 95
rect 27 47 93 61
rect 123 163 177 177
rect 123 129 133 163
rect 167 129 177 163
rect 123 95 177 129
rect 123 61 133 95
rect 167 61 177 95
rect 123 47 177 61
rect 207 95 281 177
rect 207 61 227 95
rect 261 61 281 95
rect 207 47 281 61
rect 311 163 365 177
rect 311 129 321 163
rect 355 129 365 163
rect 311 95 365 129
rect 311 61 321 95
rect 355 61 365 95
rect 311 47 365 61
rect 395 165 573 177
rect 395 131 529 165
rect 563 131 573 165
rect 395 95 573 131
rect 395 61 405 95
rect 439 93 573 95
rect 439 61 529 93
rect 395 59 529 61
rect 563 59 573 93
rect 395 47 573 59
rect 603 169 657 177
rect 603 135 613 169
rect 647 135 657 169
rect 603 101 657 135
rect 603 67 613 101
rect 647 67 657 101
rect 603 47 657 67
rect 687 101 761 177
rect 687 67 707 101
rect 741 67 761 101
rect 687 47 761 67
rect 791 169 845 177
rect 791 135 801 169
rect 835 135 845 169
rect 791 101 845 135
rect 791 67 801 101
rect 835 67 845 101
rect 791 47 845 67
rect 875 101 949 177
rect 875 67 895 101
rect 929 67 949 101
rect 875 47 949 67
rect 979 169 1033 177
rect 979 135 989 169
rect 1023 135 1033 169
rect 979 101 1033 135
rect 979 67 989 101
rect 1023 67 1033 101
rect 979 47 1033 67
rect 1063 101 1127 177
rect 1063 67 1083 101
rect 1117 67 1127 101
rect 1063 47 1127 67
<< pdiff >>
rect 27 477 85 497
rect 27 443 39 477
rect 73 443 85 477
rect 27 409 85 443
rect 27 375 39 409
rect 73 375 85 409
rect 27 341 85 375
rect 27 307 39 341
rect 73 307 85 341
rect 27 297 85 307
rect 121 485 179 497
rect 121 451 133 485
rect 167 451 179 485
rect 121 417 179 451
rect 121 383 133 417
rect 167 383 179 417
rect 121 297 179 383
rect 215 477 273 497
rect 215 443 227 477
rect 261 443 273 477
rect 215 409 273 443
rect 215 375 227 409
rect 261 375 273 409
rect 215 341 273 375
rect 215 307 227 341
rect 261 307 273 341
rect 215 297 273 307
rect 309 409 367 497
rect 309 375 321 409
rect 355 375 367 409
rect 309 341 367 375
rect 309 307 321 341
rect 355 307 367 341
rect 309 297 367 307
rect 403 485 457 497
rect 403 451 415 485
rect 449 451 457 485
rect 403 417 457 451
rect 403 383 415 417
rect 449 383 457 417
rect 403 297 457 383
rect 511 485 565 497
rect 511 451 519 485
rect 553 451 565 485
rect 511 417 565 451
rect 511 383 519 417
rect 553 383 565 417
rect 511 349 565 383
rect 511 315 519 349
rect 553 315 565 349
rect 511 297 565 315
rect 601 485 659 497
rect 601 451 613 485
rect 647 451 659 485
rect 601 417 659 451
rect 601 383 613 417
rect 647 383 659 417
rect 601 349 659 383
rect 601 315 613 349
rect 647 315 659 349
rect 601 297 659 315
rect 695 485 753 497
rect 695 451 707 485
rect 741 451 753 485
rect 695 417 753 451
rect 695 383 707 417
rect 741 383 753 417
rect 695 297 753 383
rect 789 485 847 497
rect 789 451 801 485
rect 835 451 847 485
rect 789 417 847 451
rect 789 383 801 417
rect 835 383 847 417
rect 789 349 847 383
rect 789 315 801 349
rect 835 315 847 349
rect 789 297 847 315
rect 883 485 941 497
rect 883 451 895 485
rect 929 451 941 485
rect 883 417 941 451
rect 883 383 895 417
rect 929 383 941 417
rect 883 297 941 383
rect 977 485 1035 497
rect 977 451 989 485
rect 1023 451 1035 485
rect 977 417 1035 451
rect 977 383 989 417
rect 1023 383 1035 417
rect 977 349 1035 383
rect 977 315 989 349
rect 1023 315 1035 349
rect 977 297 1035 315
rect 1071 485 1127 497
rect 1071 451 1083 485
rect 1117 451 1127 485
rect 1071 417 1127 451
rect 1071 383 1083 417
rect 1117 383 1127 417
rect 1071 297 1127 383
<< ndiffc >>
rect 39 129 73 163
rect 39 61 73 95
rect 133 129 167 163
rect 133 61 167 95
rect 227 61 261 95
rect 321 129 355 163
rect 321 61 355 95
rect 529 131 563 165
rect 405 61 439 95
rect 529 59 563 93
rect 613 135 647 169
rect 613 67 647 101
rect 707 67 741 101
rect 801 135 835 169
rect 801 67 835 101
rect 895 67 929 101
rect 989 135 1023 169
rect 989 67 1023 101
rect 1083 67 1117 101
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 133 451 167 485
rect 133 383 167 417
rect 227 443 261 477
rect 227 375 261 409
rect 227 307 261 341
rect 321 375 355 409
rect 321 307 355 341
rect 415 451 449 485
rect 415 383 449 417
rect 519 451 553 485
rect 519 383 553 417
rect 519 315 553 349
rect 613 451 647 485
rect 613 383 647 417
rect 613 315 647 349
rect 707 451 741 485
rect 707 383 741 417
rect 801 451 835 485
rect 801 383 835 417
rect 801 315 835 349
rect 895 451 929 485
rect 895 383 929 417
rect 989 451 1023 485
rect 989 383 1023 417
rect 989 315 1023 349
rect 1083 451 1117 485
rect 1083 383 1117 417
<< poly >>
rect 85 497 121 523
rect 179 497 215 523
rect 273 497 309 523
rect 367 497 403 523
rect 565 497 601 523
rect 659 497 695 523
rect 753 497 789 523
rect 847 497 883 523
rect 941 497 977 523
rect 1035 497 1071 523
rect 85 282 121 297
rect 179 282 215 297
rect 273 282 309 297
rect 367 282 403 297
rect 565 282 601 297
rect 659 282 695 297
rect 753 282 789 297
rect 847 282 883 297
rect 941 282 977 297
rect 1035 282 1071 297
rect 83 265 123 282
rect 177 265 217 282
rect 83 249 217 265
rect 83 215 99 249
rect 133 215 167 249
rect 201 215 217 249
rect 83 199 217 215
rect 271 265 311 282
rect 365 265 405 282
rect 271 249 405 265
rect 271 215 287 249
rect 321 215 355 249
rect 389 215 405 249
rect 271 199 405 215
rect 563 265 603 282
rect 657 265 697 282
rect 751 265 791 282
rect 845 265 885 282
rect 939 265 979 282
rect 1033 265 1073 282
rect 563 249 1073 265
rect 563 215 579 249
rect 613 215 647 249
rect 681 215 715 249
rect 749 215 783 249
rect 817 215 851 249
rect 885 215 919 249
rect 953 215 1073 249
rect 563 199 1073 215
rect 93 177 123 199
rect 177 177 207 199
rect 281 177 311 199
rect 365 177 395 199
rect 573 177 603 199
rect 657 177 687 199
rect 761 177 791 199
rect 845 177 875 199
rect 949 177 979 199
rect 1033 177 1063 199
rect 93 21 123 47
rect 177 21 207 47
rect 281 21 311 47
rect 365 21 395 47
rect 573 21 603 47
rect 657 21 687 47
rect 761 21 791 47
rect 845 21 875 47
rect 949 21 979 47
rect 1033 21 1063 47
<< polycont >>
rect 99 215 133 249
rect 167 215 201 249
rect 287 215 321 249
rect 355 215 389 249
rect 579 215 613 249
rect 647 215 681 249
rect 715 215 749 249
rect 783 215 817 249
rect 851 215 885 249
rect 919 215 953 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 18 477 83 493
rect 18 443 39 477
rect 73 443 83 477
rect 18 409 83 443
rect 18 375 39 409
rect 73 375 83 409
rect 18 341 83 375
rect 117 485 183 527
rect 117 451 133 485
rect 167 451 183 485
rect 117 417 183 451
rect 117 383 133 417
rect 167 383 183 417
rect 117 367 183 383
rect 217 485 465 493
rect 217 477 415 485
rect 217 443 227 477
rect 261 459 415 477
rect 261 443 271 459
rect 217 409 271 443
rect 405 451 415 459
rect 449 451 465 485
rect 217 375 227 409
rect 261 375 271 409
rect 18 307 39 341
rect 73 333 83 341
rect 217 341 271 375
rect 217 333 227 341
rect 73 307 227 333
rect 261 307 271 341
rect 18 291 271 307
rect 305 409 371 425
rect 305 375 321 409
rect 355 375 371 409
rect 305 341 371 375
rect 405 417 465 451
rect 405 383 415 417
rect 449 383 465 417
rect 405 367 465 383
rect 509 485 563 527
rect 509 451 519 485
rect 553 451 563 485
rect 509 417 563 451
rect 509 383 519 417
rect 553 383 563 417
rect 305 307 321 341
rect 355 333 371 341
rect 509 349 563 383
rect 355 307 475 333
rect 305 289 475 307
rect 509 315 519 349
rect 553 315 563 349
rect 509 299 563 315
rect 597 485 663 493
rect 597 451 613 485
rect 647 451 663 485
rect 597 417 663 451
rect 597 383 613 417
rect 647 383 663 417
rect 597 349 663 383
rect 697 485 751 527
rect 697 451 707 485
rect 741 451 751 485
rect 697 417 751 451
rect 697 383 707 417
rect 741 383 751 417
rect 697 367 751 383
rect 785 485 851 493
rect 785 451 801 485
rect 835 451 851 485
rect 785 417 851 451
rect 785 383 801 417
rect 835 383 851 417
rect 597 315 613 349
rect 647 333 663 349
rect 785 349 851 383
rect 885 485 939 527
rect 885 451 895 485
rect 929 451 939 485
rect 885 417 939 451
rect 885 383 895 417
rect 929 383 939 417
rect 885 367 939 383
rect 973 485 1039 493
rect 973 451 989 485
rect 1023 451 1039 485
rect 973 417 1039 451
rect 973 383 989 417
rect 1023 383 1039 417
rect 785 333 801 349
rect 647 315 801 333
rect 835 333 851 349
rect 973 349 1039 383
rect 1073 485 1127 527
rect 1073 451 1083 485
rect 1117 451 1127 485
rect 1073 417 1127 451
rect 1073 383 1083 417
rect 1117 383 1127 417
rect 1073 367 1127 383
rect 973 333 989 349
rect 835 315 989 333
rect 1023 333 1039 349
rect 1023 315 1083 333
rect 597 299 1083 315
rect 439 255 475 289
rect 83 249 217 255
rect 83 215 99 249
rect 133 215 167 249
rect 201 215 217 249
rect 271 249 405 255
rect 271 215 287 249
rect 321 215 355 249
rect 389 215 405 249
rect 439 249 969 255
rect 439 215 579 249
rect 613 215 647 249
rect 681 215 715 249
rect 749 215 783 249
rect 817 215 851 249
rect 885 215 919 249
rect 953 215 969 249
rect 439 181 475 215
rect 1003 181 1083 299
rect 29 163 83 181
rect 29 129 39 163
rect 73 129 83 163
rect 29 95 83 129
rect 29 61 39 95
rect 73 61 83 95
rect 29 17 83 61
rect 117 163 475 181
rect 117 129 133 163
rect 167 145 321 163
rect 167 129 183 145
rect 117 95 183 129
rect 305 129 321 145
rect 355 147 475 163
rect 509 165 563 181
rect 355 129 371 147
rect 117 61 133 95
rect 167 61 183 95
rect 117 51 183 61
rect 217 95 271 111
rect 217 61 227 95
rect 261 61 271 95
rect 217 17 271 61
rect 305 95 371 129
rect 509 131 529 165
rect 509 111 563 131
rect 305 61 321 95
rect 355 61 371 95
rect 305 51 371 61
rect 405 95 563 111
rect 439 93 563 95
rect 439 61 529 93
rect 405 59 529 61
rect 405 17 563 59
rect 597 169 1083 181
rect 597 135 613 169
rect 647 145 801 169
rect 647 135 657 145
rect 597 101 657 135
rect 791 135 801 145
rect 835 145 989 169
rect 835 135 845 145
rect 597 67 613 101
rect 647 67 657 101
rect 597 51 657 67
rect 691 101 757 111
rect 691 67 707 101
rect 741 67 757 101
rect 691 17 757 67
rect 791 101 845 135
rect 979 135 989 145
rect 1023 145 1083 169
rect 1023 135 1033 145
rect 791 67 801 101
rect 835 67 845 101
rect 791 51 845 67
rect 879 101 945 111
rect 879 67 895 101
rect 929 67 945 101
rect 879 17 945 67
rect 979 101 1033 135
rect 979 67 989 101
rect 1023 67 1033 101
rect 979 51 1033 67
rect 1067 101 1133 111
rect 1067 67 1083 101
rect 1117 67 1133 101
rect 1067 17 1133 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
flabel corelocali s 1041 221 1075 255 0 FreeSans 200 0 0 0 X
port 7 nsew
flabel corelocali s 121 221 155 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 305 221 339 255 0 FreeSans 200 0 0 0 B
port 2 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew
rlabel comment s 0 0 0 0 4 or2_6
<< properties >>
string FIXED_BBOX 0 0 1196 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 632966
string GDS_START 623536
<< end >>
