magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 940 430 994 547
rect 793 424 994 430
rect 1120 424 1186 547
rect 1310 424 1376 596
rect 1639 424 1705 596
rect 793 390 1705 424
rect 25 270 359 356
rect 505 270 743 356
rect 793 310 933 390
rect 1639 364 1705 390
rect 899 236 933 310
rect 967 270 1223 356
rect 1273 270 1558 356
rect 899 202 1619 236
rect 1381 184 1619 202
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 24 424 74 596
rect 114 458 180 649
rect 220 424 254 596
rect 294 458 360 649
rect 394 424 460 596
rect 494 581 1276 615
rect 494 458 560 581
rect 594 508 660 547
rect 728 542 794 581
rect 828 508 894 547
rect 594 474 894 508
rect 594 424 660 474
rect 1030 458 1080 581
rect 24 390 660 424
rect 1226 458 1276 581
rect 1410 458 1605 649
rect 394 364 460 390
rect 23 202 865 236
rect 23 184 461 202
rect 23 78 89 184
rect 123 17 189 150
rect 295 17 361 150
rect 395 78 461 184
rect 499 17 592 161
rect 629 78 695 202
rect 831 168 865 202
rect 729 17 795 168
rect 831 150 1155 168
rect 831 134 1361 150
rect 831 78 865 134
rect 1089 116 1361 134
rect 917 17 1053 100
rect 1089 78 1155 116
rect 1295 112 1361 116
rect 1467 112 1533 150
rect 1653 112 1705 234
rect 1191 17 1259 82
rect 1295 78 1705 112
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
<< metal1 >>
rect 0 683 1728 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 0 617 1728 649
rect 0 17 1728 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
rect 0 -49 1728 -17
<< labels >>
rlabel locali s 25 270 359 356 6 A1
port 1 nsew signal input
rlabel locali s 505 270 743 356 6 A2
port 2 nsew signal input
rlabel locali s 967 270 1223 356 6 A3
port 3 nsew signal input
rlabel locali s 1273 270 1558 356 6 B1
port 4 nsew signal input
rlabel locali s 1639 424 1705 596 6 Y
port 5 nsew signal output
rlabel locali s 1639 364 1705 390 6 Y
port 5 nsew signal output
rlabel locali s 1381 184 1619 202 6 Y
port 5 nsew signal output
rlabel locali s 1310 424 1376 596 6 Y
port 5 nsew signal output
rlabel locali s 1120 424 1186 547 6 Y
port 5 nsew signal output
rlabel locali s 940 430 994 547 6 Y
port 5 nsew signal output
rlabel locali s 899 236 933 310 6 Y
port 5 nsew signal output
rlabel locali s 899 202 1619 236 6 Y
port 5 nsew signal output
rlabel locali s 793 424 994 430 6 Y
port 5 nsew signal output
rlabel locali s 793 390 1705 424 6 Y
port 5 nsew signal output
rlabel locali s 793 310 933 390 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -49 1728 49 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1728 715 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1728 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 837174
string GDS_START 823526
<< end >>
