magic
tech sky130A
magscale 1 2
timestamp 1601050088
<< locali >>
rect 23 424 240 596
rect 374 424 440 596
rect 23 394 440 424
rect 638 424 704 596
rect 838 424 904 596
rect 1637 424 1703 547
rect 1837 424 1903 547
rect 638 394 1903 424
rect 23 390 1903 394
rect 374 360 704 390
rect 374 356 408 360
rect 25 270 270 356
rect 313 310 408 356
rect 793 326 839 356
rect 313 226 361 310
rect 442 260 839 326
rect 889 270 1223 356
rect 1257 270 1527 356
rect 1561 270 1898 356
rect 123 154 361 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 274 458 340 649
rect 474 428 604 649
rect 738 458 804 649
rect 950 492 1233 596
rect 1267 526 1317 649
rect 1357 492 1423 596
rect 1463 526 1497 649
rect 1537 581 1993 615
rect 1537 492 1603 581
rect 950 458 1603 492
rect 1737 458 1803 581
rect 1943 364 1993 581
rect 1009 226 1993 236
rect 23 120 89 226
rect 397 163 791 226
rect 837 202 1993 226
rect 837 170 1261 202
rect 837 163 903 170
rect 397 120 431 163
rect 1095 129 1161 136
rect 23 70 431 120
rect 467 70 1161 129
rect 1195 70 1261 170
rect 1295 17 1361 164
rect 1397 70 1431 202
rect 1467 17 1533 164
rect 1569 70 1619 202
rect 1653 17 1719 164
rect 1755 70 1805 202
rect 1841 17 1907 164
rect 1943 70 1993 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
rlabel locali s 1257 270 1527 356 6 A1
port 1 nsew signal input
rlabel locali s 1561 270 1898 356 6 A2
port 2 nsew signal input
rlabel locali s 889 270 1223 356 6 B1
port 3 nsew signal input
rlabel locali s 793 326 839 356 6 C1
port 4 nsew signal input
rlabel locali s 442 260 839 326 6 C1
port 4 nsew signal input
rlabel locali s 25 270 270 356 6 D1
port 5 nsew signal input
rlabel locali s 1837 424 1903 547 6 Y
port 6 nsew signal output
rlabel locali s 1637 424 1703 547 6 Y
port 6 nsew signal output
rlabel locali s 838 424 904 596 6 Y
port 6 nsew signal output
rlabel locali s 638 424 704 596 6 Y
port 6 nsew signal output
rlabel locali s 638 394 1903 424 6 Y
port 6 nsew signal output
rlabel locali s 374 424 440 596 6 Y
port 6 nsew signal output
rlabel locali s 374 360 704 390 6 Y
port 6 nsew signal output
rlabel locali s 374 356 408 360 6 Y
port 6 nsew signal output
rlabel locali s 313 310 408 356 6 Y
port 6 nsew signal output
rlabel locali s 313 226 361 310 6 Y
port 6 nsew signal output
rlabel locali s 123 154 361 226 6 Y
port 6 nsew signal output
rlabel locali s 23 424 240 596 6 Y
port 6 nsew signal output
rlabel locali s 23 394 440 424 6 Y
port 6 nsew signal output
rlabel locali s 23 390 1903 394 6 Y
port 6 nsew signal output
rlabel metal1 s 0 -49 2016 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 617 2016 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2016 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1752720
string GDS_START 1737376
<< end >>
