magic
tech sky130A
magscale 1 2
timestamp 1601050082
<< locali >>
rect 331 424 365 547
rect 331 390 619 424
rect 331 364 365 390
rect 107 294 173 360
rect 409 270 551 356
rect 585 236 619 390
rect 659 270 839 356
rect 889 270 1127 356
rect 488 202 1029 236
rect 488 192 554 202
rect 250 158 554 192
rect 250 66 316 158
rect 488 70 554 158
rect 688 70 754 202
rect 963 70 1029 202
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 23 260 73 596
rect 113 394 179 649
rect 225 581 455 615
rect 225 364 291 581
rect 405 492 455 581
rect 495 581 853 615
rect 495 526 561 581
rect 601 492 651 547
rect 405 458 651 492
rect 697 424 747 547
rect 787 458 853 581
rect 893 424 927 596
rect 967 458 1033 649
rect 1075 424 1125 596
rect 697 390 1125 424
rect 221 260 355 310
rect 23 226 355 260
rect 23 70 116 226
rect 150 17 216 192
rect 350 17 454 120
rect 588 17 654 168
rect 788 17 929 158
rect 1063 17 1129 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
rlabel locali s 889 270 1127 356 6 A
port 1 nsew signal input
rlabel locali s 659 270 839 356 6 B
port 2 nsew signal input
rlabel locali s 409 270 551 356 6 C
port 3 nsew signal input
rlabel locali s 107 294 173 360 6 D_N
port 4 nsew signal input
rlabel locali s 963 70 1029 202 6 Y
port 5 nsew signal output
rlabel locali s 688 70 754 202 6 Y
port 5 nsew signal output
rlabel locali s 585 236 619 390 6 Y
port 5 nsew signal output
rlabel locali s 488 202 1029 236 6 Y
port 5 nsew signal output
rlabel locali s 488 192 554 202 6 Y
port 5 nsew signal output
rlabel locali s 488 70 554 158 6 Y
port 5 nsew signal output
rlabel locali s 331 424 365 547 6 Y
port 5 nsew signal output
rlabel locali s 331 390 619 424 6 Y
port 5 nsew signal output
rlabel locali s 331 364 365 390 6 Y
port 5 nsew signal output
rlabel locali s 250 158 554 192 6 Y
port 5 nsew signal output
rlabel locali s 250 66 316 158 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -49 1152 49 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1152 715 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1159858
string GDS_START 1149638
<< end >>
