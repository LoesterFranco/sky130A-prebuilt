magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 2246 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 96 47 126 177
rect 190 47 220 177
rect 291 47 321 177
rect 547 47 577 177
rect 651 47 681 177
rect 755 47 785 177
rect 859 47 889 177
rect 963 47 993 177
rect 1067 47 1097 177
rect 1171 47 1201 177
rect 1275 47 1305 177
rect 1421 47 1451 177
rect 1515 47 1545 177
rect 1609 47 1639 177
rect 1703 47 1733 177
rect 1797 47 1827 177
rect 1891 47 1921 177
rect 1985 47 2015 177
rect 2089 47 2119 177
<< pmoshvt >>
rect 88 297 124 497
rect 182 297 218 497
rect 293 297 329 497
rect 491 309 527 497
rect 595 309 631 497
rect 699 309 735 497
rect 803 309 839 497
rect 907 309 943 497
rect 1011 309 1047 497
rect 1115 309 1151 497
rect 1219 309 1255 497
rect 1423 297 1459 497
rect 1517 297 1553 497
rect 1611 297 1647 497
rect 1705 297 1741 497
rect 1799 297 1835 497
rect 1893 297 1929 497
rect 1987 297 2023 497
rect 2081 297 2117 497
<< ndiff >>
rect 27 157 96 177
rect 27 123 39 157
rect 73 123 96 157
rect 27 89 96 123
rect 27 55 39 89
rect 73 55 96 89
rect 27 47 96 55
rect 126 106 190 177
rect 126 72 136 106
rect 170 72 190 106
rect 126 47 190 72
rect 220 89 291 177
rect 220 55 230 89
rect 264 55 291 89
rect 220 47 291 55
rect 321 129 383 177
rect 321 95 341 129
rect 375 95 383 129
rect 321 47 383 95
rect 485 129 547 177
rect 485 95 493 129
rect 527 95 547 129
rect 485 47 547 95
rect 577 89 651 177
rect 577 55 597 89
rect 631 55 651 89
rect 577 47 651 55
rect 681 129 755 177
rect 681 95 701 129
rect 735 95 755 129
rect 681 47 755 95
rect 785 89 859 177
rect 785 55 805 89
rect 839 55 859 89
rect 785 47 859 55
rect 889 129 963 177
rect 889 95 909 129
rect 943 95 963 129
rect 889 47 963 95
rect 993 89 1067 177
rect 993 55 1013 89
rect 1047 55 1067 89
rect 993 47 1067 55
rect 1097 129 1171 177
rect 1097 95 1117 129
rect 1151 95 1171 129
rect 1097 47 1171 95
rect 1201 89 1275 177
rect 1201 55 1221 89
rect 1255 55 1275 89
rect 1201 47 1275 55
rect 1305 129 1421 177
rect 1305 95 1352 129
rect 1386 95 1421 129
rect 1305 47 1421 95
rect 1451 169 1515 177
rect 1451 135 1471 169
rect 1505 135 1515 169
rect 1451 47 1515 135
rect 1545 89 1609 177
rect 1545 55 1565 89
rect 1599 55 1609 89
rect 1545 47 1609 55
rect 1639 169 1703 177
rect 1639 135 1659 169
rect 1693 135 1703 169
rect 1639 47 1703 135
rect 1733 89 1797 177
rect 1733 55 1753 89
rect 1787 55 1797 89
rect 1733 47 1797 55
rect 1827 169 1891 177
rect 1827 135 1847 169
rect 1881 135 1891 169
rect 1827 47 1891 135
rect 1921 89 1985 177
rect 1921 55 1941 89
rect 1975 55 1985 89
rect 1921 47 1985 55
rect 2015 169 2089 177
rect 2015 135 2035 169
rect 2069 135 2089 169
rect 2015 47 2089 135
rect 2119 89 2175 177
rect 2119 55 2129 89
rect 2163 55 2175 89
rect 2119 47 2175 55
<< pdiff >>
rect 27 489 88 497
rect 27 455 39 489
rect 73 455 88 489
rect 27 421 88 455
rect 27 387 39 421
rect 73 387 88 421
rect 27 297 88 387
rect 124 461 182 497
rect 124 427 136 461
rect 170 427 182 461
rect 124 297 182 427
rect 218 489 293 497
rect 218 455 230 489
rect 264 455 293 489
rect 218 421 293 455
rect 218 387 230 421
rect 264 387 293 421
rect 218 297 293 387
rect 329 479 383 497
rect 329 445 341 479
rect 375 445 383 479
rect 329 411 383 445
rect 329 377 341 411
rect 375 377 383 411
rect 329 343 383 377
rect 329 309 341 343
rect 375 309 383 343
rect 437 477 491 497
rect 437 443 445 477
rect 479 443 491 477
rect 437 309 491 443
rect 527 489 595 497
rect 527 455 539 489
rect 573 455 595 489
rect 527 309 595 455
rect 631 477 699 497
rect 631 443 643 477
rect 677 443 699 477
rect 631 309 699 443
rect 735 489 803 497
rect 735 455 747 489
rect 781 455 803 489
rect 735 309 803 455
rect 839 477 907 497
rect 839 443 851 477
rect 885 443 907 477
rect 839 309 907 443
rect 943 489 1011 497
rect 943 455 955 489
rect 989 455 1011 489
rect 943 309 1011 455
rect 1047 477 1115 497
rect 1047 443 1059 477
rect 1093 443 1115 477
rect 1047 309 1115 443
rect 1151 489 1219 497
rect 1151 455 1163 489
rect 1197 455 1219 489
rect 1151 309 1219 455
rect 1255 477 1423 497
rect 1255 443 1284 477
rect 1318 443 1362 477
rect 1396 443 1423 477
rect 1255 309 1423 443
rect 329 297 383 309
rect 1272 297 1423 309
rect 1459 345 1517 497
rect 1459 311 1471 345
rect 1505 311 1517 345
rect 1459 297 1517 311
rect 1553 489 1611 497
rect 1553 455 1565 489
rect 1599 455 1611 489
rect 1553 421 1611 455
rect 1553 387 1565 421
rect 1599 387 1611 421
rect 1553 297 1611 387
rect 1647 345 1705 497
rect 1647 311 1659 345
rect 1693 311 1705 345
rect 1647 297 1705 311
rect 1741 489 1799 497
rect 1741 455 1753 489
rect 1787 455 1799 489
rect 1741 421 1799 455
rect 1741 387 1753 421
rect 1787 387 1799 421
rect 1741 297 1799 387
rect 1835 345 1893 497
rect 1835 311 1847 345
rect 1881 311 1893 345
rect 1835 297 1893 311
rect 1929 489 1987 497
rect 1929 455 1941 489
rect 1975 455 1987 489
rect 1929 421 1987 455
rect 1929 387 1941 421
rect 1975 387 1987 421
rect 1929 297 1987 387
rect 2023 345 2081 497
rect 2023 311 2035 345
rect 2069 311 2081 345
rect 2023 297 2081 311
rect 2117 489 2175 497
rect 2117 455 2129 489
rect 2163 455 2175 489
rect 2117 421 2175 455
rect 2117 387 2129 421
rect 2163 387 2175 421
rect 2117 297 2175 387
<< ndiffc >>
rect 39 123 73 157
rect 39 55 73 89
rect 136 72 170 106
rect 230 55 264 89
rect 341 95 375 129
rect 493 95 527 129
rect 597 55 631 89
rect 701 95 735 129
rect 805 55 839 89
rect 909 95 943 129
rect 1013 55 1047 89
rect 1117 95 1151 129
rect 1221 55 1255 89
rect 1352 95 1386 129
rect 1471 135 1505 169
rect 1565 55 1599 89
rect 1659 135 1693 169
rect 1753 55 1787 89
rect 1847 135 1881 169
rect 1941 55 1975 89
rect 2035 135 2069 169
rect 2129 55 2163 89
<< pdiffc >>
rect 39 455 73 489
rect 39 387 73 421
rect 136 427 170 461
rect 230 455 264 489
rect 230 387 264 421
rect 341 445 375 479
rect 341 377 375 411
rect 341 309 375 343
rect 445 443 479 477
rect 539 455 573 489
rect 643 443 677 477
rect 747 455 781 489
rect 851 443 885 477
rect 955 455 989 489
rect 1059 443 1093 477
rect 1163 455 1197 489
rect 1284 443 1318 477
rect 1362 443 1396 477
rect 1471 311 1505 345
rect 1565 455 1599 489
rect 1565 387 1599 421
rect 1659 311 1693 345
rect 1753 455 1787 489
rect 1753 387 1787 421
rect 1847 311 1881 345
rect 1941 455 1975 489
rect 1941 387 1975 421
rect 2035 311 2069 345
rect 2129 455 2163 489
rect 2129 387 2163 421
<< poly >>
rect 88 497 124 523
rect 182 497 218 523
rect 293 497 329 523
rect 491 497 527 523
rect 595 497 631 523
rect 699 497 735 523
rect 803 497 839 523
rect 907 497 943 523
rect 1011 497 1047 523
rect 1115 497 1151 523
rect 1219 497 1255 523
rect 1423 497 1459 523
rect 1517 497 1553 523
rect 1611 497 1647 523
rect 1705 497 1741 523
rect 1799 497 1835 523
rect 1893 497 1929 523
rect 1987 497 2023 523
rect 2081 497 2117 523
rect 88 282 124 297
rect 182 282 218 297
rect 293 282 329 297
rect 491 294 527 309
rect 595 294 631 309
rect 699 294 735 309
rect 803 294 839 309
rect 907 294 943 309
rect 1011 294 1047 309
rect 1115 294 1151 309
rect 1219 294 1255 309
rect 86 265 126 282
rect 32 259 126 265
rect 180 259 220 282
rect 291 265 331 282
rect 414 265 1257 294
rect 1423 282 1459 297
rect 1517 282 1553 297
rect 1611 282 1647 297
rect 1705 282 1741 297
rect 1799 282 1835 297
rect 1893 282 1929 297
rect 1987 282 2023 297
rect 2081 282 2117 297
rect 32 249 220 259
rect 32 215 42 249
rect 76 215 220 249
rect 32 205 220 215
rect 32 199 126 205
rect 96 177 126 199
rect 190 177 220 205
rect 262 264 1257 265
rect 262 249 444 264
rect 1421 259 1461 282
rect 1515 259 1555 282
rect 1609 259 1649 282
rect 1703 259 1743 282
rect 1797 259 1837 282
rect 1891 259 1931 282
rect 1985 259 2025 282
rect 2079 259 2119 282
rect 262 215 272 249
rect 306 215 444 249
rect 1299 249 1375 259
rect 1299 222 1325 249
rect 262 199 444 215
rect 547 215 1325 222
rect 1359 215 1375 249
rect 291 177 321 199
rect 547 192 1375 215
rect 1421 249 2119 259
rect 1421 215 1445 249
rect 1479 215 1523 249
rect 1557 215 1601 249
rect 1635 215 1679 249
rect 1713 215 1757 249
rect 1791 215 1825 249
rect 1859 215 1903 249
rect 1937 215 1981 249
rect 2015 215 2119 249
rect 1421 205 2119 215
rect 547 177 577 192
rect 651 177 681 192
rect 755 177 785 192
rect 859 177 889 192
rect 963 177 993 192
rect 1067 177 1097 192
rect 1171 177 1201 192
rect 1275 177 1305 192
rect 1421 177 1451 205
rect 1515 177 1545 205
rect 1609 177 1639 205
rect 1703 177 1733 205
rect 1797 177 1827 205
rect 1891 177 1921 205
rect 1985 177 2015 205
rect 2089 177 2119 205
rect 96 21 126 47
rect 190 21 220 47
rect 291 21 321 47
rect 547 21 577 47
rect 651 21 681 47
rect 755 21 785 47
rect 859 21 889 47
rect 963 21 993 47
rect 1067 21 1097 47
rect 1171 21 1201 47
rect 1275 21 1305 47
rect 1421 21 1451 47
rect 1515 21 1545 47
rect 1609 21 1639 47
rect 1703 21 1733 47
rect 1797 21 1827 47
rect 1891 21 1921 47
rect 1985 21 2015 47
rect 2089 21 2119 47
<< polycont >>
rect 42 215 76 249
rect 272 215 306 249
rect 1325 215 1359 249
rect 1445 215 1479 249
rect 1523 215 1557 249
rect 1601 215 1635 249
rect 1679 215 1713 249
rect 1757 215 1791 249
rect 1825 215 1859 249
rect 1903 215 1937 249
rect 1981 215 2015 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 17 489 89 527
rect 17 455 39 489
rect 73 455 89 489
rect 17 421 89 455
rect 17 387 39 421
rect 73 387 89 421
rect 17 357 89 387
rect 133 461 170 493
rect 133 427 136 461
rect 133 323 170 427
rect 204 489 281 527
rect 204 455 230 489
rect 264 455 281 489
rect 204 421 281 455
rect 204 387 230 421
rect 264 387 281 421
rect 204 373 281 387
rect 315 479 395 493
rect 315 445 341 479
rect 375 445 395 479
rect 315 411 395 445
rect 315 377 341 411
rect 375 377 395 411
rect 429 477 479 493
rect 429 443 445 477
rect 513 489 599 527
rect 513 455 539 489
rect 573 455 599 489
rect 513 447 599 455
rect 643 477 677 493
rect 429 413 479 443
rect 721 489 807 527
rect 721 455 747 489
rect 781 455 807 489
rect 721 447 807 455
rect 851 477 885 493
rect 643 413 677 443
rect 929 489 1015 527
rect 929 455 955 489
rect 989 455 1015 489
rect 929 447 1015 455
rect 1059 477 1093 493
rect 851 413 885 443
rect 1137 489 1223 527
rect 1137 455 1163 489
rect 1197 455 1223 489
rect 1137 447 1223 455
rect 1267 489 2185 493
rect 1267 477 1565 489
rect 1059 413 1093 443
rect 1267 443 1284 477
rect 1318 443 1362 477
rect 1396 455 1565 477
rect 1599 455 1753 489
rect 1787 455 1941 489
rect 1975 455 2129 489
rect 2163 455 2185 489
rect 1396 443 2185 455
rect 1267 421 2185 443
rect 1267 413 1565 421
rect 429 387 1565 413
rect 1599 387 1753 421
rect 1787 387 1941 421
rect 1975 387 2129 421
rect 2163 387 2185 421
rect 429 379 2185 387
rect 315 343 395 377
rect 17 249 86 323
rect 17 215 42 249
rect 76 215 86 249
rect 17 199 86 215
rect 130 246 170 323
rect 130 212 131 246
rect 165 212 170 246
rect 17 157 89 165
rect 17 123 39 157
rect 73 123 89 157
rect 17 89 89 123
rect 17 55 39 89
rect 73 55 89 89
rect 130 106 170 212
rect 204 265 281 339
rect 315 309 341 343
rect 375 309 395 343
rect 315 299 395 309
rect 204 249 306 265
rect 204 215 272 249
rect 204 199 306 215
rect 350 255 395 299
rect 429 311 1471 345
rect 1505 311 1659 345
rect 1693 311 1847 345
rect 1881 311 2035 345
rect 2069 311 2185 345
rect 429 289 2185 311
rect 350 249 1375 255
rect 350 215 1325 249
rect 1359 215 1375 249
rect 350 205 1375 215
rect 1425 249 2091 255
rect 1425 215 1445 249
rect 1479 215 1523 249
rect 1557 246 1601 249
rect 1560 215 1601 246
rect 1635 215 1679 249
rect 1713 215 1757 249
rect 1791 215 1825 249
rect 1859 215 1903 249
rect 1937 215 1981 249
rect 2015 215 2091 249
rect 1425 212 1526 215
rect 1560 212 2091 215
rect 1425 205 2091 212
rect 204 124 281 199
rect 350 165 427 205
rect 2135 171 2185 289
rect 315 129 427 165
rect 130 72 136 106
rect 315 95 341 129
rect 375 95 427 129
rect 130 56 170 72
rect 17 17 89 55
rect 204 55 230 89
rect 264 55 281 89
rect 204 17 281 55
rect 315 51 427 95
rect 461 131 1411 171
rect 461 129 537 131
rect 461 95 493 129
rect 527 95 537 129
rect 701 129 745 131
rect 461 51 537 95
rect 571 89 657 97
rect 571 55 597 89
rect 631 55 657 89
rect 735 95 745 129
rect 909 129 953 131
rect 701 55 745 95
rect 779 89 865 97
rect 779 55 805 89
rect 839 55 865 89
rect 571 17 657 55
rect 779 17 865 55
rect 943 95 953 129
rect 1117 129 1161 131
rect 909 51 953 95
rect 987 89 1073 97
rect 987 55 1013 89
rect 1047 55 1073 89
rect 1151 95 1161 129
rect 1325 129 1411 131
rect 1117 55 1161 95
rect 1195 89 1281 97
rect 1195 55 1221 89
rect 1255 55 1281 89
rect 987 17 1073 55
rect 1195 17 1281 55
rect 1325 95 1352 129
rect 1386 95 1411 129
rect 1445 169 2185 171
rect 1445 135 1471 169
rect 1505 135 1659 169
rect 1693 135 1847 169
rect 1881 135 2035 169
rect 2069 135 2185 169
rect 1445 123 2185 135
rect 1325 89 1411 95
rect 1325 55 1565 89
rect 1599 55 1753 89
rect 1787 55 1941 89
rect 1975 55 2129 89
rect 2163 55 2185 89
rect 1325 51 2185 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 131 212 165 246
rect 1526 215 1557 246
rect 1557 215 1560 246
rect 1526 212 1560 215
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
<< metal1 >>
rect 0 561 2208 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 0 496 2208 527
rect 109 246 1572 252
rect 109 212 131 246
rect 165 224 1526 246
rect 165 212 177 224
rect 109 206 177 212
rect 1504 212 1526 224
rect 1560 212 1572 246
rect 1504 206 1572 212
rect 0 17 2208 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
rect 0 -48 2208 -17
<< labels >>
flabel corelocali s 29 221 63 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 29 289 63 323 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 2138 153 2172 187 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 2138 221 2172 255 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 857 289 891 323 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 969 289 1003 323 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 1080 289 1114 323 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 1211 289 1245 323 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 529 289 563 323 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 641 289 675 323 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 750 289 784 323 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 230 170 230 170 0 FreeSans 200 0 0 0 TE_B
port 2 nsew
flabel corelocali s 1323 289 1357 323 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 1414 289 1448 323 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 230 306 230 306 0 FreeSans 200 0 0 0 TE_B
port 2 nsew
flabel corelocali s 2138 289 2172 323 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 2036 289 2070 323 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 1620 289 1654 323 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 1934 289 1968 323 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 1824 289 1858 323 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 1717 289 1751 323 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew
rlabel comment s 0 0 0 0 4 ebufn_8
<< properties >>
string FIXED_BBOX 0 0 2208 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2005310
string GDS_START 1990694
<< end >>
