magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 20 199 66 323
rect 117 199 205 323
rect 471 333 531 493
rect 659 333 735 493
rect 847 333 923 493
rect 1035 333 1111 493
rect 1333 333 1409 493
rect 1521 333 1597 493
rect 1709 333 1785 493
rect 1897 333 1973 493
rect 471 289 1973 333
rect 733 181 803 289
rect 1209 215 1597 255
rect 1679 215 2068 255
rect 471 131 803 181
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 17 396 74 488
rect 108 439 163 527
rect 197 430 369 493
rect 17 357 301 396
rect 239 161 301 357
rect 17 127 301 161
rect 335 261 369 430
rect 403 299 437 527
rect 565 367 625 527
rect 779 367 813 527
rect 967 367 1001 527
rect 1165 367 1293 527
rect 1453 367 1487 527
rect 1641 367 1675 527
rect 1829 367 1863 527
rect 2017 289 2072 527
rect 335 215 405 261
rect 471 215 640 249
rect 17 51 69 127
rect 335 93 369 215
rect 837 215 1111 255
rect 103 17 179 93
rect 223 51 369 93
rect 403 97 437 181
rect 847 131 1602 181
rect 1641 131 2057 165
rect 1641 97 1675 131
rect 403 51 1205 97
rect 1253 51 1675 97
rect 1719 17 1785 97
rect 1907 17 1973 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
<< metal1 >>
rect 0 561 2116 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 0 496 2116 527
rect 0 17 2116 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
rect 0 -48 2116 -17
<< obsm1 >>
rect 347 252 405 261
rect 847 252 915 261
rect 347 224 915 252
rect 347 215 405 224
rect 847 215 915 224
<< labels >>
rlabel locali s 20 199 66 323 6 A_N
port 1 nsew signal input
rlabel locali s 117 199 205 323 6 B_N
port 2 nsew signal input
rlabel locali s 1209 215 1597 255 6 C
port 3 nsew signal input
rlabel locali s 1679 215 2068 255 6 D
port 4 nsew signal input
rlabel locali s 1897 333 1973 493 6 Y
port 5 nsew signal output
rlabel locali s 1709 333 1785 493 6 Y
port 5 nsew signal output
rlabel locali s 1521 333 1597 493 6 Y
port 5 nsew signal output
rlabel locali s 1333 333 1409 493 6 Y
port 5 nsew signal output
rlabel locali s 1035 333 1111 493 6 Y
port 5 nsew signal output
rlabel locali s 847 333 923 493 6 Y
port 5 nsew signal output
rlabel locali s 733 181 803 289 6 Y
port 5 nsew signal output
rlabel locali s 659 333 735 493 6 Y
port 5 nsew signal output
rlabel locali s 471 333 531 493 6 Y
port 5 nsew signal output
rlabel locali s 471 289 1973 333 6 Y
port 5 nsew signal output
rlabel locali s 471 131 803 181 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -48 2116 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 2116 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2116 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2380958
string GDS_START 2365442
<< end >>
