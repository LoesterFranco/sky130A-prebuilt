magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 736 561
rect 103 439 169 527
rect 311 445 445 527
rect 562 445 628 527
rect 17 199 90 335
rect 103 17 169 93
rect 304 84 360 339
rect 405 84 459 339
rect 497 133 565 339
rect 667 299 719 493
rect 685 161 719 299
rect 551 17 617 93
rect 651 68 719 161
rect 651 59 718 68
rect 0 -17 736 17
<< obsli1 >>
rect 34 403 69 493
rect 230 409 264 493
rect 488 409 522 493
rect 34 369 160 403
rect 126 265 160 369
rect 230 375 633 409
rect 126 199 196 265
rect 126 165 160 199
rect 34 131 160 165
rect 34 51 69 131
rect 230 117 264 375
rect 218 51 264 117
rect 599 265 633 375
rect 599 199 651 265
<< metal1 >>
rect 0 496 736 592
rect 0 -48 736 48
<< labels >>
rlabel locali s 17 199 90 335 6 A_N
port 1 nsew signal input
rlabel locali s 304 84 360 339 6 B
port 2 nsew signal input
rlabel locali s 405 84 459 339 6 C
port 3 nsew signal input
rlabel locali s 497 133 565 339 6 D
port 4 nsew signal input
rlabel locali s 685 161 719 299 6 X
port 5 nsew signal output
rlabel locali s 667 299 719 493 6 X
port 5 nsew signal output
rlabel locali s 651 68 719 161 6 X
port 5 nsew signal output
rlabel locali s 651 59 718 68 6 X
port 5 nsew signal output
rlabel locali s 551 17 617 93 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 103 17 169 93 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 736 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 736 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 562 445 628 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 311 445 445 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 103 439 169 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 736 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 736 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3842942
string GDS_START 3835388
<< end >>
