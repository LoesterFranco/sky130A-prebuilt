magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 108 364 359 430
rect 325 324 359 364
rect 325 272 547 324
rect 589 288 655 430
rect 313 162 418 238
rect 781 236 847 310
rect 2406 217 2472 596
rect 2406 183 2493 217
rect 2427 70 2493 183
rect 2811 70 2865 596
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 2976 683
rect 23 498 89 596
rect 123 546 280 649
rect 388 532 589 582
rect 623 532 689 649
rect 555 498 589 532
rect 723 504 799 596
rect 941 538 1007 649
rect 1142 504 1197 545
rect 723 498 1197 504
rect 23 464 521 498
rect 555 470 1197 498
rect 555 464 799 470
rect 1142 466 1197 470
rect 1232 502 1332 545
rect 1414 536 1464 649
rect 1510 502 1583 545
rect 1232 468 1583 502
rect 23 316 57 464
rect 455 366 521 464
rect 23 250 279 316
rect 23 75 73 250
rect 109 17 175 167
rect 219 85 269 167
rect 689 235 723 464
rect 757 424 833 430
rect 757 390 799 424
rect 757 364 833 390
rect 867 398 917 436
rect 1163 434 1197 466
rect 867 364 997 398
rect 1031 366 1129 432
rect 1163 400 1298 434
rect 963 332 997 364
rect 963 300 1061 332
rect 881 266 1061 300
rect 1095 300 1230 366
rect 452 201 723 235
rect 881 202 915 266
rect 1095 232 1129 300
rect 1264 258 1298 400
rect 452 119 522 201
rect 620 85 686 167
rect 219 51 686 85
rect 728 17 794 167
rect 848 70 915 202
rect 950 17 984 226
rect 1020 198 1129 232
rect 1164 224 1298 258
rect 1020 96 1086 198
rect 1164 164 1198 224
rect 1332 190 1366 468
rect 1476 464 1583 468
rect 1132 130 1198 164
rect 1232 130 1366 190
rect 1400 218 1442 355
rect 1476 315 1510 464
rect 1544 424 1604 430
rect 1544 390 1567 424
rect 1601 390 1604 424
rect 1544 359 1604 390
rect 1638 349 1688 649
rect 1728 349 1786 551
rect 1820 473 2019 539
rect 2053 532 2172 649
rect 2213 498 2279 559
rect 1476 252 1718 315
rect 1752 218 1786 349
rect 1862 373 1951 439
rect 1862 247 1928 373
rect 1400 184 1786 218
rect 1400 116 1665 150
rect 1699 119 1786 184
rect 1820 181 1928 247
rect 1985 262 2019 473
rect 2053 464 2279 498
rect 2053 330 2109 464
rect 2143 424 2279 430
rect 2177 390 2279 424
rect 2143 364 2279 390
rect 2320 364 2370 649
rect 2053 296 2372 330
rect 1985 209 2304 262
rect 1400 96 1434 116
rect 1020 62 1434 96
rect 1631 85 1665 116
rect 1820 85 1854 181
rect 1985 147 2019 209
rect 2338 175 2372 296
rect 2508 384 2566 649
rect 2613 326 2665 596
rect 2709 364 2775 649
rect 2613 260 2777 326
rect 1490 17 1597 82
rect 1631 51 1854 85
rect 1888 81 2019 147
rect 2067 17 2133 162
rect 2225 141 2372 175
rect 2225 70 2291 141
rect 2329 17 2379 107
rect 2527 17 2579 210
rect 2613 70 2665 260
rect 2734 17 2768 226
rect 2899 364 2955 649
rect 2899 17 2956 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 2976 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 799 390 833 424
rect 1567 390 1601 424
rect 2143 390 2177 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
<< metal1 >>
rect 0 683 2976 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 2976 683
rect 0 617 2976 649
rect 787 424 845 430
rect 787 390 799 424
rect 833 421 845 424
rect 1555 424 1613 430
rect 1555 421 1567 424
rect 833 393 1567 421
rect 833 390 845 393
rect 787 384 845 390
rect 1555 390 1567 393
rect 1601 421 1613 424
rect 2131 424 2189 430
rect 2131 421 2143 424
rect 1601 393 2143 421
rect 1601 390 1613 393
rect 1555 384 1613 390
rect 2131 390 2143 393
rect 2177 390 2189 424
rect 2131 384 2189 390
rect 0 17 2976 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 2976 17
rect 0 -49 2976 -17
<< labels >>
rlabel locali s 313 162 418 238 6 D
port 1 nsew signal input
rlabel locali s 2811 70 2865 596 6 Q
port 2 nsew signal output
rlabel locali s 2427 70 2493 183 6 Q_N
port 3 nsew signal output
rlabel locali s 2406 217 2472 596 6 Q_N
port 3 nsew signal output
rlabel locali s 2406 183 2493 217 6 Q_N
port 3 nsew signal output
rlabel metal1 s 2131 421 2189 430 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 2131 384 2189 393 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 1555 421 1613 430 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 1555 384 1613 393 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 787 421 845 430 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 787 393 2189 421 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 787 384 845 393 6 RESET_B
port 4 nsew signal input
rlabel locali s 589 288 655 430 6 SCD
port 5 nsew signal input
rlabel locali s 325 324 359 364 6 SCE
port 6 nsew signal input
rlabel locali s 325 272 547 324 6 SCE
port 6 nsew signal input
rlabel locali s 108 364 359 430 6 SCE
port 6 nsew signal input
rlabel locali s 781 236 847 310 6 CLK
port 7 nsew clock input
rlabel metal1 s 0 -49 2976 49 8 VGND
port 8 nsew ground bidirectional
rlabel metal1 s 0 617 2976 715 6 VPWR
port 9 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2976 666
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 21874
string GDS_START 132
<< end >>
