magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 219 393 279 425
rect 539 393 622 493
rect 219 357 622 393
rect 24 289 459 323
rect 24 211 90 289
rect 134 215 314 255
rect 350 215 459 289
rect 539 119 622 357
rect 656 153 714 280
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 21 357 87 527
rect 131 459 373 493
rect 131 357 175 459
rect 335 427 373 459
rect 412 435 488 527
rect 21 143 493 177
rect 21 51 87 143
rect 133 17 167 109
rect 203 51 279 143
rect 335 17 369 109
rect 427 85 493 143
rect 656 314 706 527
rect 656 85 706 119
rect 427 51 706 85
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel locali s 350 215 459 289 6 A1
port 1 nsew signal input
rlabel locali s 24 289 459 323 6 A1
port 1 nsew signal input
rlabel locali s 24 211 90 289 6 A1
port 1 nsew signal input
rlabel locali s 134 215 314 255 6 A2
port 2 nsew signal input
rlabel locali s 656 153 714 280 6 B1
port 3 nsew signal input
rlabel locali s 539 393 622 493 6 Y
port 4 nsew signal output
rlabel locali s 539 119 622 357 6 Y
port 4 nsew signal output
rlabel locali s 219 393 279 425 6 Y
port 4 nsew signal output
rlabel locali s 219 357 622 393 6 Y
port 4 nsew signal output
rlabel metal1 s 0 -48 736 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 736 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1009458
string GDS_START 1002726
<< end >>
