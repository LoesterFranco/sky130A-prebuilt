magic
tech sky130A
magscale 1 2
timestamp 1599588232
<< locali >>
rect 313 258 409 356
rect 511 271 579 430
rect 545 153 579 271
rect 688 326 754 392
rect 713 153 747 326
rect 881 153 919 321
rect 1175 218 1241 237
rect 1053 184 1241 218
rect 1053 153 1087 184
rect 545 119 1087 153
rect 2290 290 2375 356
rect 2517 310 2584 440
rect 2714 364 2775 596
rect 2517 70 2567 310
rect 2741 301 2775 364
rect 2741 226 2855 301
rect 2703 160 2855 226
rect 2703 71 2757 160
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2880 683
rect 21 432 72 649
rect 111 398 177 596
rect 67 364 177 398
rect 67 294 130 364
rect 218 326 268 596
rect 308 390 374 649
rect 411 578 1211 612
rect 411 403 477 578
rect 511 510 1111 544
rect 511 478 690 510
rect 25 276 130 294
rect 25 242 31 276
rect 65 242 130 276
rect 164 260 279 326
rect 25 236 130 242
rect 96 226 130 236
rect 96 192 193 226
rect 34 17 107 158
rect 141 70 193 192
rect 245 224 279 260
rect 443 237 477 403
rect 245 101 341 224
rect 443 203 511 237
rect 375 17 425 169
rect 461 85 511 203
rect 613 237 647 478
rect 724 426 822 476
rect 613 187 679 237
rect 788 282 822 426
rect 856 420 1043 470
rect 1077 454 1111 510
rect 1145 488 1211 578
rect 1253 516 1319 649
rect 1443 581 1915 615
rect 1443 482 1477 581
rect 1245 454 1477 482
rect 1077 448 1477 454
rect 1077 420 1279 448
rect 788 276 847 282
rect 788 242 799 276
rect 833 242 847 276
rect 788 237 847 242
rect 781 187 847 237
rect 953 286 987 420
rect 1343 386 1409 414
rect 1021 352 1409 386
rect 1021 320 1073 352
rect 1107 286 1309 305
rect 953 271 1309 286
rect 953 252 1141 271
rect 953 187 1019 252
rect 1275 204 1309 271
rect 1343 272 1409 352
rect 1443 392 1477 448
rect 1511 426 1662 547
rect 1443 326 1501 392
rect 1343 238 1501 272
rect 1275 170 1401 204
rect 1121 85 1187 150
rect 461 51 1187 85
rect 1267 17 1333 136
rect 1367 85 1401 170
rect 1435 126 1501 238
rect 1535 255 1594 389
rect 1535 85 1569 255
rect 1628 208 1662 426
rect 1696 245 1747 581
rect 1781 426 1847 547
rect 1781 211 1815 426
rect 1881 392 1915 581
rect 1628 202 1711 208
rect 1628 168 1663 202
rect 1697 168 1711 202
rect 1628 128 1711 168
rect 1367 51 1569 85
rect 1603 78 1711 128
rect 1749 85 1815 211
rect 1849 326 1915 392
rect 1949 554 2015 596
rect 2203 588 2279 649
rect 1949 520 2394 554
rect 2428 542 2494 649
rect 2608 542 2674 649
rect 1949 420 2015 520
rect 2360 508 2394 520
rect 2062 426 2162 486
rect 2360 474 2680 508
rect 1849 153 1883 326
rect 1949 237 1983 420
rect 1917 187 1983 237
rect 2017 271 2094 337
rect 2017 153 2051 271
rect 2128 237 2162 426
rect 1849 119 2051 153
rect 2085 203 2162 237
rect 2196 390 2386 440
rect 2196 211 2248 390
rect 2646 326 2680 474
rect 2809 364 2859 649
rect 2085 119 2119 203
rect 2196 169 2373 211
rect 2153 135 2373 169
rect 2417 202 2483 310
rect 2417 168 2431 202
rect 2465 168 2483 202
rect 2417 162 2483 168
rect 2153 85 2187 135
rect 1749 51 2187 85
rect 2221 17 2271 101
rect 2307 75 2373 135
rect 2415 17 2481 128
rect 2646 260 2707 326
rect 2603 17 2669 226
rect 2791 17 2857 126
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2880 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 31 242 65 276
rect 799 242 833 276
rect 1663 168 1697 202
rect 2431 168 2465 202
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
<< metal1 >>
rect 0 683 2880 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2880 683
rect 0 617 2880 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 2880 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2880 17
rect 0 -49 2880 -17
<< obsm1 >>
rect 19 276 77 282
rect 19 242 31 276
rect 65 273 77 276
rect 787 276 845 282
rect 787 273 799 276
rect 65 245 799 273
rect 65 242 77 245
rect 19 236 77 242
rect 787 242 799 245
rect 833 242 845 276
rect 787 236 845 242
rect 1651 202 1709 208
rect 1651 168 1663 202
rect 1697 199 1709 202
rect 2419 202 2477 208
rect 2419 199 2431 202
rect 1697 171 2431 199
rect 1697 168 1709 171
rect 1651 162 1709 168
rect 2419 168 2431 171
rect 2465 168 2477 202
rect 2419 162 2477 168
<< labels >>
rlabel locali s 313 258 409 356 6 A
port 1 nsew signal input
rlabel locali s 1175 218 1241 237 6 B
port 2 nsew signal input
rlabel locali s 1053 184 1241 218 6 B
port 2 nsew signal input
rlabel locali s 1053 153 1087 184 6 B
port 2 nsew signal input
rlabel locali s 881 153 919 321 6 B
port 2 nsew signal input
rlabel locali s 713 153 747 326 6 B
port 2 nsew signal input
rlabel locali s 688 326 754 392 6 B
port 2 nsew signal input
rlabel locali s 545 153 579 271 6 B
port 2 nsew signal input
rlabel locali s 545 119 1087 153 6 B
port 2 nsew signal input
rlabel locali s 511 271 579 430 6 B
port 2 nsew signal input
rlabel locali s 2290 290 2375 356 6 CI
port 3 nsew signal input
rlabel locali s 2517 310 2584 440 6 COUT
port 4 nsew signal output
rlabel locali s 2517 70 2567 310 6 COUT
port 4 nsew signal output
rlabel locali s 2741 301 2775 364 6 SUM
port 5 nsew signal output
rlabel locali s 2741 226 2855 301 6 SUM
port 5 nsew signal output
rlabel locali s 2714 364 2775 596 6 SUM
port 5 nsew signal output
rlabel locali s 2703 160 2855 226 6 SUM
port 5 nsew signal output
rlabel locali s 2703 71 2757 160 6 SUM
port 5 nsew signal output
rlabel metal1 s 0 -49 2880 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 7 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 617 2880 715 6 VPWR
port 9 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2880 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 2552342
string GDS_START 2532674
<< end >>
