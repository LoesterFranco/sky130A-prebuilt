magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 90 47 120 131
rect 185 47 215 131
rect 289 47 319 131
<< pmoshvt >>
rect 82 297 118 497
rect 187 297 223 497
rect 281 297 317 497
<< ndiff >>
rect 27 101 90 131
rect 27 67 35 101
rect 69 67 90 101
rect 27 47 90 67
rect 120 97 185 131
rect 120 63 131 97
rect 165 63 185 97
rect 120 47 185 63
rect 215 101 289 131
rect 215 67 235 101
rect 269 67 289 101
rect 215 47 289 67
rect 319 97 371 131
rect 319 63 329 97
rect 363 63 371 97
rect 319 47 371 63
<< pdiff >>
rect 27 471 82 497
rect 27 437 35 471
rect 69 437 82 471
rect 27 366 82 437
rect 27 332 35 366
rect 69 332 82 366
rect 27 297 82 332
rect 118 473 187 497
rect 118 439 131 473
rect 165 439 187 473
rect 118 405 187 439
rect 118 371 131 405
rect 165 371 187 405
rect 118 297 187 371
rect 223 471 281 497
rect 223 437 235 471
rect 269 437 281 471
rect 223 297 281 437
rect 317 476 371 497
rect 317 442 329 476
rect 363 442 371 476
rect 317 297 371 442
<< ndiffc >>
rect 35 67 69 101
rect 131 63 165 97
rect 235 67 269 101
rect 329 63 363 97
<< pdiffc >>
rect 35 437 69 471
rect 35 332 69 366
rect 131 439 165 473
rect 131 371 165 405
rect 235 437 269 471
rect 329 442 363 476
<< poly >>
rect 82 497 118 523
rect 187 497 223 523
rect 281 497 317 523
rect 82 282 118 297
rect 187 282 223 297
rect 281 282 317 297
rect 80 279 120 282
rect 185 279 225 282
rect 279 279 319 282
rect 69 249 143 279
rect 69 215 89 249
rect 123 215 143 249
rect 69 196 143 215
rect 185 249 319 279
rect 185 215 203 249
rect 237 215 319 249
rect 69 195 120 196
rect 90 131 120 195
rect 185 149 319 215
rect 185 131 215 149
rect 289 131 319 149
rect 90 21 120 47
rect 185 21 215 47
rect 289 21 319 47
<< polycont >>
rect 89 215 123 249
rect 203 215 237 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 17 471 71 487
rect 17 437 35 471
rect 69 437 71 471
rect 17 366 71 437
rect 105 473 181 527
rect 105 439 131 473
rect 165 439 181 473
rect 105 405 181 439
rect 105 371 131 405
rect 165 371 181 405
rect 232 471 269 487
rect 232 437 235 471
rect 303 476 380 527
rect 303 442 329 476
rect 363 442 380 476
rect 232 406 269 437
rect 232 371 375 406
rect 17 332 35 366
rect 69 333 71 366
rect 69 332 263 333
rect 17 299 263 332
rect 17 117 51 299
rect 85 249 167 265
rect 85 215 89 249
rect 123 215 167 249
rect 85 149 167 215
rect 203 249 263 299
rect 237 215 263 249
rect 203 199 263 215
rect 297 165 375 371
rect 228 131 375 165
rect 17 101 69 117
rect 17 67 35 101
rect 17 51 69 67
rect 121 97 176 113
rect 121 63 131 97
rect 165 63 176 97
rect 121 17 176 63
rect 228 101 269 131
rect 228 67 235 101
rect 228 51 269 67
rect 303 63 329 97
rect 363 63 380 97
rect 303 17 380 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew
flabel corelocali s 131 153 165 187 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 131 221 165 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 322 238 322 238 0 FreeSans 200 0 0 0 X
port 6 nsew
flabel corelocali s 322 170 322 170 0 FreeSans 200 0 0 0 X
port 6 nsew
flabel corelocali s 322 306 322 306 0 FreeSans 200 0 0 0 X
port 6 nsew
flabel corelocali s 322 374 322 374 0 FreeSans 200 0 0 0 X
port 6 nsew
rlabel comment s 0 0 0 0 4 clkbuf_2
<< properties >>
string FIXED_BBOX 0 0 460 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1765424
string GDS_START 1760910
<< end >>
