magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1196 561
rect 225 325 291 425
rect 29 291 291 325
rect 393 383 459 527
rect 561 383 627 527
rect 751 383 885 527
rect 1001 383 1067 527
rect 29 163 63 291
rect 109 215 311 256
rect 357 215 491 259
rect 533 215 673 257
rect 709 215 915 259
rect 951 215 1179 259
rect 29 129 459 163
rect 37 17 103 93
rect 137 51 171 129
rect 205 17 275 93
rect 1001 17 1067 93
rect 0 -17 1196 17
<< obsli1 >>
rect 157 459 359 493
rect 157 359 191 459
rect 325 341 359 459
rect 493 341 527 493
rect 665 341 699 493
rect 933 341 967 493
rect 1101 341 1135 493
rect 325 307 1152 341
rect 493 129 711 163
rect 749 129 1135 163
rect 493 93 527 129
rect 309 59 527 93
rect 561 59 899 93
rect 1101 51 1135 129
<< metal1 >>
rect 0 496 1196 592
rect 0 -48 1196 48
<< labels >>
rlabel locali s 357 215 491 259 6 A1
port 1 nsew signal input
rlabel locali s 533 215 673 257 6 A2
port 2 nsew signal input
rlabel locali s 709 215 915 259 6 A3
port 3 nsew signal input
rlabel locali s 951 215 1179 259 6 A4
port 4 nsew signal input
rlabel locali s 109 215 311 256 6 B1
port 5 nsew signal input
rlabel locali s 225 325 291 425 6 Y
port 6 nsew signal output
rlabel locali s 137 51 171 129 6 Y
port 6 nsew signal output
rlabel locali s 29 291 291 325 6 Y
port 6 nsew signal output
rlabel locali s 29 163 63 291 6 Y
port 6 nsew signal output
rlabel locali s 29 129 459 163 6 Y
port 6 nsew signal output
rlabel locali s 1001 17 1067 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 205 17 275 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 37 17 103 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 1196 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1196 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1001 383 1067 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 751 383 885 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 561 383 627 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 393 383 459 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 1196 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 1196 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3720546
string GDS_START 3710476
<< end >>
