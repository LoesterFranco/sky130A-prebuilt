magic
tech sky130A
magscale 1 2
timestamp 1604502729
<< locali >>
rect 109 270 167 356
rect 975 236 1041 317
rect 1364 467 1523 533
rect 1380 262 1414 467
rect 1328 197 1414 262
rect 1741 231 1807 297
rect 1328 88 1607 197
rect 2519 168 2569 596
rect 2503 88 2569 168
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2592 683
rect 24 236 75 596
rect 115 390 165 649
rect 201 581 787 615
rect 201 326 235 581
rect 269 513 596 547
rect 269 364 367 513
rect 409 414 497 479
rect 409 378 483 414
rect 531 409 596 513
rect 201 260 289 326
rect 201 236 258 260
rect 24 202 258 236
rect 323 204 367 364
rect 24 70 90 202
rect 124 17 190 168
rect 224 85 258 202
rect 295 123 367 204
rect 433 123 483 378
rect 562 218 596 409
rect 637 410 703 547
rect 737 450 787 581
rect 821 581 1009 615
rect 821 410 855 581
rect 637 376 855 410
rect 637 375 703 376
rect 889 375 941 547
rect 975 512 1009 581
rect 1081 546 1153 649
rect 1230 581 1743 615
rect 1230 512 1330 581
rect 975 478 1330 512
rect 562 184 635 218
rect 517 85 567 150
rect 224 51 567 85
rect 601 85 635 184
rect 669 119 703 375
rect 737 310 798 342
rect 737 276 857 310
rect 739 85 789 225
rect 601 51 789 85
rect 823 85 857 276
rect 891 134 941 375
rect 991 398 1057 444
rect 991 364 1160 398
rect 1194 364 1262 444
rect 1126 317 1160 364
rect 1126 251 1194 317
rect 1126 202 1160 251
rect 993 168 1160 202
rect 1228 213 1262 364
rect 1296 368 1330 478
rect 1296 302 1346 368
rect 993 85 1059 168
rect 823 51 1059 85
rect 1093 17 1194 127
rect 1228 77 1294 213
rect 1448 234 1511 430
rect 1557 297 1591 581
rect 1625 364 1675 547
rect 1549 231 1607 297
rect 1641 213 1675 364
rect 1709 365 1743 581
rect 1777 399 1811 649
rect 1851 581 2395 615
rect 1851 399 1945 581
rect 2160 548 2231 581
rect 1709 331 1877 365
rect 1641 77 1707 213
rect 1741 17 1809 197
rect 1843 114 1877 331
rect 1911 268 1945 399
rect 1979 514 2013 547
rect 2277 514 2327 547
rect 1979 480 2327 514
rect 1979 380 2013 480
rect 1911 148 1977 268
rect 2053 252 2103 446
rect 2137 286 2203 430
rect 2239 370 2327 480
rect 2014 148 2183 252
rect 2239 250 2273 370
rect 2361 336 2395 581
rect 2429 370 2479 649
rect 2307 270 2395 336
rect 1843 51 2115 114
rect 2149 98 2183 148
rect 2217 244 2273 250
rect 2217 132 2283 244
rect 2429 236 2485 336
rect 2317 202 2485 236
rect 2317 98 2351 202
rect 2149 64 2351 98
rect 2385 17 2469 162
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2592 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
<< metal1 >>
rect 0 683 2592 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2592 683
rect 0 617 2592 649
rect 0 17 2592 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2592 17
rect 0 -49 2592 -17
<< obsm1 >>
rect 403 421 461 430
rect 883 421 941 430
rect 1459 421 1517 430
rect 2131 421 2189 430
rect 403 393 2189 421
rect 403 384 461 393
rect 883 384 941 393
rect 1459 384 1517 393
rect 2131 384 2189 393
<< labels >>
rlabel locali s 109 270 167 356 6 A
port 1 nsew signal input
rlabel locali s 975 236 1041 317 6 B
port 2 nsew signal input
rlabel locali s 1741 231 1807 297 6 CIN
port 3 nsew signal input
rlabel locali s 1380 262 1414 467 6 COUT
port 4 nsew signal output
rlabel locali s 1364 467 1523 533 6 COUT
port 4 nsew signal output
rlabel locali s 1328 197 1414 262 6 COUT
port 4 nsew signal output
rlabel locali s 1328 88 1607 197 6 COUT
port 4 nsew signal output
rlabel locali s 2519 168 2569 596 6 SUM
port 5 nsew signal output
rlabel locali s 2503 88 2569 168 6 SUM
port 5 nsew signal output
rlabel metal1 s 0 -49 2592 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 2592 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2592 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 2593892
string GDS_START 2574762
<< end >>
