magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 2392 561
rect 104 427 170 527
rect 19 195 89 325
rect 103 17 169 93
rect 376 449 442 527
rect 356 157 390 337
rect 752 433 786 527
rect 492 271 559 337
rect 617 157 651 223
rect 707 207 807 331
rect 356 123 651 157
rect 1185 367 1219 527
rect 395 17 461 89
rect 495 61 530 123
rect 1561 427 1622 527
rect 1779 325 1815 527
rect 753 17 793 105
rect 1143 17 1217 117
rect 1851 306 1917 486
rect 1953 323 1987 527
rect 1851 299 1923 306
rect 1882 286 1923 299
rect 1889 178 1923 286
rect 1882 165 1923 178
rect 1548 17 1622 123
rect 1851 158 1923 165
rect 2143 299 2204 527
rect 2238 289 2288 465
rect 1779 17 1817 139
rect 1851 51 1917 158
rect 1951 17 1997 138
rect 2138 17 2204 161
rect 2247 159 2288 289
rect 2322 279 2356 527
rect 2238 53 2288 159
rect 2322 17 2356 191
rect 0 -17 2392 17
<< obsli1 >>
rect 36 393 70 493
rect 36 391 169 393
rect 36 359 129 391
rect 123 357 129 359
rect 163 357 169 391
rect 123 194 169 357
rect 123 161 162 194
rect 35 127 162 161
rect 204 187 249 493
rect 204 153 210 187
rect 244 153 249 187
rect 204 143 249 153
rect 35 69 69 127
rect 203 69 249 143
rect 287 415 342 489
rect 539 449 718 483
rect 287 372 650 415
rect 287 89 321 372
rect 424 225 458 372
rect 616 337 650 372
rect 684 399 718 449
rect 841 413 897 488
rect 937 438 1151 472
rect 841 399 875 413
rect 684 365 875 399
rect 995 391 1083 402
rect 616 271 655 337
rect 424 191 493 225
rect 841 173 875 365
rect 685 139 875 173
rect 909 207 957 381
rect 995 357 1041 391
rect 1075 357 1083 391
rect 995 331 1083 357
rect 1117 315 1151 438
rect 1253 427 1303 493
rect 1348 433 1525 467
rect 1117 297 1219 315
rect 1059 263 1219 297
rect 909 187 1025 207
rect 909 153 949 187
rect 983 153 1025 187
rect 909 141 1025 153
rect 287 55 361 89
rect 685 89 719 139
rect 841 107 875 139
rect 1059 107 1093 263
rect 1185 249 1219 263
rect 1127 213 1161 219
rect 1253 213 1287 427
rect 1321 391 1359 393
rect 1321 357 1325 391
rect 1321 249 1359 357
rect 1393 315 1457 381
rect 1127 153 1287 213
rect 1393 207 1431 315
rect 1491 281 1525 433
rect 1679 381 1745 491
rect 1559 315 1745 381
rect 564 55 719 89
rect 841 73 911 107
rect 945 73 1093 107
rect 1253 107 1287 153
rect 1321 187 1431 207
rect 1321 153 1328 187
rect 1362 153 1431 187
rect 1321 141 1431 153
rect 1465 265 1525 281
rect 1708 265 1745 315
rect 1465 199 1674 265
rect 1708 199 1855 265
rect 1465 107 1499 199
rect 1708 165 1745 199
rect 1253 73 1345 107
rect 1391 73 1499 107
rect 1672 60 1745 165
rect 2041 265 2107 485
rect 2041 199 2213 265
rect 2041 69 2091 199
<< obsli1c >>
rect 129 357 163 391
rect 210 153 244 187
rect 1041 357 1075 391
rect 949 153 983 187
rect 1325 357 1359 391
rect 1328 153 1362 187
<< metal1 >>
rect 0 496 2392 592
rect 0 -48 2392 48
<< obsm1 >>
rect 117 391 175 397
rect 117 357 129 391
rect 163 388 175 391
rect 1029 391 1087 397
rect 1029 388 1041 391
rect 163 360 1041 388
rect 163 357 175 360
rect 117 351 175 357
rect 1029 357 1041 360
rect 1075 388 1087 391
rect 1313 391 1371 397
rect 1313 388 1325 391
rect 1075 360 1325 388
rect 1075 357 1087 360
rect 1029 351 1087 357
rect 1313 357 1325 360
rect 1359 357 1371 391
rect 1313 351 1371 357
rect 198 187 256 193
rect 198 153 210 187
rect 244 184 256 187
rect 937 187 995 193
rect 937 184 949 187
rect 244 156 949 184
rect 244 153 256 156
rect 198 147 256 153
rect 937 153 949 156
rect 983 184 995 187
rect 1316 187 1374 193
rect 1316 184 1328 187
rect 983 156 1328 184
rect 983 153 995 156
rect 937 147 995 153
rect 1316 153 1328 156
rect 1362 153 1374 187
rect 1316 147 1374 153
<< labels >>
rlabel locali s 492 271 559 337 6 D
port 1 nsew signal input
rlabel locali s 1889 178 1923 286 6 Q
port 2 nsew signal output
rlabel locali s 1882 286 1923 299 6 Q
port 2 nsew signal output
rlabel locali s 1882 165 1923 178 6 Q
port 2 nsew signal output
rlabel locali s 1851 306 1917 486 6 Q
port 2 nsew signal output
rlabel locali s 1851 299 1923 306 6 Q
port 2 nsew signal output
rlabel locali s 1851 158 1923 165 6 Q
port 2 nsew signal output
rlabel locali s 1851 51 1917 158 6 Q
port 2 nsew signal output
rlabel locali s 2247 159 2288 289 6 Q_N
port 3 nsew signal output
rlabel locali s 2238 289 2288 465 6 Q_N
port 3 nsew signal output
rlabel locali s 2238 53 2288 159 6 Q_N
port 3 nsew signal output
rlabel locali s 707 207 807 331 6 SCD
port 4 nsew signal input
rlabel locali s 617 157 651 223 6 SCE
port 5 nsew signal input
rlabel locali s 495 61 530 123 6 SCE
port 5 nsew signal input
rlabel locali s 356 157 390 337 6 SCE
port 5 nsew signal input
rlabel locali s 356 123 651 157 6 SCE
port 5 nsew signal input
rlabel locali s 19 195 89 325 6 CLK
port 6 nsew clock input
rlabel locali s 2322 17 2356 191 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 2138 17 2204 161 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1951 17 1997 138 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1779 17 1817 139 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1548 17 1622 123 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1143 17 1217 117 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 753 17 793 105 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 395 17 461 89 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 103 17 169 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 2392 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 2392 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 2322 279 2356 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 2143 299 2204 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1953 323 1987 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1779 325 1815 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1561 427 1622 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1185 367 1219 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 752 433 786 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 376 449 442 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 104 427 170 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 2392 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 2392 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2392 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 361040
string GDS_START 343158
<< end >>
