magic
tech sky130A
magscale 1 2
timestamp 1604502705
<< nwell >>
rect -38 332 1094 704
<< pwell >>
rect 0 0 1056 49
<< scnmos >>
rect 84 74 114 222
rect 338 74 368 222
rect 424 74 454 222
rect 510 74 540 222
rect 596 74 626 222
rect 682 74 712 222
rect 768 74 798 222
rect 856 74 886 222
rect 942 74 972 222
<< pmoshvt >>
rect 98 368 128 592
rect 300 368 330 592
rect 390 368 420 592
rect 480 368 510 592
rect 580 368 610 592
rect 670 368 700 592
rect 760 368 790 592
rect 850 368 880 592
rect 940 368 970 592
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 210 171 222
rect 114 176 125 210
rect 159 176 171 210
rect 114 120 171 176
rect 114 86 125 120
rect 159 86 171 120
rect 114 74 171 86
rect 281 210 338 222
rect 281 176 293 210
rect 327 176 338 210
rect 281 120 338 176
rect 281 86 293 120
rect 327 86 338 120
rect 281 74 338 86
rect 368 193 424 222
rect 368 159 379 193
rect 413 159 424 193
rect 368 120 424 159
rect 368 86 379 120
rect 413 86 424 120
rect 368 74 424 86
rect 454 210 510 222
rect 454 176 465 210
rect 499 176 510 210
rect 454 120 510 176
rect 454 86 465 120
rect 499 86 510 120
rect 454 74 510 86
rect 540 193 596 222
rect 540 159 551 193
rect 585 159 596 193
rect 540 120 596 159
rect 540 86 551 120
rect 585 86 596 120
rect 540 74 596 86
rect 626 210 682 222
rect 626 176 637 210
rect 671 176 682 210
rect 626 120 682 176
rect 626 86 637 120
rect 671 86 682 120
rect 626 74 682 86
rect 712 207 768 222
rect 712 173 723 207
rect 757 173 768 207
rect 712 74 768 173
rect 798 120 856 222
rect 798 86 810 120
rect 844 86 856 120
rect 798 74 856 86
rect 886 177 942 222
rect 886 143 897 177
rect 931 143 942 177
rect 886 74 942 143
rect 972 153 1029 222
rect 972 119 983 153
rect 1017 119 1029 153
rect 972 74 1029 119
<< pdiff >>
rect 39 580 98 592
rect 39 546 51 580
rect 85 546 98 580
rect 39 510 98 546
rect 39 476 51 510
rect 85 476 98 510
rect 39 440 98 476
rect 39 406 51 440
rect 85 406 98 440
rect 39 368 98 406
rect 128 580 187 592
rect 128 546 141 580
rect 175 546 187 580
rect 128 497 187 546
rect 128 463 141 497
rect 175 463 187 497
rect 128 414 187 463
rect 128 380 141 414
rect 175 380 187 414
rect 128 368 187 380
rect 241 580 300 592
rect 241 546 253 580
rect 287 546 300 580
rect 241 497 300 546
rect 241 463 253 497
rect 287 463 300 497
rect 241 414 300 463
rect 241 380 253 414
rect 287 380 300 414
rect 241 368 300 380
rect 330 580 390 592
rect 330 546 343 580
rect 377 546 390 580
rect 330 497 390 546
rect 330 463 343 497
rect 377 463 390 497
rect 330 414 390 463
rect 330 380 343 414
rect 377 380 390 414
rect 330 368 390 380
rect 420 580 480 592
rect 420 546 433 580
rect 467 546 480 580
rect 420 497 480 546
rect 420 463 433 497
rect 467 463 480 497
rect 420 414 480 463
rect 420 380 433 414
rect 467 380 480 414
rect 420 368 480 380
rect 510 580 580 592
rect 510 546 523 580
rect 557 546 580 580
rect 510 497 580 546
rect 510 463 523 497
rect 557 463 580 497
rect 510 414 580 463
rect 510 380 523 414
rect 557 380 580 414
rect 510 368 580 380
rect 610 580 670 592
rect 610 546 623 580
rect 657 546 670 580
rect 610 497 670 546
rect 610 463 623 497
rect 657 463 670 497
rect 610 414 670 463
rect 610 380 623 414
rect 657 380 670 414
rect 610 368 670 380
rect 700 547 760 592
rect 700 513 713 547
rect 747 513 760 547
rect 700 479 760 513
rect 700 445 713 479
rect 747 445 760 479
rect 700 411 760 445
rect 700 377 713 411
rect 747 377 760 411
rect 700 368 760 377
rect 790 580 850 592
rect 790 546 803 580
rect 837 546 850 580
rect 790 462 850 546
rect 790 428 803 462
rect 837 428 850 462
rect 790 368 850 428
rect 880 547 940 592
rect 880 513 893 547
rect 927 513 940 547
rect 880 479 940 513
rect 880 445 893 479
rect 927 445 940 479
rect 880 411 940 445
rect 880 377 893 411
rect 927 377 940 411
rect 880 368 940 377
rect 970 580 1029 592
rect 970 546 983 580
rect 1017 546 1029 580
rect 970 497 1029 546
rect 970 463 983 497
rect 1017 463 1029 497
rect 970 414 1029 463
rect 970 380 983 414
rect 1017 380 1029 414
rect 970 368 1029 380
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 125 176 159 210
rect 125 86 159 120
rect 293 176 327 210
rect 293 86 327 120
rect 379 159 413 193
rect 379 86 413 120
rect 465 176 499 210
rect 465 86 499 120
rect 551 159 585 193
rect 551 86 585 120
rect 637 176 671 210
rect 637 86 671 120
rect 723 173 757 207
rect 810 86 844 120
rect 897 143 931 177
rect 983 119 1017 153
<< pdiffc >>
rect 51 546 85 580
rect 51 476 85 510
rect 51 406 85 440
rect 141 546 175 580
rect 141 463 175 497
rect 141 380 175 414
rect 253 546 287 580
rect 253 463 287 497
rect 253 380 287 414
rect 343 546 377 580
rect 343 463 377 497
rect 343 380 377 414
rect 433 546 467 580
rect 433 463 467 497
rect 433 380 467 414
rect 523 546 557 580
rect 523 463 557 497
rect 523 380 557 414
rect 623 546 657 580
rect 623 463 657 497
rect 623 380 657 414
rect 713 513 747 547
rect 713 445 747 479
rect 713 377 747 411
rect 803 546 837 580
rect 803 428 837 462
rect 893 513 927 547
rect 893 445 927 479
rect 893 377 927 411
rect 983 546 1017 580
rect 983 463 1017 497
rect 983 380 1017 414
<< poly >>
rect 98 592 128 618
rect 300 592 330 618
rect 390 592 420 618
rect 480 592 510 618
rect 580 592 610 618
rect 670 592 700 618
rect 760 592 790 618
rect 850 592 880 618
rect 940 592 970 618
rect 98 353 128 368
rect 300 353 330 368
rect 390 353 420 368
rect 480 353 510 368
rect 580 353 610 368
rect 670 353 700 368
rect 760 353 790 368
rect 850 353 880 368
rect 940 353 970 368
rect 95 345 131 353
rect 297 345 333 353
rect 387 345 423 353
rect 477 345 513 353
rect 577 345 613 353
rect 25 315 613 345
rect 667 345 703 353
rect 757 345 793 353
rect 847 345 883 353
rect 937 345 973 353
rect 667 315 1009 345
rect 25 310 131 315
rect 25 276 41 310
rect 75 276 131 310
rect 25 260 131 276
rect 682 294 1009 315
rect 84 222 114 260
rect 193 246 626 267
rect 193 212 209 246
rect 243 237 626 246
rect 243 212 259 237
rect 338 222 368 237
rect 424 222 454 237
rect 510 222 540 237
rect 596 222 626 237
rect 682 260 823 294
rect 857 260 891 294
rect 925 260 959 294
rect 993 260 1009 294
rect 682 244 1009 260
rect 682 222 712 244
rect 768 222 798 244
rect 856 222 886 244
rect 942 222 972 244
rect 193 178 259 212
rect 193 144 209 178
rect 243 144 259 178
rect 193 110 259 144
rect 193 76 209 110
rect 243 76 259 110
rect 84 48 114 74
rect 193 60 259 76
rect 338 48 368 74
rect 424 48 454 74
rect 510 48 540 74
rect 596 48 626 74
rect 682 48 712 74
rect 768 48 798 74
rect 856 48 886 74
rect 942 48 972 74
<< polycont >>
rect 41 276 75 310
rect 209 212 243 246
rect 823 260 857 294
rect 891 260 925 294
rect 959 260 993 294
rect 209 144 243 178
rect 209 76 243 110
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 35 580 85 649
rect 35 546 51 580
rect 35 510 85 546
rect 35 476 51 510
rect 35 440 85 476
rect 35 406 51 440
rect 35 390 85 406
rect 125 580 191 596
rect 125 546 141 580
rect 175 546 191 580
rect 125 497 191 546
rect 125 463 141 497
rect 175 463 191 497
rect 125 414 191 463
rect 125 380 141 414
rect 175 380 191 414
rect 25 310 91 356
rect 25 276 41 310
rect 75 276 91 310
rect 25 260 91 276
rect 125 262 191 380
rect 237 580 287 596
rect 237 546 253 580
rect 237 497 287 546
rect 237 463 253 497
rect 237 414 287 463
rect 237 380 253 414
rect 237 330 287 380
rect 327 580 377 649
rect 327 546 343 580
rect 327 497 377 546
rect 327 463 343 497
rect 327 414 377 463
rect 327 380 343 414
rect 327 364 377 380
rect 417 580 467 596
rect 417 546 433 580
rect 417 497 467 546
rect 417 463 433 497
rect 417 414 467 463
rect 417 380 433 414
rect 417 330 467 380
rect 507 580 573 649
rect 507 546 523 580
rect 557 546 573 580
rect 507 497 573 546
rect 507 463 523 497
rect 557 463 573 497
rect 507 414 573 463
rect 507 380 523 414
rect 557 380 573 414
rect 507 364 573 380
rect 607 581 1033 615
rect 607 580 657 581
rect 607 546 623 580
rect 803 580 837 581
rect 607 497 657 546
rect 607 463 623 497
rect 607 414 657 463
rect 607 380 623 414
rect 607 330 657 380
rect 237 296 657 330
rect 697 513 713 547
rect 747 513 763 547
rect 697 479 763 513
rect 697 445 713 479
rect 747 445 763 479
rect 697 411 763 445
rect 983 580 1033 581
rect 803 462 837 546
rect 803 412 837 428
rect 877 513 893 547
rect 927 513 943 547
rect 877 479 943 513
rect 877 445 893 479
rect 927 445 943 479
rect 697 377 713 411
rect 747 378 763 411
rect 877 411 943 445
rect 877 378 893 411
rect 747 377 893 378
rect 927 377 943 411
rect 697 344 943 377
rect 1017 546 1033 580
rect 983 497 1033 546
rect 1017 463 1033 497
rect 983 414 1033 463
rect 1017 380 1033 414
rect 983 364 1033 380
rect 697 310 763 344
rect 125 246 259 262
rect 125 226 209 246
rect 23 210 73 226
rect 23 176 39 210
rect 23 120 73 176
rect 23 86 39 120
rect 23 17 73 86
rect 109 212 209 226
rect 243 212 259 246
rect 109 210 259 212
rect 109 176 125 210
rect 159 178 259 210
rect 159 176 209 178
rect 109 144 209 176
rect 243 144 259 178
rect 109 120 259 144
rect 109 86 125 120
rect 159 110 259 120
rect 159 86 209 110
rect 109 76 209 86
rect 243 76 259 110
rect 109 60 259 76
rect 293 228 687 262
rect 293 210 327 228
rect 465 210 499 228
rect 293 120 327 176
rect 293 70 327 86
rect 363 193 429 194
rect 363 159 379 193
rect 413 159 429 193
rect 363 120 429 159
rect 363 86 379 120
rect 413 86 429 120
rect 363 17 429 86
rect 637 210 687 228
rect 465 120 499 176
rect 465 70 499 86
rect 535 193 601 194
rect 535 159 551 193
rect 585 159 601 193
rect 535 120 601 159
rect 535 86 551 120
rect 585 86 601 120
rect 535 17 601 86
rect 671 176 687 210
rect 637 120 687 176
rect 723 226 763 310
rect 807 294 1031 310
rect 807 260 823 294
rect 857 260 891 294
rect 925 260 959 294
rect 993 260 1031 294
rect 807 236 1031 260
rect 723 207 773 226
rect 757 202 773 207
rect 757 177 931 202
rect 757 173 897 177
rect 723 154 897 173
rect 671 86 810 120
rect 844 86 861 120
rect 897 119 931 143
rect 967 153 1033 202
rect 967 119 983 153
rect 1017 119 1033 153
rect 637 85 861 86
rect 967 85 1033 119
rect 637 51 1033 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 683 1056 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 0 617 1056 649
rect 0 17 1056 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -49 1056 -17
<< labels >>
rlabel comment s 0 0 0 0 4 einvn_4
flabel pwell s 0 0 1056 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 0 617 1056 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 0 617 1056 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 1056 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 TE_B
port 2 nsew
flabel corelocali s 895 242 929 276 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 991 242 1025 276 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 Z
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 1056 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2119416
string GDS_START 2110256
<< end >>
