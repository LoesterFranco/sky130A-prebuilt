magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 22 215 88 255
rect 696 323 772 493
rect 884 323 960 493
rect 1072 323 1148 493
rect 1260 323 1336 493
rect 696 289 1448 323
rect 1372 181 1448 289
rect 696 147 1448 181
rect 696 52 772 147
rect 884 52 960 147
rect 1072 52 1148 147
rect 1260 52 1336 147
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 19 323 85 432
rect 129 357 163 527
rect 19 289 166 323
rect 210 309 296 493
rect 132 265 166 289
rect 132 199 228 265
rect 262 255 296 309
rect 330 323 396 493
rect 440 357 474 527
rect 508 323 584 493
rect 628 357 662 527
rect 816 367 850 527
rect 1004 367 1038 527
rect 1192 367 1226 527
rect 1380 367 1414 527
rect 330 289 662 323
rect 628 255 662 289
rect 262 215 584 255
rect 628 215 1182 255
rect 132 181 166 199
rect 19 147 166 181
rect 262 165 296 215
rect 628 181 662 215
rect 19 52 85 147
rect 129 17 163 113
rect 210 52 296 165
rect 330 147 662 181
rect 330 52 396 147
rect 440 17 474 113
rect 508 52 584 147
rect 628 17 662 113
rect 816 17 850 113
rect 1004 17 1038 113
rect 1192 17 1226 113
rect 1380 17 1414 113
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< labels >>
rlabel locali s 22 215 88 255 6 A
port 1 nsew signal input
rlabel locali s 1372 181 1448 289 6 X
port 2 nsew signal output
rlabel locali s 1260 323 1336 493 6 X
port 2 nsew signal output
rlabel locali s 1260 52 1336 147 6 X
port 2 nsew signal output
rlabel locali s 1072 323 1148 493 6 X
port 2 nsew signal output
rlabel locali s 1072 52 1148 147 6 X
port 2 nsew signal output
rlabel locali s 884 323 960 493 6 X
port 2 nsew signal output
rlabel locali s 884 52 960 147 6 X
port 2 nsew signal output
rlabel locali s 696 323 772 493 6 X
port 2 nsew signal output
rlabel locali s 696 289 1448 323 6 X
port 2 nsew signal output
rlabel locali s 696 147 1448 181 6 X
port 2 nsew signal output
rlabel locali s 696 52 772 147 6 X
port 2 nsew signal output
rlabel metal1 s 0 -48 1472 48 8 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 496 1472 592 6 VPWR
port 4 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1472 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1714314
string GDS_START 1703340
<< end >>
