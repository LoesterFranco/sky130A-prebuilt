magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 301 333 377 493
rect 489 401 565 493
rect 677 401 753 493
rect 489 333 753 401
rect 865 333 941 493
rect 1157 333 1233 493
rect 1345 333 1421 493
rect 301 289 1421 333
rect 86 215 166 255
rect 609 215 711 289
rect 745 215 986 255
rect 1037 215 1420 255
rect 609 181 643 215
rect 301 127 643 181
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 17 289 85 493
rect 129 289 267 527
rect 421 367 455 527
rect 609 435 643 527
rect 797 367 831 527
rect 985 367 1123 527
rect 1277 367 1311 527
rect 1465 289 1531 527
rect 17 181 52 289
rect 211 215 565 255
rect 211 181 267 215
rect 17 143 267 181
rect 17 51 85 143
rect 677 143 1421 181
rect 677 127 1035 143
rect 129 17 179 109
rect 217 51 1035 93
rect 1073 17 1123 109
rect 1157 51 1233 143
rect 1277 17 1311 109
rect 1345 51 1421 143
rect 1465 17 1531 181
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
<< metal1 >>
rect 0 561 1564 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 0 496 1564 527
rect 0 17 1564 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
rect 0 -48 1564 -17
<< labels >>
rlabel locali s 86 215 166 255 6 A_N
port 1 nsew signal input
rlabel locali s 745 215 986 255 6 B
port 2 nsew signal input
rlabel locali s 1037 215 1420 255 6 C
port 3 nsew signal input
rlabel locali s 1345 333 1421 493 6 Y
port 4 nsew signal output
rlabel locali s 1157 333 1233 493 6 Y
port 4 nsew signal output
rlabel locali s 865 333 941 493 6 Y
port 4 nsew signal output
rlabel locali s 677 401 753 493 6 Y
port 4 nsew signal output
rlabel locali s 609 215 711 289 6 Y
port 4 nsew signal output
rlabel locali s 609 181 643 215 6 Y
port 4 nsew signal output
rlabel locali s 489 401 565 493 6 Y
port 4 nsew signal output
rlabel locali s 489 333 753 401 6 Y
port 4 nsew signal output
rlabel locali s 301 333 377 493 6 Y
port 4 nsew signal output
rlabel locali s 301 289 1421 333 6 Y
port 4 nsew signal output
rlabel locali s 301 127 643 181 6 Y
port 4 nsew signal output
rlabel metal1 s 0 -48 1564 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 1564 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1564 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2287458
string GDS_START 2275096
<< end >>
