magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 1382 704
<< pwell >>
rect 0 0 1344 49
<< scnmos >>
rect 87 74 117 202
rect 201 74 231 202
rect 439 74 469 222
rect 530 74 560 222
rect 648 74 678 222
rect 734 74 764 222
rect 943 74 973 222
rect 1043 74 1073 222
rect 1129 74 1159 222
rect 1229 74 1259 222
<< pmoshvt >>
rect 86 368 116 568
rect 210 368 240 568
rect 442 368 472 592
rect 532 368 562 592
rect 642 368 672 592
rect 732 368 762 592
rect 928 368 958 592
rect 1018 368 1048 592
rect 1128 368 1158 592
rect 1226 368 1256 592
<< ndiff >>
rect 30 190 87 202
rect 30 156 42 190
rect 76 156 87 190
rect 30 120 87 156
rect 30 86 42 120
rect 76 86 87 120
rect 30 74 87 86
rect 117 190 201 202
rect 117 156 142 190
rect 176 156 201 190
rect 117 120 201 156
rect 117 86 142 120
rect 176 86 201 120
rect 117 74 201 86
rect 231 190 288 202
rect 231 156 242 190
rect 276 156 288 190
rect 231 120 288 156
rect 231 86 242 120
rect 276 86 288 120
rect 231 74 288 86
rect 373 136 439 222
rect 373 102 385 136
rect 419 102 439 136
rect 373 74 439 102
rect 469 168 530 222
rect 469 134 485 168
rect 519 134 530 168
rect 469 74 530 134
rect 560 100 648 222
rect 560 74 587 100
rect 575 66 587 74
rect 621 74 648 100
rect 678 116 734 222
rect 678 82 689 116
rect 723 82 734 116
rect 678 74 734 82
rect 764 184 832 222
rect 764 150 780 184
rect 814 150 832 184
rect 764 74 832 150
rect 886 174 943 222
rect 886 140 898 174
rect 932 140 943 174
rect 886 74 943 140
rect 973 147 1043 222
rect 973 113 998 147
rect 1032 113 1043 147
rect 973 74 1043 113
rect 1073 210 1129 222
rect 1073 176 1084 210
rect 1118 176 1129 210
rect 1073 120 1129 176
rect 1073 86 1084 120
rect 1118 86 1129 120
rect 1073 74 1129 86
rect 1159 147 1229 222
rect 1159 113 1184 147
rect 1218 113 1229 147
rect 1159 74 1229 113
rect 1259 210 1316 222
rect 1259 176 1270 210
rect 1304 176 1316 210
rect 1259 120 1316 176
rect 1259 86 1270 120
rect 1304 86 1316 120
rect 1259 74 1316 86
rect 621 66 633 74
rect 575 54 633 66
<< pdiff >>
rect 134 568 192 578
rect 373 573 442 592
rect 27 560 86 568
rect 27 526 39 560
rect 73 526 86 560
rect 27 492 86 526
rect 27 458 39 492
rect 73 458 86 492
rect 27 424 86 458
rect 27 390 39 424
rect 73 390 86 424
rect 27 368 86 390
rect 116 566 210 568
rect 116 532 146 566
rect 180 532 210 566
rect 116 368 210 532
rect 240 414 319 568
rect 240 380 263 414
rect 297 380 319 414
rect 240 368 319 380
rect 373 539 385 573
rect 419 539 442 573
rect 373 368 442 539
rect 472 580 532 592
rect 472 546 485 580
rect 519 546 532 580
rect 472 497 532 546
rect 472 463 485 497
rect 519 463 532 497
rect 472 414 532 463
rect 472 380 485 414
rect 519 380 532 414
rect 472 368 532 380
rect 562 580 642 592
rect 562 546 585 580
rect 619 546 642 580
rect 562 488 642 546
rect 562 454 585 488
rect 619 454 642 488
rect 562 368 642 454
rect 672 580 732 592
rect 672 546 685 580
rect 719 546 732 580
rect 672 500 732 546
rect 672 466 685 500
rect 719 466 732 500
rect 672 420 732 466
rect 672 386 685 420
rect 719 386 732 420
rect 672 368 732 386
rect 762 580 928 592
rect 762 546 775 580
rect 809 546 881 580
rect 915 546 928 580
rect 762 508 928 546
rect 762 474 775 508
rect 809 474 881 508
rect 915 474 928 508
rect 762 368 928 474
rect 958 580 1018 592
rect 958 546 971 580
rect 1005 546 1018 580
rect 958 510 1018 546
rect 958 476 971 510
rect 1005 476 1018 510
rect 958 440 1018 476
rect 958 406 971 440
rect 1005 406 1018 440
rect 958 368 1018 406
rect 1048 580 1128 592
rect 1048 546 1071 580
rect 1105 546 1128 580
rect 1048 508 1128 546
rect 1048 474 1071 508
rect 1105 474 1128 508
rect 1048 368 1128 474
rect 1158 580 1226 592
rect 1158 546 1171 580
rect 1205 546 1226 580
rect 1158 500 1226 546
rect 1158 466 1171 500
rect 1205 466 1226 500
rect 1158 420 1226 466
rect 1158 386 1171 420
rect 1205 386 1226 420
rect 1158 368 1226 386
rect 1256 580 1317 592
rect 1256 546 1271 580
rect 1305 546 1317 580
rect 1256 510 1317 546
rect 1256 476 1271 510
rect 1305 476 1317 510
rect 1256 440 1317 476
rect 1256 406 1271 440
rect 1305 406 1317 440
rect 1256 368 1317 406
<< ndiffc >>
rect 42 156 76 190
rect 42 86 76 120
rect 142 156 176 190
rect 142 86 176 120
rect 242 156 276 190
rect 242 86 276 120
rect 385 102 419 136
rect 485 134 519 168
rect 587 66 621 100
rect 689 82 723 116
rect 780 150 814 184
rect 898 140 932 174
rect 998 113 1032 147
rect 1084 176 1118 210
rect 1084 86 1118 120
rect 1184 113 1218 147
rect 1270 176 1304 210
rect 1270 86 1304 120
<< pdiffc >>
rect 39 526 73 560
rect 39 458 73 492
rect 39 390 73 424
rect 146 532 180 566
rect 263 380 297 414
rect 385 539 419 573
rect 485 546 519 580
rect 485 463 519 497
rect 485 380 519 414
rect 585 546 619 580
rect 585 454 619 488
rect 685 546 719 580
rect 685 466 719 500
rect 685 386 719 420
rect 775 546 809 580
rect 881 546 915 580
rect 775 474 809 508
rect 881 474 915 508
rect 971 546 1005 580
rect 971 476 1005 510
rect 971 406 1005 440
rect 1071 546 1105 580
rect 1071 474 1105 508
rect 1171 546 1205 580
rect 1171 466 1205 500
rect 1171 386 1205 420
rect 1271 546 1305 580
rect 1271 476 1305 510
rect 1271 406 1305 440
<< poly >>
rect 86 568 116 594
rect 210 568 240 594
rect 442 592 472 618
rect 532 592 562 618
rect 642 592 672 618
rect 732 592 762 618
rect 928 592 958 618
rect 1018 592 1048 618
rect 1128 592 1158 618
rect 1226 592 1256 618
rect 86 353 116 368
rect 210 353 240 368
rect 442 353 472 368
rect 532 353 562 368
rect 642 353 672 368
rect 732 353 762 368
rect 928 353 958 368
rect 1018 353 1048 368
rect 1128 353 1158 368
rect 1226 353 1256 368
rect 83 326 119 353
rect 83 310 153 326
rect 83 276 103 310
rect 137 276 153 310
rect 207 302 243 353
rect 439 336 475 353
rect 369 324 475 336
rect 529 324 565 353
rect 639 336 675 353
rect 729 336 765 353
rect 369 320 565 324
rect 83 260 153 276
rect 201 286 267 302
rect 87 202 117 260
rect 201 252 217 286
rect 251 252 267 286
rect 369 286 385 320
rect 419 286 565 320
rect 369 270 565 286
rect 625 320 765 336
rect 625 286 641 320
rect 675 286 709 320
rect 743 286 765 320
rect 625 270 765 286
rect 925 336 961 353
rect 1015 336 1051 353
rect 1125 336 1161 353
rect 1223 336 1259 353
rect 925 320 1077 336
rect 925 286 959 320
rect 993 286 1027 320
rect 1061 286 1077 320
rect 925 270 1077 286
rect 1125 320 1259 336
rect 1125 286 1141 320
rect 1175 286 1209 320
rect 1243 286 1259 320
rect 1125 270 1259 286
rect 201 236 267 252
rect 439 237 565 270
rect 201 202 231 236
rect 439 222 469 237
rect 530 222 560 237
rect 648 222 678 270
rect 734 222 764 270
rect 943 222 973 270
rect 1043 222 1073 270
rect 1129 222 1159 270
rect 1229 222 1259 270
rect 87 48 117 74
rect 201 48 231 74
rect 439 48 469 74
rect 530 48 560 74
rect 648 48 678 74
rect 734 48 764 74
rect 943 48 973 74
rect 1043 48 1073 74
rect 1129 48 1159 74
rect 1229 48 1259 74
<< polycont >>
rect 103 276 137 310
rect 217 252 251 286
rect 385 286 419 320
rect 641 286 675 320
rect 709 286 743 320
rect 959 286 993 320
rect 1027 286 1061 320
rect 1141 286 1175 320
rect 1209 286 1243 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 19 560 89 572
rect 19 526 39 560
rect 73 526 89 560
rect 19 492 89 526
rect 130 566 196 649
rect 130 532 146 566
rect 180 532 196 566
rect 130 516 196 532
rect 369 573 435 649
rect 369 539 385 573
rect 419 539 435 573
rect 369 516 435 539
rect 469 580 535 596
rect 469 546 485 580
rect 519 546 535 580
rect 19 458 39 492
rect 73 482 89 492
rect 469 497 535 546
rect 73 458 435 482
rect 19 448 435 458
rect 19 424 89 448
rect 19 390 39 424
rect 73 390 89 424
rect 19 206 53 390
rect 237 380 263 414
rect 297 380 335 414
rect 237 364 335 380
rect 87 310 167 356
rect 87 276 103 310
rect 137 276 167 310
rect 87 260 167 276
rect 201 286 267 302
rect 201 252 217 286
rect 251 252 267 286
rect 201 236 267 252
rect 301 236 335 364
rect 369 320 435 448
rect 469 463 485 497
rect 519 463 535 497
rect 469 414 535 463
rect 569 580 635 649
rect 569 546 585 580
rect 619 546 635 580
rect 569 488 635 546
rect 569 454 585 488
rect 619 454 635 488
rect 569 438 635 454
rect 669 580 735 596
rect 669 546 685 580
rect 719 546 735 580
rect 669 500 735 546
rect 669 466 685 500
rect 719 466 735 500
rect 469 380 485 414
rect 519 404 535 414
rect 669 424 735 466
rect 769 580 921 649
rect 769 546 775 580
rect 809 546 881 580
rect 915 546 921 580
rect 769 508 921 546
rect 769 474 775 508
rect 809 474 881 508
rect 915 474 921 508
rect 769 458 921 474
rect 955 580 1021 596
rect 955 546 971 580
rect 1005 546 1021 580
rect 955 510 1021 546
rect 955 476 971 510
rect 1005 476 1021 510
rect 955 440 1021 476
rect 1055 580 1121 649
rect 1055 546 1071 580
rect 1105 546 1121 580
rect 1055 508 1121 546
rect 1055 474 1071 508
rect 1105 474 1121 508
rect 1055 458 1121 474
rect 1155 580 1221 596
rect 1155 546 1171 580
rect 1205 546 1221 580
rect 1155 500 1221 546
rect 1155 466 1171 500
rect 1205 466 1221 500
rect 955 424 971 440
rect 669 420 971 424
rect 669 404 685 420
rect 519 386 685 404
rect 719 406 971 420
rect 1005 424 1021 440
rect 1155 424 1221 466
rect 1005 420 1221 424
rect 1005 406 1171 420
rect 719 390 1171 406
rect 719 386 839 390
rect 519 380 839 386
rect 469 370 839 380
rect 1155 386 1171 390
rect 1205 386 1221 420
rect 1255 580 1321 649
rect 1255 546 1271 580
rect 1305 546 1321 580
rect 1255 510 1321 546
rect 1255 476 1271 510
rect 1305 476 1321 510
rect 1255 440 1321 476
rect 1255 406 1271 440
rect 1305 406 1321 440
rect 1255 390 1321 406
rect 1155 370 1221 386
rect 469 364 535 370
rect 625 320 759 336
rect 369 286 385 320
rect 419 286 435 320
rect 369 270 435 286
rect 469 286 641 320
rect 675 286 709 320
rect 743 286 759 320
rect 469 236 503 286
rect 793 252 839 370
rect 889 320 1077 356
rect 1273 336 1319 356
rect 889 286 959 320
rect 993 286 1027 320
rect 1061 286 1077 320
rect 889 270 1077 286
rect 1125 320 1319 336
rect 1125 286 1141 320
rect 1175 286 1209 320
rect 1243 286 1319 320
rect 1125 270 1319 286
rect 19 190 92 206
rect 301 202 503 236
rect 537 218 839 252
rect 19 156 42 190
rect 76 156 92 190
rect 19 120 92 156
rect 19 86 42 120
rect 76 86 92 120
rect 19 70 92 86
rect 126 190 192 202
rect 126 156 142 190
rect 176 156 192 190
rect 126 120 192 156
rect 126 86 142 120
rect 176 86 192 120
rect 126 17 192 86
rect 226 190 335 202
rect 226 156 242 190
rect 276 156 335 190
rect 537 168 571 218
rect 882 210 1320 236
rect 882 202 1084 210
rect 226 120 335 156
rect 226 86 242 120
rect 276 86 335 120
rect 226 70 335 86
rect 369 136 435 168
rect 369 102 385 136
rect 419 102 435 136
rect 469 134 485 168
rect 519 134 571 168
rect 605 150 780 184
rect 814 150 836 184
rect 882 174 948 202
rect 369 100 435 102
rect 605 100 639 150
rect 882 140 898 174
rect 932 140 948 174
rect 1118 202 1270 210
rect 1118 176 1134 202
rect 882 124 948 140
rect 982 147 1048 163
rect 369 66 587 100
rect 621 66 639 100
rect 673 82 689 116
rect 723 85 739 116
rect 982 113 998 147
rect 1032 113 1048 147
rect 982 85 1048 113
rect 723 82 1048 85
rect 673 51 1048 82
rect 1084 120 1134 176
rect 1304 176 1320 210
rect 1118 86 1134 120
rect 1084 70 1134 86
rect 1168 147 1234 163
rect 1168 113 1184 147
rect 1218 113 1234 147
rect 1168 17 1234 113
rect 1270 120 1320 176
rect 1304 86 1320 120
rect 1270 70 1320 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
<< metal1 >>
rect 0 683 1344 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 0 617 1344 649
rect 0 17 1344 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
rect 0 -49 1344 -17
<< labels >>
rlabel comment s 0 0 0 0 4 nand4bb_2
flabel pwell s 0 0 1344 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 1344 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 1344 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 1344 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew
flabel corelocali s 799 242 833 276 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 1279 316 1313 350 0 FreeSans 340 0 0 0 D
port 4 nsew
flabel corelocali s 223 242 257 276 0 FreeSans 340 0 0 0 B_N
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 1344 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1866798
string GDS_START 1856182
<< end >>
