magic
tech sky130A
magscale 1 2
timestamp 1601050088
<< locali >>
rect 91 332 359 367
rect 91 298 545 332
rect 313 162 420 253
rect 469 252 545 298
rect 589 288 655 430
rect 867 332 928 355
rect 757 252 928 332
rect 757 184 839 252
rect 2614 226 2665 596
rect 2599 70 2665 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2688 683
rect 23 435 89 596
rect 123 469 189 649
rect 297 503 511 596
rect 619 537 685 649
rect 733 526 799 596
rect 941 560 1007 649
rect 1165 526 1215 545
rect 733 503 1215 526
rect 297 491 1215 503
rect 297 478 799 491
rect 297 469 757 478
rect 689 466 757 469
rect 23 401 541 435
rect 23 253 57 401
rect 407 366 541 401
rect 23 210 275 253
rect 23 84 73 210
rect 209 187 275 210
rect 109 17 175 176
rect 689 218 723 466
rect 784 432 833 444
rect 757 424 833 432
rect 757 390 799 424
rect 867 434 917 457
rect 867 390 996 434
rect 1031 394 1126 457
rect 1165 443 1215 491
rect 1250 498 1376 545
rect 1441 532 1508 649
rect 1549 498 1615 549
rect 1250 477 1615 498
rect 1342 464 1615 477
rect 1165 409 1308 443
rect 757 366 833 390
rect 962 360 996 390
rect 1090 375 1126 394
rect 454 184 723 218
rect 962 289 1056 360
rect 1090 309 1240 375
rect 962 218 1009 289
rect 1090 253 1126 309
rect 1274 274 1308 409
rect 873 184 1009 218
rect 1043 222 1126 253
rect 1160 240 1308 274
rect 221 85 287 128
rect 454 119 520 184
rect 873 150 907 184
rect 612 85 682 150
rect 221 51 682 85
rect 718 17 776 150
rect 827 100 907 150
rect 941 17 1007 150
rect 1043 85 1124 222
rect 1160 207 1195 240
rect 1159 119 1195 207
rect 1342 206 1376 464
rect 1229 172 1376 206
rect 1410 218 1465 361
rect 1499 315 1533 464
rect 1567 424 1633 430
rect 1601 390 1633 424
rect 1567 363 1633 390
rect 1677 349 1711 649
rect 1745 343 1801 551
rect 1858 510 2063 576
rect 1849 425 1995 476
rect 1499 252 1663 315
rect 1745 218 1779 343
rect 1849 254 1883 425
rect 2029 391 2063 510
rect 2097 504 2147 649
rect 2189 504 2262 596
rect 1410 184 1779 218
rect 1813 188 1883 254
rect 1917 357 2063 391
rect 2128 424 2194 430
rect 2128 390 2143 424
rect 2177 390 2194 424
rect 2128 364 2194 390
rect 1917 253 1951 357
rect 2228 323 2262 504
rect 2296 420 2362 649
rect 2396 420 2462 596
rect 2417 326 2462 420
rect 2508 364 2574 649
rect 1997 289 2347 323
rect 1997 287 2063 289
rect 2213 253 2279 255
rect 1917 219 2279 253
rect 1229 119 1294 172
rect 1410 116 1620 150
rect 1654 119 1731 184
rect 1410 85 1444 116
rect 1043 51 1444 85
rect 1586 85 1620 116
rect 1813 85 1847 188
rect 1917 154 1951 219
rect 2313 185 2347 289
rect 1486 17 1552 82
rect 1586 51 1847 85
rect 1881 70 1951 154
rect 2039 17 2105 162
rect 2202 151 2347 185
rect 2417 260 2574 326
rect 2202 70 2268 151
rect 2314 17 2381 117
rect 2417 70 2467 260
rect 2513 17 2563 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2688 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 799 390 833 424
rect 1567 390 1601 424
rect 2143 390 2177 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
<< metal1 >>
rect 0 683 2688 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2688 683
rect 0 617 2688 649
rect 787 424 845 430
rect 787 390 799 424
rect 833 421 845 424
rect 1555 424 1613 430
rect 1555 421 1567 424
rect 833 393 1567 421
rect 833 390 845 393
rect 787 384 845 390
rect 1555 390 1567 393
rect 1601 421 1613 424
rect 2131 424 2189 430
rect 2131 421 2143 424
rect 1601 393 2143 421
rect 1601 390 1613 393
rect 1555 384 1613 390
rect 2131 390 2143 393
rect 2177 390 2189 424
rect 2131 384 2189 390
rect 0 17 2688 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2688 17
rect 0 -49 2688 -17
<< labels >>
rlabel locali s 313 162 420 253 6 D
port 1 nsew signal input
rlabel locali s 2614 226 2665 596 6 Q
port 2 nsew signal output
rlabel locali s 2599 70 2665 226 6 Q
port 2 nsew signal output
rlabel metal1 s 2131 421 2189 430 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 2131 384 2189 393 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 1555 421 1613 430 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 1555 384 1613 393 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 787 421 845 430 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 787 393 2189 421 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 787 384 845 393 6 RESET_B
port 3 nsew signal input
rlabel locali s 589 288 655 430 6 SCD
port 4 nsew signal input
rlabel locali s 469 252 545 298 6 SCE
port 5 nsew signal input
rlabel locali s 91 332 359 367 6 SCE
port 5 nsew signal input
rlabel locali s 91 298 545 332 6 SCE
port 5 nsew signal input
rlabel locali s 867 332 928 355 6 CLK
port 6 nsew clock input
rlabel locali s 757 252 928 332 6 CLK
port 6 nsew clock input
rlabel locali s 757 184 839 252 6 CLK
port 6 nsew clock input
rlabel metal1 s 0 -49 2688 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 617 2688 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2688 666
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 231846
string GDS_START 210444
<< end >>
