magic
tech sky130A
magscale 1 2
timestamp 1601050082
<< locali >>
rect 495 378 561 547
rect 21 252 87 310
rect 121 286 309 356
rect 495 344 667 378
rect 357 252 423 310
rect 21 218 423 252
rect 465 236 599 310
rect 633 252 667 344
rect 701 286 839 356
rect 633 218 841 252
rect 509 85 652 116
rect 775 85 841 218
rect 509 51 841 85
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 23 424 73 596
rect 113 458 179 649
rect 213 424 279 596
rect 319 458 369 649
rect 403 581 651 615
rect 403 424 455 581
rect 23 390 455 424
rect 23 364 73 390
rect 595 446 651 581
rect 685 480 751 649
rect 785 446 841 596
rect 595 412 841 446
rect 775 390 841 412
rect 23 17 73 184
rect 109 85 175 184
rect 209 150 741 184
rect 209 119 275 150
rect 686 134 741 150
rect 309 85 375 116
rect 109 51 375 85
rect 409 17 475 116
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel locali s 701 286 839 356 6 A1
port 1 nsew signal input
rlabel locali s 121 286 309 356 6 A2
port 2 nsew signal input
rlabel locali s 357 252 423 310 6 A3
port 3 nsew signal input
rlabel locali s 21 252 87 310 6 A3
port 3 nsew signal input
rlabel locali s 21 218 423 252 6 A3
port 3 nsew signal input
rlabel locali s 465 236 599 310 6 B1
port 4 nsew signal input
rlabel locali s 775 85 841 218 6 Y
port 5 nsew signal output
rlabel locali s 633 252 667 344 6 Y
port 5 nsew signal output
rlabel locali s 633 218 841 252 6 Y
port 5 nsew signal output
rlabel locali s 509 85 652 116 6 Y
port 5 nsew signal output
rlabel locali s 509 51 841 85 6 Y
port 5 nsew signal output
rlabel locali s 495 378 561 547 6 Y
port 5 nsew signal output
rlabel locali s 495 344 667 378 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -49 864 49 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 617 864 715 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3666150
string GDS_START 3657910
<< end >>
