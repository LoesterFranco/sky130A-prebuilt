magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 736 561
rect 17 296 85 493
rect 119 441 201 527
rect 350 443 416 527
rect 17 165 68 296
rect 206 199 272 265
rect 17 90 89 165
rect 142 17 176 165
rect 610 307 676 527
rect 442 215 556 257
rect 590 215 719 257
rect 554 17 588 111
rect 0 -17 736 17
<< obsli1 >>
rect 450 407 515 493
rect 119 373 515 407
rect 119 265 172 373
rect 215 305 340 339
rect 102 199 172 265
rect 306 165 340 305
rect 232 131 340 165
rect 374 291 515 373
rect 232 90 266 131
rect 374 51 408 291
rect 454 147 688 181
rect 454 51 520 147
rect 622 54 688 147
<< metal1 >>
rect 0 496 736 592
rect 0 -48 736 48
<< labels >>
rlabel locali s 590 215 719 257 6 A1
port 1 nsew signal input
rlabel locali s 442 215 556 257 6 A2
port 2 nsew signal input
rlabel locali s 206 199 272 265 6 B1_N
port 3 nsew signal input
rlabel locali s 17 296 85 493 6 X
port 4 nsew signal output
rlabel locali s 17 165 68 296 6 X
port 4 nsew signal output
rlabel locali s 17 90 89 165 6 X
port 4 nsew signal output
rlabel locali s 554 17 588 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 142 17 176 165 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 736 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 736 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 610 307 676 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 350 443 416 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 119 441 201 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 736 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 736 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1373440
string GDS_START 1367336
<< end >>
