magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 3166 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 89 47 119 131
rect 183 47 213 131
rect 381 47 411 131
rect 453 47 483 131
rect 688 47 718 131
rect 794 47 824 131
rect 876 47 906 131
rect 973 47 1003 119
rect 1091 47 1121 119
rect 1197 47 1227 131
rect 1323 47 1353 131
rect 1441 47 1471 175
rect 1525 47 1555 175
rect 1739 47 1769 175
rect 1834 47 1864 119
rect 1962 47 1992 119
rect 2058 47 2088 131
rect 2186 47 2216 131
rect 2292 47 2322 175
rect 2385 47 2415 175
rect 2583 47 2613 131
rect 2690 47 2720 177
rect 2907 47 2937 131
rect 3012 47 3042 177
<< pmoshvt >>
rect 81 363 117 491
rect 175 363 211 491
rect 373 363 409 491
rect 455 363 491 491
rect 680 413 716 497
rect 774 413 810 497
rect 868 413 904 497
rect 975 413 1011 497
rect 1069 413 1105 497
rect 1199 413 1235 497
rect 1315 413 1351 497
rect 1433 329 1469 497
rect 1527 329 1563 497
rect 1674 329 1710 497
rect 1838 413 1874 497
rect 1932 413 1968 497
rect 2060 413 2096 497
rect 2178 413 2214 497
rect 2284 329 2320 497
rect 2366 329 2402 497
rect 2575 301 2611 429
rect 2682 297 2718 497
rect 2899 353 2935 481
rect 3004 297 3040 497
<< ndiff >>
rect 27 119 89 131
rect 27 85 35 119
rect 69 85 89 119
rect 27 47 89 85
rect 119 93 183 131
rect 119 59 129 93
rect 163 59 183 93
rect 119 47 183 59
rect 213 119 265 131
rect 213 85 223 119
rect 257 85 265 119
rect 213 47 265 85
rect 319 111 381 131
rect 319 77 327 111
rect 361 77 381 111
rect 319 47 381 77
rect 411 47 453 131
rect 483 103 552 131
rect 483 69 510 103
rect 544 69 552 103
rect 483 47 552 69
rect 623 111 688 131
rect 623 77 631 111
rect 665 77 688 111
rect 623 47 688 77
rect 718 89 794 131
rect 718 55 740 89
rect 774 55 794 89
rect 718 47 794 55
rect 824 47 876 131
rect 906 119 956 131
rect 1376 131 1441 175
rect 1146 119 1197 131
rect 906 111 973 119
rect 906 77 929 111
rect 963 77 973 111
rect 906 47 973 77
rect 1003 93 1091 119
rect 1003 59 1036 93
rect 1070 59 1091 93
rect 1003 47 1091 59
rect 1121 47 1197 119
rect 1227 89 1323 131
rect 1227 55 1277 89
rect 1311 55 1323 89
rect 1227 47 1323 55
rect 1353 93 1441 131
rect 1353 59 1371 93
rect 1405 59 1441 93
rect 1353 47 1441 59
rect 1471 153 1525 175
rect 1471 119 1481 153
rect 1515 119 1525 153
rect 1471 47 1525 119
rect 1555 127 1612 175
rect 1555 93 1570 127
rect 1604 93 1612 127
rect 1555 47 1612 93
rect 1666 93 1739 175
rect 1666 59 1674 93
rect 1708 59 1739 93
rect 1666 47 1739 59
rect 1769 119 1819 175
rect 2231 131 2292 175
rect 2007 119 2058 131
rect 1769 47 1834 119
rect 1864 93 1962 119
rect 1864 59 1899 93
rect 1933 59 1962 93
rect 1864 47 1962 59
rect 1992 47 2058 119
rect 2088 89 2186 131
rect 2088 55 2110 89
rect 2144 55 2186 89
rect 2088 47 2186 55
rect 2216 93 2292 131
rect 2216 59 2226 93
rect 2260 59 2292 93
rect 2216 47 2292 59
rect 2322 163 2385 175
rect 2322 129 2333 163
rect 2367 129 2385 163
rect 2322 47 2385 129
rect 2415 101 2467 175
rect 2628 161 2690 177
rect 2628 131 2636 161
rect 2415 67 2425 101
rect 2459 67 2467 101
rect 2415 47 2467 67
rect 2521 103 2583 131
rect 2521 69 2529 103
rect 2563 69 2583 103
rect 2521 47 2583 69
rect 2613 127 2636 131
rect 2670 127 2690 161
rect 2613 93 2690 127
rect 2613 59 2636 93
rect 2670 59 2690 93
rect 2613 47 2690 59
rect 2720 127 2791 177
rect 2952 131 3012 177
rect 2720 93 2749 127
rect 2783 93 2791 127
rect 2720 47 2791 93
rect 2845 119 2907 131
rect 2845 85 2863 119
rect 2897 85 2907 119
rect 2845 47 2907 85
rect 2937 93 3012 131
rect 2937 59 2958 93
rect 2992 59 3012 93
rect 2937 47 3012 59
rect 3042 129 3094 177
rect 3042 95 3052 129
rect 3086 95 3094 129
rect 3042 47 3094 95
<< pdiff >>
rect 27 477 81 491
rect 27 443 35 477
rect 69 443 81 477
rect 27 409 81 443
rect 27 375 35 409
rect 69 375 81 409
rect 27 363 81 375
rect 117 461 175 491
rect 117 427 129 461
rect 163 427 175 461
rect 117 363 175 427
rect 211 477 265 491
rect 211 443 223 477
rect 257 443 265 477
rect 211 409 265 443
rect 211 375 223 409
rect 257 375 265 409
rect 211 363 265 375
rect 319 479 373 491
rect 319 445 327 479
rect 361 445 373 479
rect 319 411 373 445
rect 319 377 327 411
rect 361 377 373 411
rect 319 363 373 377
rect 409 363 455 491
rect 491 477 545 491
rect 491 443 503 477
rect 537 443 545 477
rect 491 409 545 443
rect 611 477 680 497
rect 611 443 619 477
rect 653 443 680 477
rect 611 413 680 443
rect 716 477 774 497
rect 716 443 728 477
rect 762 443 774 477
rect 716 413 774 443
rect 810 413 868 497
rect 904 477 975 497
rect 904 443 929 477
rect 963 443 975 477
rect 904 413 975 443
rect 1011 484 1069 497
rect 1011 450 1023 484
rect 1057 450 1069 484
rect 1011 413 1069 450
rect 1105 413 1199 497
rect 1235 475 1315 497
rect 1235 441 1257 475
rect 1291 441 1315 475
rect 1235 413 1315 441
rect 1351 459 1433 497
rect 1351 425 1387 459
rect 1421 425 1433 459
rect 1351 413 1433 425
rect 491 375 503 409
rect 537 375 545 409
rect 491 363 545 375
rect 1369 391 1433 413
rect 1369 357 1387 391
rect 1421 357 1433 391
rect 1369 329 1433 357
rect 1469 329 1527 497
rect 1563 485 1674 497
rect 1563 451 1581 485
rect 1615 451 1674 485
rect 1563 417 1674 451
rect 1563 383 1581 417
rect 1615 383 1674 417
rect 1563 329 1674 383
rect 1710 413 1838 497
rect 1874 484 1932 497
rect 1874 450 1886 484
rect 1920 450 1932 484
rect 1874 413 1932 450
rect 1968 413 2060 497
rect 2096 485 2178 497
rect 2096 451 2120 485
rect 2154 451 2178 485
rect 2096 413 2178 451
rect 2214 459 2284 497
rect 2214 425 2238 459
rect 2272 425 2284 459
rect 2214 413 2284 425
rect 1710 329 1774 413
rect 2231 329 2284 413
rect 2320 329 2366 497
rect 2402 485 2456 497
rect 2402 451 2414 485
rect 2448 451 2456 485
rect 2628 485 2682 497
rect 2402 329 2456 451
rect 2628 451 2636 485
rect 2670 451 2682 485
rect 2628 429 2682 451
rect 2521 349 2575 429
rect 2521 315 2529 349
rect 2563 315 2575 349
rect 2521 301 2575 315
rect 2611 301 2682 429
rect 2630 297 2682 301
rect 2718 448 2791 497
rect 2952 481 3004 497
rect 2718 414 2749 448
rect 2783 414 2791 448
rect 2718 380 2791 414
rect 2718 346 2749 380
rect 2783 346 2791 380
rect 2845 467 2899 481
rect 2845 433 2853 467
rect 2887 433 2899 467
rect 2845 399 2899 433
rect 2845 365 2853 399
rect 2887 365 2899 399
rect 2845 353 2899 365
rect 2935 473 3004 481
rect 2935 439 2958 473
rect 2992 439 3004 473
rect 2935 405 3004 439
rect 2935 371 2958 405
rect 2992 371 3004 405
rect 2935 353 3004 371
rect 2718 297 2791 346
rect 2952 297 3004 353
rect 3040 449 3094 497
rect 3040 415 3052 449
rect 3086 415 3094 449
rect 3040 381 3094 415
rect 3040 347 3052 381
rect 3086 347 3094 381
rect 3040 297 3094 347
<< ndiffc >>
rect 35 85 69 119
rect 129 59 163 93
rect 223 85 257 119
rect 327 77 361 111
rect 510 69 544 103
rect 631 77 665 111
rect 740 55 774 89
rect 929 77 963 111
rect 1036 59 1070 93
rect 1277 55 1311 89
rect 1371 59 1405 93
rect 1481 119 1515 153
rect 1570 93 1604 127
rect 1674 59 1708 93
rect 1899 59 1933 93
rect 2110 55 2144 89
rect 2226 59 2260 93
rect 2333 129 2367 163
rect 2425 67 2459 101
rect 2529 69 2563 103
rect 2636 127 2670 161
rect 2636 59 2670 93
rect 2749 93 2783 127
rect 2863 85 2897 119
rect 2958 59 2992 93
rect 3052 95 3086 129
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 129 427 163 461
rect 223 443 257 477
rect 223 375 257 409
rect 327 445 361 479
rect 327 377 361 411
rect 503 443 537 477
rect 619 443 653 477
rect 728 443 762 477
rect 929 443 963 477
rect 1023 450 1057 484
rect 1257 441 1291 475
rect 1387 425 1421 459
rect 503 375 537 409
rect 1387 357 1421 391
rect 1581 451 1615 485
rect 1581 383 1615 417
rect 1886 450 1920 484
rect 2120 451 2154 485
rect 2238 425 2272 459
rect 2414 451 2448 485
rect 2636 451 2670 485
rect 2529 315 2563 349
rect 2749 414 2783 448
rect 2749 346 2783 380
rect 2853 433 2887 467
rect 2853 365 2887 399
rect 2958 439 2992 473
rect 2958 371 2992 405
rect 3052 415 3086 449
rect 3052 347 3086 381
<< poly >>
rect 81 491 117 517
rect 175 491 211 517
rect 373 491 409 517
rect 455 491 491 517
rect 680 497 716 523
rect 774 497 810 523
rect 868 497 904 523
rect 975 497 1011 523
rect 1069 497 1105 523
rect 1199 497 1235 523
rect 1315 497 1351 523
rect 1433 497 1469 523
rect 1527 497 1563 523
rect 1674 497 1710 523
rect 1838 497 1874 523
rect 1932 497 1968 523
rect 2060 497 2096 523
rect 2178 497 2214 523
rect 2284 497 2320 523
rect 2366 497 2402 523
rect 2682 497 2718 523
rect 680 398 716 413
rect 774 398 810 413
rect 868 398 904 413
rect 975 398 1011 413
rect 1069 398 1105 413
rect 1199 398 1235 413
rect 1315 398 1351 413
rect 678 397 718 398
rect 772 397 812 398
rect 579 365 636 381
rect 81 348 117 363
rect 175 348 211 363
rect 373 348 409 363
rect 455 348 491 363
rect 45 318 119 348
rect 45 280 75 318
rect 21 264 75 280
rect 173 274 213 348
rect 371 331 411 348
rect 21 230 31 264
rect 65 230 75 264
rect 21 214 75 230
rect 127 264 213 274
rect 309 315 411 331
rect 453 345 493 348
rect 579 345 592 365
rect 453 331 592 345
rect 626 331 636 365
rect 453 315 636 331
rect 678 367 812 397
rect 309 281 319 315
rect 353 281 411 315
rect 309 265 411 281
rect 127 230 143 264
rect 177 230 213 264
rect 127 220 213 230
rect 45 176 75 214
rect 45 146 119 176
rect 89 131 119 146
rect 183 131 213 220
rect 381 131 411 265
rect 453 203 517 219
rect 453 169 463 203
rect 497 177 517 203
rect 678 177 718 367
rect 866 325 906 398
rect 815 315 906 325
rect 815 281 831 315
rect 865 281 906 315
rect 815 271 906 281
rect 497 169 718 177
rect 453 147 718 169
rect 760 203 824 219
rect 760 169 770 203
rect 804 169 824 203
rect 760 153 824 169
rect 453 131 483 147
rect 688 131 718 147
rect 794 131 824 153
rect 876 131 906 271
rect 973 279 1013 398
rect 1067 375 1107 398
rect 1197 381 1237 398
rect 1055 365 1131 375
rect 1055 331 1071 365
rect 1105 331 1131 365
rect 1055 321 1131 331
rect 1197 365 1271 381
rect 1197 331 1217 365
rect 1251 331 1271 365
rect 1197 315 1271 331
rect 973 249 1131 279
rect 1091 219 1131 249
rect 973 191 1049 207
rect 973 157 997 191
rect 1031 157 1049 191
rect 973 141 1049 157
rect 1091 203 1155 219
rect 1091 169 1111 203
rect 1145 169 1155 203
rect 1091 153 1155 169
rect 973 119 1003 141
rect 1091 119 1121 153
rect 1197 131 1227 315
rect 1313 229 1353 398
rect 1838 398 1874 413
rect 1932 398 1968 413
rect 2060 398 2096 413
rect 2178 398 2214 413
rect 1836 381 1876 398
rect 1812 365 1876 381
rect 1930 375 1970 398
rect 2058 381 2098 398
rect 1812 331 1822 365
rect 1856 331 1876 365
rect 1433 314 1469 329
rect 1527 314 1563 329
rect 1674 314 1710 329
rect 1812 315 1876 331
rect 1918 365 1994 375
rect 1918 331 1934 365
rect 1968 331 1994 365
rect 1918 321 1994 331
rect 2058 365 2134 381
rect 2058 331 2080 365
rect 2114 331 2134 365
rect 1431 297 1471 314
rect 1395 281 1471 297
rect 1395 247 1405 281
rect 1439 247 1471 281
rect 1395 231 1471 247
rect 1283 213 1353 229
rect 1283 179 1293 213
rect 1327 179 1353 213
rect 1283 163 1353 179
rect 1441 175 1471 231
rect 1525 297 1565 314
rect 1525 281 1621 297
rect 1525 247 1577 281
rect 1611 247 1621 281
rect 1525 231 1621 247
rect 1672 263 1712 314
rect 1836 279 1876 315
rect 2058 315 2134 331
rect 1672 247 1769 263
rect 1836 249 1992 279
rect 1525 175 1555 231
rect 1672 213 1715 247
rect 1749 213 1769 247
rect 1672 197 1769 213
rect 1739 175 1769 197
rect 1834 191 1911 207
rect 1323 131 1353 163
rect 1834 157 1857 191
rect 1891 157 1911 191
rect 1834 141 1911 157
rect 1834 119 1864 141
rect 1962 119 1992 249
rect 2058 131 2088 315
rect 2176 229 2216 398
rect 2575 429 2611 455
rect 2284 314 2320 329
rect 2366 314 2402 329
rect 2282 281 2322 314
rect 2139 213 2216 229
rect 2258 265 2322 281
rect 2364 297 2404 314
rect 2364 281 2470 297
rect 2575 286 2611 301
rect 2899 481 2935 507
rect 3004 497 3040 523
rect 2899 338 2935 353
rect 2897 337 2937 338
rect 2872 307 2937 337
rect 2364 267 2426 281
rect 2258 231 2268 265
rect 2302 231 2322 265
rect 2258 215 2322 231
rect 2139 179 2149 213
rect 2183 179 2216 213
rect 2139 163 2216 179
rect 2292 175 2322 215
rect 2385 247 2426 267
rect 2460 247 2470 281
rect 2573 269 2613 286
rect 2682 282 2718 297
rect 2385 231 2470 247
rect 2523 253 2613 269
rect 2680 265 2720 282
rect 2385 175 2415 231
rect 2523 219 2533 253
rect 2567 219 2613 253
rect 2523 203 2613 219
rect 2186 131 2216 163
rect 2583 131 2613 203
rect 2661 259 2720 265
rect 2872 259 2902 307
rect 3004 282 3040 297
rect 3002 265 3042 282
rect 2661 249 2902 259
rect 2661 215 2671 249
rect 2705 215 2902 249
rect 2661 205 2902 215
rect 2661 199 2720 205
rect 2690 177 2720 199
rect 2872 176 2902 205
rect 2974 249 3042 265
rect 2974 215 2984 249
rect 3018 215 3042 249
rect 2974 199 3042 215
rect 3012 177 3042 199
rect 2872 146 2937 176
rect 2907 131 2937 146
rect 89 21 119 47
rect 183 21 213 47
rect 381 21 411 47
rect 453 21 483 47
rect 688 21 718 47
rect 794 21 824 47
rect 876 21 906 47
rect 973 21 1003 47
rect 1091 21 1121 47
rect 1197 21 1227 47
rect 1323 21 1353 47
rect 1441 21 1471 47
rect 1525 21 1555 47
rect 1739 21 1769 47
rect 1834 21 1864 47
rect 1962 21 1992 47
rect 2058 21 2088 47
rect 2186 21 2216 47
rect 2292 21 2322 47
rect 2385 21 2415 47
rect 2583 21 2613 47
rect 2690 21 2720 47
rect 2907 21 2937 47
rect 3012 21 3042 47
<< polycont >>
rect 31 230 65 264
rect 592 331 626 365
rect 319 281 353 315
rect 143 230 177 264
rect 463 169 497 203
rect 831 281 865 315
rect 770 169 804 203
rect 1071 331 1105 365
rect 1217 331 1251 365
rect 997 157 1031 191
rect 1111 169 1145 203
rect 1822 331 1856 365
rect 1934 331 1968 365
rect 2080 331 2114 365
rect 1405 247 1439 281
rect 1293 179 1327 213
rect 1577 247 1611 281
rect 1715 213 1749 247
rect 1857 157 1891 191
rect 2268 231 2302 265
rect 2149 179 2183 213
rect 2426 247 2460 281
rect 2533 219 2567 253
rect 2671 215 2705 249
rect 2984 215 3018 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3128 561
rect 34 477 69 493
rect 34 443 35 477
rect 34 409 69 443
rect 103 461 179 527
rect 103 427 129 461
rect 163 427 179 461
rect 223 477 264 493
rect 257 443 264 477
rect 34 375 35 409
rect 223 409 264 443
rect 69 391 177 393
rect 69 375 131 391
rect 34 359 131 375
rect 165 357 177 391
rect 17 264 87 325
rect 17 230 31 264
rect 65 230 87 264
rect 17 195 87 230
rect 131 264 177 357
rect 131 230 143 264
rect 131 161 177 230
rect 34 127 177 161
rect 257 375 264 409
rect 311 479 377 527
rect 311 445 327 479
rect 361 445 377 479
rect 619 477 653 493
rect 311 411 377 445
rect 311 377 327 411
rect 361 377 377 411
rect 477 443 503 477
rect 537 443 553 477
rect 477 409 553 443
rect 477 375 503 409
rect 537 375 553 409
rect 702 477 778 527
rect 702 443 728 477
rect 762 443 778 477
rect 929 477 963 493
rect 619 381 653 443
rect 223 187 264 375
rect 298 315 353 337
rect 298 281 319 315
rect 298 205 353 281
rect 223 153 230 187
rect 34 119 69 127
rect 34 85 35 119
rect 223 119 264 153
rect 387 203 451 339
rect 510 273 553 375
rect 589 365 653 381
rect 589 331 592 365
rect 626 349 653 365
rect 626 331 779 349
rect 589 315 779 331
rect 510 255 655 273
rect 510 237 621 255
rect 557 221 621 237
rect 557 215 655 221
rect 745 219 779 315
rect 831 315 895 475
rect 865 281 895 315
rect 831 265 895 281
rect 1007 450 1023 484
rect 1057 450 1183 484
rect 929 255 963 443
rect 387 169 463 203
rect 497 169 521 203
rect 387 153 521 169
rect 387 152 451 153
rect 34 69 69 85
rect 103 59 129 93
rect 163 59 179 93
rect 257 85 264 119
rect 223 69 264 85
rect 311 111 361 127
rect 311 77 327 111
rect 103 17 179 59
rect 311 17 361 77
rect 395 69 451 152
rect 557 119 591 215
rect 745 203 814 219
rect 745 169 770 203
rect 804 169 814 203
rect 745 159 814 169
rect 510 103 591 119
rect 544 69 591 103
rect 510 53 591 69
rect 625 153 814 159
rect 625 125 779 153
rect 625 111 665 125
rect 625 77 631 111
rect 929 111 963 221
rect 997 357 1029 391
rect 1063 365 1115 391
rect 1063 357 1071 365
rect 997 331 1071 357
rect 1105 331 1115 365
rect 997 315 1115 331
rect 997 191 1049 315
rect 1149 281 1183 450
rect 1241 475 1317 527
rect 1565 485 1631 527
rect 1241 441 1257 475
rect 1291 441 1317 475
rect 1387 459 1421 475
rect 1387 407 1421 425
rect 1565 451 1581 485
rect 1615 451 1631 485
rect 2104 485 2180 527
rect 1565 417 1631 451
rect 1860 450 1886 484
rect 1920 450 2046 484
rect 2104 451 2120 485
rect 2154 451 2180 485
rect 2388 485 2686 527
rect 2238 459 2272 475
rect 1217 391 1517 407
rect 1217 365 1387 391
rect 1251 357 1387 365
rect 1421 357 1517 391
rect 1565 383 1581 417
rect 1615 383 1631 417
rect 1822 391 1869 397
rect 1251 331 1277 357
rect 1217 315 1277 331
rect 1389 281 1439 297
rect 1149 247 1405 281
rect 1149 239 1243 247
rect 1031 157 1049 191
rect 997 141 1049 157
rect 1085 169 1111 203
rect 1145 187 1165 203
rect 1085 153 1131 169
rect 1085 129 1165 153
rect 625 61 665 77
rect 724 55 740 89
rect 774 55 790 89
rect 1199 93 1243 239
rect 1395 231 1439 247
rect 1483 213 1517 357
rect 1822 365 1835 391
rect 1856 331 1869 357
rect 1561 323 1782 331
rect 1561 289 1743 323
rect 1777 289 1782 323
rect 1822 315 1869 331
rect 1927 365 1978 381
rect 1927 331 1934 365
rect 1968 331 1978 365
rect 1561 283 1782 289
rect 1561 281 1627 283
rect 1561 247 1577 281
rect 1611 247 1627 281
rect 1927 261 1978 331
rect 1834 255 1978 261
rect 1689 213 1715 247
rect 1749 213 1775 247
rect 1277 179 1293 213
rect 1327 187 1359 213
rect 1277 153 1317 179
rect 1351 153 1359 187
rect 1483 179 1775 213
rect 1834 221 1835 255
rect 1869 225 1978 255
rect 2012 281 2046 450
rect 2388 451 2414 485
rect 2448 451 2636 485
rect 2670 451 2686 485
rect 2238 417 2272 425
rect 2743 448 2819 493
rect 2080 383 2686 417
rect 2080 365 2140 383
rect 2114 331 2140 365
rect 2080 315 2140 331
rect 2012 265 2302 281
rect 2012 247 2268 265
rect 1869 221 1902 225
rect 1834 191 1902 221
rect 1483 153 1531 179
rect 1277 147 1359 153
rect 1455 119 1481 153
rect 1515 119 1531 153
rect 1834 157 1857 191
rect 1891 157 1902 191
rect 1570 127 1609 143
rect 1834 141 1902 157
rect 929 61 963 77
rect 724 17 790 55
rect 1020 59 1036 93
rect 1070 59 1243 93
rect 1020 53 1243 59
rect 1277 89 1311 105
rect 1604 93 1609 127
rect 2012 93 2046 247
rect 2258 231 2268 247
rect 2258 215 2302 231
rect 2131 187 2149 213
rect 2131 153 2143 187
rect 2183 179 2216 213
rect 2177 153 2216 179
rect 2346 163 2383 383
rect 2131 147 2216 153
rect 2307 129 2333 163
rect 2367 129 2383 163
rect 2426 323 2529 349
rect 2426 289 2433 323
rect 2467 315 2529 323
rect 2563 315 2581 349
rect 2467 289 2469 315
rect 2426 281 2469 289
rect 2460 247 2469 281
rect 2652 265 2686 383
rect 2743 414 2749 448
rect 2783 414 2819 448
rect 2743 380 2819 414
rect 2743 346 2749 380
rect 2783 346 2819 380
rect 2743 326 2819 346
rect 2853 467 2904 483
rect 2887 433 2904 467
rect 2853 399 2904 433
rect 2887 365 2904 399
rect 2853 345 2904 365
rect 2949 473 3008 527
rect 2949 439 2958 473
rect 2992 439 3008 473
rect 2949 405 3008 439
rect 2949 371 2958 405
rect 2992 371 3008 405
rect 2949 353 3008 371
rect 3052 449 3109 493
rect 3086 415 3109 449
rect 3052 381 3109 415
rect 2764 304 2819 326
rect 2426 185 2469 247
rect 2503 253 2618 265
rect 2503 219 2533 253
rect 2567 219 2618 253
rect 2652 249 2705 265
rect 2652 215 2671 249
rect 2652 199 2705 215
rect 2426 151 2563 185
rect 1277 17 1311 55
rect 1355 59 1371 93
rect 1405 85 1421 93
rect 1570 85 1609 93
rect 1405 59 1609 85
rect 1355 51 1609 59
rect 1658 59 1674 93
rect 1708 59 1735 93
rect 1658 17 1735 59
rect 1883 59 1899 93
rect 1933 59 2046 93
rect 1883 53 2046 59
rect 2082 89 2144 105
rect 2425 101 2460 117
rect 2082 55 2110 89
rect 2082 17 2144 55
rect 2196 59 2226 93
rect 2260 85 2276 93
rect 2260 67 2425 85
rect 2459 67 2460 101
rect 2260 59 2460 67
rect 2196 51 2460 59
rect 2523 103 2563 151
rect 2523 69 2529 103
rect 2523 53 2563 69
rect 2620 127 2636 161
rect 2670 127 2686 161
rect 2764 143 2823 304
rect 2620 93 2686 127
rect 2620 59 2636 93
rect 2670 59 2686 93
rect 2620 17 2686 59
rect 2743 127 2823 143
rect 2743 93 2749 127
rect 2783 93 2823 127
rect 2743 51 2823 93
rect 2863 265 2904 345
rect 3086 347 3109 381
rect 3052 321 3109 347
rect 2863 249 3018 265
rect 2863 215 2984 249
rect 2863 199 3018 215
rect 2863 119 2904 199
rect 3062 165 3109 321
rect 2897 85 2904 119
rect 3052 129 3109 165
rect 2863 51 2904 85
rect 2950 93 3008 109
rect 2950 59 2958 93
rect 2992 59 3008 93
rect 2950 17 3008 59
rect 3086 95 3109 129
rect 3052 51 3109 95
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3128 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 2881 527 2915 561
rect 2973 527 3007 561
rect 3065 527 3099 561
rect 131 357 165 391
rect 230 153 264 187
rect 621 221 655 255
rect 929 221 963 255
rect 1029 357 1063 391
rect 1131 169 1145 187
rect 1145 169 1165 187
rect 1131 153 1165 169
rect 1835 365 1869 391
rect 1835 357 1856 365
rect 1856 357 1869 365
rect 1743 289 1777 323
rect 1317 179 1327 187
rect 1327 179 1351 187
rect 1317 153 1351 179
rect 1835 221 1869 255
rect 2143 179 2149 187
rect 2149 179 2177 187
rect 2143 153 2177 179
rect 2433 289 2467 323
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
rect 2881 -17 2915 17
rect 2973 -17 3007 17
rect 3065 -17 3099 17
<< metal1 >>
rect 0 561 3128 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3128 561
rect 0 496 3128 527
rect 119 391 177 397
rect 119 357 131 391
rect 165 388 177 391
rect 1017 391 1075 397
rect 1017 388 1029 391
rect 165 360 1029 388
rect 165 357 177 360
rect 119 351 177 357
rect 1017 357 1029 360
rect 1063 388 1075 391
rect 1823 391 1881 397
rect 1823 388 1835 391
rect 1063 360 1835 388
rect 1063 357 1075 360
rect 1017 351 1075 357
rect 1823 357 1835 360
rect 1869 357 1881 391
rect 1823 351 1881 357
rect 1731 323 1789 329
rect 1731 289 1743 323
rect 1777 320 1789 323
rect 2421 323 2479 329
rect 2421 320 2433 323
rect 1777 292 2433 320
rect 1777 289 1789 292
rect 1731 283 1789 289
rect 2421 289 2433 292
rect 2467 289 2479 323
rect 2421 283 2479 289
rect 609 255 667 261
rect 609 221 621 255
rect 655 252 667 255
rect 917 255 975 261
rect 917 252 929 255
rect 655 224 929 252
rect 655 221 667 224
rect 609 215 667 221
rect 917 221 929 224
rect 963 221 975 255
rect 1823 255 1881 261
rect 1823 252 1835 255
rect 917 215 975 221
rect 1134 224 1835 252
rect 1134 193 1177 224
rect 1823 221 1835 224
rect 1869 221 1881 255
rect 1823 215 1881 221
rect 218 187 276 193
rect 218 153 230 187
rect 264 184 276 187
rect 1119 187 1177 193
rect 1119 184 1131 187
rect 264 156 1131 184
rect 264 153 276 156
rect 218 147 276 153
rect 1119 153 1131 156
rect 1165 153 1177 187
rect 1119 147 1177 153
rect 1305 187 1363 193
rect 1305 153 1317 187
rect 1351 184 1363 187
rect 2131 187 2189 193
rect 2131 184 2143 187
rect 1351 156 2143 184
rect 1351 153 1363 156
rect 1305 147 1363 153
rect 2131 153 2143 156
rect 2177 153 2189 187
rect 2131 147 2189 153
rect 0 17 3128 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3128 17
rect 0 -48 3128 -17
<< labels >>
flabel corelocali s 305 289 339 323 0 FreeSans 200 0 0 0 SCD
port 4 nsew
flabel corelocali s 305 221 339 255 0 FreeSans 200 0 0 0 SCD
port 4 nsew
flabel corelocali s 397 289 431 323 0 FreeSans 200 0 0 0 SCE
port 5 nsew
flabel corelocali s 397 221 431 255 0 FreeSans 200 0 0 0 SCE
port 5 nsew
flabel corelocali s 397 85 431 119 0 FreeSans 400 0 0 0 SCE
port 5 nsew
flabel corelocali s 2513 221 2547 255 0 FreeSans 200 0 0 0 RESET_B
port 3 nsew
flabel corelocali s 29 -17 63 17 3 FreeSans 400 0 0 0 VGND
port 7 nsew
flabel corelocali s 29 221 63 255 0 FreeSans 400 0 0 0 CLK
port 1 nsew
flabel corelocali s 29 289 63 323 0 FreeSans 400 0 0 0 CLK
port 1 nsew
flabel corelocali s 3065 85 3099 119 0 FreeSans 400 0 0 0 Q
port 11 nsew
flabel corelocali s 3065 357 3099 391 0 FreeSans 400 0 0 0 Q
port 11 nsew
flabel corelocali s 3065 425 3099 459 0 FreeSans 400 0 0 0 Q
port 11 nsew
flabel corelocali s 29 527 63 561 3 FreeSans 400 0 0 0 VPWR
port 10 nsew
flabel corelocali s 857 289 891 323 0 FreeSans 200 0 0 0 D
port 2 nsew
flabel corelocali s 857 425 891 459 0 FreeSans 200 0 0 0 D
port 2 nsew
flabel corelocali s 2789 221 2823 255 0 FreeSans 400 0 0 0 Q_N
port 12 nsew
flabel corelocali s 2789 153 2823 187 0 FreeSans 400 0 0 0 Q_N
port 12 nsew
flabel corelocali s 2789 85 2823 119 0 FreeSans 400 0 0 0 Q_N
port 12 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 7 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 10 nsew
flabel metal1 s 1317 153 1351 187 0 FreeSans 200 0 0 0 SET_B
port 6 nsew
flabel nbase s 29 527 63 561 3 FreeSans 400 0 0 0 VPB
port 9 nsew
flabel nbase s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
port 9 nsew
flabel pwell s 29 -17 63 17 3 FreeSans 400 0 0 0 VNB
port 8 nsew
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
port 8 nsew
rlabel comment s 0 0 0 0 4 sdfbbp_1
<< properties >>
string FIXED_BBOX 0 0 3128 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 146246
string GDS_START 122988
<< end >>
