magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 1418 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 89 47 119 177
rect 277 47 307 177
rect 371 47 401 177
rect 475 47 505 177
rect 559 47 589 177
rect 653 47 683 177
rect 747 47 777 177
rect 841 47 871 177
rect 935 47 965 177
rect 1029 47 1059 177
rect 1123 47 1153 177
rect 1227 47 1257 177
<< pmoshvt >>
rect 81 297 117 497
rect 279 297 315 497
rect 373 297 409 497
rect 467 297 503 497
rect 561 297 597 497
rect 655 297 691 497
rect 749 297 785 497
rect 843 297 879 497
rect 937 297 973 497
rect 1031 297 1067 497
rect 1125 297 1161 497
rect 1219 297 1255 497
<< ndiff >>
rect 27 165 89 177
rect 27 131 35 165
rect 69 131 89 165
rect 27 97 89 131
rect 27 63 35 97
rect 69 63 89 97
rect 27 47 89 63
rect 119 165 171 177
rect 119 131 129 165
rect 163 131 171 165
rect 119 97 171 131
rect 119 63 129 97
rect 163 63 171 97
rect 119 47 171 63
rect 225 165 277 177
rect 225 131 233 165
rect 267 131 277 165
rect 225 97 277 131
rect 225 63 233 97
rect 267 63 277 97
rect 225 47 277 63
rect 307 97 371 177
rect 307 63 327 97
rect 361 63 371 97
rect 307 47 371 63
rect 401 165 475 177
rect 401 131 421 165
rect 455 131 475 165
rect 401 97 475 131
rect 401 63 421 97
rect 455 63 475 97
rect 401 47 475 63
rect 505 97 559 177
rect 505 63 515 97
rect 549 63 559 97
rect 505 47 559 63
rect 589 165 653 177
rect 589 131 609 165
rect 643 131 653 165
rect 589 97 653 131
rect 589 63 609 97
rect 643 63 653 97
rect 589 47 653 63
rect 683 97 747 177
rect 683 63 703 97
rect 737 63 747 97
rect 683 47 747 63
rect 777 165 841 177
rect 777 131 797 165
rect 831 131 841 165
rect 777 97 841 131
rect 777 63 797 97
rect 831 63 841 97
rect 777 47 841 63
rect 871 97 935 177
rect 871 63 891 97
rect 925 63 935 97
rect 871 47 935 63
rect 965 165 1029 177
rect 965 131 985 165
rect 1019 131 1029 165
rect 965 97 1029 131
rect 965 63 985 97
rect 1019 63 1029 97
rect 965 47 1029 63
rect 1059 97 1123 177
rect 1059 63 1079 97
rect 1113 63 1123 97
rect 1059 47 1123 63
rect 1153 165 1227 177
rect 1153 131 1173 165
rect 1207 131 1227 165
rect 1153 97 1227 131
rect 1153 63 1173 97
rect 1207 63 1227 97
rect 1153 47 1227 63
rect 1257 97 1309 177
rect 1257 63 1267 97
rect 1301 63 1309 97
rect 1257 47 1309 63
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 479 171 497
rect 117 445 129 479
rect 163 445 171 479
rect 117 411 171 445
rect 117 377 129 411
rect 163 377 171 411
rect 117 343 171 377
rect 117 309 129 343
rect 163 309 171 343
rect 117 297 171 309
rect 225 479 279 497
rect 225 445 233 479
rect 267 445 279 479
rect 225 411 279 445
rect 225 377 233 411
rect 267 377 279 411
rect 225 343 279 377
rect 225 309 233 343
rect 267 309 279 343
rect 225 297 279 309
rect 315 485 373 497
rect 315 451 327 485
rect 361 451 373 485
rect 315 417 373 451
rect 315 383 327 417
rect 361 383 373 417
rect 315 297 373 383
rect 409 479 467 497
rect 409 445 421 479
rect 455 445 467 479
rect 409 411 467 445
rect 409 377 421 411
rect 455 377 467 411
rect 409 343 467 377
rect 409 309 421 343
rect 455 309 467 343
rect 409 297 467 309
rect 503 485 561 497
rect 503 451 515 485
rect 549 451 561 485
rect 503 417 561 451
rect 503 383 515 417
rect 549 383 561 417
rect 503 297 561 383
rect 597 479 655 497
rect 597 445 609 479
rect 643 445 655 479
rect 597 411 655 445
rect 597 377 609 411
rect 643 377 655 411
rect 597 343 655 377
rect 597 309 609 343
rect 643 309 655 343
rect 597 297 655 309
rect 691 485 749 497
rect 691 451 703 485
rect 737 451 749 485
rect 691 417 749 451
rect 691 383 703 417
rect 737 383 749 417
rect 691 297 749 383
rect 785 479 843 497
rect 785 445 797 479
rect 831 445 843 479
rect 785 411 843 445
rect 785 377 797 411
rect 831 377 843 411
rect 785 343 843 377
rect 785 309 797 343
rect 831 309 843 343
rect 785 297 843 309
rect 879 485 937 497
rect 879 451 891 485
rect 925 451 937 485
rect 879 417 937 451
rect 879 383 891 417
rect 925 383 937 417
rect 879 297 937 383
rect 973 479 1031 497
rect 973 445 985 479
rect 1019 445 1031 479
rect 973 411 1031 445
rect 973 377 985 411
rect 1019 377 1031 411
rect 973 343 1031 377
rect 973 309 985 343
rect 1019 309 1031 343
rect 973 297 1031 309
rect 1067 485 1125 497
rect 1067 451 1079 485
rect 1113 451 1125 485
rect 1067 417 1125 451
rect 1067 383 1079 417
rect 1113 383 1125 417
rect 1067 297 1125 383
rect 1161 479 1219 497
rect 1161 445 1173 479
rect 1207 445 1219 479
rect 1161 411 1219 445
rect 1161 377 1173 411
rect 1207 377 1219 411
rect 1161 343 1219 377
rect 1161 309 1173 343
rect 1207 309 1219 343
rect 1161 297 1219 309
rect 1255 485 1309 497
rect 1255 451 1267 485
rect 1301 451 1309 485
rect 1255 417 1309 451
rect 1255 383 1267 417
rect 1301 383 1309 417
rect 1255 297 1309 383
<< ndiffc >>
rect 35 131 69 165
rect 35 63 69 97
rect 129 131 163 165
rect 129 63 163 97
rect 233 131 267 165
rect 233 63 267 97
rect 327 63 361 97
rect 421 131 455 165
rect 421 63 455 97
rect 515 63 549 97
rect 609 131 643 165
rect 609 63 643 97
rect 703 63 737 97
rect 797 131 831 165
rect 797 63 831 97
rect 891 63 925 97
rect 985 131 1019 165
rect 985 63 1019 97
rect 1079 63 1113 97
rect 1173 131 1207 165
rect 1173 63 1207 97
rect 1267 63 1301 97
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 445 163 479
rect 129 377 163 411
rect 129 309 163 343
rect 233 445 267 479
rect 233 377 267 411
rect 233 309 267 343
rect 327 451 361 485
rect 327 383 361 417
rect 421 445 455 479
rect 421 377 455 411
rect 421 309 455 343
rect 515 451 549 485
rect 515 383 549 417
rect 609 445 643 479
rect 609 377 643 411
rect 609 309 643 343
rect 703 451 737 485
rect 703 383 737 417
rect 797 445 831 479
rect 797 377 831 411
rect 797 309 831 343
rect 891 451 925 485
rect 891 383 925 417
rect 985 445 1019 479
rect 985 377 1019 411
rect 985 309 1019 343
rect 1079 451 1113 485
rect 1079 383 1113 417
rect 1173 445 1207 479
rect 1173 377 1207 411
rect 1173 309 1207 343
rect 1267 451 1301 485
rect 1267 383 1301 417
<< poly >>
rect 81 497 117 523
rect 279 497 315 523
rect 373 497 409 523
rect 467 497 503 523
rect 561 497 597 523
rect 655 497 691 523
rect 749 497 785 523
rect 843 497 879 523
rect 937 497 973 523
rect 1031 497 1067 523
rect 1125 497 1161 523
rect 1219 497 1255 523
rect 81 282 117 297
rect 279 282 315 297
rect 373 282 409 297
rect 467 282 503 297
rect 561 282 597 297
rect 655 282 691 297
rect 749 282 785 297
rect 843 282 879 297
rect 937 282 973 297
rect 1031 282 1067 297
rect 1125 282 1161 297
rect 1219 282 1255 297
rect 79 265 119 282
rect 21 249 119 265
rect 21 215 38 249
rect 72 215 119 249
rect 21 199 119 215
rect 89 177 119 199
rect 277 259 317 282
rect 371 259 411 282
rect 465 259 505 282
rect 277 249 505 259
rect 277 215 327 249
rect 361 215 395 249
rect 429 215 505 249
rect 277 205 505 215
rect 277 177 307 205
rect 371 177 401 205
rect 475 177 505 205
rect 559 259 599 282
rect 653 259 693 282
rect 747 259 787 282
rect 841 259 881 282
rect 935 259 975 282
rect 1029 259 1069 282
rect 1123 259 1163 282
rect 1217 259 1257 282
rect 559 249 1257 259
rect 559 215 583 249
rect 617 215 661 249
rect 695 215 739 249
rect 773 215 817 249
rect 851 215 895 249
rect 929 215 963 249
rect 997 215 1041 249
rect 1075 215 1119 249
rect 1153 215 1197 249
rect 1231 215 1257 249
rect 559 205 1257 215
rect 559 177 589 205
rect 653 177 683 205
rect 747 177 777 205
rect 841 177 871 205
rect 935 177 965 205
rect 1029 177 1059 205
rect 1123 177 1153 205
rect 1227 177 1257 205
rect 89 21 119 47
rect 277 21 307 47
rect 371 21 401 47
rect 475 21 505 47
rect 559 21 589 47
rect 653 21 683 47
rect 747 21 777 47
rect 841 21 871 47
rect 935 21 965 47
rect 1029 21 1059 47
rect 1123 21 1153 47
rect 1227 21 1257 47
<< polycont >>
rect 38 215 72 249
rect 327 215 361 249
rect 395 215 429 249
rect 583 215 617 249
rect 661 215 695 249
rect 739 215 773 249
rect 817 215 851 249
rect 895 215 929 249
rect 963 215 997 249
rect 1041 215 1075 249
rect 1119 215 1153 249
rect 1197 215 1231 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 35 485 69 527
rect 35 417 69 451
rect 35 349 69 383
rect 35 289 69 315
rect 103 479 179 493
rect 103 445 129 479
rect 163 445 179 479
rect 103 411 179 445
rect 103 377 129 411
rect 163 377 179 411
rect 103 343 179 377
rect 103 309 129 343
rect 163 309 179 343
rect 145 255 179 309
rect 217 479 283 493
rect 217 445 233 479
rect 267 445 283 479
rect 217 411 283 445
rect 217 377 233 411
rect 267 377 283 411
rect 217 343 283 377
rect 327 485 361 527
rect 327 417 361 451
rect 327 357 361 383
rect 395 479 471 493
rect 395 445 421 479
rect 455 445 471 479
rect 395 411 471 445
rect 395 377 421 411
rect 455 377 471 411
rect 217 309 233 343
rect 267 323 283 343
rect 395 343 471 377
rect 515 485 549 527
rect 515 417 549 451
rect 515 357 549 383
rect 583 479 659 493
rect 583 445 609 479
rect 643 445 659 479
rect 583 411 659 445
rect 583 377 609 411
rect 643 377 659 411
rect 395 323 421 343
rect 267 309 421 323
rect 455 323 471 343
rect 583 343 659 377
rect 703 485 737 527
rect 703 417 737 451
rect 703 367 737 383
rect 771 479 847 493
rect 771 445 797 479
rect 831 445 847 479
rect 771 411 847 445
rect 771 377 797 411
rect 831 377 847 411
rect 455 309 549 323
rect 217 289 549 309
rect 583 309 609 343
rect 643 323 659 343
rect 771 343 847 377
rect 891 485 925 527
rect 891 417 925 451
rect 891 367 925 383
rect 959 479 1035 493
rect 959 445 985 479
rect 1019 445 1035 479
rect 959 411 1035 445
rect 959 377 985 411
rect 1019 377 1035 411
rect 771 323 797 343
rect 643 309 797 323
rect 831 323 847 343
rect 959 343 1035 377
rect 1079 485 1113 527
rect 1079 417 1113 451
rect 1079 367 1113 383
rect 1147 479 1223 493
rect 1147 445 1173 479
rect 1207 445 1223 479
rect 1147 411 1223 445
rect 1147 377 1173 411
rect 1207 377 1223 411
rect 959 323 985 343
rect 831 309 985 323
rect 1019 323 1035 343
rect 1147 343 1223 377
rect 1267 485 1301 527
rect 1267 417 1301 451
rect 1267 367 1301 383
rect 1147 323 1173 343
rect 1019 309 1173 323
rect 1207 323 1223 343
rect 1207 309 1361 323
rect 583 289 1361 309
rect 515 255 549 289
rect 17 249 101 255
rect 17 215 38 249
rect 72 215 101 249
rect 145 249 471 255
rect 145 215 327 249
rect 361 215 395 249
rect 429 215 471 249
rect 515 249 1249 255
rect 515 215 583 249
rect 617 215 661 249
rect 695 215 739 249
rect 773 215 817 249
rect 851 215 895 249
rect 929 215 963 249
rect 997 215 1041 249
rect 1075 215 1119 249
rect 1153 215 1197 249
rect 1231 215 1249 249
rect 145 181 179 215
rect 515 181 549 215
rect 1283 181 1361 289
rect 35 165 69 181
rect 35 97 69 131
rect 35 17 69 63
rect 103 165 179 181
rect 103 131 129 165
rect 163 131 179 165
rect 103 97 179 131
rect 103 63 129 97
rect 163 63 179 97
rect 103 52 179 63
rect 217 165 549 181
rect 217 131 233 165
rect 267 147 421 165
rect 267 131 283 147
rect 217 97 283 131
rect 395 131 421 147
rect 455 147 549 165
rect 583 165 1361 181
rect 455 131 471 147
rect 217 63 233 97
rect 267 63 283 97
rect 217 52 283 63
rect 327 97 361 113
rect 327 17 361 63
rect 395 97 471 131
rect 583 131 609 165
rect 643 147 797 165
rect 643 131 659 147
rect 395 63 421 97
rect 455 63 471 97
rect 395 52 471 63
rect 515 97 549 113
rect 515 17 549 63
rect 583 97 659 131
rect 771 131 797 147
rect 831 147 985 165
rect 831 131 847 147
rect 583 63 609 97
rect 643 63 659 97
rect 583 52 659 63
rect 703 97 737 113
rect 703 17 737 63
rect 771 97 847 131
rect 959 131 985 147
rect 1019 147 1173 165
rect 1019 131 1035 147
rect 771 63 797 97
rect 831 63 847 97
rect 771 52 847 63
rect 891 97 925 113
rect 891 17 925 63
rect 959 97 1035 131
rect 1147 131 1173 147
rect 1207 147 1361 165
rect 1207 131 1223 147
rect 959 63 985 97
rect 1019 63 1035 97
rect 959 52 1035 63
rect 1079 97 1113 113
rect 1079 17 1113 63
rect 1147 97 1223 131
rect 1147 63 1173 97
rect 1207 63 1223 97
rect 1147 52 1223 63
rect 1267 97 1301 113
rect 1267 17 1301 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
<< metal1 >>
rect 0 561 1380 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 0 496 1380 527
rect 0 17 1380 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
rect 0 -48 1380 -17
<< labels >>
flabel corelocali s 30 221 64 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 1317 221 1351 255 0 FreeSans 200 0 0 0 Y
port 6 nsew
flabel corelocali s 1317 289 1351 323 0 FreeSans 200 0 0 0 Y
port 6 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew
rlabel comment s 0 0 0 0 4 bufinv_8
<< properties >>
string FIXED_BBOX 0 0 1380 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1743172
string GDS_START 1732476
<< end >>
