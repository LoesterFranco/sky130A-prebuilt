magic
tech sky130A
magscale 1 2
timestamp 1604502701
<< nwell >>
rect -38 332 710 704
<< pwell >>
rect 0 0 672 49
<< scpmos >>
rect 108 385 138 553
rect 198 385 228 553
rect 346 368 376 592
rect 430 368 460 592
rect 544 368 574 592
<< nmoslvt >>
rect 82 119 112 247
rect 154 119 184 247
rect 348 74 378 222
rect 463 74 493 222
rect 549 74 579 222
<< ndiff >>
rect 27 235 82 247
rect 27 201 37 235
rect 71 201 82 235
rect 27 165 82 201
rect 27 131 37 165
rect 71 131 82 165
rect 27 119 82 131
rect 112 119 154 247
rect 184 235 239 247
rect 184 201 195 235
rect 229 201 239 235
rect 184 165 239 201
rect 184 131 195 165
rect 229 131 239 165
rect 184 119 239 131
rect 293 152 348 222
rect 293 118 303 152
rect 337 118 348 152
rect 293 74 348 118
rect 378 91 463 222
rect 378 74 403 91
rect 393 57 403 74
rect 437 74 463 91
rect 493 152 549 222
rect 493 118 504 152
rect 538 118 549 152
rect 493 74 549 118
rect 579 210 641 222
rect 579 176 595 210
rect 629 176 641 210
rect 579 120 641 176
rect 579 86 595 120
rect 629 86 641 120
rect 579 74 641 86
rect 437 57 448 74
rect 393 38 448 57
<< pdiff >>
rect 287 580 346 592
rect 287 553 299 580
rect 39 524 108 553
rect 39 490 51 524
rect 85 490 108 524
rect 39 431 108 490
rect 39 397 51 431
rect 85 397 108 431
rect 39 385 108 397
rect 138 541 198 553
rect 138 507 151 541
rect 185 507 198 541
rect 138 440 198 507
rect 138 406 151 440
rect 185 406 198 440
rect 138 385 198 406
rect 228 546 299 553
rect 333 546 346 580
rect 228 500 346 546
rect 228 466 299 500
rect 333 466 346 500
rect 228 385 346 466
rect 293 368 346 385
rect 376 368 430 592
rect 460 580 544 592
rect 460 546 487 580
rect 521 546 544 580
rect 460 500 544 546
rect 460 466 487 500
rect 521 466 544 500
rect 460 420 544 466
rect 460 386 487 420
rect 521 386 544 420
rect 460 368 544 386
rect 574 580 633 592
rect 574 546 587 580
rect 621 546 633 580
rect 574 477 633 546
rect 574 443 587 477
rect 621 443 633 477
rect 574 368 633 443
<< ndiffc >>
rect 37 201 71 235
rect 37 131 71 165
rect 195 201 229 235
rect 195 131 229 165
rect 303 118 337 152
rect 403 57 437 91
rect 504 118 538 152
rect 595 176 629 210
rect 595 86 629 120
<< pdiffc >>
rect 51 490 85 524
rect 51 397 85 431
rect 151 507 185 541
rect 151 406 185 440
rect 299 546 333 580
rect 299 466 333 500
rect 487 546 521 580
rect 487 466 521 500
rect 487 386 521 420
rect 587 546 621 580
rect 587 443 621 477
<< poly >>
rect 346 592 376 618
rect 430 592 460 618
rect 544 592 574 618
rect 108 553 138 579
rect 198 553 228 579
rect 108 370 138 385
rect 198 370 228 385
rect 82 340 141 370
rect 195 353 231 370
rect 346 353 376 368
rect 430 353 460 368
rect 544 353 574 368
rect 82 247 112 340
rect 189 337 255 353
rect 189 303 205 337
rect 239 303 255 337
rect 343 336 379 353
rect 189 292 255 303
rect 154 262 255 292
rect 303 320 379 336
rect 303 286 319 320
rect 353 286 379 320
rect 303 270 379 286
rect 427 336 463 353
rect 427 320 493 336
rect 541 326 577 353
rect 427 286 443 320
rect 477 286 493 320
rect 427 270 493 286
rect 154 247 184 262
rect 348 222 378 270
rect 463 222 493 270
rect 535 310 601 326
rect 535 276 551 310
rect 585 276 601 310
rect 535 260 601 276
rect 549 222 579 260
rect 82 51 112 119
rect 154 93 184 119
rect 348 51 378 74
rect 82 21 378 51
rect 463 48 493 74
rect 549 48 579 74
<< polycont >>
rect 205 303 239 337
rect 319 286 353 320
rect 443 286 477 320
rect 551 276 585 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 35 524 101 649
rect 283 580 349 649
rect 35 490 51 524
rect 85 490 101 524
rect 35 458 101 490
rect 135 541 201 557
rect 135 507 151 541
rect 185 507 201 541
rect 35 431 85 458
rect 35 397 51 431
rect 135 440 201 507
rect 283 546 299 580
rect 333 546 349 580
rect 283 500 349 546
rect 283 466 299 500
rect 333 466 349 500
rect 283 458 349 466
rect 409 580 537 596
rect 409 546 487 580
rect 521 546 537 580
rect 409 500 537 546
rect 409 466 487 500
rect 521 466 537 500
rect 409 458 537 466
rect 135 424 151 440
rect 35 381 85 397
rect 121 406 151 424
rect 185 406 201 440
rect 121 390 201 406
rect 235 390 437 424
rect 121 251 155 390
rect 235 356 269 390
rect 189 337 269 356
rect 189 303 205 337
rect 239 303 269 337
rect 189 287 269 303
rect 303 320 369 356
rect 303 286 319 320
rect 353 286 369 320
rect 303 270 369 286
rect 403 336 437 390
rect 471 420 537 458
rect 571 580 637 649
rect 571 546 587 580
rect 621 546 637 580
rect 571 477 637 546
rect 571 443 587 477
rect 621 443 637 477
rect 571 438 637 443
rect 471 386 487 420
rect 521 404 537 420
rect 521 386 655 404
rect 471 370 655 386
rect 403 320 493 336
rect 403 286 443 320
rect 477 286 493 320
rect 403 270 493 286
rect 527 310 587 326
rect 527 276 551 310
rect 585 276 587 310
rect 527 260 587 276
rect 21 235 87 251
rect 21 201 37 235
rect 71 201 87 235
rect 121 236 245 251
rect 527 236 561 260
rect 121 235 561 236
rect 121 217 195 235
rect 21 165 87 201
rect 21 131 37 165
rect 71 131 87 165
rect 21 17 87 131
rect 179 201 195 217
rect 229 202 561 235
rect 621 226 655 370
rect 595 210 655 226
rect 229 201 245 202
rect 179 165 245 201
rect 629 176 655 210
rect 179 131 195 165
rect 229 131 245 165
rect 179 115 245 131
rect 287 152 554 168
rect 287 118 303 152
rect 337 134 504 152
rect 337 118 353 134
rect 287 102 353 118
rect 488 118 504 134
rect 538 118 554 152
rect 488 102 554 118
rect 595 120 655 176
rect 387 91 453 100
rect 387 57 403 91
rect 437 57 453 91
rect 629 86 655 120
rect 595 70 655 86
rect 387 17 453 57
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel comment s 0 0 0 0 4 xnor2_1
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 415 464 449 498 0 FreeSans 340 0 0 0 Y
port 7 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 B
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 672 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 464242
string GDS_START 458282
<< end >>
