magic
tech sky130A
magscale 1 2
timestamp 1601050082
<< locali >>
rect 201 290 267 356
rect 910 289 1044 356
rect 1361 88 1427 596
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 19 364 89 596
rect 137 458 215 649
rect 307 510 481 576
rect 589 530 697 649
rect 307 424 341 510
rect 445 444 511 476
rect 123 390 341 424
rect 375 410 665 444
rect 19 188 53 364
rect 123 310 157 390
rect 87 256 157 310
rect 375 290 409 410
rect 631 377 665 410
rect 731 420 797 596
rect 87 222 312 256
rect 346 224 409 290
rect 451 277 517 368
rect 631 311 697 377
rect 731 277 765 420
rect 842 415 909 591
rect 943 415 1009 649
rect 842 377 876 415
rect 1043 390 1112 591
rect 1146 390 1327 649
rect 799 311 876 377
rect 451 243 807 277
rect 278 190 312 222
rect 19 154 244 188
rect 19 70 73 154
rect 109 17 176 120
rect 210 85 244 154
rect 278 124 449 190
rect 584 151 707 201
rect 566 85 632 117
rect 210 51 632 85
rect 668 17 707 151
rect 741 121 807 243
rect 842 255 876 311
rect 1078 322 1112 390
rect 842 115 919 255
rect 953 17 1019 255
rect 1078 188 1261 322
rect 1111 115 1177 188
rect 1261 17 1327 154
rect 1463 364 1513 649
rect 1463 17 1513 244
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
rlabel locali s 201 290 267 356 6 GATE
port 1 nsew signal input
rlabel locali s 1361 88 1427 596 6 GCLK
port 2 nsew signal output
rlabel locali s 910 289 1044 356 6 CLK
port 3 nsew clock input
rlabel metal1 s 0 -49 1536 49 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1536 715 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1536 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2909356
string GDS_START 2896962
<< end >>
