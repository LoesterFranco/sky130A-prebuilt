magic
tech sky130A
magscale 1 2
timestamp 1604502697
<< nwell >>
rect -38 261 5190 827
<< pwell >>
rect 29 1071 63 1105
rect 1225 1071 1259 1105
rect 1317 1071 1351 1105
rect 2513 1071 2547 1105
rect 2605 1071 2639 1105
rect 3801 1071 3835 1105
rect 3893 1071 3927 1105
rect 5089 1071 5123 1105
rect 29 -17 63 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 3801 -17 3835 17
rect 3893 -17 3927 17
rect 5089 -17 5123 17
<< scnmos >>
rect 89 911 119 1041
rect 173 911 203 1041
rect 277 915 307 1019
rect 361 915 391 1019
rect 587 937 617 1041
rect 671 937 701 1041
rect 897 915 927 1019
rect 981 915 1011 1019
rect 1085 911 1115 1041
rect 1169 911 1199 1041
rect 1377 911 1407 1041
rect 1461 911 1491 1041
rect 1565 915 1595 1019
rect 1649 915 1679 1019
rect 1875 937 1905 1041
rect 1959 937 1989 1041
rect 2185 915 2215 1019
rect 2269 915 2299 1019
rect 2373 911 2403 1041
rect 2457 911 2487 1041
rect 2665 911 2695 1041
rect 2749 911 2779 1041
rect 2853 915 2883 1019
rect 2937 915 2967 1019
rect 3163 937 3193 1041
rect 3247 937 3277 1041
rect 3473 915 3503 1019
rect 3557 915 3587 1019
rect 3661 911 3691 1041
rect 3745 911 3775 1041
rect 3953 911 3983 1041
rect 4037 911 4067 1041
rect 4141 915 4171 1019
rect 4225 915 4255 1019
rect 4451 937 4481 1041
rect 4535 937 4565 1041
rect 4761 915 4791 1019
rect 4845 915 4875 1019
rect 4949 911 4979 1041
rect 5033 911 5063 1041
rect 89 47 119 177
rect 173 47 203 177
rect 277 69 307 173
rect 361 69 391 173
rect 587 47 617 151
rect 671 47 701 151
rect 897 69 927 173
rect 981 69 1011 173
rect 1085 47 1115 177
rect 1169 47 1199 177
rect 1377 47 1407 177
rect 1461 47 1491 177
rect 1565 69 1595 173
rect 1649 69 1679 173
rect 1875 47 1905 151
rect 1959 47 1989 151
rect 2185 69 2215 173
rect 2269 69 2299 173
rect 2373 47 2403 177
rect 2457 47 2487 177
rect 2665 47 2695 177
rect 2749 47 2779 177
rect 2853 69 2883 173
rect 2937 69 2967 173
rect 3163 47 3193 151
rect 3247 47 3277 151
rect 3473 69 3503 173
rect 3557 69 3587 173
rect 3661 47 3691 177
rect 3745 47 3775 177
rect 3953 47 3983 177
rect 4037 47 4067 177
rect 4141 69 4171 173
rect 4225 69 4255 173
rect 4451 47 4481 151
rect 4535 47 4565 151
rect 4761 69 4791 173
rect 4845 69 4875 173
rect 4949 47 4979 177
rect 5033 47 5063 177
<< pmoshvt >>
rect 81 591 117 791
rect 175 591 211 791
rect 280 591 316 755
rect 374 591 410 755
rect 572 591 608 791
rect 680 591 716 791
rect 878 591 914 755
rect 972 591 1008 755
rect 1077 591 1113 791
rect 1171 591 1207 791
rect 1369 591 1405 791
rect 1463 591 1499 791
rect 1568 591 1604 755
rect 1662 591 1698 755
rect 1860 591 1896 791
rect 1968 591 2004 791
rect 2166 591 2202 755
rect 2260 591 2296 755
rect 2365 591 2401 791
rect 2459 591 2495 791
rect 2657 591 2693 791
rect 2751 591 2787 791
rect 2856 591 2892 755
rect 2950 591 2986 755
rect 3148 591 3184 791
rect 3256 591 3292 791
rect 3454 591 3490 755
rect 3548 591 3584 755
rect 3653 591 3689 791
rect 3747 591 3783 791
rect 3945 591 3981 791
rect 4039 591 4075 791
rect 4144 591 4180 755
rect 4238 591 4274 755
rect 4436 591 4472 791
rect 4544 591 4580 791
rect 4742 591 4778 755
rect 4836 591 4872 755
rect 4941 591 4977 791
rect 5035 591 5071 791
rect 81 297 117 497
rect 175 297 211 497
rect 280 333 316 497
rect 374 333 410 497
rect 572 297 608 497
rect 680 297 716 497
rect 878 333 914 497
rect 972 333 1008 497
rect 1077 297 1113 497
rect 1171 297 1207 497
rect 1369 297 1405 497
rect 1463 297 1499 497
rect 1568 333 1604 497
rect 1662 333 1698 497
rect 1860 297 1896 497
rect 1968 297 2004 497
rect 2166 333 2202 497
rect 2260 333 2296 497
rect 2365 297 2401 497
rect 2459 297 2495 497
rect 2657 297 2693 497
rect 2751 297 2787 497
rect 2856 333 2892 497
rect 2950 333 2986 497
rect 3148 297 3184 497
rect 3256 297 3292 497
rect 3454 333 3490 497
rect 3548 333 3584 497
rect 3653 297 3689 497
rect 3747 297 3783 497
rect 3945 297 3981 497
rect 4039 297 4075 497
rect 4144 333 4180 497
rect 4238 333 4274 497
rect 4436 297 4472 497
rect 4544 297 4580 497
rect 4742 333 4778 497
rect 4836 333 4872 497
rect 4941 297 4977 497
rect 5035 297 5071 497
<< ndiff >>
rect 27 1029 89 1041
rect 27 995 45 1029
rect 79 995 89 1029
rect 27 961 89 995
rect 27 927 45 961
rect 79 927 89 961
rect 27 911 89 927
rect 119 1029 173 1041
rect 119 995 129 1029
rect 163 995 173 1029
rect 119 911 173 995
rect 203 1021 262 1041
rect 203 987 218 1021
rect 252 1019 262 1021
rect 252 987 277 1019
rect 203 953 277 987
rect 203 919 218 953
rect 252 919 277 953
rect 203 915 277 919
rect 307 969 361 1019
rect 307 935 317 969
rect 351 935 361 969
rect 307 915 361 935
rect 391 984 443 1019
rect 391 950 401 984
rect 435 950 443 984
rect 391 915 443 950
rect 535 1006 587 1041
rect 535 972 543 1006
rect 577 972 587 1006
rect 535 937 587 972
rect 617 1006 671 1041
rect 617 972 627 1006
rect 661 972 671 1006
rect 617 937 671 972
rect 701 1006 753 1041
rect 701 972 711 1006
rect 745 972 753 1006
rect 701 937 753 972
rect 203 911 262 915
rect 1026 1021 1085 1041
rect 1026 1019 1036 1021
rect 845 984 897 1019
rect 845 950 853 984
rect 887 950 897 984
rect 845 915 897 950
rect 927 969 981 1019
rect 927 935 937 969
rect 971 935 981 969
rect 927 915 981 935
rect 1011 987 1036 1019
rect 1070 987 1085 1021
rect 1011 953 1085 987
rect 1011 919 1036 953
rect 1070 919 1085 953
rect 1011 915 1085 919
rect 1026 911 1085 915
rect 1115 1029 1169 1041
rect 1115 995 1125 1029
rect 1159 995 1169 1029
rect 1115 911 1169 995
rect 1199 1029 1261 1041
rect 1199 995 1209 1029
rect 1243 995 1261 1029
rect 1199 961 1261 995
rect 1199 927 1209 961
rect 1243 927 1261 961
rect 1199 911 1261 927
rect 1315 1029 1377 1041
rect 1315 995 1333 1029
rect 1367 995 1377 1029
rect 1315 961 1377 995
rect 1315 927 1333 961
rect 1367 927 1377 961
rect 1315 911 1377 927
rect 1407 1029 1461 1041
rect 1407 995 1417 1029
rect 1451 995 1461 1029
rect 1407 911 1461 995
rect 1491 1021 1550 1041
rect 1491 987 1506 1021
rect 1540 1019 1550 1021
rect 1540 987 1565 1019
rect 1491 953 1565 987
rect 1491 919 1506 953
rect 1540 919 1565 953
rect 1491 915 1565 919
rect 1595 969 1649 1019
rect 1595 935 1605 969
rect 1639 935 1649 969
rect 1595 915 1649 935
rect 1679 984 1731 1019
rect 1679 950 1689 984
rect 1723 950 1731 984
rect 1679 915 1731 950
rect 1823 1006 1875 1041
rect 1823 972 1831 1006
rect 1865 972 1875 1006
rect 1823 937 1875 972
rect 1905 1006 1959 1041
rect 1905 972 1915 1006
rect 1949 972 1959 1006
rect 1905 937 1959 972
rect 1989 1006 2041 1041
rect 1989 972 1999 1006
rect 2033 972 2041 1006
rect 1989 937 2041 972
rect 1491 911 1550 915
rect 2314 1021 2373 1041
rect 2314 1019 2324 1021
rect 2133 984 2185 1019
rect 2133 950 2141 984
rect 2175 950 2185 984
rect 2133 915 2185 950
rect 2215 969 2269 1019
rect 2215 935 2225 969
rect 2259 935 2269 969
rect 2215 915 2269 935
rect 2299 987 2324 1019
rect 2358 987 2373 1021
rect 2299 953 2373 987
rect 2299 919 2324 953
rect 2358 919 2373 953
rect 2299 915 2373 919
rect 2314 911 2373 915
rect 2403 1029 2457 1041
rect 2403 995 2413 1029
rect 2447 995 2457 1029
rect 2403 911 2457 995
rect 2487 1029 2549 1041
rect 2487 995 2497 1029
rect 2531 995 2549 1029
rect 2487 961 2549 995
rect 2487 927 2497 961
rect 2531 927 2549 961
rect 2487 911 2549 927
rect 2603 1029 2665 1041
rect 2603 995 2621 1029
rect 2655 995 2665 1029
rect 2603 961 2665 995
rect 2603 927 2621 961
rect 2655 927 2665 961
rect 2603 911 2665 927
rect 2695 1029 2749 1041
rect 2695 995 2705 1029
rect 2739 995 2749 1029
rect 2695 911 2749 995
rect 2779 1021 2838 1041
rect 2779 987 2794 1021
rect 2828 1019 2838 1021
rect 2828 987 2853 1019
rect 2779 953 2853 987
rect 2779 919 2794 953
rect 2828 919 2853 953
rect 2779 915 2853 919
rect 2883 969 2937 1019
rect 2883 935 2893 969
rect 2927 935 2937 969
rect 2883 915 2937 935
rect 2967 984 3019 1019
rect 2967 950 2977 984
rect 3011 950 3019 984
rect 2967 915 3019 950
rect 3111 1006 3163 1041
rect 3111 972 3119 1006
rect 3153 972 3163 1006
rect 3111 937 3163 972
rect 3193 1006 3247 1041
rect 3193 972 3203 1006
rect 3237 972 3247 1006
rect 3193 937 3247 972
rect 3277 1006 3329 1041
rect 3277 972 3287 1006
rect 3321 972 3329 1006
rect 3277 937 3329 972
rect 2779 911 2838 915
rect 3602 1021 3661 1041
rect 3602 1019 3612 1021
rect 3421 984 3473 1019
rect 3421 950 3429 984
rect 3463 950 3473 984
rect 3421 915 3473 950
rect 3503 969 3557 1019
rect 3503 935 3513 969
rect 3547 935 3557 969
rect 3503 915 3557 935
rect 3587 987 3612 1019
rect 3646 987 3661 1021
rect 3587 953 3661 987
rect 3587 919 3612 953
rect 3646 919 3661 953
rect 3587 915 3661 919
rect 3602 911 3661 915
rect 3691 1029 3745 1041
rect 3691 995 3701 1029
rect 3735 995 3745 1029
rect 3691 911 3745 995
rect 3775 1029 3837 1041
rect 3775 995 3785 1029
rect 3819 995 3837 1029
rect 3775 961 3837 995
rect 3775 927 3785 961
rect 3819 927 3837 961
rect 3775 911 3837 927
rect 3891 1029 3953 1041
rect 3891 995 3909 1029
rect 3943 995 3953 1029
rect 3891 961 3953 995
rect 3891 927 3909 961
rect 3943 927 3953 961
rect 3891 911 3953 927
rect 3983 1029 4037 1041
rect 3983 995 3993 1029
rect 4027 995 4037 1029
rect 3983 911 4037 995
rect 4067 1021 4126 1041
rect 4067 987 4082 1021
rect 4116 1019 4126 1021
rect 4116 987 4141 1019
rect 4067 953 4141 987
rect 4067 919 4082 953
rect 4116 919 4141 953
rect 4067 915 4141 919
rect 4171 969 4225 1019
rect 4171 935 4181 969
rect 4215 935 4225 969
rect 4171 915 4225 935
rect 4255 984 4307 1019
rect 4255 950 4265 984
rect 4299 950 4307 984
rect 4255 915 4307 950
rect 4399 1006 4451 1041
rect 4399 972 4407 1006
rect 4441 972 4451 1006
rect 4399 937 4451 972
rect 4481 1006 4535 1041
rect 4481 972 4491 1006
rect 4525 972 4535 1006
rect 4481 937 4535 972
rect 4565 1006 4617 1041
rect 4565 972 4575 1006
rect 4609 972 4617 1006
rect 4565 937 4617 972
rect 4067 911 4126 915
rect 4890 1021 4949 1041
rect 4890 1019 4900 1021
rect 4709 984 4761 1019
rect 4709 950 4717 984
rect 4751 950 4761 984
rect 4709 915 4761 950
rect 4791 969 4845 1019
rect 4791 935 4801 969
rect 4835 935 4845 969
rect 4791 915 4845 935
rect 4875 987 4900 1019
rect 4934 987 4949 1021
rect 4875 953 4949 987
rect 4875 919 4900 953
rect 4934 919 4949 953
rect 4875 915 4949 919
rect 4890 911 4949 915
rect 4979 1029 5033 1041
rect 4979 995 4989 1029
rect 5023 995 5033 1029
rect 4979 911 5033 995
rect 5063 1029 5125 1041
rect 5063 995 5073 1029
rect 5107 995 5125 1029
rect 5063 961 5125 995
rect 5063 927 5073 961
rect 5107 927 5125 961
rect 5063 911 5125 927
rect 27 161 89 177
rect 27 127 45 161
rect 79 127 89 161
rect 27 93 89 127
rect 27 59 45 93
rect 79 59 89 93
rect 27 47 89 59
rect 119 93 173 177
rect 119 59 129 93
rect 163 59 173 93
rect 119 47 173 59
rect 203 173 262 177
rect 203 169 277 173
rect 203 135 218 169
rect 252 135 277 169
rect 203 101 277 135
rect 203 67 218 101
rect 252 69 277 101
rect 307 153 361 173
rect 307 119 317 153
rect 351 119 361 153
rect 307 69 361 119
rect 391 138 443 173
rect 391 104 401 138
rect 435 104 443 138
rect 391 69 443 104
rect 252 67 262 69
rect 203 47 262 67
rect 1026 173 1085 177
rect 535 116 587 151
rect 535 82 543 116
rect 577 82 587 116
rect 535 47 587 82
rect 617 116 671 151
rect 617 82 627 116
rect 661 82 671 116
rect 617 47 671 82
rect 701 116 753 151
rect 701 82 711 116
rect 745 82 753 116
rect 701 47 753 82
rect 845 138 897 173
rect 845 104 853 138
rect 887 104 897 138
rect 845 69 897 104
rect 927 153 981 173
rect 927 119 937 153
rect 971 119 981 153
rect 927 69 981 119
rect 1011 169 1085 173
rect 1011 135 1036 169
rect 1070 135 1085 169
rect 1011 101 1085 135
rect 1011 69 1036 101
rect 1026 67 1036 69
rect 1070 67 1085 101
rect 1026 47 1085 67
rect 1115 93 1169 177
rect 1115 59 1125 93
rect 1159 59 1169 93
rect 1115 47 1169 59
rect 1199 161 1261 177
rect 1199 127 1209 161
rect 1243 127 1261 161
rect 1199 93 1261 127
rect 1199 59 1209 93
rect 1243 59 1261 93
rect 1199 47 1261 59
rect 1315 161 1377 177
rect 1315 127 1333 161
rect 1367 127 1377 161
rect 1315 93 1377 127
rect 1315 59 1333 93
rect 1367 59 1377 93
rect 1315 47 1377 59
rect 1407 93 1461 177
rect 1407 59 1417 93
rect 1451 59 1461 93
rect 1407 47 1461 59
rect 1491 173 1550 177
rect 1491 169 1565 173
rect 1491 135 1506 169
rect 1540 135 1565 169
rect 1491 101 1565 135
rect 1491 67 1506 101
rect 1540 69 1565 101
rect 1595 153 1649 173
rect 1595 119 1605 153
rect 1639 119 1649 153
rect 1595 69 1649 119
rect 1679 138 1731 173
rect 1679 104 1689 138
rect 1723 104 1731 138
rect 1679 69 1731 104
rect 1540 67 1550 69
rect 1491 47 1550 67
rect 2314 173 2373 177
rect 1823 116 1875 151
rect 1823 82 1831 116
rect 1865 82 1875 116
rect 1823 47 1875 82
rect 1905 116 1959 151
rect 1905 82 1915 116
rect 1949 82 1959 116
rect 1905 47 1959 82
rect 1989 116 2041 151
rect 1989 82 1999 116
rect 2033 82 2041 116
rect 1989 47 2041 82
rect 2133 138 2185 173
rect 2133 104 2141 138
rect 2175 104 2185 138
rect 2133 69 2185 104
rect 2215 153 2269 173
rect 2215 119 2225 153
rect 2259 119 2269 153
rect 2215 69 2269 119
rect 2299 169 2373 173
rect 2299 135 2324 169
rect 2358 135 2373 169
rect 2299 101 2373 135
rect 2299 69 2324 101
rect 2314 67 2324 69
rect 2358 67 2373 101
rect 2314 47 2373 67
rect 2403 93 2457 177
rect 2403 59 2413 93
rect 2447 59 2457 93
rect 2403 47 2457 59
rect 2487 161 2549 177
rect 2487 127 2497 161
rect 2531 127 2549 161
rect 2487 93 2549 127
rect 2487 59 2497 93
rect 2531 59 2549 93
rect 2487 47 2549 59
rect 2603 161 2665 177
rect 2603 127 2621 161
rect 2655 127 2665 161
rect 2603 93 2665 127
rect 2603 59 2621 93
rect 2655 59 2665 93
rect 2603 47 2665 59
rect 2695 93 2749 177
rect 2695 59 2705 93
rect 2739 59 2749 93
rect 2695 47 2749 59
rect 2779 173 2838 177
rect 2779 169 2853 173
rect 2779 135 2794 169
rect 2828 135 2853 169
rect 2779 101 2853 135
rect 2779 67 2794 101
rect 2828 69 2853 101
rect 2883 153 2937 173
rect 2883 119 2893 153
rect 2927 119 2937 153
rect 2883 69 2937 119
rect 2967 138 3019 173
rect 2967 104 2977 138
rect 3011 104 3019 138
rect 2967 69 3019 104
rect 2828 67 2838 69
rect 2779 47 2838 67
rect 3602 173 3661 177
rect 3111 116 3163 151
rect 3111 82 3119 116
rect 3153 82 3163 116
rect 3111 47 3163 82
rect 3193 116 3247 151
rect 3193 82 3203 116
rect 3237 82 3247 116
rect 3193 47 3247 82
rect 3277 116 3329 151
rect 3277 82 3287 116
rect 3321 82 3329 116
rect 3277 47 3329 82
rect 3421 138 3473 173
rect 3421 104 3429 138
rect 3463 104 3473 138
rect 3421 69 3473 104
rect 3503 153 3557 173
rect 3503 119 3513 153
rect 3547 119 3557 153
rect 3503 69 3557 119
rect 3587 169 3661 173
rect 3587 135 3612 169
rect 3646 135 3661 169
rect 3587 101 3661 135
rect 3587 69 3612 101
rect 3602 67 3612 69
rect 3646 67 3661 101
rect 3602 47 3661 67
rect 3691 93 3745 177
rect 3691 59 3701 93
rect 3735 59 3745 93
rect 3691 47 3745 59
rect 3775 161 3837 177
rect 3775 127 3785 161
rect 3819 127 3837 161
rect 3775 93 3837 127
rect 3775 59 3785 93
rect 3819 59 3837 93
rect 3775 47 3837 59
rect 3891 161 3953 177
rect 3891 127 3909 161
rect 3943 127 3953 161
rect 3891 93 3953 127
rect 3891 59 3909 93
rect 3943 59 3953 93
rect 3891 47 3953 59
rect 3983 93 4037 177
rect 3983 59 3993 93
rect 4027 59 4037 93
rect 3983 47 4037 59
rect 4067 173 4126 177
rect 4067 169 4141 173
rect 4067 135 4082 169
rect 4116 135 4141 169
rect 4067 101 4141 135
rect 4067 67 4082 101
rect 4116 69 4141 101
rect 4171 153 4225 173
rect 4171 119 4181 153
rect 4215 119 4225 153
rect 4171 69 4225 119
rect 4255 138 4307 173
rect 4255 104 4265 138
rect 4299 104 4307 138
rect 4255 69 4307 104
rect 4116 67 4126 69
rect 4067 47 4126 67
rect 4890 173 4949 177
rect 4399 116 4451 151
rect 4399 82 4407 116
rect 4441 82 4451 116
rect 4399 47 4451 82
rect 4481 116 4535 151
rect 4481 82 4491 116
rect 4525 82 4535 116
rect 4481 47 4535 82
rect 4565 116 4617 151
rect 4565 82 4575 116
rect 4609 82 4617 116
rect 4565 47 4617 82
rect 4709 138 4761 173
rect 4709 104 4717 138
rect 4751 104 4761 138
rect 4709 69 4761 104
rect 4791 153 4845 173
rect 4791 119 4801 153
rect 4835 119 4845 153
rect 4791 69 4845 119
rect 4875 169 4949 173
rect 4875 135 4900 169
rect 4934 135 4949 169
rect 4875 101 4949 135
rect 4875 69 4900 101
rect 4890 67 4900 69
rect 4934 67 4949 101
rect 4890 47 4949 67
rect 4979 93 5033 177
rect 4979 59 4989 93
rect 5023 59 5033 93
rect 4979 47 5033 59
rect 5063 161 5125 177
rect 5063 127 5073 161
rect 5107 127 5125 161
rect 5063 93 5125 127
rect 5063 59 5073 93
rect 5107 59 5125 93
rect 5063 47 5125 59
<< pdiff >>
rect 27 773 81 791
rect 27 739 35 773
rect 69 739 81 773
rect 27 705 81 739
rect 27 671 35 705
rect 69 671 81 705
rect 27 637 81 671
rect 27 603 35 637
rect 69 603 81 637
rect 27 591 81 603
rect 117 717 175 791
rect 117 683 129 717
rect 163 683 175 717
rect 117 637 175 683
rect 117 603 129 637
rect 163 603 175 637
rect 117 591 175 603
rect 211 755 263 791
rect 518 779 572 791
rect 211 749 280 755
rect 211 715 223 749
rect 257 715 280 749
rect 211 645 280 715
rect 211 611 223 645
rect 257 611 280 645
rect 211 591 280 611
rect 316 701 374 755
rect 316 667 328 701
rect 362 667 374 701
rect 316 591 374 667
rect 410 743 464 755
rect 410 709 422 743
rect 456 709 464 743
rect 410 645 464 709
rect 410 611 422 645
rect 456 611 464 645
rect 410 591 464 611
rect 518 745 526 779
rect 560 745 572 779
rect 518 711 572 745
rect 518 677 526 711
rect 560 677 572 711
rect 518 643 572 677
rect 518 609 526 643
rect 560 609 572 643
rect 518 591 572 609
rect 608 779 680 791
rect 608 745 627 779
rect 661 745 680 779
rect 608 711 680 745
rect 608 677 627 711
rect 661 677 680 711
rect 608 643 680 677
rect 608 609 627 643
rect 661 609 680 643
rect 608 591 680 609
rect 716 779 770 791
rect 716 745 728 779
rect 762 745 770 779
rect 1025 755 1077 791
rect 716 711 770 745
rect 716 677 728 711
rect 762 677 770 711
rect 716 643 770 677
rect 716 609 728 643
rect 762 609 770 643
rect 716 591 770 609
rect 824 743 878 755
rect 824 709 832 743
rect 866 709 878 743
rect 824 645 878 709
rect 824 611 832 645
rect 866 611 878 645
rect 824 591 878 611
rect 914 701 972 755
rect 914 667 926 701
rect 960 667 972 701
rect 914 591 972 667
rect 1008 749 1077 755
rect 1008 715 1031 749
rect 1065 715 1077 749
rect 1008 645 1077 715
rect 1008 611 1031 645
rect 1065 611 1077 645
rect 1008 591 1077 611
rect 1113 717 1171 791
rect 1113 683 1125 717
rect 1159 683 1171 717
rect 1113 637 1171 683
rect 1113 603 1125 637
rect 1159 603 1171 637
rect 1113 591 1171 603
rect 1207 773 1261 791
rect 1207 739 1219 773
rect 1253 739 1261 773
rect 1207 705 1261 739
rect 1207 671 1219 705
rect 1253 671 1261 705
rect 1207 637 1261 671
rect 1207 603 1219 637
rect 1253 603 1261 637
rect 1207 591 1261 603
rect 1315 773 1369 791
rect 1315 739 1323 773
rect 1357 739 1369 773
rect 1315 705 1369 739
rect 1315 671 1323 705
rect 1357 671 1369 705
rect 1315 637 1369 671
rect 1315 603 1323 637
rect 1357 603 1369 637
rect 1315 591 1369 603
rect 1405 717 1463 791
rect 1405 683 1417 717
rect 1451 683 1463 717
rect 1405 637 1463 683
rect 1405 603 1417 637
rect 1451 603 1463 637
rect 1405 591 1463 603
rect 1499 755 1551 791
rect 1806 779 1860 791
rect 1499 749 1568 755
rect 1499 715 1511 749
rect 1545 715 1568 749
rect 1499 645 1568 715
rect 1499 611 1511 645
rect 1545 611 1568 645
rect 1499 591 1568 611
rect 1604 701 1662 755
rect 1604 667 1616 701
rect 1650 667 1662 701
rect 1604 591 1662 667
rect 1698 743 1752 755
rect 1698 709 1710 743
rect 1744 709 1752 743
rect 1698 645 1752 709
rect 1698 611 1710 645
rect 1744 611 1752 645
rect 1698 591 1752 611
rect 1806 745 1814 779
rect 1848 745 1860 779
rect 1806 711 1860 745
rect 1806 677 1814 711
rect 1848 677 1860 711
rect 1806 643 1860 677
rect 1806 609 1814 643
rect 1848 609 1860 643
rect 1806 591 1860 609
rect 1896 779 1968 791
rect 1896 745 1915 779
rect 1949 745 1968 779
rect 1896 711 1968 745
rect 1896 677 1915 711
rect 1949 677 1968 711
rect 1896 643 1968 677
rect 1896 609 1915 643
rect 1949 609 1968 643
rect 1896 591 1968 609
rect 2004 779 2058 791
rect 2004 745 2016 779
rect 2050 745 2058 779
rect 2313 755 2365 791
rect 2004 711 2058 745
rect 2004 677 2016 711
rect 2050 677 2058 711
rect 2004 643 2058 677
rect 2004 609 2016 643
rect 2050 609 2058 643
rect 2004 591 2058 609
rect 2112 743 2166 755
rect 2112 709 2120 743
rect 2154 709 2166 743
rect 2112 645 2166 709
rect 2112 611 2120 645
rect 2154 611 2166 645
rect 2112 591 2166 611
rect 2202 701 2260 755
rect 2202 667 2214 701
rect 2248 667 2260 701
rect 2202 591 2260 667
rect 2296 749 2365 755
rect 2296 715 2319 749
rect 2353 715 2365 749
rect 2296 645 2365 715
rect 2296 611 2319 645
rect 2353 611 2365 645
rect 2296 591 2365 611
rect 2401 717 2459 791
rect 2401 683 2413 717
rect 2447 683 2459 717
rect 2401 637 2459 683
rect 2401 603 2413 637
rect 2447 603 2459 637
rect 2401 591 2459 603
rect 2495 773 2549 791
rect 2495 739 2507 773
rect 2541 739 2549 773
rect 2495 705 2549 739
rect 2495 671 2507 705
rect 2541 671 2549 705
rect 2495 637 2549 671
rect 2495 603 2507 637
rect 2541 603 2549 637
rect 2495 591 2549 603
rect 2603 773 2657 791
rect 2603 739 2611 773
rect 2645 739 2657 773
rect 2603 705 2657 739
rect 2603 671 2611 705
rect 2645 671 2657 705
rect 2603 637 2657 671
rect 2603 603 2611 637
rect 2645 603 2657 637
rect 2603 591 2657 603
rect 2693 717 2751 791
rect 2693 683 2705 717
rect 2739 683 2751 717
rect 2693 637 2751 683
rect 2693 603 2705 637
rect 2739 603 2751 637
rect 2693 591 2751 603
rect 2787 755 2839 791
rect 3094 779 3148 791
rect 2787 749 2856 755
rect 2787 715 2799 749
rect 2833 715 2856 749
rect 2787 645 2856 715
rect 2787 611 2799 645
rect 2833 611 2856 645
rect 2787 591 2856 611
rect 2892 701 2950 755
rect 2892 667 2904 701
rect 2938 667 2950 701
rect 2892 591 2950 667
rect 2986 743 3040 755
rect 2986 709 2998 743
rect 3032 709 3040 743
rect 2986 645 3040 709
rect 2986 611 2998 645
rect 3032 611 3040 645
rect 2986 591 3040 611
rect 3094 745 3102 779
rect 3136 745 3148 779
rect 3094 711 3148 745
rect 3094 677 3102 711
rect 3136 677 3148 711
rect 3094 643 3148 677
rect 3094 609 3102 643
rect 3136 609 3148 643
rect 3094 591 3148 609
rect 3184 779 3256 791
rect 3184 745 3203 779
rect 3237 745 3256 779
rect 3184 711 3256 745
rect 3184 677 3203 711
rect 3237 677 3256 711
rect 3184 643 3256 677
rect 3184 609 3203 643
rect 3237 609 3256 643
rect 3184 591 3256 609
rect 3292 779 3346 791
rect 3292 745 3304 779
rect 3338 745 3346 779
rect 3601 755 3653 791
rect 3292 711 3346 745
rect 3292 677 3304 711
rect 3338 677 3346 711
rect 3292 643 3346 677
rect 3292 609 3304 643
rect 3338 609 3346 643
rect 3292 591 3346 609
rect 3400 743 3454 755
rect 3400 709 3408 743
rect 3442 709 3454 743
rect 3400 645 3454 709
rect 3400 611 3408 645
rect 3442 611 3454 645
rect 3400 591 3454 611
rect 3490 701 3548 755
rect 3490 667 3502 701
rect 3536 667 3548 701
rect 3490 591 3548 667
rect 3584 749 3653 755
rect 3584 715 3607 749
rect 3641 715 3653 749
rect 3584 645 3653 715
rect 3584 611 3607 645
rect 3641 611 3653 645
rect 3584 591 3653 611
rect 3689 717 3747 791
rect 3689 683 3701 717
rect 3735 683 3747 717
rect 3689 637 3747 683
rect 3689 603 3701 637
rect 3735 603 3747 637
rect 3689 591 3747 603
rect 3783 773 3837 791
rect 3783 739 3795 773
rect 3829 739 3837 773
rect 3783 705 3837 739
rect 3783 671 3795 705
rect 3829 671 3837 705
rect 3783 637 3837 671
rect 3783 603 3795 637
rect 3829 603 3837 637
rect 3783 591 3837 603
rect 3891 773 3945 791
rect 3891 739 3899 773
rect 3933 739 3945 773
rect 3891 705 3945 739
rect 3891 671 3899 705
rect 3933 671 3945 705
rect 3891 637 3945 671
rect 3891 603 3899 637
rect 3933 603 3945 637
rect 3891 591 3945 603
rect 3981 717 4039 791
rect 3981 683 3993 717
rect 4027 683 4039 717
rect 3981 637 4039 683
rect 3981 603 3993 637
rect 4027 603 4039 637
rect 3981 591 4039 603
rect 4075 755 4127 791
rect 4382 779 4436 791
rect 4075 749 4144 755
rect 4075 715 4087 749
rect 4121 715 4144 749
rect 4075 645 4144 715
rect 4075 611 4087 645
rect 4121 611 4144 645
rect 4075 591 4144 611
rect 4180 701 4238 755
rect 4180 667 4192 701
rect 4226 667 4238 701
rect 4180 591 4238 667
rect 4274 743 4328 755
rect 4274 709 4286 743
rect 4320 709 4328 743
rect 4274 645 4328 709
rect 4274 611 4286 645
rect 4320 611 4328 645
rect 4274 591 4328 611
rect 4382 745 4390 779
rect 4424 745 4436 779
rect 4382 711 4436 745
rect 4382 677 4390 711
rect 4424 677 4436 711
rect 4382 643 4436 677
rect 4382 609 4390 643
rect 4424 609 4436 643
rect 4382 591 4436 609
rect 4472 779 4544 791
rect 4472 745 4491 779
rect 4525 745 4544 779
rect 4472 711 4544 745
rect 4472 677 4491 711
rect 4525 677 4544 711
rect 4472 643 4544 677
rect 4472 609 4491 643
rect 4525 609 4544 643
rect 4472 591 4544 609
rect 4580 779 4634 791
rect 4580 745 4592 779
rect 4626 745 4634 779
rect 4889 755 4941 791
rect 4580 711 4634 745
rect 4580 677 4592 711
rect 4626 677 4634 711
rect 4580 643 4634 677
rect 4580 609 4592 643
rect 4626 609 4634 643
rect 4580 591 4634 609
rect 4688 743 4742 755
rect 4688 709 4696 743
rect 4730 709 4742 743
rect 4688 645 4742 709
rect 4688 611 4696 645
rect 4730 611 4742 645
rect 4688 591 4742 611
rect 4778 701 4836 755
rect 4778 667 4790 701
rect 4824 667 4836 701
rect 4778 591 4836 667
rect 4872 749 4941 755
rect 4872 715 4895 749
rect 4929 715 4941 749
rect 4872 645 4941 715
rect 4872 611 4895 645
rect 4929 611 4941 645
rect 4872 591 4941 611
rect 4977 717 5035 791
rect 4977 683 4989 717
rect 5023 683 5035 717
rect 4977 637 5035 683
rect 4977 603 4989 637
rect 5023 603 5035 637
rect 4977 591 5035 603
rect 5071 773 5125 791
rect 5071 739 5083 773
rect 5117 739 5125 773
rect 5071 705 5125 739
rect 5071 671 5083 705
rect 5117 671 5125 705
rect 5071 637 5125 671
rect 5071 603 5083 637
rect 5117 603 5125 637
rect 5071 591 5125 603
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 485 175 497
rect 117 451 129 485
rect 163 451 175 485
rect 117 405 175 451
rect 117 371 129 405
rect 163 371 175 405
rect 117 297 175 371
rect 211 477 280 497
rect 211 443 223 477
rect 257 443 280 477
rect 211 373 280 443
rect 211 339 223 373
rect 257 339 280 373
rect 211 333 280 339
rect 316 421 374 497
rect 316 387 328 421
rect 362 387 374 421
rect 316 333 374 387
rect 410 477 464 497
rect 410 443 422 477
rect 456 443 464 477
rect 410 379 464 443
rect 410 345 422 379
rect 456 345 464 379
rect 410 333 464 345
rect 518 479 572 497
rect 518 445 526 479
rect 560 445 572 479
rect 518 411 572 445
rect 518 377 526 411
rect 560 377 572 411
rect 518 343 572 377
rect 211 297 263 333
rect 518 309 526 343
rect 560 309 572 343
rect 518 297 572 309
rect 608 479 680 497
rect 608 445 627 479
rect 661 445 680 479
rect 608 411 680 445
rect 608 377 627 411
rect 661 377 680 411
rect 608 343 680 377
rect 608 309 627 343
rect 661 309 680 343
rect 608 297 680 309
rect 716 479 770 497
rect 716 445 728 479
rect 762 445 770 479
rect 716 411 770 445
rect 716 377 728 411
rect 762 377 770 411
rect 716 343 770 377
rect 716 309 728 343
rect 762 309 770 343
rect 824 477 878 497
rect 824 443 832 477
rect 866 443 878 477
rect 824 379 878 443
rect 824 345 832 379
rect 866 345 878 379
rect 824 333 878 345
rect 914 421 972 497
rect 914 387 926 421
rect 960 387 972 421
rect 914 333 972 387
rect 1008 477 1077 497
rect 1008 443 1031 477
rect 1065 443 1077 477
rect 1008 373 1077 443
rect 1008 339 1031 373
rect 1065 339 1077 373
rect 1008 333 1077 339
rect 716 297 770 309
rect 1025 297 1077 333
rect 1113 485 1171 497
rect 1113 451 1125 485
rect 1159 451 1171 485
rect 1113 405 1171 451
rect 1113 371 1125 405
rect 1159 371 1171 405
rect 1113 297 1171 371
rect 1207 485 1261 497
rect 1207 451 1219 485
rect 1253 451 1261 485
rect 1207 417 1261 451
rect 1207 383 1219 417
rect 1253 383 1261 417
rect 1207 349 1261 383
rect 1207 315 1219 349
rect 1253 315 1261 349
rect 1207 297 1261 315
rect 1315 485 1369 497
rect 1315 451 1323 485
rect 1357 451 1369 485
rect 1315 417 1369 451
rect 1315 383 1323 417
rect 1357 383 1369 417
rect 1315 349 1369 383
rect 1315 315 1323 349
rect 1357 315 1369 349
rect 1315 297 1369 315
rect 1405 485 1463 497
rect 1405 451 1417 485
rect 1451 451 1463 485
rect 1405 405 1463 451
rect 1405 371 1417 405
rect 1451 371 1463 405
rect 1405 297 1463 371
rect 1499 477 1568 497
rect 1499 443 1511 477
rect 1545 443 1568 477
rect 1499 373 1568 443
rect 1499 339 1511 373
rect 1545 339 1568 373
rect 1499 333 1568 339
rect 1604 421 1662 497
rect 1604 387 1616 421
rect 1650 387 1662 421
rect 1604 333 1662 387
rect 1698 477 1752 497
rect 1698 443 1710 477
rect 1744 443 1752 477
rect 1698 379 1752 443
rect 1698 345 1710 379
rect 1744 345 1752 379
rect 1698 333 1752 345
rect 1806 479 1860 497
rect 1806 445 1814 479
rect 1848 445 1860 479
rect 1806 411 1860 445
rect 1806 377 1814 411
rect 1848 377 1860 411
rect 1806 343 1860 377
rect 1499 297 1551 333
rect 1806 309 1814 343
rect 1848 309 1860 343
rect 1806 297 1860 309
rect 1896 479 1968 497
rect 1896 445 1915 479
rect 1949 445 1968 479
rect 1896 411 1968 445
rect 1896 377 1915 411
rect 1949 377 1968 411
rect 1896 343 1968 377
rect 1896 309 1915 343
rect 1949 309 1968 343
rect 1896 297 1968 309
rect 2004 479 2058 497
rect 2004 445 2016 479
rect 2050 445 2058 479
rect 2004 411 2058 445
rect 2004 377 2016 411
rect 2050 377 2058 411
rect 2004 343 2058 377
rect 2004 309 2016 343
rect 2050 309 2058 343
rect 2112 477 2166 497
rect 2112 443 2120 477
rect 2154 443 2166 477
rect 2112 379 2166 443
rect 2112 345 2120 379
rect 2154 345 2166 379
rect 2112 333 2166 345
rect 2202 421 2260 497
rect 2202 387 2214 421
rect 2248 387 2260 421
rect 2202 333 2260 387
rect 2296 477 2365 497
rect 2296 443 2319 477
rect 2353 443 2365 477
rect 2296 373 2365 443
rect 2296 339 2319 373
rect 2353 339 2365 373
rect 2296 333 2365 339
rect 2004 297 2058 309
rect 2313 297 2365 333
rect 2401 485 2459 497
rect 2401 451 2413 485
rect 2447 451 2459 485
rect 2401 405 2459 451
rect 2401 371 2413 405
rect 2447 371 2459 405
rect 2401 297 2459 371
rect 2495 485 2549 497
rect 2495 451 2507 485
rect 2541 451 2549 485
rect 2495 417 2549 451
rect 2495 383 2507 417
rect 2541 383 2549 417
rect 2495 349 2549 383
rect 2495 315 2507 349
rect 2541 315 2549 349
rect 2495 297 2549 315
rect 2603 485 2657 497
rect 2603 451 2611 485
rect 2645 451 2657 485
rect 2603 417 2657 451
rect 2603 383 2611 417
rect 2645 383 2657 417
rect 2603 349 2657 383
rect 2603 315 2611 349
rect 2645 315 2657 349
rect 2603 297 2657 315
rect 2693 485 2751 497
rect 2693 451 2705 485
rect 2739 451 2751 485
rect 2693 405 2751 451
rect 2693 371 2705 405
rect 2739 371 2751 405
rect 2693 297 2751 371
rect 2787 477 2856 497
rect 2787 443 2799 477
rect 2833 443 2856 477
rect 2787 373 2856 443
rect 2787 339 2799 373
rect 2833 339 2856 373
rect 2787 333 2856 339
rect 2892 421 2950 497
rect 2892 387 2904 421
rect 2938 387 2950 421
rect 2892 333 2950 387
rect 2986 477 3040 497
rect 2986 443 2998 477
rect 3032 443 3040 477
rect 2986 379 3040 443
rect 2986 345 2998 379
rect 3032 345 3040 379
rect 2986 333 3040 345
rect 3094 479 3148 497
rect 3094 445 3102 479
rect 3136 445 3148 479
rect 3094 411 3148 445
rect 3094 377 3102 411
rect 3136 377 3148 411
rect 3094 343 3148 377
rect 2787 297 2839 333
rect 3094 309 3102 343
rect 3136 309 3148 343
rect 3094 297 3148 309
rect 3184 479 3256 497
rect 3184 445 3203 479
rect 3237 445 3256 479
rect 3184 411 3256 445
rect 3184 377 3203 411
rect 3237 377 3256 411
rect 3184 343 3256 377
rect 3184 309 3203 343
rect 3237 309 3256 343
rect 3184 297 3256 309
rect 3292 479 3346 497
rect 3292 445 3304 479
rect 3338 445 3346 479
rect 3292 411 3346 445
rect 3292 377 3304 411
rect 3338 377 3346 411
rect 3292 343 3346 377
rect 3292 309 3304 343
rect 3338 309 3346 343
rect 3400 477 3454 497
rect 3400 443 3408 477
rect 3442 443 3454 477
rect 3400 379 3454 443
rect 3400 345 3408 379
rect 3442 345 3454 379
rect 3400 333 3454 345
rect 3490 421 3548 497
rect 3490 387 3502 421
rect 3536 387 3548 421
rect 3490 333 3548 387
rect 3584 477 3653 497
rect 3584 443 3607 477
rect 3641 443 3653 477
rect 3584 373 3653 443
rect 3584 339 3607 373
rect 3641 339 3653 373
rect 3584 333 3653 339
rect 3292 297 3346 309
rect 3601 297 3653 333
rect 3689 485 3747 497
rect 3689 451 3701 485
rect 3735 451 3747 485
rect 3689 405 3747 451
rect 3689 371 3701 405
rect 3735 371 3747 405
rect 3689 297 3747 371
rect 3783 485 3837 497
rect 3783 451 3795 485
rect 3829 451 3837 485
rect 3783 417 3837 451
rect 3783 383 3795 417
rect 3829 383 3837 417
rect 3783 349 3837 383
rect 3783 315 3795 349
rect 3829 315 3837 349
rect 3783 297 3837 315
rect 3891 485 3945 497
rect 3891 451 3899 485
rect 3933 451 3945 485
rect 3891 417 3945 451
rect 3891 383 3899 417
rect 3933 383 3945 417
rect 3891 349 3945 383
rect 3891 315 3899 349
rect 3933 315 3945 349
rect 3891 297 3945 315
rect 3981 485 4039 497
rect 3981 451 3993 485
rect 4027 451 4039 485
rect 3981 405 4039 451
rect 3981 371 3993 405
rect 4027 371 4039 405
rect 3981 297 4039 371
rect 4075 477 4144 497
rect 4075 443 4087 477
rect 4121 443 4144 477
rect 4075 373 4144 443
rect 4075 339 4087 373
rect 4121 339 4144 373
rect 4075 333 4144 339
rect 4180 421 4238 497
rect 4180 387 4192 421
rect 4226 387 4238 421
rect 4180 333 4238 387
rect 4274 477 4328 497
rect 4274 443 4286 477
rect 4320 443 4328 477
rect 4274 379 4328 443
rect 4274 345 4286 379
rect 4320 345 4328 379
rect 4274 333 4328 345
rect 4382 479 4436 497
rect 4382 445 4390 479
rect 4424 445 4436 479
rect 4382 411 4436 445
rect 4382 377 4390 411
rect 4424 377 4436 411
rect 4382 343 4436 377
rect 4075 297 4127 333
rect 4382 309 4390 343
rect 4424 309 4436 343
rect 4382 297 4436 309
rect 4472 479 4544 497
rect 4472 445 4491 479
rect 4525 445 4544 479
rect 4472 411 4544 445
rect 4472 377 4491 411
rect 4525 377 4544 411
rect 4472 343 4544 377
rect 4472 309 4491 343
rect 4525 309 4544 343
rect 4472 297 4544 309
rect 4580 479 4634 497
rect 4580 445 4592 479
rect 4626 445 4634 479
rect 4580 411 4634 445
rect 4580 377 4592 411
rect 4626 377 4634 411
rect 4580 343 4634 377
rect 4580 309 4592 343
rect 4626 309 4634 343
rect 4688 477 4742 497
rect 4688 443 4696 477
rect 4730 443 4742 477
rect 4688 379 4742 443
rect 4688 345 4696 379
rect 4730 345 4742 379
rect 4688 333 4742 345
rect 4778 421 4836 497
rect 4778 387 4790 421
rect 4824 387 4836 421
rect 4778 333 4836 387
rect 4872 477 4941 497
rect 4872 443 4895 477
rect 4929 443 4941 477
rect 4872 373 4941 443
rect 4872 339 4895 373
rect 4929 339 4941 373
rect 4872 333 4941 339
rect 4580 297 4634 309
rect 4889 297 4941 333
rect 4977 485 5035 497
rect 4977 451 4989 485
rect 5023 451 5035 485
rect 4977 405 5035 451
rect 4977 371 4989 405
rect 5023 371 5035 405
rect 4977 297 5035 371
rect 5071 485 5125 497
rect 5071 451 5083 485
rect 5117 451 5125 485
rect 5071 417 5125 451
rect 5071 383 5083 417
rect 5117 383 5125 417
rect 5071 349 5125 383
rect 5071 315 5083 349
rect 5117 315 5125 349
rect 5071 297 5125 315
<< ndiffc >>
rect 45 995 79 1029
rect 45 927 79 961
rect 129 995 163 1029
rect 218 987 252 1021
rect 218 919 252 953
rect 317 935 351 969
rect 401 950 435 984
rect 543 972 577 1006
rect 627 972 661 1006
rect 711 972 745 1006
rect 853 950 887 984
rect 937 935 971 969
rect 1036 987 1070 1021
rect 1036 919 1070 953
rect 1125 995 1159 1029
rect 1209 995 1243 1029
rect 1209 927 1243 961
rect 1333 995 1367 1029
rect 1333 927 1367 961
rect 1417 995 1451 1029
rect 1506 987 1540 1021
rect 1506 919 1540 953
rect 1605 935 1639 969
rect 1689 950 1723 984
rect 1831 972 1865 1006
rect 1915 972 1949 1006
rect 1999 972 2033 1006
rect 2141 950 2175 984
rect 2225 935 2259 969
rect 2324 987 2358 1021
rect 2324 919 2358 953
rect 2413 995 2447 1029
rect 2497 995 2531 1029
rect 2497 927 2531 961
rect 2621 995 2655 1029
rect 2621 927 2655 961
rect 2705 995 2739 1029
rect 2794 987 2828 1021
rect 2794 919 2828 953
rect 2893 935 2927 969
rect 2977 950 3011 984
rect 3119 972 3153 1006
rect 3203 972 3237 1006
rect 3287 972 3321 1006
rect 3429 950 3463 984
rect 3513 935 3547 969
rect 3612 987 3646 1021
rect 3612 919 3646 953
rect 3701 995 3735 1029
rect 3785 995 3819 1029
rect 3785 927 3819 961
rect 3909 995 3943 1029
rect 3909 927 3943 961
rect 3993 995 4027 1029
rect 4082 987 4116 1021
rect 4082 919 4116 953
rect 4181 935 4215 969
rect 4265 950 4299 984
rect 4407 972 4441 1006
rect 4491 972 4525 1006
rect 4575 972 4609 1006
rect 4717 950 4751 984
rect 4801 935 4835 969
rect 4900 987 4934 1021
rect 4900 919 4934 953
rect 4989 995 5023 1029
rect 5073 995 5107 1029
rect 5073 927 5107 961
rect 45 127 79 161
rect 45 59 79 93
rect 129 59 163 93
rect 218 135 252 169
rect 218 67 252 101
rect 317 119 351 153
rect 401 104 435 138
rect 543 82 577 116
rect 627 82 661 116
rect 711 82 745 116
rect 853 104 887 138
rect 937 119 971 153
rect 1036 135 1070 169
rect 1036 67 1070 101
rect 1125 59 1159 93
rect 1209 127 1243 161
rect 1209 59 1243 93
rect 1333 127 1367 161
rect 1333 59 1367 93
rect 1417 59 1451 93
rect 1506 135 1540 169
rect 1506 67 1540 101
rect 1605 119 1639 153
rect 1689 104 1723 138
rect 1831 82 1865 116
rect 1915 82 1949 116
rect 1999 82 2033 116
rect 2141 104 2175 138
rect 2225 119 2259 153
rect 2324 135 2358 169
rect 2324 67 2358 101
rect 2413 59 2447 93
rect 2497 127 2531 161
rect 2497 59 2531 93
rect 2621 127 2655 161
rect 2621 59 2655 93
rect 2705 59 2739 93
rect 2794 135 2828 169
rect 2794 67 2828 101
rect 2893 119 2927 153
rect 2977 104 3011 138
rect 3119 82 3153 116
rect 3203 82 3237 116
rect 3287 82 3321 116
rect 3429 104 3463 138
rect 3513 119 3547 153
rect 3612 135 3646 169
rect 3612 67 3646 101
rect 3701 59 3735 93
rect 3785 127 3819 161
rect 3785 59 3819 93
rect 3909 127 3943 161
rect 3909 59 3943 93
rect 3993 59 4027 93
rect 4082 135 4116 169
rect 4082 67 4116 101
rect 4181 119 4215 153
rect 4265 104 4299 138
rect 4407 82 4441 116
rect 4491 82 4525 116
rect 4575 82 4609 116
rect 4717 104 4751 138
rect 4801 119 4835 153
rect 4900 135 4934 169
rect 4900 67 4934 101
rect 4989 59 5023 93
rect 5073 127 5107 161
rect 5073 59 5107 93
<< pdiffc >>
rect 35 739 69 773
rect 35 671 69 705
rect 35 603 69 637
rect 129 683 163 717
rect 129 603 163 637
rect 223 715 257 749
rect 223 611 257 645
rect 328 667 362 701
rect 422 709 456 743
rect 422 611 456 645
rect 526 745 560 779
rect 526 677 560 711
rect 526 609 560 643
rect 627 745 661 779
rect 627 677 661 711
rect 627 609 661 643
rect 728 745 762 779
rect 728 677 762 711
rect 728 609 762 643
rect 832 709 866 743
rect 832 611 866 645
rect 926 667 960 701
rect 1031 715 1065 749
rect 1031 611 1065 645
rect 1125 683 1159 717
rect 1125 603 1159 637
rect 1219 739 1253 773
rect 1219 671 1253 705
rect 1219 603 1253 637
rect 1323 739 1357 773
rect 1323 671 1357 705
rect 1323 603 1357 637
rect 1417 683 1451 717
rect 1417 603 1451 637
rect 1511 715 1545 749
rect 1511 611 1545 645
rect 1616 667 1650 701
rect 1710 709 1744 743
rect 1710 611 1744 645
rect 1814 745 1848 779
rect 1814 677 1848 711
rect 1814 609 1848 643
rect 1915 745 1949 779
rect 1915 677 1949 711
rect 1915 609 1949 643
rect 2016 745 2050 779
rect 2016 677 2050 711
rect 2016 609 2050 643
rect 2120 709 2154 743
rect 2120 611 2154 645
rect 2214 667 2248 701
rect 2319 715 2353 749
rect 2319 611 2353 645
rect 2413 683 2447 717
rect 2413 603 2447 637
rect 2507 739 2541 773
rect 2507 671 2541 705
rect 2507 603 2541 637
rect 2611 739 2645 773
rect 2611 671 2645 705
rect 2611 603 2645 637
rect 2705 683 2739 717
rect 2705 603 2739 637
rect 2799 715 2833 749
rect 2799 611 2833 645
rect 2904 667 2938 701
rect 2998 709 3032 743
rect 2998 611 3032 645
rect 3102 745 3136 779
rect 3102 677 3136 711
rect 3102 609 3136 643
rect 3203 745 3237 779
rect 3203 677 3237 711
rect 3203 609 3237 643
rect 3304 745 3338 779
rect 3304 677 3338 711
rect 3304 609 3338 643
rect 3408 709 3442 743
rect 3408 611 3442 645
rect 3502 667 3536 701
rect 3607 715 3641 749
rect 3607 611 3641 645
rect 3701 683 3735 717
rect 3701 603 3735 637
rect 3795 739 3829 773
rect 3795 671 3829 705
rect 3795 603 3829 637
rect 3899 739 3933 773
rect 3899 671 3933 705
rect 3899 603 3933 637
rect 3993 683 4027 717
rect 3993 603 4027 637
rect 4087 715 4121 749
rect 4087 611 4121 645
rect 4192 667 4226 701
rect 4286 709 4320 743
rect 4286 611 4320 645
rect 4390 745 4424 779
rect 4390 677 4424 711
rect 4390 609 4424 643
rect 4491 745 4525 779
rect 4491 677 4525 711
rect 4491 609 4525 643
rect 4592 745 4626 779
rect 4592 677 4626 711
rect 4592 609 4626 643
rect 4696 709 4730 743
rect 4696 611 4730 645
rect 4790 667 4824 701
rect 4895 715 4929 749
rect 4895 611 4929 645
rect 4989 683 5023 717
rect 4989 603 5023 637
rect 5083 739 5117 773
rect 5083 671 5117 705
rect 5083 603 5117 637
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 451 163 485
rect 129 371 163 405
rect 223 443 257 477
rect 223 339 257 373
rect 328 387 362 421
rect 422 443 456 477
rect 422 345 456 379
rect 526 445 560 479
rect 526 377 560 411
rect 526 309 560 343
rect 627 445 661 479
rect 627 377 661 411
rect 627 309 661 343
rect 728 445 762 479
rect 728 377 762 411
rect 728 309 762 343
rect 832 443 866 477
rect 832 345 866 379
rect 926 387 960 421
rect 1031 443 1065 477
rect 1031 339 1065 373
rect 1125 451 1159 485
rect 1125 371 1159 405
rect 1219 451 1253 485
rect 1219 383 1253 417
rect 1219 315 1253 349
rect 1323 451 1357 485
rect 1323 383 1357 417
rect 1323 315 1357 349
rect 1417 451 1451 485
rect 1417 371 1451 405
rect 1511 443 1545 477
rect 1511 339 1545 373
rect 1616 387 1650 421
rect 1710 443 1744 477
rect 1710 345 1744 379
rect 1814 445 1848 479
rect 1814 377 1848 411
rect 1814 309 1848 343
rect 1915 445 1949 479
rect 1915 377 1949 411
rect 1915 309 1949 343
rect 2016 445 2050 479
rect 2016 377 2050 411
rect 2016 309 2050 343
rect 2120 443 2154 477
rect 2120 345 2154 379
rect 2214 387 2248 421
rect 2319 443 2353 477
rect 2319 339 2353 373
rect 2413 451 2447 485
rect 2413 371 2447 405
rect 2507 451 2541 485
rect 2507 383 2541 417
rect 2507 315 2541 349
rect 2611 451 2645 485
rect 2611 383 2645 417
rect 2611 315 2645 349
rect 2705 451 2739 485
rect 2705 371 2739 405
rect 2799 443 2833 477
rect 2799 339 2833 373
rect 2904 387 2938 421
rect 2998 443 3032 477
rect 2998 345 3032 379
rect 3102 445 3136 479
rect 3102 377 3136 411
rect 3102 309 3136 343
rect 3203 445 3237 479
rect 3203 377 3237 411
rect 3203 309 3237 343
rect 3304 445 3338 479
rect 3304 377 3338 411
rect 3304 309 3338 343
rect 3408 443 3442 477
rect 3408 345 3442 379
rect 3502 387 3536 421
rect 3607 443 3641 477
rect 3607 339 3641 373
rect 3701 451 3735 485
rect 3701 371 3735 405
rect 3795 451 3829 485
rect 3795 383 3829 417
rect 3795 315 3829 349
rect 3899 451 3933 485
rect 3899 383 3933 417
rect 3899 315 3933 349
rect 3993 451 4027 485
rect 3993 371 4027 405
rect 4087 443 4121 477
rect 4087 339 4121 373
rect 4192 387 4226 421
rect 4286 443 4320 477
rect 4286 345 4320 379
rect 4390 445 4424 479
rect 4390 377 4424 411
rect 4390 309 4424 343
rect 4491 445 4525 479
rect 4491 377 4525 411
rect 4491 309 4525 343
rect 4592 445 4626 479
rect 4592 377 4626 411
rect 4592 309 4626 343
rect 4696 443 4730 477
rect 4696 345 4730 379
rect 4790 387 4824 421
rect 4895 443 4929 477
rect 4895 339 4929 373
rect 4989 451 5023 485
rect 4989 371 5023 405
rect 5083 451 5117 485
rect 5083 383 5117 417
rect 5083 315 5117 349
<< poly >>
rect 89 1041 119 1069
rect 173 1041 203 1067
rect 277 1037 488 1067
rect 587 1041 617 1067
rect 671 1041 701 1067
rect 277 1019 307 1037
rect 361 1019 391 1037
rect 458 919 488 1037
rect 800 1037 1011 1067
rect 1085 1041 1115 1067
rect 1169 1041 1199 1069
rect 1377 1041 1407 1069
rect 1461 1041 1491 1067
rect 587 919 617 937
rect 89 883 119 911
rect 173 883 203 911
rect 277 889 307 915
rect 361 889 391 915
rect 458 889 617 919
rect 671 919 701 937
rect 800 919 830 1037
rect 897 1019 927 1037
rect 981 1019 1011 1037
rect 671 889 830 919
rect 897 889 927 915
rect 981 889 1011 915
rect 1565 1037 1776 1067
rect 1875 1041 1905 1067
rect 1959 1041 1989 1067
rect 1565 1019 1595 1037
rect 1649 1019 1679 1037
rect 1746 919 1776 1037
rect 2088 1037 2299 1067
rect 2373 1041 2403 1067
rect 2457 1041 2487 1069
rect 2665 1041 2695 1069
rect 2749 1041 2779 1067
rect 1875 919 1905 937
rect 49 873 213 883
rect 49 839 65 873
rect 99 839 133 873
rect 167 839 213 873
rect 564 873 618 889
rect 49 829 213 839
rect 420 837 486 847
rect 81 791 117 829
rect 175 791 211 829
rect 420 823 436 837
rect 278 803 436 823
rect 470 803 486 837
rect 564 839 574 873
rect 608 839 618 873
rect 564 823 618 839
rect 670 873 724 889
rect 1085 883 1115 911
rect 1169 883 1199 911
rect 1377 883 1407 911
rect 1461 883 1491 911
rect 1565 889 1595 915
rect 1649 889 1679 915
rect 1746 889 1905 919
rect 1959 919 1989 937
rect 2088 919 2118 1037
rect 2185 1019 2215 1037
rect 2269 1019 2299 1037
rect 1959 889 2118 919
rect 2185 889 2215 915
rect 2269 889 2299 915
rect 2853 1037 3064 1067
rect 3163 1041 3193 1067
rect 3247 1041 3277 1067
rect 2853 1019 2883 1037
rect 2937 1019 2967 1037
rect 3034 919 3064 1037
rect 3376 1037 3587 1067
rect 3661 1041 3691 1067
rect 3745 1041 3775 1069
rect 3953 1041 3983 1069
rect 4037 1041 4067 1067
rect 3163 919 3193 937
rect 670 839 680 873
rect 714 839 724 873
rect 1075 873 1239 883
rect 670 823 724 839
rect 802 837 868 847
rect 570 806 610 823
rect 678 806 718 823
rect 278 793 486 803
rect 280 755 316 793
rect 374 755 410 793
rect 572 791 608 806
rect 680 791 716 806
rect 802 803 818 837
rect 852 823 868 837
rect 1075 839 1121 873
rect 1155 839 1189 873
rect 1223 839 1239 873
rect 1075 829 1239 839
rect 1337 873 1501 883
rect 1337 839 1353 873
rect 1387 839 1421 873
rect 1455 839 1501 873
rect 1852 873 1906 889
rect 1337 829 1501 839
rect 1708 837 1774 847
rect 852 803 1010 823
rect 802 793 1010 803
rect 878 755 914 793
rect 972 755 1008 793
rect 1077 791 1113 829
rect 1171 791 1207 829
rect 1369 791 1405 829
rect 1463 791 1499 829
rect 1708 823 1724 837
rect 1566 803 1724 823
rect 1758 803 1774 837
rect 1852 839 1862 873
rect 1896 839 1906 873
rect 1852 823 1906 839
rect 1958 873 2012 889
rect 2373 883 2403 911
rect 2457 883 2487 911
rect 2665 883 2695 911
rect 2749 883 2779 911
rect 2853 889 2883 915
rect 2937 889 2967 915
rect 3034 889 3193 919
rect 3247 919 3277 937
rect 3376 919 3406 1037
rect 3473 1019 3503 1037
rect 3557 1019 3587 1037
rect 3247 889 3406 919
rect 3473 889 3503 915
rect 3557 889 3587 915
rect 4141 1037 4352 1067
rect 4451 1041 4481 1067
rect 4535 1041 4565 1067
rect 4141 1019 4171 1037
rect 4225 1019 4255 1037
rect 4322 919 4352 1037
rect 4664 1037 4875 1067
rect 4949 1041 4979 1067
rect 5033 1041 5063 1069
rect 4451 919 4481 937
rect 1958 839 1968 873
rect 2002 839 2012 873
rect 2363 873 2527 883
rect 1958 823 2012 839
rect 2090 837 2156 847
rect 1858 806 1898 823
rect 1966 806 2006 823
rect 1566 793 1774 803
rect 1568 755 1604 793
rect 1662 755 1698 793
rect 1860 791 1896 806
rect 1968 791 2004 806
rect 2090 803 2106 837
rect 2140 823 2156 837
rect 2363 839 2409 873
rect 2443 839 2477 873
rect 2511 839 2527 873
rect 2363 829 2527 839
rect 2625 873 2789 883
rect 2625 839 2641 873
rect 2675 839 2709 873
rect 2743 839 2789 873
rect 3140 873 3194 889
rect 2625 829 2789 839
rect 2996 837 3062 847
rect 2140 803 2298 823
rect 2090 793 2298 803
rect 2166 755 2202 793
rect 2260 755 2296 793
rect 2365 791 2401 829
rect 2459 791 2495 829
rect 2657 791 2693 829
rect 2751 791 2787 829
rect 2996 823 3012 837
rect 2854 803 3012 823
rect 3046 803 3062 837
rect 3140 839 3150 873
rect 3184 839 3194 873
rect 3140 823 3194 839
rect 3246 873 3300 889
rect 3661 883 3691 911
rect 3745 883 3775 911
rect 3953 883 3983 911
rect 4037 883 4067 911
rect 4141 889 4171 915
rect 4225 889 4255 915
rect 4322 889 4481 919
rect 4535 919 4565 937
rect 4664 919 4694 1037
rect 4761 1019 4791 1037
rect 4845 1019 4875 1037
rect 4535 889 4694 919
rect 4761 889 4791 915
rect 4845 889 4875 915
rect 3246 839 3256 873
rect 3290 839 3300 873
rect 3651 873 3815 883
rect 3246 823 3300 839
rect 3378 837 3444 847
rect 3146 806 3186 823
rect 3254 806 3294 823
rect 2854 793 3062 803
rect 2856 755 2892 793
rect 2950 755 2986 793
rect 3148 791 3184 806
rect 3256 791 3292 806
rect 3378 803 3394 837
rect 3428 823 3444 837
rect 3651 839 3697 873
rect 3731 839 3765 873
rect 3799 839 3815 873
rect 3651 829 3815 839
rect 3913 873 4077 883
rect 3913 839 3929 873
rect 3963 839 3997 873
rect 4031 839 4077 873
rect 4428 873 4482 889
rect 3913 829 4077 839
rect 4284 837 4350 847
rect 3428 803 3586 823
rect 3378 793 3586 803
rect 3454 755 3490 793
rect 3548 755 3584 793
rect 3653 791 3689 829
rect 3747 791 3783 829
rect 3945 791 3981 829
rect 4039 791 4075 829
rect 4284 823 4300 837
rect 4142 803 4300 823
rect 4334 803 4350 837
rect 4428 839 4438 873
rect 4472 839 4482 873
rect 4428 823 4482 839
rect 4534 873 4588 889
rect 4949 883 4979 911
rect 5033 883 5063 911
rect 4534 839 4544 873
rect 4578 839 4588 873
rect 4939 873 5103 883
rect 4534 823 4588 839
rect 4666 837 4732 847
rect 4434 806 4474 823
rect 4542 806 4582 823
rect 4142 793 4350 803
rect 4144 755 4180 793
rect 4238 755 4274 793
rect 4436 791 4472 806
rect 4544 791 4580 806
rect 4666 803 4682 837
rect 4716 823 4732 837
rect 4939 839 4985 873
rect 5019 839 5053 873
rect 5087 839 5103 873
rect 4939 829 5103 839
rect 4716 803 4874 823
rect 4666 793 4874 803
rect 4742 755 4778 793
rect 4836 755 4872 793
rect 4941 791 4977 829
rect 5035 791 5071 829
rect 81 565 117 591
rect 175 565 211 591
rect 280 565 316 591
rect 374 565 410 591
rect 572 565 608 591
rect 680 565 716 591
rect 878 565 914 591
rect 972 565 1008 591
rect 1077 565 1113 591
rect 1171 565 1207 591
rect 1369 565 1405 591
rect 1463 565 1499 591
rect 1568 565 1604 591
rect 1662 565 1698 591
rect 1860 565 1896 591
rect 1968 565 2004 591
rect 2166 565 2202 591
rect 2260 565 2296 591
rect 2365 565 2401 591
rect 2459 565 2495 591
rect 2657 565 2693 591
rect 2751 565 2787 591
rect 2856 565 2892 591
rect 2950 565 2986 591
rect 3148 565 3184 591
rect 3256 565 3292 591
rect 3454 565 3490 591
rect 3548 565 3584 591
rect 3653 565 3689 591
rect 3747 565 3783 591
rect 3945 565 3981 591
rect 4039 565 4075 591
rect 4144 565 4180 591
rect 4238 565 4274 591
rect 4436 565 4472 591
rect 4544 565 4580 591
rect 4742 565 4778 591
rect 4836 565 4872 591
rect 4941 565 4977 591
rect 5035 565 5071 591
rect 81 497 117 523
rect 175 497 211 523
rect 280 497 316 523
rect 374 497 410 523
rect 572 497 608 523
rect 680 497 716 523
rect 878 497 914 523
rect 972 497 1008 523
rect 1077 497 1113 523
rect 1171 497 1207 523
rect 1369 497 1405 523
rect 1463 497 1499 523
rect 1568 497 1604 523
rect 1662 497 1698 523
rect 1860 497 1896 523
rect 1968 497 2004 523
rect 2166 497 2202 523
rect 2260 497 2296 523
rect 2365 497 2401 523
rect 2459 497 2495 523
rect 2657 497 2693 523
rect 2751 497 2787 523
rect 2856 497 2892 523
rect 2950 497 2986 523
rect 3148 497 3184 523
rect 3256 497 3292 523
rect 3454 497 3490 523
rect 3548 497 3584 523
rect 3653 497 3689 523
rect 3747 497 3783 523
rect 3945 497 3981 523
rect 4039 497 4075 523
rect 4144 497 4180 523
rect 4238 497 4274 523
rect 4436 497 4472 523
rect 4544 497 4580 523
rect 4742 497 4778 523
rect 4836 497 4872 523
rect 4941 497 4977 523
rect 5035 497 5071 523
rect 81 259 117 297
rect 175 259 211 297
rect 280 295 316 333
rect 374 295 410 333
rect 278 285 486 295
rect 278 265 436 285
rect 49 249 213 259
rect 49 215 65 249
rect 99 215 133 249
rect 167 215 213 249
rect 420 251 436 265
rect 470 251 486 285
rect 572 282 608 297
rect 680 282 716 297
rect 878 295 914 333
rect 972 295 1008 333
rect 802 285 1010 295
rect 570 265 610 282
rect 678 265 718 282
rect 420 241 486 251
rect 564 249 618 265
rect 49 205 213 215
rect 564 215 574 249
rect 608 215 618 249
rect 89 177 119 205
rect 173 177 203 205
rect 564 199 618 215
rect 670 249 724 265
rect 670 215 680 249
rect 714 215 724 249
rect 802 251 818 285
rect 852 265 1010 285
rect 852 251 868 265
rect 1077 259 1113 297
rect 1171 259 1207 297
rect 1369 259 1405 297
rect 1463 259 1499 297
rect 1568 295 1604 333
rect 1662 295 1698 333
rect 1566 285 1774 295
rect 1566 265 1724 285
rect 802 241 868 251
rect 1075 249 1239 259
rect 670 199 724 215
rect 1075 215 1121 249
rect 1155 215 1189 249
rect 1223 215 1239 249
rect 1075 205 1239 215
rect 1337 249 1501 259
rect 1337 215 1353 249
rect 1387 215 1421 249
rect 1455 215 1501 249
rect 1708 251 1724 265
rect 1758 251 1774 285
rect 1860 282 1896 297
rect 1968 282 2004 297
rect 2166 295 2202 333
rect 2260 295 2296 333
rect 2090 285 2298 295
rect 1858 265 1898 282
rect 1966 265 2006 282
rect 1708 241 1774 251
rect 1852 249 1906 265
rect 1337 205 1501 215
rect 1852 215 1862 249
rect 1896 215 1906 249
rect 277 173 307 199
rect 361 173 391 199
rect 458 169 617 199
rect 277 51 307 69
rect 361 51 391 69
rect 458 51 488 169
rect 587 151 617 169
rect 671 169 830 199
rect 897 173 927 199
rect 981 173 1011 199
rect 1085 177 1115 205
rect 1169 177 1199 205
rect 1377 177 1407 205
rect 1461 177 1491 205
rect 1852 199 1906 215
rect 1958 249 2012 265
rect 1958 215 1968 249
rect 2002 215 2012 249
rect 2090 251 2106 285
rect 2140 265 2298 285
rect 2140 251 2156 265
rect 2365 259 2401 297
rect 2459 259 2495 297
rect 2657 259 2693 297
rect 2751 259 2787 297
rect 2856 295 2892 333
rect 2950 295 2986 333
rect 2854 285 3062 295
rect 2854 265 3012 285
rect 2090 241 2156 251
rect 2363 249 2527 259
rect 1958 199 2012 215
rect 2363 215 2409 249
rect 2443 215 2477 249
rect 2511 215 2527 249
rect 2363 205 2527 215
rect 2625 249 2789 259
rect 2625 215 2641 249
rect 2675 215 2709 249
rect 2743 215 2789 249
rect 2996 251 3012 265
rect 3046 251 3062 285
rect 3148 282 3184 297
rect 3256 282 3292 297
rect 3454 295 3490 333
rect 3548 295 3584 333
rect 3378 285 3586 295
rect 3146 265 3186 282
rect 3254 265 3294 282
rect 2996 241 3062 251
rect 3140 249 3194 265
rect 2625 205 2789 215
rect 3140 215 3150 249
rect 3184 215 3194 249
rect 671 151 701 169
rect 89 19 119 47
rect 173 21 203 47
rect 277 21 488 51
rect 800 51 830 169
rect 897 51 927 69
rect 981 51 1011 69
rect 587 21 617 47
rect 671 21 701 47
rect 800 21 1011 51
rect 1565 173 1595 199
rect 1649 173 1679 199
rect 1746 169 1905 199
rect 1565 51 1595 69
rect 1649 51 1679 69
rect 1746 51 1776 169
rect 1875 151 1905 169
rect 1959 169 2118 199
rect 2185 173 2215 199
rect 2269 173 2299 199
rect 2373 177 2403 205
rect 2457 177 2487 205
rect 2665 177 2695 205
rect 2749 177 2779 205
rect 3140 199 3194 215
rect 3246 249 3300 265
rect 3246 215 3256 249
rect 3290 215 3300 249
rect 3378 251 3394 285
rect 3428 265 3586 285
rect 3428 251 3444 265
rect 3653 259 3689 297
rect 3747 259 3783 297
rect 3945 259 3981 297
rect 4039 259 4075 297
rect 4144 295 4180 333
rect 4238 295 4274 333
rect 4142 285 4350 295
rect 4142 265 4300 285
rect 3378 241 3444 251
rect 3651 249 3815 259
rect 3246 199 3300 215
rect 3651 215 3697 249
rect 3731 215 3765 249
rect 3799 215 3815 249
rect 3651 205 3815 215
rect 3913 249 4077 259
rect 3913 215 3929 249
rect 3963 215 3997 249
rect 4031 215 4077 249
rect 4284 251 4300 265
rect 4334 251 4350 285
rect 4436 282 4472 297
rect 4544 282 4580 297
rect 4742 295 4778 333
rect 4836 295 4872 333
rect 4666 285 4874 295
rect 4434 265 4474 282
rect 4542 265 4582 282
rect 4284 241 4350 251
rect 4428 249 4482 265
rect 3913 205 4077 215
rect 4428 215 4438 249
rect 4472 215 4482 249
rect 1959 151 1989 169
rect 1085 21 1115 47
rect 1169 19 1199 47
rect 1377 19 1407 47
rect 1461 21 1491 47
rect 1565 21 1776 51
rect 2088 51 2118 169
rect 2185 51 2215 69
rect 2269 51 2299 69
rect 1875 21 1905 47
rect 1959 21 1989 47
rect 2088 21 2299 51
rect 2853 173 2883 199
rect 2937 173 2967 199
rect 3034 169 3193 199
rect 2853 51 2883 69
rect 2937 51 2967 69
rect 3034 51 3064 169
rect 3163 151 3193 169
rect 3247 169 3406 199
rect 3473 173 3503 199
rect 3557 173 3587 199
rect 3661 177 3691 205
rect 3745 177 3775 205
rect 3953 177 3983 205
rect 4037 177 4067 205
rect 4428 199 4482 215
rect 4534 249 4588 265
rect 4534 215 4544 249
rect 4578 215 4588 249
rect 4666 251 4682 285
rect 4716 265 4874 285
rect 4716 251 4732 265
rect 4941 259 4977 297
rect 5035 259 5071 297
rect 4666 241 4732 251
rect 4939 249 5103 259
rect 4534 199 4588 215
rect 4939 215 4985 249
rect 5019 215 5053 249
rect 5087 215 5103 249
rect 4939 205 5103 215
rect 3247 151 3277 169
rect 2373 21 2403 47
rect 2457 19 2487 47
rect 2665 19 2695 47
rect 2749 21 2779 47
rect 2853 21 3064 51
rect 3376 51 3406 169
rect 3473 51 3503 69
rect 3557 51 3587 69
rect 3163 21 3193 47
rect 3247 21 3277 47
rect 3376 21 3587 51
rect 4141 173 4171 199
rect 4225 173 4255 199
rect 4322 169 4481 199
rect 4141 51 4171 69
rect 4225 51 4255 69
rect 4322 51 4352 169
rect 4451 151 4481 169
rect 4535 169 4694 199
rect 4761 173 4791 199
rect 4845 173 4875 199
rect 4949 177 4979 205
rect 5033 177 5063 205
rect 4535 151 4565 169
rect 3661 21 3691 47
rect 3745 19 3775 47
rect 3953 19 3983 47
rect 4037 21 4067 47
rect 4141 21 4352 51
rect 4664 51 4694 169
rect 4761 51 4791 69
rect 4845 51 4875 69
rect 4451 21 4481 47
rect 4535 21 4565 47
rect 4664 21 4875 51
rect 4949 21 4979 47
rect 5033 19 5063 47
<< polycont >>
rect 65 839 99 873
rect 133 839 167 873
rect 436 803 470 837
rect 574 839 608 873
rect 680 839 714 873
rect 818 803 852 837
rect 1121 839 1155 873
rect 1189 839 1223 873
rect 1353 839 1387 873
rect 1421 839 1455 873
rect 1724 803 1758 837
rect 1862 839 1896 873
rect 1968 839 2002 873
rect 2106 803 2140 837
rect 2409 839 2443 873
rect 2477 839 2511 873
rect 2641 839 2675 873
rect 2709 839 2743 873
rect 3012 803 3046 837
rect 3150 839 3184 873
rect 3256 839 3290 873
rect 3394 803 3428 837
rect 3697 839 3731 873
rect 3765 839 3799 873
rect 3929 839 3963 873
rect 3997 839 4031 873
rect 4300 803 4334 837
rect 4438 839 4472 873
rect 4544 839 4578 873
rect 4682 803 4716 837
rect 4985 839 5019 873
rect 5053 839 5087 873
rect 65 215 99 249
rect 133 215 167 249
rect 436 251 470 285
rect 574 215 608 249
rect 680 215 714 249
rect 818 251 852 285
rect 1121 215 1155 249
rect 1189 215 1223 249
rect 1353 215 1387 249
rect 1421 215 1455 249
rect 1724 251 1758 285
rect 1862 215 1896 249
rect 1968 215 2002 249
rect 2106 251 2140 285
rect 2409 215 2443 249
rect 2477 215 2511 249
rect 2641 215 2675 249
rect 2709 215 2743 249
rect 3012 251 3046 285
rect 3150 215 3184 249
rect 3256 215 3290 249
rect 3394 251 3428 285
rect 3697 215 3731 249
rect 3765 215 3799 249
rect 3929 215 3963 249
rect 3997 215 4031 249
rect 4300 251 4334 285
rect 4438 215 4472 249
rect 4544 215 4578 249
rect 4682 251 4716 285
rect 4985 215 5019 249
rect 5053 215 5087 249
<< locali >>
rect 0 1071 29 1105
rect 63 1071 121 1105
rect 155 1071 213 1105
rect 247 1071 305 1105
rect 339 1071 397 1105
rect 431 1071 489 1105
rect 523 1071 581 1105
rect 615 1071 673 1105
rect 707 1071 765 1105
rect 799 1071 857 1105
rect 891 1071 949 1105
rect 983 1071 1041 1105
rect 1075 1071 1133 1105
rect 1167 1071 1225 1105
rect 1259 1071 1317 1105
rect 1351 1071 1409 1105
rect 1443 1071 1501 1105
rect 1535 1071 1593 1105
rect 1627 1071 1685 1105
rect 1719 1071 1777 1105
rect 1811 1071 1869 1105
rect 1903 1071 1961 1105
rect 1995 1071 2053 1105
rect 2087 1071 2145 1105
rect 2179 1071 2237 1105
rect 2271 1071 2329 1105
rect 2363 1071 2421 1105
rect 2455 1071 2513 1105
rect 2547 1071 2605 1105
rect 2639 1071 2697 1105
rect 2731 1071 2789 1105
rect 2823 1071 2881 1105
rect 2915 1071 2973 1105
rect 3007 1071 3065 1105
rect 3099 1071 3157 1105
rect 3191 1071 3249 1105
rect 3283 1071 3341 1105
rect 3375 1071 3433 1105
rect 3467 1071 3525 1105
rect 3559 1071 3617 1105
rect 3651 1071 3709 1105
rect 3743 1071 3801 1105
rect 3835 1071 3893 1105
rect 3927 1071 3985 1105
rect 4019 1071 4077 1105
rect 4111 1071 4169 1105
rect 4203 1071 4261 1105
rect 4295 1071 4353 1105
rect 4387 1071 4445 1105
rect 4479 1071 4537 1105
rect 4571 1071 4629 1105
rect 4663 1071 4721 1105
rect 4755 1071 4813 1105
rect 4847 1071 4905 1105
rect 4939 1071 4997 1105
rect 5031 1071 5089 1105
rect 5123 1071 5152 1105
rect 29 1029 95 1037
rect 29 995 45 1029
rect 79 995 95 1029
rect 29 961 95 995
rect 129 1029 172 1071
rect 163 995 172 1029
rect 129 979 172 995
rect 206 1021 435 1037
rect 206 987 218 1021
rect 252 1003 435 1021
rect 252 987 267 1003
rect 29 927 45 961
rect 79 945 95 961
rect 206 953 267 987
rect 401 984 435 1003
rect 206 945 218 953
rect 79 927 218 945
rect 29 919 218 927
rect 252 919 267 953
rect 29 911 267 919
rect 301 935 317 969
rect 351 935 367 969
rect 301 911 367 935
rect 535 1006 585 1022
rect 535 972 543 1006
rect 577 972 585 1006
rect 535 971 585 972
rect 401 934 435 950
rect 469 937 585 971
rect 619 1006 669 1071
rect 619 972 627 1006
rect 661 972 669 1006
rect 619 956 669 972
rect 703 1006 753 1022
rect 703 972 711 1006
rect 745 972 753 1006
rect 703 971 753 972
rect 853 1021 1082 1037
rect 853 1003 1036 1021
rect 853 984 887 1003
rect 703 937 819 971
rect 206 903 267 911
rect 19 873 183 877
rect 19 839 65 873
rect 99 839 133 873
rect 167 839 183 873
rect 19 823 183 839
rect 19 773 257 789
rect 19 739 35 773
rect 69 755 257 773
rect 69 739 79 755
rect 19 705 79 739
rect 223 749 257 755
rect 19 671 35 705
rect 69 671 79 705
rect 19 660 79 671
rect 113 717 179 721
rect 113 683 129 717
rect 163 683 179 717
rect 113 667 179 683
rect 19 603 35 660
rect 69 646 79 660
rect 69 603 85 646
rect 19 595 85 603
rect 119 637 179 667
rect 119 603 129 637
rect 163 603 179 637
rect 119 561 179 603
rect 317 737 351 911
rect 469 847 503 937
rect 420 837 503 847
rect 420 803 436 837
rect 470 827 503 837
rect 558 873 625 883
rect 558 839 574 873
rect 608 839 625 873
rect 558 829 625 839
rect 663 873 730 883
rect 663 839 680 873
rect 714 839 730 873
rect 663 829 730 839
rect 785 847 819 937
rect 1021 987 1036 1003
rect 1070 987 1082 1021
rect 853 934 887 950
rect 921 935 937 969
rect 971 935 987 969
rect 921 911 987 935
rect 1021 953 1082 987
rect 1116 1029 1159 1071
rect 1116 995 1125 1029
rect 1116 979 1159 995
rect 1193 1029 1259 1037
rect 1193 995 1209 1029
rect 1243 995 1259 1029
rect 1021 919 1036 953
rect 1070 945 1082 953
rect 1193 961 1259 995
rect 1193 945 1209 961
rect 1070 927 1209 945
rect 1243 927 1259 961
rect 1070 919 1259 927
rect 1021 911 1259 919
rect 1317 1029 1383 1037
rect 1317 995 1333 1029
rect 1367 995 1383 1029
rect 1317 961 1383 995
rect 1417 1029 1460 1071
rect 1451 995 1460 1029
rect 1417 979 1460 995
rect 1494 1021 1723 1037
rect 1494 987 1506 1021
rect 1540 1003 1723 1021
rect 1540 987 1555 1003
rect 1317 927 1333 961
rect 1367 945 1383 961
rect 1494 953 1555 987
rect 1689 984 1723 1003
rect 1494 945 1506 953
rect 1367 927 1506 945
rect 1317 919 1506 927
rect 1540 919 1555 953
rect 1317 911 1555 919
rect 1589 935 1605 969
rect 1639 935 1655 969
rect 1589 911 1655 935
rect 1823 1006 1873 1022
rect 1823 972 1831 1006
rect 1865 972 1873 1006
rect 1823 971 1873 972
rect 1689 934 1723 950
rect 1757 937 1873 971
rect 1907 1006 1957 1071
rect 1907 972 1915 1006
rect 1949 972 1957 1006
rect 1907 956 1957 972
rect 1991 1006 2041 1022
rect 1991 972 1999 1006
rect 2033 972 2041 1006
rect 1991 971 2041 972
rect 2141 1021 2370 1037
rect 2141 1003 2324 1021
rect 2141 984 2175 1003
rect 1991 937 2107 971
rect 785 837 868 847
rect 785 827 818 837
rect 470 803 524 827
rect 420 795 524 803
rect 764 803 818 827
rect 852 803 868 837
rect 764 795 868 803
rect 420 793 576 795
rect 490 779 576 793
rect 490 761 526 779
rect 422 743 456 759
rect 223 660 257 715
rect 293 731 379 737
rect 293 697 305 731
rect 339 701 379 731
rect 293 667 328 697
rect 362 667 379 701
rect 293 663 379 667
rect 257 611 283 629
rect 223 595 283 611
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 283 561
rect 19 485 85 493
rect 19 428 35 485
rect 69 442 85 485
rect 119 485 179 527
rect 119 451 129 485
rect 163 451 179 485
rect 69 428 79 442
rect 19 417 79 428
rect 119 421 179 451
rect 19 383 35 417
rect 69 383 79 417
rect 19 349 79 383
rect 113 405 179 421
rect 113 371 129 405
rect 163 371 179 405
rect 113 367 179 371
rect 223 477 283 493
rect 257 459 283 477
rect 223 373 257 428
rect 317 425 351 663
rect 422 660 456 709
rect 385 611 422 629
rect 385 595 456 611
rect 510 745 526 761
rect 560 745 576 779
rect 510 711 576 745
rect 510 677 526 711
rect 560 677 576 711
rect 510 643 576 677
rect 510 609 526 643
rect 560 609 576 643
rect 510 595 576 609
rect 611 779 677 795
rect 611 745 627 779
rect 661 745 677 779
rect 611 711 677 745
rect 611 677 627 711
rect 661 677 677 711
rect 611 643 677 677
rect 611 609 627 643
rect 661 609 677 643
rect 611 561 677 609
rect 712 793 868 795
rect 712 779 798 793
rect 712 745 728 779
rect 762 761 798 779
rect 762 745 778 761
rect 712 711 778 745
rect 712 677 728 711
rect 762 677 778 711
rect 712 643 778 677
rect 712 609 728 643
rect 762 609 778 643
rect 712 595 778 609
rect 832 743 866 759
rect 937 737 971 911
rect 1021 903 1082 911
rect 1494 903 1555 911
rect 1105 873 1269 877
rect 1105 839 1121 873
rect 1155 839 1189 873
rect 1223 839 1269 873
rect 1105 823 1269 839
rect 1307 873 1471 877
rect 1307 839 1353 873
rect 1387 839 1421 873
rect 1455 839 1471 873
rect 1307 823 1471 839
rect 1031 773 1269 789
rect 1031 755 1219 773
rect 1031 749 1065 755
rect 832 660 866 709
rect 909 731 995 737
rect 909 701 949 731
rect 909 667 926 701
rect 983 697 995 731
rect 960 667 995 697
rect 909 663 995 667
rect 1209 739 1219 755
rect 1253 739 1269 773
rect 866 611 903 629
rect 832 595 903 611
rect 385 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 903 561
rect 385 477 456 493
rect 385 459 422 477
rect 19 315 35 349
rect 69 333 79 349
rect 293 421 379 425
rect 293 391 328 421
rect 293 357 305 391
rect 362 387 379 421
rect 339 357 379 387
rect 293 351 379 357
rect 422 379 456 428
rect 223 333 257 339
rect 69 315 257 333
rect 19 299 257 315
rect 19 249 183 265
rect 19 215 65 249
rect 99 215 133 249
rect 167 215 183 249
rect 19 211 183 215
rect 206 177 267 185
rect 317 177 351 351
rect 422 329 456 345
rect 510 479 576 493
rect 510 445 526 479
rect 560 445 576 479
rect 510 411 576 445
rect 510 377 526 411
rect 560 377 576 411
rect 510 343 576 377
rect 510 327 526 343
rect 490 309 526 327
rect 560 309 576 343
rect 490 295 576 309
rect 420 293 576 295
rect 611 479 677 527
rect 611 445 627 479
rect 661 445 677 479
rect 611 411 677 445
rect 611 377 627 411
rect 661 377 677 411
rect 611 343 677 377
rect 611 309 627 343
rect 661 309 677 343
rect 611 293 677 309
rect 712 479 778 493
rect 712 445 728 479
rect 762 445 778 479
rect 712 411 778 445
rect 712 377 728 411
rect 762 377 778 411
rect 712 343 778 377
rect 712 309 728 343
rect 762 327 778 343
rect 832 477 903 493
rect 866 459 903 477
rect 832 379 866 428
rect 937 425 971 663
rect 1031 660 1065 715
rect 1005 611 1031 629
rect 1005 595 1065 611
rect 1109 717 1175 721
rect 1109 683 1125 717
rect 1159 683 1175 717
rect 1109 667 1175 683
rect 1209 705 1269 739
rect 1209 671 1219 705
rect 1253 671 1269 705
rect 1109 637 1169 667
rect 1209 660 1269 671
rect 1209 646 1219 660
rect 1109 603 1125 637
rect 1159 603 1169 637
rect 1109 561 1169 603
rect 1203 603 1219 646
rect 1253 603 1269 660
rect 1203 595 1269 603
rect 1307 773 1545 789
rect 1307 739 1323 773
rect 1357 755 1545 773
rect 1357 739 1367 755
rect 1307 705 1367 739
rect 1511 749 1545 755
rect 1307 671 1323 705
rect 1357 671 1367 705
rect 1307 660 1367 671
rect 1401 717 1467 721
rect 1401 683 1417 717
rect 1451 683 1467 717
rect 1401 667 1467 683
rect 1307 603 1323 660
rect 1357 646 1367 660
rect 1357 603 1373 646
rect 1307 595 1373 603
rect 1407 637 1467 667
rect 1407 603 1417 637
rect 1451 603 1467 637
rect 1407 561 1467 603
rect 1605 737 1639 911
rect 1757 847 1791 937
rect 1708 837 1791 847
rect 1708 803 1724 837
rect 1758 827 1791 837
rect 1846 873 1913 883
rect 1846 839 1862 873
rect 1896 839 1913 873
rect 1846 829 1913 839
rect 1951 873 2018 883
rect 1951 839 1968 873
rect 2002 839 2018 873
rect 1951 829 2018 839
rect 2073 847 2107 937
rect 2309 987 2324 1003
rect 2358 987 2370 1021
rect 2141 934 2175 950
rect 2209 935 2225 969
rect 2259 935 2275 969
rect 2209 911 2275 935
rect 2309 953 2370 987
rect 2404 1029 2447 1071
rect 2404 995 2413 1029
rect 2404 979 2447 995
rect 2481 1029 2547 1037
rect 2481 995 2497 1029
rect 2531 995 2547 1029
rect 2309 919 2324 953
rect 2358 945 2370 953
rect 2481 961 2547 995
rect 2481 945 2497 961
rect 2358 927 2497 945
rect 2531 927 2547 961
rect 2358 919 2547 927
rect 2309 911 2547 919
rect 2605 1029 2671 1037
rect 2605 995 2621 1029
rect 2655 995 2671 1029
rect 2605 961 2671 995
rect 2705 1029 2748 1071
rect 2739 995 2748 1029
rect 2705 979 2748 995
rect 2782 1021 3011 1037
rect 2782 987 2794 1021
rect 2828 1003 3011 1021
rect 2828 987 2843 1003
rect 2605 927 2621 961
rect 2655 945 2671 961
rect 2782 953 2843 987
rect 2977 984 3011 1003
rect 2782 945 2794 953
rect 2655 927 2794 945
rect 2605 919 2794 927
rect 2828 919 2843 953
rect 2605 911 2843 919
rect 2877 935 2893 969
rect 2927 935 2943 969
rect 2877 911 2943 935
rect 3111 1006 3161 1022
rect 3111 972 3119 1006
rect 3153 972 3161 1006
rect 3111 971 3161 972
rect 2977 934 3011 950
rect 3045 937 3161 971
rect 3195 1006 3245 1071
rect 3195 972 3203 1006
rect 3237 972 3245 1006
rect 3195 956 3245 972
rect 3279 1006 3329 1022
rect 3279 972 3287 1006
rect 3321 972 3329 1006
rect 3279 971 3329 972
rect 3429 1021 3658 1037
rect 3429 1003 3612 1021
rect 3429 984 3463 1003
rect 3279 937 3395 971
rect 2073 837 2156 847
rect 2073 827 2106 837
rect 1758 803 1812 827
rect 1708 795 1812 803
rect 2052 803 2106 827
rect 2140 803 2156 837
rect 2052 795 2156 803
rect 1708 793 1864 795
rect 1778 779 1864 793
rect 1778 761 1814 779
rect 1710 743 1744 759
rect 1511 660 1545 715
rect 1581 731 1667 737
rect 1581 697 1593 731
rect 1627 701 1667 731
rect 1581 667 1616 697
rect 1650 667 1667 701
rect 1581 663 1667 667
rect 1545 611 1571 629
rect 1511 595 1571 611
rect 1005 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1571 561
rect 1005 477 1065 493
rect 1005 459 1031 477
rect 909 421 995 425
rect 909 387 926 421
rect 960 391 995 421
rect 909 357 949 387
rect 983 357 995 391
rect 909 351 995 357
rect 1031 373 1065 428
rect 832 329 866 345
rect 762 309 798 327
rect 712 295 798 309
rect 712 293 868 295
rect 420 285 524 293
rect 420 251 436 285
rect 470 261 524 285
rect 764 285 868 293
rect 764 261 818 285
rect 470 251 503 261
rect 420 241 503 251
rect 29 169 267 177
rect 29 161 218 169
rect 29 127 45 161
rect 79 143 218 161
rect 79 127 95 143
rect 29 93 95 127
rect 206 135 218 143
rect 252 135 267 169
rect 29 59 45 93
rect 79 59 95 93
rect 29 51 95 59
rect 129 93 172 109
rect 163 59 172 93
rect 129 17 172 59
rect 206 101 267 135
rect 301 153 367 177
rect 301 119 317 153
rect 351 119 367 153
rect 401 138 435 154
rect 206 67 218 101
rect 252 85 267 101
rect 469 151 503 241
rect 558 249 625 259
rect 558 215 574 249
rect 608 215 625 249
rect 558 205 625 215
rect 663 249 730 259
rect 663 215 680 249
rect 714 215 730 249
rect 663 205 730 215
rect 785 251 818 261
rect 852 251 868 285
rect 785 241 868 251
rect 785 151 819 241
rect 937 177 971 351
rect 1109 485 1169 527
rect 1109 451 1125 485
rect 1159 451 1169 485
rect 1109 421 1169 451
rect 1203 485 1269 493
rect 1203 442 1219 485
rect 1209 428 1219 442
rect 1253 428 1269 485
rect 1109 405 1175 421
rect 1109 371 1125 405
rect 1159 371 1175 405
rect 1109 367 1175 371
rect 1209 417 1269 428
rect 1209 383 1219 417
rect 1253 383 1269 417
rect 1031 333 1065 339
rect 1209 349 1269 383
rect 1209 333 1219 349
rect 1031 315 1219 333
rect 1253 315 1269 349
rect 1031 299 1269 315
rect 1307 485 1373 493
rect 1307 428 1323 485
rect 1357 442 1373 485
rect 1407 485 1467 527
rect 1407 451 1417 485
rect 1451 451 1467 485
rect 1357 428 1367 442
rect 1307 417 1367 428
rect 1407 421 1467 451
rect 1307 383 1323 417
rect 1357 383 1367 417
rect 1307 349 1367 383
rect 1401 405 1467 421
rect 1401 371 1417 405
rect 1451 371 1467 405
rect 1401 367 1467 371
rect 1511 477 1571 493
rect 1545 459 1571 477
rect 1511 373 1545 428
rect 1605 425 1639 663
rect 1710 660 1744 709
rect 1673 611 1710 629
rect 1673 595 1744 611
rect 1798 745 1814 761
rect 1848 745 1864 779
rect 1798 711 1864 745
rect 1798 677 1814 711
rect 1848 677 1864 711
rect 1798 643 1864 677
rect 1798 609 1814 643
rect 1848 609 1864 643
rect 1798 595 1864 609
rect 1899 779 1965 795
rect 1899 745 1915 779
rect 1949 745 1965 779
rect 1899 711 1965 745
rect 1899 677 1915 711
rect 1949 677 1965 711
rect 1899 643 1965 677
rect 1899 609 1915 643
rect 1949 609 1965 643
rect 1899 561 1965 609
rect 2000 793 2156 795
rect 2000 779 2086 793
rect 2000 745 2016 779
rect 2050 761 2086 779
rect 2050 745 2066 761
rect 2000 711 2066 745
rect 2000 677 2016 711
rect 2050 677 2066 711
rect 2000 643 2066 677
rect 2000 609 2016 643
rect 2050 609 2066 643
rect 2000 595 2066 609
rect 2120 743 2154 759
rect 2225 737 2259 911
rect 2309 903 2370 911
rect 2782 903 2843 911
rect 2393 873 2557 877
rect 2393 839 2409 873
rect 2443 839 2477 873
rect 2511 839 2557 873
rect 2393 823 2557 839
rect 2595 873 2759 877
rect 2595 839 2641 873
rect 2675 839 2709 873
rect 2743 839 2759 873
rect 2595 823 2759 839
rect 2319 773 2557 789
rect 2319 755 2507 773
rect 2319 749 2353 755
rect 2120 660 2154 709
rect 2197 731 2283 737
rect 2197 701 2237 731
rect 2197 667 2214 701
rect 2271 697 2283 731
rect 2248 667 2283 697
rect 2197 663 2283 667
rect 2497 739 2507 755
rect 2541 739 2557 773
rect 2154 611 2191 629
rect 2120 595 2191 611
rect 1673 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2191 561
rect 1673 477 1744 493
rect 1673 459 1710 477
rect 1307 315 1323 349
rect 1357 333 1367 349
rect 1581 421 1667 425
rect 1581 391 1616 421
rect 1581 357 1593 391
rect 1650 387 1667 421
rect 1627 357 1667 387
rect 1581 351 1667 357
rect 1710 379 1744 428
rect 1511 333 1545 339
rect 1357 315 1545 333
rect 1307 299 1545 315
rect 1105 249 1269 265
rect 1105 215 1121 249
rect 1155 215 1189 249
rect 1223 215 1269 249
rect 1105 211 1269 215
rect 1307 249 1471 265
rect 1307 215 1353 249
rect 1387 215 1421 249
rect 1455 215 1471 249
rect 1307 211 1471 215
rect 1021 177 1082 185
rect 1494 177 1555 185
rect 1605 177 1639 351
rect 1710 329 1744 345
rect 1798 479 1864 493
rect 1798 445 1814 479
rect 1848 445 1864 479
rect 1798 411 1864 445
rect 1798 377 1814 411
rect 1848 377 1864 411
rect 1798 343 1864 377
rect 1798 327 1814 343
rect 1778 309 1814 327
rect 1848 309 1864 343
rect 1778 295 1864 309
rect 1708 293 1864 295
rect 1899 479 1965 527
rect 1899 445 1915 479
rect 1949 445 1965 479
rect 1899 411 1965 445
rect 1899 377 1915 411
rect 1949 377 1965 411
rect 1899 343 1965 377
rect 1899 309 1915 343
rect 1949 309 1965 343
rect 1899 293 1965 309
rect 2000 479 2066 493
rect 2000 445 2016 479
rect 2050 445 2066 479
rect 2000 411 2066 445
rect 2000 377 2016 411
rect 2050 377 2066 411
rect 2000 343 2066 377
rect 2000 309 2016 343
rect 2050 327 2066 343
rect 2120 477 2191 493
rect 2154 459 2191 477
rect 2120 379 2154 428
rect 2225 425 2259 663
rect 2319 660 2353 715
rect 2293 611 2319 629
rect 2293 595 2353 611
rect 2397 717 2463 721
rect 2397 683 2413 717
rect 2447 683 2463 717
rect 2397 667 2463 683
rect 2497 705 2557 739
rect 2497 671 2507 705
rect 2541 671 2557 705
rect 2397 637 2457 667
rect 2497 660 2557 671
rect 2497 646 2507 660
rect 2397 603 2413 637
rect 2447 603 2457 637
rect 2397 561 2457 603
rect 2491 603 2507 646
rect 2541 603 2557 660
rect 2491 595 2557 603
rect 2595 773 2833 789
rect 2595 739 2611 773
rect 2645 755 2833 773
rect 2645 739 2655 755
rect 2595 705 2655 739
rect 2799 749 2833 755
rect 2595 671 2611 705
rect 2645 671 2655 705
rect 2595 660 2655 671
rect 2689 717 2755 721
rect 2689 683 2705 717
rect 2739 683 2755 717
rect 2689 667 2755 683
rect 2595 603 2611 660
rect 2645 646 2655 660
rect 2645 603 2661 646
rect 2595 595 2661 603
rect 2695 637 2755 667
rect 2695 603 2705 637
rect 2739 603 2755 637
rect 2695 561 2755 603
rect 2893 737 2927 911
rect 3045 847 3079 937
rect 2996 837 3079 847
rect 2996 803 3012 837
rect 3046 827 3079 837
rect 3134 873 3201 883
rect 3134 839 3150 873
rect 3184 839 3201 873
rect 3134 829 3201 839
rect 3239 873 3306 883
rect 3239 839 3256 873
rect 3290 839 3306 873
rect 3239 829 3306 839
rect 3361 847 3395 937
rect 3597 987 3612 1003
rect 3646 987 3658 1021
rect 3429 934 3463 950
rect 3497 935 3513 969
rect 3547 935 3563 969
rect 3497 911 3563 935
rect 3597 953 3658 987
rect 3692 1029 3735 1071
rect 3692 995 3701 1029
rect 3692 979 3735 995
rect 3769 1029 3835 1037
rect 3769 995 3785 1029
rect 3819 995 3835 1029
rect 3597 919 3612 953
rect 3646 945 3658 953
rect 3769 961 3835 995
rect 3769 945 3785 961
rect 3646 927 3785 945
rect 3819 927 3835 961
rect 3646 919 3835 927
rect 3597 911 3835 919
rect 3893 1029 3959 1037
rect 3893 995 3909 1029
rect 3943 995 3959 1029
rect 3893 961 3959 995
rect 3993 1029 4036 1071
rect 4027 995 4036 1029
rect 3993 979 4036 995
rect 4070 1021 4299 1037
rect 4070 987 4082 1021
rect 4116 1003 4299 1021
rect 4116 987 4131 1003
rect 3893 927 3909 961
rect 3943 945 3959 961
rect 4070 953 4131 987
rect 4265 984 4299 1003
rect 4070 945 4082 953
rect 3943 927 4082 945
rect 3893 919 4082 927
rect 4116 919 4131 953
rect 3893 911 4131 919
rect 4165 935 4181 969
rect 4215 935 4231 969
rect 4165 911 4231 935
rect 4399 1006 4449 1022
rect 4399 972 4407 1006
rect 4441 972 4449 1006
rect 4399 971 4449 972
rect 4265 934 4299 950
rect 4333 937 4449 971
rect 4483 1006 4533 1071
rect 4483 972 4491 1006
rect 4525 972 4533 1006
rect 4483 956 4533 972
rect 4567 1006 4617 1022
rect 4567 972 4575 1006
rect 4609 972 4617 1006
rect 4567 971 4617 972
rect 4717 1021 4946 1037
rect 4717 1003 4900 1021
rect 4717 984 4751 1003
rect 4567 937 4683 971
rect 3361 837 3444 847
rect 3361 827 3394 837
rect 3046 803 3100 827
rect 2996 795 3100 803
rect 3340 803 3394 827
rect 3428 803 3444 837
rect 3340 795 3444 803
rect 2996 793 3152 795
rect 3066 779 3152 793
rect 3066 761 3102 779
rect 2998 743 3032 759
rect 2799 660 2833 715
rect 2869 731 2955 737
rect 2869 697 2881 731
rect 2915 701 2955 731
rect 2869 667 2904 697
rect 2938 667 2955 701
rect 2869 663 2955 667
rect 2833 611 2859 629
rect 2799 595 2859 611
rect 2293 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2859 561
rect 2293 477 2353 493
rect 2293 459 2319 477
rect 2197 421 2283 425
rect 2197 387 2214 421
rect 2248 391 2283 421
rect 2197 357 2237 387
rect 2271 357 2283 391
rect 2197 351 2283 357
rect 2319 373 2353 428
rect 2120 329 2154 345
rect 2050 309 2086 327
rect 2000 295 2086 309
rect 2000 293 2156 295
rect 1708 285 1812 293
rect 1708 251 1724 285
rect 1758 261 1812 285
rect 2052 285 2156 293
rect 2052 261 2106 285
rect 1758 251 1791 261
rect 1708 241 1791 251
rect 469 117 585 151
rect 401 85 435 104
rect 252 67 435 85
rect 206 51 435 67
rect 535 116 585 117
rect 535 82 543 116
rect 577 82 585 116
rect 535 66 585 82
rect 619 116 669 132
rect 619 82 627 116
rect 661 82 669 116
rect 619 17 669 82
rect 703 117 819 151
rect 853 138 887 154
rect 703 116 753 117
rect 703 82 711 116
rect 745 82 753 116
rect 703 66 753 82
rect 921 153 987 177
rect 921 119 937 153
rect 971 119 987 153
rect 1021 169 1259 177
rect 1021 135 1036 169
rect 1070 161 1259 169
rect 1070 143 1209 161
rect 1070 135 1082 143
rect 853 85 887 104
rect 1021 101 1082 135
rect 1193 127 1209 143
rect 1243 127 1259 161
rect 1021 85 1036 101
rect 853 67 1036 85
rect 1070 67 1082 101
rect 853 51 1082 67
rect 1116 93 1159 109
rect 1116 59 1125 93
rect 1116 17 1159 59
rect 1193 93 1259 127
rect 1193 59 1209 93
rect 1243 59 1259 93
rect 1193 51 1259 59
rect 1317 169 1555 177
rect 1317 161 1506 169
rect 1317 127 1333 161
rect 1367 143 1506 161
rect 1367 127 1383 143
rect 1317 93 1383 127
rect 1494 135 1506 143
rect 1540 135 1555 169
rect 1317 59 1333 93
rect 1367 59 1383 93
rect 1317 51 1383 59
rect 1417 93 1460 109
rect 1451 59 1460 93
rect 1417 17 1460 59
rect 1494 101 1555 135
rect 1589 153 1655 177
rect 1589 119 1605 153
rect 1639 119 1655 153
rect 1689 138 1723 154
rect 1494 67 1506 101
rect 1540 85 1555 101
rect 1757 151 1791 241
rect 1846 249 1913 259
rect 1846 215 1862 249
rect 1896 215 1913 249
rect 1846 205 1913 215
rect 1951 249 2018 259
rect 1951 215 1968 249
rect 2002 215 2018 249
rect 1951 205 2018 215
rect 2073 251 2106 261
rect 2140 251 2156 285
rect 2073 241 2156 251
rect 2073 151 2107 241
rect 2225 177 2259 351
rect 2397 485 2457 527
rect 2397 451 2413 485
rect 2447 451 2457 485
rect 2397 421 2457 451
rect 2491 485 2557 493
rect 2491 442 2507 485
rect 2497 428 2507 442
rect 2541 428 2557 485
rect 2397 405 2463 421
rect 2397 371 2413 405
rect 2447 371 2463 405
rect 2397 367 2463 371
rect 2497 417 2557 428
rect 2497 383 2507 417
rect 2541 383 2557 417
rect 2319 333 2353 339
rect 2497 349 2557 383
rect 2497 333 2507 349
rect 2319 315 2507 333
rect 2541 315 2557 349
rect 2319 299 2557 315
rect 2595 485 2661 493
rect 2595 428 2611 485
rect 2645 442 2661 485
rect 2695 485 2755 527
rect 2695 451 2705 485
rect 2739 451 2755 485
rect 2645 428 2655 442
rect 2595 417 2655 428
rect 2695 421 2755 451
rect 2595 383 2611 417
rect 2645 383 2655 417
rect 2595 349 2655 383
rect 2689 405 2755 421
rect 2689 371 2705 405
rect 2739 371 2755 405
rect 2689 367 2755 371
rect 2799 477 2859 493
rect 2833 459 2859 477
rect 2799 373 2833 428
rect 2893 425 2927 663
rect 2998 660 3032 709
rect 2961 611 2998 629
rect 2961 595 3032 611
rect 3086 745 3102 761
rect 3136 745 3152 779
rect 3086 711 3152 745
rect 3086 677 3102 711
rect 3136 677 3152 711
rect 3086 643 3152 677
rect 3086 609 3102 643
rect 3136 609 3152 643
rect 3086 595 3152 609
rect 3187 779 3253 795
rect 3187 745 3203 779
rect 3237 745 3253 779
rect 3187 711 3253 745
rect 3187 677 3203 711
rect 3237 677 3253 711
rect 3187 643 3253 677
rect 3187 609 3203 643
rect 3237 609 3253 643
rect 3187 561 3253 609
rect 3288 793 3444 795
rect 3288 779 3374 793
rect 3288 745 3304 779
rect 3338 761 3374 779
rect 3338 745 3354 761
rect 3288 711 3354 745
rect 3288 677 3304 711
rect 3338 677 3354 711
rect 3288 643 3354 677
rect 3288 609 3304 643
rect 3338 609 3354 643
rect 3288 595 3354 609
rect 3408 743 3442 759
rect 3513 737 3547 911
rect 3597 903 3658 911
rect 4070 903 4131 911
rect 3681 873 3845 877
rect 3681 839 3697 873
rect 3731 839 3765 873
rect 3799 839 3845 873
rect 3681 823 3845 839
rect 3883 873 4047 877
rect 3883 839 3929 873
rect 3963 839 3997 873
rect 4031 839 4047 873
rect 3883 823 4047 839
rect 3607 773 3845 789
rect 3607 755 3795 773
rect 3607 749 3641 755
rect 3408 660 3442 709
rect 3485 731 3571 737
rect 3485 701 3525 731
rect 3485 667 3502 701
rect 3559 697 3571 731
rect 3536 667 3571 697
rect 3485 663 3571 667
rect 3785 739 3795 755
rect 3829 739 3845 773
rect 3442 611 3479 629
rect 3408 595 3479 611
rect 2961 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3157 561
rect 3191 527 3249 561
rect 3283 527 3341 561
rect 3375 527 3433 561
rect 3467 527 3479 561
rect 2961 477 3032 493
rect 2961 459 2998 477
rect 2595 315 2611 349
rect 2645 333 2655 349
rect 2869 421 2955 425
rect 2869 391 2904 421
rect 2869 357 2881 391
rect 2938 387 2955 421
rect 2915 357 2955 387
rect 2869 351 2955 357
rect 2998 379 3032 428
rect 2799 333 2833 339
rect 2645 315 2833 333
rect 2595 299 2833 315
rect 2393 249 2557 265
rect 2393 215 2409 249
rect 2443 215 2477 249
rect 2511 215 2557 249
rect 2393 211 2557 215
rect 2595 249 2759 265
rect 2595 215 2641 249
rect 2675 215 2709 249
rect 2743 215 2759 249
rect 2595 211 2759 215
rect 2309 177 2370 185
rect 2782 177 2843 185
rect 2893 177 2927 351
rect 2998 329 3032 345
rect 3086 479 3152 493
rect 3086 445 3102 479
rect 3136 445 3152 479
rect 3086 411 3152 445
rect 3086 377 3102 411
rect 3136 377 3152 411
rect 3086 343 3152 377
rect 3086 327 3102 343
rect 3066 309 3102 327
rect 3136 309 3152 343
rect 3066 295 3152 309
rect 2996 293 3152 295
rect 3187 479 3253 527
rect 3187 445 3203 479
rect 3237 445 3253 479
rect 3187 411 3253 445
rect 3187 377 3203 411
rect 3237 377 3253 411
rect 3187 343 3253 377
rect 3187 309 3203 343
rect 3237 309 3253 343
rect 3187 293 3253 309
rect 3288 479 3354 493
rect 3288 445 3304 479
rect 3338 445 3354 479
rect 3288 411 3354 445
rect 3288 377 3304 411
rect 3338 377 3354 411
rect 3288 343 3354 377
rect 3288 309 3304 343
rect 3338 327 3354 343
rect 3408 477 3479 493
rect 3442 459 3479 477
rect 3408 379 3442 428
rect 3513 425 3547 663
rect 3607 660 3641 715
rect 3581 611 3607 629
rect 3581 595 3641 611
rect 3685 717 3751 721
rect 3685 683 3701 717
rect 3735 683 3751 717
rect 3685 667 3751 683
rect 3785 705 3845 739
rect 3785 671 3795 705
rect 3829 671 3845 705
rect 3685 637 3745 667
rect 3785 660 3845 671
rect 3785 646 3795 660
rect 3685 603 3701 637
rect 3735 603 3745 637
rect 3685 561 3745 603
rect 3779 603 3795 646
rect 3829 603 3845 660
rect 3779 595 3845 603
rect 3883 773 4121 789
rect 3883 739 3899 773
rect 3933 755 4121 773
rect 3933 739 3943 755
rect 3883 705 3943 739
rect 4087 749 4121 755
rect 3883 671 3899 705
rect 3933 671 3943 705
rect 3883 660 3943 671
rect 3977 717 4043 721
rect 3977 683 3993 717
rect 4027 683 4043 717
rect 3977 667 4043 683
rect 3883 603 3899 660
rect 3933 646 3943 660
rect 3933 603 3949 646
rect 3883 595 3949 603
rect 3983 637 4043 667
rect 3983 603 3993 637
rect 4027 603 4043 637
rect 3983 561 4043 603
rect 4181 737 4215 911
rect 4333 847 4367 937
rect 4284 837 4367 847
rect 4284 803 4300 837
rect 4334 827 4367 837
rect 4422 873 4489 883
rect 4422 839 4438 873
rect 4472 839 4489 873
rect 4422 829 4489 839
rect 4527 873 4594 883
rect 4527 839 4544 873
rect 4578 839 4594 873
rect 4527 829 4594 839
rect 4649 847 4683 937
rect 4885 987 4900 1003
rect 4934 987 4946 1021
rect 4717 934 4751 950
rect 4785 935 4801 969
rect 4835 935 4851 969
rect 4785 911 4851 935
rect 4885 953 4946 987
rect 4980 1029 5023 1071
rect 4980 995 4989 1029
rect 4980 979 5023 995
rect 5057 1029 5123 1037
rect 5057 995 5073 1029
rect 5107 995 5123 1029
rect 4885 919 4900 953
rect 4934 945 4946 953
rect 5057 961 5123 995
rect 5057 945 5073 961
rect 4934 927 5073 945
rect 5107 927 5123 961
rect 4934 919 5123 927
rect 4885 911 5123 919
rect 4649 837 4732 847
rect 4649 827 4682 837
rect 4334 803 4388 827
rect 4284 795 4388 803
rect 4628 803 4682 827
rect 4716 803 4732 837
rect 4628 795 4732 803
rect 4284 793 4440 795
rect 4354 779 4440 793
rect 4354 761 4390 779
rect 4286 743 4320 759
rect 4087 660 4121 715
rect 4157 731 4243 737
rect 4157 697 4169 731
rect 4203 701 4243 731
rect 4157 667 4192 697
rect 4226 667 4243 701
rect 4157 663 4243 667
rect 4121 611 4147 629
rect 4087 595 4147 611
rect 3581 527 3617 561
rect 3651 527 3709 561
rect 3743 527 3801 561
rect 3835 527 3893 561
rect 3927 527 3985 561
rect 4019 527 4077 561
rect 4111 527 4147 561
rect 3581 477 3641 493
rect 3581 459 3607 477
rect 3485 421 3571 425
rect 3485 387 3502 421
rect 3536 391 3571 421
rect 3485 357 3525 387
rect 3559 357 3571 391
rect 3485 351 3571 357
rect 3607 373 3641 428
rect 3408 329 3442 345
rect 3338 309 3374 327
rect 3288 295 3374 309
rect 3288 293 3444 295
rect 2996 285 3100 293
rect 2996 251 3012 285
rect 3046 261 3100 285
rect 3340 285 3444 293
rect 3340 261 3394 285
rect 3046 251 3079 261
rect 2996 241 3079 251
rect 1757 117 1873 151
rect 1689 85 1723 104
rect 1540 67 1723 85
rect 1494 51 1723 67
rect 1823 116 1873 117
rect 1823 82 1831 116
rect 1865 82 1873 116
rect 1823 66 1873 82
rect 1907 116 1957 132
rect 1907 82 1915 116
rect 1949 82 1957 116
rect 1907 17 1957 82
rect 1991 117 2107 151
rect 2141 138 2175 154
rect 1991 116 2041 117
rect 1991 82 1999 116
rect 2033 82 2041 116
rect 1991 66 2041 82
rect 2209 153 2275 177
rect 2209 119 2225 153
rect 2259 119 2275 153
rect 2309 169 2547 177
rect 2309 135 2324 169
rect 2358 161 2547 169
rect 2358 143 2497 161
rect 2358 135 2370 143
rect 2141 85 2175 104
rect 2309 101 2370 135
rect 2481 127 2497 143
rect 2531 127 2547 161
rect 2309 85 2324 101
rect 2141 67 2324 85
rect 2358 67 2370 101
rect 2141 51 2370 67
rect 2404 93 2447 109
rect 2404 59 2413 93
rect 2404 17 2447 59
rect 2481 93 2547 127
rect 2481 59 2497 93
rect 2531 59 2547 93
rect 2481 51 2547 59
rect 2605 169 2843 177
rect 2605 161 2794 169
rect 2605 127 2621 161
rect 2655 143 2794 161
rect 2655 127 2671 143
rect 2605 93 2671 127
rect 2782 135 2794 143
rect 2828 135 2843 169
rect 2605 59 2621 93
rect 2655 59 2671 93
rect 2605 51 2671 59
rect 2705 93 2748 109
rect 2739 59 2748 93
rect 2705 17 2748 59
rect 2782 101 2843 135
rect 2877 153 2943 177
rect 2877 119 2893 153
rect 2927 119 2943 153
rect 2977 138 3011 154
rect 2782 67 2794 101
rect 2828 85 2843 101
rect 3045 151 3079 241
rect 3134 249 3201 259
rect 3134 215 3150 249
rect 3184 215 3201 249
rect 3134 205 3201 215
rect 3239 249 3306 259
rect 3239 215 3256 249
rect 3290 215 3306 249
rect 3239 205 3306 215
rect 3361 251 3394 261
rect 3428 251 3444 285
rect 3361 241 3444 251
rect 3361 151 3395 241
rect 3513 177 3547 351
rect 3685 485 3745 527
rect 3685 451 3701 485
rect 3735 451 3745 485
rect 3685 421 3745 451
rect 3779 485 3845 493
rect 3779 442 3795 485
rect 3785 428 3795 442
rect 3829 428 3845 485
rect 3685 405 3751 421
rect 3685 371 3701 405
rect 3735 371 3751 405
rect 3685 367 3751 371
rect 3785 417 3845 428
rect 3785 383 3795 417
rect 3829 383 3845 417
rect 3607 333 3641 339
rect 3785 349 3845 383
rect 3785 333 3795 349
rect 3607 315 3795 333
rect 3829 315 3845 349
rect 3607 299 3845 315
rect 3883 485 3949 493
rect 3883 428 3899 485
rect 3933 442 3949 485
rect 3983 485 4043 527
rect 3983 451 3993 485
rect 4027 451 4043 485
rect 3933 428 3943 442
rect 3883 417 3943 428
rect 3983 421 4043 451
rect 3883 383 3899 417
rect 3933 383 3943 417
rect 3883 349 3943 383
rect 3977 405 4043 421
rect 3977 371 3993 405
rect 4027 371 4043 405
rect 3977 367 4043 371
rect 4087 477 4147 493
rect 4121 459 4147 477
rect 4087 373 4121 428
rect 4181 425 4215 663
rect 4286 660 4320 709
rect 4249 611 4286 629
rect 4249 595 4320 611
rect 4374 745 4390 761
rect 4424 745 4440 779
rect 4374 711 4440 745
rect 4374 677 4390 711
rect 4424 677 4440 711
rect 4374 643 4440 677
rect 4374 609 4390 643
rect 4424 609 4440 643
rect 4374 595 4440 609
rect 4475 779 4541 795
rect 4475 745 4491 779
rect 4525 745 4541 779
rect 4475 711 4541 745
rect 4475 677 4491 711
rect 4525 677 4541 711
rect 4475 643 4541 677
rect 4475 609 4491 643
rect 4525 609 4541 643
rect 4475 561 4541 609
rect 4576 793 4732 795
rect 4576 779 4662 793
rect 4576 745 4592 779
rect 4626 761 4662 779
rect 4626 745 4642 761
rect 4576 711 4642 745
rect 4576 677 4592 711
rect 4626 677 4642 711
rect 4576 643 4642 677
rect 4576 609 4592 643
rect 4626 609 4642 643
rect 4576 595 4642 609
rect 4696 743 4730 759
rect 4801 737 4835 911
rect 4885 903 4946 911
rect 4969 873 5133 877
rect 4969 839 4985 873
rect 5019 839 5053 873
rect 5087 839 5133 873
rect 4969 823 5133 839
rect 4895 773 5133 789
rect 4895 755 5083 773
rect 4895 749 4929 755
rect 4696 660 4730 709
rect 4773 731 4859 737
rect 4773 701 4813 731
rect 4773 667 4790 701
rect 4847 697 4859 731
rect 4824 667 4859 697
rect 4773 663 4859 667
rect 5073 739 5083 755
rect 5117 739 5133 773
rect 4730 611 4767 629
rect 4696 595 4767 611
rect 4249 527 4261 561
rect 4295 527 4353 561
rect 4387 527 4445 561
rect 4479 527 4537 561
rect 4571 527 4629 561
rect 4663 527 4721 561
rect 4755 527 4767 561
rect 4249 477 4320 493
rect 4249 459 4286 477
rect 3883 315 3899 349
rect 3933 333 3943 349
rect 4157 421 4243 425
rect 4157 391 4192 421
rect 4157 357 4169 391
rect 4226 387 4243 421
rect 4203 357 4243 387
rect 4157 351 4243 357
rect 4286 379 4320 428
rect 4087 333 4121 339
rect 3933 315 4121 333
rect 3883 299 4121 315
rect 3681 249 3845 265
rect 3681 215 3697 249
rect 3731 215 3765 249
rect 3799 215 3845 249
rect 3681 211 3845 215
rect 3883 249 4047 265
rect 3883 215 3929 249
rect 3963 215 3997 249
rect 4031 215 4047 249
rect 3883 211 4047 215
rect 3597 177 3658 185
rect 4070 177 4131 185
rect 4181 177 4215 351
rect 4286 329 4320 345
rect 4374 479 4440 493
rect 4374 445 4390 479
rect 4424 445 4440 479
rect 4374 411 4440 445
rect 4374 377 4390 411
rect 4424 377 4440 411
rect 4374 343 4440 377
rect 4374 327 4390 343
rect 4354 309 4390 327
rect 4424 309 4440 343
rect 4354 295 4440 309
rect 4284 293 4440 295
rect 4475 479 4541 527
rect 4475 445 4491 479
rect 4525 445 4541 479
rect 4475 411 4541 445
rect 4475 377 4491 411
rect 4525 377 4541 411
rect 4475 343 4541 377
rect 4475 309 4491 343
rect 4525 309 4541 343
rect 4475 293 4541 309
rect 4576 479 4642 493
rect 4576 445 4592 479
rect 4626 445 4642 479
rect 4576 411 4642 445
rect 4576 377 4592 411
rect 4626 377 4642 411
rect 4576 343 4642 377
rect 4576 309 4592 343
rect 4626 327 4642 343
rect 4696 477 4767 493
rect 4730 459 4767 477
rect 4696 379 4730 428
rect 4801 425 4835 663
rect 4895 660 4929 715
rect 4869 611 4895 629
rect 4869 595 4929 611
rect 4973 717 5039 721
rect 4973 683 4989 717
rect 5023 683 5039 717
rect 4973 667 5039 683
rect 5073 705 5133 739
rect 5073 671 5083 705
rect 5117 671 5133 705
rect 4973 637 5033 667
rect 5073 660 5133 671
rect 5073 646 5083 660
rect 4973 603 4989 637
rect 5023 603 5033 637
rect 4973 561 5033 603
rect 5067 603 5083 646
rect 5117 603 5133 660
rect 5067 595 5133 603
rect 4869 527 4905 561
rect 4939 527 4997 561
rect 5031 527 5089 561
rect 5123 527 5152 561
rect 4869 477 4929 493
rect 4869 459 4895 477
rect 4773 421 4859 425
rect 4773 387 4790 421
rect 4824 391 4859 421
rect 4773 357 4813 387
rect 4847 357 4859 391
rect 4773 351 4859 357
rect 4895 373 4929 428
rect 4696 329 4730 345
rect 4626 309 4662 327
rect 4576 295 4662 309
rect 4576 293 4732 295
rect 4284 285 4388 293
rect 4284 251 4300 285
rect 4334 261 4388 285
rect 4628 285 4732 293
rect 4628 261 4682 285
rect 4334 251 4367 261
rect 4284 241 4367 251
rect 3045 117 3161 151
rect 2977 85 3011 104
rect 2828 67 3011 85
rect 2782 51 3011 67
rect 3111 116 3161 117
rect 3111 82 3119 116
rect 3153 82 3161 116
rect 3111 66 3161 82
rect 3195 116 3245 132
rect 3195 82 3203 116
rect 3237 82 3245 116
rect 3195 17 3245 82
rect 3279 117 3395 151
rect 3429 138 3463 154
rect 3279 116 3329 117
rect 3279 82 3287 116
rect 3321 82 3329 116
rect 3279 66 3329 82
rect 3497 153 3563 177
rect 3497 119 3513 153
rect 3547 119 3563 153
rect 3597 169 3835 177
rect 3597 135 3612 169
rect 3646 161 3835 169
rect 3646 143 3785 161
rect 3646 135 3658 143
rect 3429 85 3463 104
rect 3597 101 3658 135
rect 3769 127 3785 143
rect 3819 127 3835 161
rect 3597 85 3612 101
rect 3429 67 3612 85
rect 3646 67 3658 101
rect 3429 51 3658 67
rect 3692 93 3735 109
rect 3692 59 3701 93
rect 3692 17 3735 59
rect 3769 93 3835 127
rect 3769 59 3785 93
rect 3819 59 3835 93
rect 3769 51 3835 59
rect 3893 169 4131 177
rect 3893 161 4082 169
rect 3893 127 3909 161
rect 3943 143 4082 161
rect 3943 127 3959 143
rect 3893 93 3959 127
rect 4070 135 4082 143
rect 4116 135 4131 169
rect 3893 59 3909 93
rect 3943 59 3959 93
rect 3893 51 3959 59
rect 3993 93 4036 109
rect 4027 59 4036 93
rect 3993 17 4036 59
rect 4070 101 4131 135
rect 4165 153 4231 177
rect 4165 119 4181 153
rect 4215 119 4231 153
rect 4265 138 4299 154
rect 4070 67 4082 101
rect 4116 85 4131 101
rect 4333 151 4367 241
rect 4422 249 4489 259
rect 4422 215 4438 249
rect 4472 215 4489 249
rect 4422 205 4489 215
rect 4527 249 4594 259
rect 4527 215 4544 249
rect 4578 215 4594 249
rect 4527 205 4594 215
rect 4649 251 4682 261
rect 4716 251 4732 285
rect 4649 241 4732 251
rect 4649 151 4683 241
rect 4801 177 4835 351
rect 4973 485 5033 527
rect 4973 451 4989 485
rect 5023 451 5033 485
rect 4973 421 5033 451
rect 5067 485 5133 493
rect 5067 442 5083 485
rect 5073 428 5083 442
rect 5117 428 5133 485
rect 4973 405 5039 421
rect 4973 371 4989 405
rect 5023 371 5039 405
rect 4973 367 5039 371
rect 5073 417 5133 428
rect 5073 383 5083 417
rect 5117 383 5133 417
rect 4895 333 4929 339
rect 5073 349 5133 383
rect 5073 333 5083 349
rect 4895 315 5083 333
rect 5117 315 5133 349
rect 4895 299 5133 315
rect 4969 249 5133 265
rect 4969 215 4985 249
rect 5019 215 5053 249
rect 5087 215 5133 249
rect 4969 211 5133 215
rect 4885 177 4946 185
rect 4333 117 4449 151
rect 4265 85 4299 104
rect 4116 67 4299 85
rect 4070 51 4299 67
rect 4399 116 4449 117
rect 4399 82 4407 116
rect 4441 82 4449 116
rect 4399 66 4449 82
rect 4483 116 4533 132
rect 4483 82 4491 116
rect 4525 82 4533 116
rect 4483 17 4533 82
rect 4567 117 4683 151
rect 4717 138 4751 154
rect 4567 116 4617 117
rect 4567 82 4575 116
rect 4609 82 4617 116
rect 4567 66 4617 82
rect 4785 153 4851 177
rect 4785 119 4801 153
rect 4835 119 4851 153
rect 4885 169 5123 177
rect 4885 135 4900 169
rect 4934 161 5123 169
rect 4934 143 5073 161
rect 4934 135 4946 143
rect 4717 85 4751 104
rect 4885 101 4946 135
rect 5057 127 5073 143
rect 5107 127 5123 161
rect 4885 85 4900 101
rect 4717 67 4900 85
rect 4934 67 4946 101
rect 4717 51 4946 67
rect 4980 93 5023 109
rect 4980 59 4989 93
rect 4980 17 5023 59
rect 5057 93 5123 127
rect 5057 59 5073 93
rect 5107 59 5123 93
rect 5057 51 5123 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3341 17
rect 3375 -17 3433 17
rect 3467 -17 3525 17
rect 3559 -17 3617 17
rect 3651 -17 3709 17
rect 3743 -17 3801 17
rect 3835 -17 3893 17
rect 3927 -17 3985 17
rect 4019 -17 4077 17
rect 4111 -17 4169 17
rect 4203 -17 4261 17
rect 4295 -17 4353 17
rect 4387 -17 4445 17
rect 4479 -17 4537 17
rect 4571 -17 4629 17
rect 4663 -17 4721 17
rect 4755 -17 4813 17
rect 4847 -17 4905 17
rect 4939 -17 4997 17
rect 5031 -17 5089 17
rect 5123 -17 5152 17
<< viali >>
rect 29 1071 63 1105
rect 121 1071 155 1105
rect 213 1071 247 1105
rect 305 1071 339 1105
rect 397 1071 431 1105
rect 489 1071 523 1105
rect 581 1071 615 1105
rect 673 1071 707 1105
rect 765 1071 799 1105
rect 857 1071 891 1105
rect 949 1071 983 1105
rect 1041 1071 1075 1105
rect 1133 1071 1167 1105
rect 1225 1071 1259 1105
rect 1317 1071 1351 1105
rect 1409 1071 1443 1105
rect 1501 1071 1535 1105
rect 1593 1071 1627 1105
rect 1685 1071 1719 1105
rect 1777 1071 1811 1105
rect 1869 1071 1903 1105
rect 1961 1071 1995 1105
rect 2053 1071 2087 1105
rect 2145 1071 2179 1105
rect 2237 1071 2271 1105
rect 2329 1071 2363 1105
rect 2421 1071 2455 1105
rect 2513 1071 2547 1105
rect 2605 1071 2639 1105
rect 2697 1071 2731 1105
rect 2789 1071 2823 1105
rect 2881 1071 2915 1105
rect 2973 1071 3007 1105
rect 3065 1071 3099 1105
rect 3157 1071 3191 1105
rect 3249 1071 3283 1105
rect 3341 1071 3375 1105
rect 3433 1071 3467 1105
rect 3525 1071 3559 1105
rect 3617 1071 3651 1105
rect 3709 1071 3743 1105
rect 3801 1071 3835 1105
rect 3893 1071 3927 1105
rect 3985 1071 4019 1105
rect 4077 1071 4111 1105
rect 4169 1071 4203 1105
rect 4261 1071 4295 1105
rect 4353 1071 4387 1105
rect 4445 1071 4479 1105
rect 4537 1071 4571 1105
rect 4629 1071 4663 1105
rect 4721 1071 4755 1105
rect 4813 1071 4847 1105
rect 4905 1071 4939 1105
rect 4997 1071 5031 1105
rect 5089 1071 5123 1105
rect 35 637 69 660
rect 35 626 69 637
rect 305 701 339 731
rect 305 697 328 701
rect 328 697 339 701
rect 223 645 257 660
rect 223 626 257 645
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 35 451 69 462
rect 35 428 69 451
rect 223 443 257 462
rect 223 428 257 443
rect 422 645 456 660
rect 422 626 456 645
rect 949 701 983 731
rect 949 697 960 701
rect 960 697 983 701
rect 832 645 866 660
rect 832 626 866 645
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 422 443 456 462
rect 422 428 456 443
rect 305 387 328 391
rect 328 387 339 391
rect 305 357 339 387
rect 832 443 866 462
rect 832 428 866 443
rect 1031 645 1065 660
rect 1031 626 1065 645
rect 1219 637 1253 660
rect 1219 626 1253 637
rect 1323 637 1357 660
rect 1323 626 1357 637
rect 1593 701 1627 731
rect 1593 697 1616 701
rect 1616 697 1627 701
rect 1511 645 1545 660
rect 1511 626 1545 645
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1031 443 1065 462
rect 1031 428 1065 443
rect 949 387 960 391
rect 960 387 983 391
rect 949 357 983 387
rect 1219 451 1253 462
rect 1219 428 1253 451
rect 1323 451 1357 462
rect 1323 428 1357 451
rect 1511 443 1545 462
rect 1511 428 1545 443
rect 1710 645 1744 660
rect 1710 626 1744 645
rect 2237 701 2271 731
rect 2237 697 2248 701
rect 2248 697 2271 701
rect 2120 645 2154 660
rect 2120 626 2154 645
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 1710 443 1744 462
rect 1710 428 1744 443
rect 1593 387 1616 391
rect 1616 387 1627 391
rect 1593 357 1627 387
rect 2120 443 2154 462
rect 2120 428 2154 443
rect 2319 645 2353 660
rect 2319 626 2353 645
rect 2507 637 2541 660
rect 2507 626 2541 637
rect 2611 637 2645 660
rect 2611 626 2645 637
rect 2881 701 2915 731
rect 2881 697 2904 701
rect 2904 697 2915 701
rect 2799 645 2833 660
rect 2799 626 2833 645
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 2319 443 2353 462
rect 2319 428 2353 443
rect 2237 387 2248 391
rect 2248 387 2271 391
rect 2237 357 2271 387
rect 2507 451 2541 462
rect 2507 428 2541 451
rect 2611 451 2645 462
rect 2611 428 2645 451
rect 2799 443 2833 462
rect 2799 428 2833 443
rect 2998 645 3032 660
rect 2998 626 3032 645
rect 3525 701 3559 731
rect 3525 697 3536 701
rect 3536 697 3559 701
rect 3408 645 3442 660
rect 3408 626 3442 645
rect 2973 527 3007 561
rect 3065 527 3099 561
rect 3157 527 3191 561
rect 3249 527 3283 561
rect 3341 527 3375 561
rect 3433 527 3467 561
rect 2998 443 3032 462
rect 2998 428 3032 443
rect 2881 387 2904 391
rect 2904 387 2915 391
rect 2881 357 2915 387
rect 3408 443 3442 462
rect 3408 428 3442 443
rect 3607 645 3641 660
rect 3607 626 3641 645
rect 3795 637 3829 660
rect 3795 626 3829 637
rect 3899 637 3933 660
rect 3899 626 3933 637
rect 4169 701 4203 731
rect 4169 697 4192 701
rect 4192 697 4203 701
rect 4087 645 4121 660
rect 4087 626 4121 645
rect 3617 527 3651 561
rect 3709 527 3743 561
rect 3801 527 3835 561
rect 3893 527 3927 561
rect 3985 527 4019 561
rect 4077 527 4111 561
rect 3607 443 3641 462
rect 3607 428 3641 443
rect 3525 387 3536 391
rect 3536 387 3559 391
rect 3525 357 3559 387
rect 3795 451 3829 462
rect 3795 428 3829 451
rect 3899 451 3933 462
rect 3899 428 3933 451
rect 4087 443 4121 462
rect 4087 428 4121 443
rect 4286 645 4320 660
rect 4286 626 4320 645
rect 4813 701 4847 731
rect 4813 697 4824 701
rect 4824 697 4847 701
rect 4696 645 4730 660
rect 4696 626 4730 645
rect 4261 527 4295 561
rect 4353 527 4387 561
rect 4445 527 4479 561
rect 4537 527 4571 561
rect 4629 527 4663 561
rect 4721 527 4755 561
rect 4286 443 4320 462
rect 4286 428 4320 443
rect 4169 387 4192 391
rect 4192 387 4203 391
rect 4169 357 4203 387
rect 4696 443 4730 462
rect 4696 428 4730 443
rect 4895 645 4929 660
rect 4895 626 4929 645
rect 5083 637 5117 660
rect 5083 626 5117 637
rect 4905 527 4939 561
rect 4997 527 5031 561
rect 5089 527 5123 561
rect 4895 443 4929 462
rect 4895 428 4929 443
rect 4813 387 4824 391
rect 4824 387 4847 391
rect 4813 357 4847 387
rect 5083 451 5117 462
rect 5083 428 5117 451
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
rect 2881 -17 2915 17
rect 2973 -17 3007 17
rect 3065 -17 3099 17
rect 3157 -17 3191 17
rect 3249 -17 3283 17
rect 3341 -17 3375 17
rect 3433 -17 3467 17
rect 3525 -17 3559 17
rect 3617 -17 3651 17
rect 3709 -17 3743 17
rect 3801 -17 3835 17
rect 3893 -17 3927 17
rect 3985 -17 4019 17
rect 4077 -17 4111 17
rect 4169 -17 4203 17
rect 4261 -17 4295 17
rect 4353 -17 4387 17
rect 4445 -17 4479 17
rect 4537 -17 4571 17
rect 4629 -17 4663 17
rect 4721 -17 4755 17
rect 4813 -17 4847 17
rect 4905 -17 4939 17
rect 4997 -17 5031 17
rect 5089 -17 5123 17
<< metal1 >>
rect 0 1105 5152 1136
rect 0 1071 29 1105
rect 63 1071 121 1105
rect 155 1071 213 1105
rect 247 1071 305 1105
rect 339 1071 397 1105
rect 431 1071 489 1105
rect 523 1071 581 1105
rect 615 1071 673 1105
rect 707 1071 765 1105
rect 799 1071 857 1105
rect 891 1071 949 1105
rect 983 1071 1041 1105
rect 1075 1071 1133 1105
rect 1167 1071 1225 1105
rect 1259 1071 1317 1105
rect 1351 1071 1409 1105
rect 1443 1071 1501 1105
rect 1535 1071 1593 1105
rect 1627 1071 1685 1105
rect 1719 1071 1777 1105
rect 1811 1071 1869 1105
rect 1903 1071 1961 1105
rect 1995 1071 2053 1105
rect 2087 1071 2145 1105
rect 2179 1071 2237 1105
rect 2271 1071 2329 1105
rect 2363 1071 2421 1105
rect 2455 1071 2513 1105
rect 2547 1071 2605 1105
rect 2639 1071 2697 1105
rect 2731 1071 2789 1105
rect 2823 1071 2881 1105
rect 2915 1071 2973 1105
rect 3007 1071 3065 1105
rect 3099 1071 3157 1105
rect 3191 1071 3249 1105
rect 3283 1071 3341 1105
rect 3375 1071 3433 1105
rect 3467 1071 3525 1105
rect 3559 1071 3617 1105
rect 3651 1071 3709 1105
rect 3743 1071 3801 1105
rect 3835 1071 3893 1105
rect 3927 1071 3985 1105
rect 4019 1071 4077 1105
rect 4111 1071 4169 1105
rect 4203 1071 4261 1105
rect 4295 1071 4353 1105
rect 4387 1071 4445 1105
rect 4479 1071 4537 1105
rect 4571 1071 4629 1105
rect 4663 1071 4721 1105
rect 4755 1071 4813 1105
rect 4847 1071 4905 1105
rect 4939 1071 4997 1105
rect 5031 1071 5089 1105
rect 5123 1071 5152 1105
rect 0 1040 5152 1071
rect 293 731 351 737
rect 293 697 305 731
rect 339 728 351 731
rect 937 731 995 737
rect 937 728 949 731
rect 339 700 949 728
rect 339 697 351 700
rect 293 691 351 697
rect 937 697 949 700
rect 983 728 995 731
rect 1581 731 1639 737
rect 1581 728 1593 731
rect 983 700 1593 728
rect 983 697 995 700
rect 937 691 995 697
rect 1581 697 1593 700
rect 1627 728 1639 731
rect 2225 731 2283 737
rect 2225 728 2237 731
rect 1627 700 2237 728
rect 1627 697 1639 700
rect 1581 691 1639 697
rect 2225 697 2237 700
rect 2271 728 2283 731
rect 2869 731 2927 737
rect 2869 728 2881 731
rect 2271 700 2881 728
rect 2271 697 2283 700
rect 2225 691 2283 697
rect 2869 697 2881 700
rect 2915 728 2927 731
rect 3513 731 3571 737
rect 3513 728 3525 731
rect 2915 700 3525 728
rect 2915 697 2927 700
rect 2869 691 2927 697
rect 3513 697 3525 700
rect 3559 728 3571 731
rect 4157 731 4215 737
rect 4157 728 4169 731
rect 3559 700 4169 728
rect 3559 697 3571 700
rect 3513 691 3571 697
rect 4157 697 4169 700
rect 4203 728 4215 731
rect 4801 731 4859 737
rect 4801 728 4813 731
rect 4203 700 4813 728
rect 4203 697 4215 700
rect 4157 691 4215 697
rect 4801 697 4813 700
rect 4847 697 4859 731
rect 4801 691 4859 697
rect 23 660 81 666
rect 23 626 35 660
rect 69 657 81 660
rect 211 660 269 666
rect 211 657 223 660
rect 69 629 223 657
rect 69 626 81 629
rect 23 620 81 626
rect 211 626 223 629
rect 257 657 269 660
rect 410 660 468 666
rect 410 657 422 660
rect 257 629 422 657
rect 257 626 269 629
rect 211 620 269 626
rect 410 626 422 629
rect 456 626 468 660
rect 410 620 468 626
rect 820 660 878 666
rect 820 626 832 660
rect 866 657 878 660
rect 1019 660 1077 666
rect 1019 657 1031 660
rect 866 629 1031 657
rect 866 626 878 629
rect 820 620 878 626
rect 1019 626 1031 629
rect 1065 657 1077 660
rect 1207 660 1265 666
rect 1207 657 1219 660
rect 1065 629 1219 657
rect 1065 626 1077 629
rect 1019 620 1077 626
rect 1207 626 1219 629
rect 1253 626 1265 660
rect 1207 620 1265 626
rect 1311 660 1369 666
rect 1311 626 1323 660
rect 1357 657 1369 660
rect 1499 660 1557 666
rect 1499 657 1511 660
rect 1357 629 1511 657
rect 1357 626 1369 629
rect 1311 620 1369 626
rect 1499 626 1511 629
rect 1545 657 1557 660
rect 1698 660 1756 666
rect 1698 657 1710 660
rect 1545 629 1710 657
rect 1545 626 1557 629
rect 1499 620 1557 626
rect 1698 626 1710 629
rect 1744 626 1756 660
rect 1698 620 1756 626
rect 2108 660 2166 666
rect 2108 626 2120 660
rect 2154 657 2166 660
rect 2307 660 2365 666
rect 2307 657 2319 660
rect 2154 629 2319 657
rect 2154 626 2166 629
rect 2108 620 2166 626
rect 2307 626 2319 629
rect 2353 657 2365 660
rect 2495 660 2553 666
rect 2495 657 2507 660
rect 2353 629 2507 657
rect 2353 626 2365 629
rect 2307 620 2365 626
rect 2495 626 2507 629
rect 2541 626 2553 660
rect 2495 620 2553 626
rect 2599 660 2657 666
rect 2599 626 2611 660
rect 2645 657 2657 660
rect 2787 660 2845 666
rect 2787 657 2799 660
rect 2645 629 2799 657
rect 2645 626 2657 629
rect 2599 620 2657 626
rect 2787 626 2799 629
rect 2833 657 2845 660
rect 2986 660 3044 666
rect 2986 657 2998 660
rect 2833 629 2998 657
rect 2833 626 2845 629
rect 2787 620 2845 626
rect 2986 626 2998 629
rect 3032 626 3044 660
rect 2986 620 3044 626
rect 3396 660 3454 666
rect 3396 626 3408 660
rect 3442 657 3454 660
rect 3595 660 3653 666
rect 3595 657 3607 660
rect 3442 629 3607 657
rect 3442 626 3454 629
rect 3396 620 3454 626
rect 3595 626 3607 629
rect 3641 657 3653 660
rect 3783 660 3841 666
rect 3783 657 3795 660
rect 3641 629 3795 657
rect 3641 626 3653 629
rect 3595 620 3653 626
rect 3783 626 3795 629
rect 3829 626 3841 660
rect 3783 620 3841 626
rect 3887 660 3945 666
rect 3887 626 3899 660
rect 3933 657 3945 660
rect 4075 660 4133 666
rect 4075 657 4087 660
rect 3933 629 4087 657
rect 3933 626 3945 629
rect 3887 620 3945 626
rect 4075 626 4087 629
rect 4121 657 4133 660
rect 4274 660 4332 666
rect 4274 657 4286 660
rect 4121 629 4286 657
rect 4121 626 4133 629
rect 4075 620 4133 626
rect 4274 626 4286 629
rect 4320 626 4332 660
rect 4274 620 4332 626
rect 4684 660 4742 666
rect 4684 626 4696 660
rect 4730 657 4742 660
rect 4883 660 4941 666
rect 4883 657 4895 660
rect 4730 629 4895 657
rect 4730 626 4742 629
rect 4684 620 4742 626
rect 4883 626 4895 629
rect 4929 657 4941 660
rect 5071 660 5129 666
rect 5071 657 5083 660
rect 4929 629 5083 657
rect 4929 626 4941 629
rect 4883 620 4941 626
rect 5071 626 5083 629
rect 5117 626 5129 660
rect 5071 620 5129 626
rect 0 561 5152 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3157 561
rect 3191 527 3249 561
rect 3283 527 3341 561
rect 3375 527 3433 561
rect 3467 527 3617 561
rect 3651 527 3709 561
rect 3743 527 3801 561
rect 3835 527 3893 561
rect 3927 527 3985 561
rect 4019 527 4077 561
rect 4111 527 4261 561
rect 4295 527 4353 561
rect 4387 527 4445 561
rect 4479 527 4537 561
rect 4571 527 4629 561
rect 4663 527 4721 561
rect 4755 527 4905 561
rect 4939 527 4997 561
rect 5031 527 5089 561
rect 5123 527 5152 561
rect 0 496 5152 527
rect 23 462 81 468
rect 23 428 35 462
rect 69 459 81 462
rect 211 462 269 468
rect 211 459 223 462
rect 69 431 223 459
rect 69 428 81 431
rect 23 422 81 428
rect 211 428 223 431
rect 257 459 269 462
rect 410 462 468 468
rect 410 459 422 462
rect 257 431 422 459
rect 257 428 269 431
rect 211 422 269 428
rect 410 428 422 431
rect 456 428 468 462
rect 410 422 468 428
rect 820 462 878 468
rect 820 428 832 462
rect 866 459 878 462
rect 1019 462 1077 468
rect 1019 459 1031 462
rect 866 431 1031 459
rect 866 428 878 431
rect 820 422 878 428
rect 1019 428 1031 431
rect 1065 459 1077 462
rect 1207 462 1265 468
rect 1207 459 1219 462
rect 1065 431 1219 459
rect 1065 428 1077 431
rect 1019 422 1077 428
rect 1207 428 1219 431
rect 1253 428 1265 462
rect 1207 422 1265 428
rect 1311 462 1369 468
rect 1311 428 1323 462
rect 1357 459 1369 462
rect 1499 462 1557 468
rect 1499 459 1511 462
rect 1357 431 1511 459
rect 1357 428 1369 431
rect 1311 422 1369 428
rect 1499 428 1511 431
rect 1545 459 1557 462
rect 1698 462 1756 468
rect 1698 459 1710 462
rect 1545 431 1710 459
rect 1545 428 1557 431
rect 1499 422 1557 428
rect 1698 428 1710 431
rect 1744 428 1756 462
rect 1698 422 1756 428
rect 2108 462 2166 468
rect 2108 428 2120 462
rect 2154 459 2166 462
rect 2307 462 2365 468
rect 2307 459 2319 462
rect 2154 431 2319 459
rect 2154 428 2166 431
rect 2108 422 2166 428
rect 2307 428 2319 431
rect 2353 459 2365 462
rect 2495 462 2553 468
rect 2495 459 2507 462
rect 2353 431 2507 459
rect 2353 428 2365 431
rect 2307 422 2365 428
rect 2495 428 2507 431
rect 2541 428 2553 462
rect 2495 422 2553 428
rect 2599 462 2657 468
rect 2599 428 2611 462
rect 2645 459 2657 462
rect 2787 462 2845 468
rect 2787 459 2799 462
rect 2645 431 2799 459
rect 2645 428 2657 431
rect 2599 422 2657 428
rect 2787 428 2799 431
rect 2833 459 2845 462
rect 2986 462 3044 468
rect 2986 459 2998 462
rect 2833 431 2998 459
rect 2833 428 2845 431
rect 2787 422 2845 428
rect 2986 428 2998 431
rect 3032 428 3044 462
rect 2986 422 3044 428
rect 3396 462 3454 468
rect 3396 428 3408 462
rect 3442 459 3454 462
rect 3595 462 3653 468
rect 3595 459 3607 462
rect 3442 431 3607 459
rect 3442 428 3454 431
rect 3396 422 3454 428
rect 3595 428 3607 431
rect 3641 459 3653 462
rect 3783 462 3841 468
rect 3783 459 3795 462
rect 3641 431 3795 459
rect 3641 428 3653 431
rect 3595 422 3653 428
rect 3783 428 3795 431
rect 3829 428 3841 462
rect 3783 422 3841 428
rect 3887 462 3945 468
rect 3887 428 3899 462
rect 3933 459 3945 462
rect 4075 462 4133 468
rect 4075 459 4087 462
rect 3933 431 4087 459
rect 3933 428 3945 431
rect 3887 422 3945 428
rect 4075 428 4087 431
rect 4121 459 4133 462
rect 4274 462 4332 468
rect 4274 459 4286 462
rect 4121 431 4286 459
rect 4121 428 4133 431
rect 4075 422 4133 428
rect 4274 428 4286 431
rect 4320 428 4332 462
rect 4274 422 4332 428
rect 4684 462 4742 468
rect 4684 428 4696 462
rect 4730 459 4742 462
rect 4883 462 4941 468
rect 4883 459 4895 462
rect 4730 431 4895 459
rect 4730 428 4742 431
rect 4684 422 4742 428
rect 4883 428 4895 431
rect 4929 459 4941 462
rect 5071 462 5129 468
rect 5071 459 5083 462
rect 4929 431 5083 459
rect 4929 428 4941 431
rect 4883 422 4941 428
rect 5071 428 5083 431
rect 5117 428 5129 462
rect 5071 422 5129 428
rect 293 391 351 397
rect 293 357 305 391
rect 339 388 351 391
rect 937 391 995 397
rect 937 388 949 391
rect 339 360 949 388
rect 339 357 351 360
rect 293 351 351 357
rect 937 357 949 360
rect 983 388 995 391
rect 1581 391 1639 397
rect 1581 388 1593 391
rect 983 360 1593 388
rect 983 357 995 360
rect 937 351 995 357
rect 1581 357 1593 360
rect 1627 388 1639 391
rect 2225 391 2283 397
rect 2225 388 2237 391
rect 1627 360 2237 388
rect 1627 357 1639 360
rect 1581 351 1639 357
rect 2225 357 2237 360
rect 2271 388 2283 391
rect 2869 391 2927 397
rect 2869 388 2881 391
rect 2271 360 2881 388
rect 2271 357 2283 360
rect 2225 351 2283 357
rect 2869 357 2881 360
rect 2915 388 2927 391
rect 3513 391 3571 397
rect 3513 388 3525 391
rect 2915 360 3525 388
rect 2915 357 2927 360
rect 2869 351 2927 357
rect 3513 357 3525 360
rect 3559 388 3571 391
rect 4157 391 4215 397
rect 4157 388 4169 391
rect 3559 360 4169 388
rect 3559 357 3571 360
rect 3513 351 3571 357
rect 4157 357 4169 360
rect 4203 388 4215 391
rect 4801 391 4859 397
rect 4801 388 4813 391
rect 4203 360 4813 388
rect 4203 357 4215 360
rect 4157 351 4215 357
rect 4801 357 4813 360
rect 4847 357 4859 391
rect 4801 351 4859 357
rect 0 17 5152 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3341 17
rect 3375 -17 3433 17
rect 3467 -17 3525 17
rect 3559 -17 3617 17
rect 3651 -17 3709 17
rect 3743 -17 3801 17
rect 3835 -17 3893 17
rect 3927 -17 3985 17
rect 4019 -17 4077 17
rect 4111 -17 4169 17
rect 4203 -17 4261 17
rect 4295 -17 4353 17
rect 4387 -17 4445 17
rect 4479 -17 4537 17
rect 4571 -17 4629 17
rect 4663 -17 4721 17
rect 4755 -17 4813 17
rect 4847 -17 4905 17
rect 4939 -17 4997 17
rect 5031 -17 5089 17
rect 5123 -17 5152 17
rect 0 -48 5152 -17
<< labels >>
rlabel comment s 0 0 0 0 4 muxb16to1_2
flabel metal1 s 305 357 339 391 0 FreeSans 200 0 0 0 Z
port 37 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 33 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 36 nsew
flabel metal1 s 29 1071 63 1105 0 FreeSans 200 0 0 0 VGND
port 33 nsew
flabel metal1 s 305 697 339 731 0 FreeSans 200 0 0 0 Z
port 37 nsew
flabel metal1 s 1225 -17 1259 17 0 FreeSans 200 180 0 0 VGND
port 33 nsew
flabel metal1 s 1225 527 1259 561 0 FreeSans 200 180 0 0 VPWR
port 36 nsew
flabel metal1 s 3893 527 3927 561 0 FreeSans 200 0 0 0 VPWR
port 36 nsew
flabel metal1 s 3893 -17 3927 17 0 FreeSans 200 0 0 0 VGND
port 33 nsew
flabel metal1 s 1225 1071 1259 1105 0 FreeSans 200 180 0 0 VGND
port 33 nsew
flabel metal1 s 1242 544 1242 544 0 FreeSans 200 180 0 0 VPWR
port 36 nsew
flabel metal1 s 3910 544 3910 544 0 FreeSans 200 0 0 0 VPWR
port 36 nsew
flabel metal1 s 3893 1071 3927 1105 0 FreeSans 200 0 0 0 VGND
port 33 nsew
flabel metal1 s 3801 527 3835 561 0 FreeSans 200 180 0 0 VPWR
port 36 nsew
flabel metal1 s 3801 -17 3835 17 0 FreeSans 200 180 0 0 VGND
port 33 nsew
flabel metal1 s 46 1088 46 1088 0 FreeSans 200 0 0 0 VGND
port 33 nsew
flabel metal1 s 46 544 46 544 0 FreeSans 200 0 0 0 VPWR
port 36 nsew
flabel metal1 s 2605 527 2639 561 0 FreeSans 200 0 0 0 VPWR
port 36 nsew
flabel metal1 s 2605 -17 2639 17 0 FreeSans 200 0 0 0 VGND
port 33 nsew
flabel metal1 s 3818 544 3818 544 0 FreeSans 200 180 0 0 VPWR
port 36 nsew
flabel metal1 s 3801 1071 3835 1105 0 FreeSans 200 180 0 0 VGND
port 33 nsew
flabel metal1 s 46 0 46 0 0 FreeSans 200 0 0 0 VGND
port 33 nsew
flabel metal1 s 46 544 46 544 0 FreeSans 200 0 0 0 VPWR
port 36 nsew
flabel metal1 s 2622 544 2622 544 0 FreeSans 200 0 0 0 VPWR
port 36 nsew
flabel metal1 s 2605 1071 2639 1105 0 FreeSans 200 0 0 0 VGND
port 33 nsew
flabel metal1 s 1317 527 1351 561 0 FreeSans 200 0 0 0 VPWR
port 36 nsew
flabel metal1 s 1317 1071 1351 1105 0 FreeSans 200 0 0 0 VGND
port 33 nsew
flabel metal1 s 1334 544 1334 544 0 FreeSans 200 0 0 0 VPWR
port 36 nsew
flabel metal1 s 1317 -17 1351 17 0 FreeSans 200 0 0 0 VGND
port 33 nsew
flabel metal1 s 2513 527 2547 561 0 FreeSans 200 180 0 0 VPWR
port 36 nsew
flabel metal1 s 2513 1071 2547 1105 0 FreeSans 200 180 0 0 VGND
port 33 nsew
flabel metal1 s 2530 544 2530 544 0 FreeSans 200 180 0 0 VPWR
port 36 nsew
flabel metal1 s 2513 -17 2547 17 0 FreeSans 200 180 0 0 VGND
port 33 nsew
flabel metal1 s 5089 527 5123 561 0 FreeSans 200 180 0 0 VPWR
port 36 nsew
flabel metal1 s 5089 1071 5123 1105 0 FreeSans 200 180 0 0 VGND
port 33 nsew
flabel metal1 s 5106 544 5106 544 0 FreeSans 200 180 0 0 VPWR
port 36 nsew
flabel metal1 s 5089 -17 5123 17 0 FreeSans 200 180 0 0 VGND
port 33 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 34 nsew
flabel pwell s 29 1071 63 1105 0 FreeSans 200 0 0 0 VNB
port 34 nsew
flabel pwell s 1225 -17 1259 17 0 FreeSans 200 180 0 0 VNB
port 34 nsew
flabel pwell s 3893 -17 3927 17 0 FreeSans 200 0 0 0 VNB
port 34 nsew
flabel pwell s 1225 1071 1259 1105 0 FreeSans 200 180 0 0 VNB
port 34 nsew
flabel pwell s 3893 1071 3927 1105 0 FreeSans 200 0 0 0 VNB
port 34 nsew
flabel pwell s 3801 -17 3835 17 0 FreeSans 200 180 0 0 VNB
port 34 nsew
flabel pwell s 46 1088 46 1088 0 FreeSans 200 0 0 0 VNB
port 34 nsew
flabel pwell s 2605 -17 2639 17 0 FreeSans 200 0 0 0 VNB
port 34 nsew
flabel pwell s 3801 1071 3835 1105 0 FreeSans 200 180 0 0 VNB
port 34 nsew
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
port 34 nsew
flabel pwell s 2605 1071 2639 1105 0 FreeSans 200 0 0 0 VNB
port 34 nsew
flabel pwell s 1317 1071 1351 1105 0 FreeSans 200 0 0 0 VNB
port 34 nsew
flabel pwell s 1317 -17 1351 17 0 FreeSans 200 0 0 0 VNB
port 34 nsew
flabel pwell s 2513 1071 2547 1105 0 FreeSans 200 180 0 0 VNB
port 34 nsew
flabel pwell s 2513 -17 2547 17 0 FreeSans 200 180 0 0 VNB
port 34 nsew
flabel pwell s 5089 1071 5123 1105 0 FreeSans 200 180 0 0 VNB
port 34 nsew
flabel pwell s 5089 -17 5123 17 0 FreeSans 200 180 0 0 VNB
port 34 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 35 nsew
flabel nbase s 1225 527 1259 561 0 FreeSans 200 180 0 0 VPB
port 35 nsew
flabel nbase s 3893 527 3927 561 0 FreeSans 200 0 0 0 VPB
port 35 nsew
flabel nbase s 1242 544 1242 544 0 FreeSans 200 180 0 0 VPB
port 35 nsew
flabel nbase s 3910 544 3910 544 0 FreeSans 200 0 0 0 VPB
port 35 nsew
flabel nbase s 3801 527 3835 561 0 FreeSans 200 180 0 0 VPB
port 35 nsew
flabel nbase s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
port 35 nsew
flabel nbase s 2605 527 2639 561 0 FreeSans 200 0 0 0 VPB
port 35 nsew
flabel nbase s 3818 544 3818 544 0 FreeSans 200 180 0 0 VPB
port 35 nsew
flabel nbase s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
port 35 nsew
flabel nbase s 2622 544 2622 544 0 FreeSans 200 0 0 0 VPB
port 35 nsew
flabel nbase s 1317 527 1351 561 0 FreeSans 200 0 0 0 VPB
port 35 nsew
flabel nbase s 1334 544 1334 544 0 FreeSans 200 0 0 0 VPB
port 35 nsew
flabel nbase s 2513 527 2547 561 0 FreeSans 200 180 0 0 VPB
port 35 nsew
flabel nbase s 2530 544 2530 544 0 FreeSans 200 180 0 0 VPB
port 35 nsew
flabel nbase s 5089 527 5123 561 0 FreeSans 200 180 0 0 VPB
port 35 nsew
flabel nbase s 5106 544 5106 544 0 FreeSans 200 180 0 0 VPB
port 35 nsew
flabel corelocali s 1317 221 1351 255 0 FreeSans 200 0 0 0 D[2]
port 14 nsew
flabel corelocali s 1225 221 1259 255 0 FreeSans 200 0 0 0 D[1]
port 15 nsew
flabel corelocali s 4537 221 4571 255 0 FreeSans 200 0 0 0 S[7]
port 25 nsew
flabel corelocali s 4445 221 4479 255 0 FreeSans 200 0 0 0 S[6]
port 26 nsew
flabel corelocali s 3249 221 3283 255 0 FreeSans 200 0 0 0 S[5]
port 27 nsew
flabel corelocali s 1225 833 1259 867 0 FreeSans 200 0 0 0 D[9]
port 7 nsew
flabel corelocali s 29 833 63 867 0 FreeSans 200 0 0 0 D[8]
port 8 nsew
flabel corelocali s 4445 833 4479 867 0 FreeSans 200 0 0 0 S[14]
port 18 nsew
flabel corelocali s 3249 833 3283 867 0 FreeSans 200 0 0 0 S[13]
port 19 nsew
flabel corelocali s 3157 833 3191 867 0 FreeSans 200 0 0 0 S[12]
port 20 nsew
flabel corelocali s 1961 833 1995 867 0 FreeSans 200 0 0 0 S[11]
port 21 nsew
flabel corelocali s 1869 833 1903 867 0 FreeSans 200 0 0 0 S[10]
port 22 nsew
flabel corelocali s 673 833 707 867 0 FreeSans 200 0 0 0 S[9]
port 23 nsew
flabel corelocali s 581 833 615 867 0 FreeSans 200 0 0 0 S[8]
port 24 nsew
flabel corelocali s 5089 833 5123 867 0 FreeSans 200 0 0 0 D[15]
port 1 nsew
flabel corelocali s 3893 833 3927 867 0 FreeSans 200 0 0 0 D[14]
port 2 nsew
flabel corelocali s 3801 833 3835 867 0 FreeSans 200 0 0 0 D[13]
port 3 nsew
flabel corelocali s 2605 833 2639 867 0 FreeSans 200 0 0 0 D[12]
port 4 nsew
flabel corelocali s 2513 833 2547 867 0 FreeSans 200 0 0 0 D[11]
port 5 nsew
flabel corelocali s 1317 833 1351 867 0 FreeSans 200 0 0 0 D[10]
port 6 nsew
flabel corelocali s 4537 833 4571 867 0 FreeSans 200 0 0 0 S[15]
port 17 nsew
flabel corelocali s 3157 221 3191 255 0 FreeSans 200 0 0 0 S[4]
port 28 nsew
flabel corelocali s 1961 221 1995 255 0 FreeSans 200 0 0 0 S[3]
port 29 nsew
flabel corelocali s 1869 221 1903 255 0 FreeSans 200 0 0 0 S[2]
port 30 nsew
flabel corelocali s 673 221 707 255 0 FreeSans 200 0 0 0 S[1]
port 31 nsew
flabel corelocali s 581 221 615 255 0 FreeSans 200 0 0 0 S[0]
port 32 nsew
flabel corelocali s 5089 221 5123 255 0 FreeSans 200 0 0 0 D[7]
port 9 nsew
flabel corelocali s 3893 221 3927 255 0 FreeSans 200 0 0 0 D[6]
port 10 nsew
flabel corelocali s 3801 221 3835 255 0 FreeSans 200 0 0 0 D[5]
port 11 nsew
flabel corelocali s 2605 221 2639 255 0 FreeSans 200 0 0 0 D[4]
port 12 nsew
flabel corelocali s 2513 221 2547 255 0 FreeSans 200 0 0 0 D[3]
port 13 nsew
flabel corelocali s 29 221 63 255 0 FreeSans 200 0 0 0 D[0]
port 16 nsew
<< properties >>
string FIXED_BBOX 0 0 5152 1088
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3118222
string GDS_START 3026152
<< end >>
