magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1564 561
rect 18 333 77 527
rect 191 455 257 527
rect 723 439 777 527
rect 887 455 953 527
rect 1056 455 1122 527
rect 1224 455 1291 527
rect 1471 455 1537 527
rect 361 405 694 421
rect 809 405 1536 421
rect 361 371 1536 405
rect 193 303 726 337
rect 193 266 282 303
rect 80 215 282 266
rect 341 215 636 269
rect 670 199 726 303
rect 852 303 1400 337
rect 852 282 995 303
rect 760 199 995 282
rect 1074 215 1288 269
rect 1366 199 1400 303
rect 1434 268 1536 371
rect 1434 165 1470 268
rect 1313 131 1470 165
rect 105 17 171 89
rect 293 17 327 105
rect 449 17 515 89
rect 621 17 687 89
rect 1313 90 1347 131
rect 1056 54 1347 90
rect 0 -17 1564 17
<< obsli1 >>
rect 291 455 687 493
rect 111 421 155 438
rect 291 421 327 455
rect 111 387 327 421
rect 111 372 155 387
rect 31 173 359 181
rect 31 159 626 173
rect 31 139 767 159
rect 31 125 248 139
rect 355 125 767 139
rect 801 127 1234 163
rect 31 107 71 125
rect 205 119 248 125
rect 205 85 214 119
rect 721 91 767 125
rect 721 51 984 91
rect 1396 85 1502 96
rect 1396 62 1536 85
<< obsli1c >>
rect 214 85 248 119
rect 1502 85 1536 119
<< metal1 >>
rect 0 496 1564 592
rect 0 -48 1564 48
<< obsm1 >>
rect 202 119 260 125
rect 202 85 214 119
rect 248 116 260 119
rect 1490 119 1548 125
rect 1490 116 1502 119
rect 248 88 1502 116
rect 248 85 260 88
rect 202 79 260 85
rect 1490 85 1502 88
rect 1536 85 1548 119
rect 1490 79 1548 85
<< labels >>
rlabel locali s 670 199 726 303 6 A1
port 1 nsew signal input
rlabel locali s 193 303 726 337 6 A1
port 1 nsew signal input
rlabel locali s 193 266 282 303 6 A1
port 1 nsew signal input
rlabel locali s 80 215 282 266 6 A1
port 1 nsew signal input
rlabel locali s 341 215 636 269 6 A2
port 2 nsew signal input
rlabel locali s 1366 199 1400 303 6 B1
port 3 nsew signal input
rlabel locali s 852 303 1400 337 6 B1
port 3 nsew signal input
rlabel locali s 852 282 995 303 6 B1
port 3 nsew signal input
rlabel locali s 760 199 995 282 6 B1
port 3 nsew signal input
rlabel locali s 1074 215 1288 269 6 C1
port 4 nsew signal input
rlabel locali s 1434 268 1536 371 6 Y
port 5 nsew signal output
rlabel locali s 1434 165 1470 268 6 Y
port 5 nsew signal output
rlabel locali s 1313 131 1470 165 6 Y
port 5 nsew signal output
rlabel locali s 1313 90 1347 131 6 Y
port 5 nsew signal output
rlabel locali s 1056 54 1347 90 6 Y
port 5 nsew signal output
rlabel locali s 809 405 1536 421 6 Y
port 5 nsew signal output
rlabel locali s 361 405 694 421 6 Y
port 5 nsew signal output
rlabel locali s 361 371 1536 405 6 Y
port 5 nsew signal output
rlabel locali s 621 17 687 89 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 449 17 515 89 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 293 17 327 105 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 105 17 171 89 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 1564 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1564 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1471 455 1537 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1224 455 1291 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1056 455 1122 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 887 455 953 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 723 439 777 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 191 455 257 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 18 333 77 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 1564 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 1564 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1564 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1308074
string GDS_START 1298054
<< end >>
