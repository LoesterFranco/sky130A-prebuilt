magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 614 704
<< pwell >>
rect 0 0 576 49
<< scnmos >>
rect 84 116 114 226
rect 239 78 269 226
rect 317 78 347 226
rect 425 78 455 226
<< pmoshvt >>
rect 117 368 147 536
rect 234 368 264 592
rect 324 368 354 592
rect 434 368 464 592
<< ndiff >>
rect 27 188 84 226
rect 27 154 39 188
rect 73 154 84 188
rect 27 116 84 154
rect 114 162 239 226
rect 114 128 125 162
rect 159 128 194 162
rect 228 128 239 162
rect 114 116 239 128
rect 129 78 239 116
rect 269 78 317 226
rect 347 78 425 226
rect 455 214 547 226
rect 455 180 501 214
rect 535 180 547 214
rect 455 124 547 180
rect 455 90 466 124
rect 500 90 547 124
rect 455 78 547 90
<< pdiff >>
rect 165 580 234 592
rect 165 546 177 580
rect 211 546 234 580
rect 165 536 234 546
rect 58 524 117 536
rect 58 490 70 524
rect 104 490 117 524
rect 58 440 117 490
rect 58 406 70 440
rect 104 406 117 440
rect 58 368 117 406
rect 147 508 234 536
rect 147 474 177 508
rect 211 474 234 508
rect 147 424 234 474
rect 147 390 177 424
rect 211 390 234 424
rect 147 368 234 390
rect 264 580 324 592
rect 264 546 277 580
rect 311 546 324 580
rect 264 510 324 546
rect 264 476 277 510
rect 311 476 324 510
rect 264 440 324 476
rect 264 406 277 440
rect 311 406 324 440
rect 264 368 324 406
rect 354 580 434 592
rect 354 546 377 580
rect 411 546 434 580
rect 354 508 434 546
rect 354 474 377 508
rect 411 474 434 508
rect 354 368 434 474
rect 464 580 523 592
rect 464 546 477 580
rect 511 546 523 580
rect 464 497 523 546
rect 464 463 477 497
rect 511 463 523 497
rect 464 414 523 463
rect 464 380 477 414
rect 511 380 523 414
rect 464 368 523 380
<< ndiffc >>
rect 39 154 73 188
rect 125 128 159 162
rect 194 128 228 162
rect 501 180 535 214
rect 466 90 500 124
<< pdiffc >>
rect 177 546 211 580
rect 70 490 104 524
rect 70 406 104 440
rect 177 474 211 508
rect 177 390 211 424
rect 277 546 311 580
rect 277 476 311 510
rect 277 406 311 440
rect 377 546 411 580
rect 377 474 411 508
rect 477 546 511 580
rect 477 463 511 497
rect 477 380 511 414
<< poly >>
rect 234 592 264 618
rect 324 592 354 618
rect 434 592 464 618
rect 117 536 147 562
rect 117 353 147 368
rect 234 353 264 368
rect 324 353 354 368
rect 434 353 464 368
rect 114 336 150 353
rect 231 336 267 353
rect 321 336 357 353
rect 84 320 155 336
rect 84 286 105 320
rect 139 286 155 320
rect 84 270 155 286
rect 203 320 269 336
rect 203 286 219 320
rect 253 286 269 320
rect 203 270 269 286
rect 84 226 114 270
rect 239 226 269 270
rect 317 320 383 336
rect 431 330 467 353
rect 317 286 333 320
rect 367 286 383 320
rect 317 270 383 286
rect 425 314 491 330
rect 425 280 441 314
rect 475 280 491 314
rect 317 226 347 270
rect 425 264 491 280
rect 425 226 455 264
rect 84 90 114 116
rect 239 52 269 78
rect 317 52 347 78
rect 425 52 455 78
<< polycont >>
rect 105 286 139 320
rect 219 286 253 320
rect 333 286 367 320
rect 441 280 475 314
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 161 580 227 649
rect 161 546 177 580
rect 211 546 227 580
rect 21 524 120 540
rect 21 490 70 524
rect 104 490 120 524
rect 21 440 120 490
rect 21 406 70 440
rect 104 406 120 440
rect 21 390 120 406
rect 161 508 227 546
rect 161 474 177 508
rect 211 474 227 508
rect 161 424 227 474
rect 161 390 177 424
rect 211 390 227 424
rect 261 580 327 596
rect 261 546 277 580
rect 311 546 327 580
rect 261 510 327 546
rect 261 476 277 510
rect 311 476 327 510
rect 261 440 327 476
rect 361 580 427 649
rect 361 546 377 580
rect 411 546 427 580
rect 361 508 427 546
rect 361 474 377 508
rect 411 474 427 508
rect 361 458 427 474
rect 461 580 559 596
rect 461 546 477 580
rect 511 546 559 580
rect 461 497 559 546
rect 461 463 477 497
rect 511 463 559 497
rect 261 406 277 440
rect 311 424 327 440
rect 461 424 559 463
rect 311 414 559 424
rect 311 406 477 414
rect 261 390 477 406
rect 21 230 55 390
rect 461 380 477 390
rect 511 380 559 414
rect 461 364 559 380
rect 89 320 167 356
rect 89 286 105 320
rect 139 286 167 320
rect 89 270 167 286
rect 203 320 269 356
rect 203 286 219 320
rect 253 286 269 320
rect 203 270 269 286
rect 313 320 383 356
rect 313 286 333 320
rect 367 286 383 320
rect 313 270 383 286
rect 417 314 491 330
rect 417 280 441 314
rect 475 280 491 314
rect 417 264 491 280
rect 417 230 451 264
rect 525 230 559 364
rect 21 196 451 230
rect 485 214 559 230
rect 21 188 75 196
rect 21 154 39 188
rect 73 154 75 188
rect 485 180 501 214
rect 535 180 559 214
rect 21 112 75 154
rect 109 128 125 162
rect 159 128 194 162
rect 228 128 244 162
rect 485 158 559 180
rect 109 17 244 128
rect 450 124 559 158
rect 450 90 466 124
rect 500 90 559 124
rect 450 74 559 90
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
rlabel comment s 0 0 0 0 4 nand3b_1
flabel pwell s 0 0 576 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 0 617 576 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 576 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 576 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 511 390 545 424 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 511 464 545 498 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 511 538 545 572 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 B
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 576 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1731184
string GDS_START 1725580
<< end >>
