magic
tech sky130A
magscale 1 2
timestamp 1599588244
<< locali >>
rect 87 290 167 356
rect 201 290 267 356
rect 1351 364 1423 596
rect 1177 236 1247 310
rect 1389 226 1423 364
rect 1346 70 1423 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 19 390 90 566
rect 131 390 197 649
rect 460 572 526 649
rect 238 538 335 566
rect 238 504 849 538
rect 927 506 1086 649
rect 238 390 335 504
rect 19 250 53 390
rect 301 334 335 390
rect 369 402 449 470
rect 651 436 749 470
rect 369 368 681 402
rect 301 268 381 334
rect 301 250 335 268
rect 19 150 89 250
rect 213 184 335 250
rect 415 234 449 368
rect 369 184 449 234
rect 507 150 573 318
rect 615 304 681 368
rect 715 372 749 436
rect 783 406 849 504
rect 1127 472 1193 572
rect 897 406 1193 472
rect 1251 412 1317 649
rect 1093 378 1193 406
rect 715 338 1014 372
rect 980 326 1014 338
rect 1093 344 1317 378
rect 615 238 867 304
rect 980 260 1059 326
rect 980 204 1014 260
rect 1093 226 1127 344
rect 1283 330 1317 344
rect 1283 264 1355 330
rect 19 116 573 150
rect 763 170 1014 204
rect 125 17 191 82
rect 471 17 640 82
rect 763 70 829 170
rect 934 17 1002 136
rect 1048 70 1127 226
rect 1228 17 1294 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 683 1440 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 0 617 1440 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 1440 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -49 1440 -17
<< labels >>
rlabel locali s 87 290 167 356 6 D
port 1 nsew signal input
rlabel locali s 1389 226 1423 364 6 Q
port 2 nsew signal output
rlabel locali s 1351 364 1423 596 6 Q
port 2 nsew signal output
rlabel locali s 1346 70 1423 226 6 Q
port 2 nsew signal output
rlabel locali s 1177 236 1247 310 6 RESET_B
port 3 nsew signal input
rlabel locali s 201 290 267 356 6 GATE_N
port 4 nsew clock input
rlabel metal1 s 0 -49 1440 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 6 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 617 1440 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1440 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3059618
string GDS_START 3048966
<< end >>
