magic
tech sky130A
magscale 1 2
timestamp 1599588232
<< locali >>
rect 85 290 161 356
rect 195 324 517 358
rect 195 287 261 324
rect 409 236 517 324
rect 619 398 653 596
rect 799 398 833 596
rect 619 364 833 398
rect 799 330 833 364
rect 799 296 935 330
rect 889 230 935 296
rect 619 196 935 230
rect 619 70 653 196
rect 782 70 832 196
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 17 390 71 596
rect 111 420 177 649
rect 215 426 281 596
rect 321 460 371 649
rect 409 426 475 596
rect 513 460 579 649
rect 215 392 585 426
rect 17 253 51 390
rect 303 253 369 290
rect 17 219 369 253
rect 551 330 585 392
rect 693 432 759 649
rect 873 364 939 649
rect 551 264 765 330
rect 17 70 108 219
rect 551 185 585 264
rect 142 17 208 185
rect 242 117 294 185
rect 328 151 585 185
rect 242 67 480 117
rect 514 17 580 117
rect 689 17 739 162
rect 868 17 934 162
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
rlabel locali s 85 290 161 356 6 A_N
port 1 nsew signal input
rlabel locali s 409 236 517 324 6 B
port 2 nsew signal input
rlabel locali s 195 324 517 358 6 B
port 2 nsew signal input
rlabel locali s 195 287 261 324 6 B
port 2 nsew signal input
rlabel locali s 889 230 935 296 6 X
port 3 nsew signal output
rlabel locali s 799 398 833 596 6 X
port 3 nsew signal output
rlabel locali s 799 330 833 364 6 X
port 3 nsew signal output
rlabel locali s 799 296 935 330 6 X
port 3 nsew signal output
rlabel locali s 782 70 832 196 6 X
port 3 nsew signal output
rlabel locali s 619 398 653 596 6 X
port 3 nsew signal output
rlabel locali s 619 364 833 398 6 X
port 3 nsew signal output
rlabel locali s 619 196 935 230 6 X
port 3 nsew signal output
rlabel locali s 619 70 653 196 6 X
port 3 nsew signal output
rlabel metal1 s 0 -49 960 49 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 5 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 617 960 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3212828
string GDS_START 3204404
<< end >>
