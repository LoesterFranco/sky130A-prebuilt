magic
tech sky130A
magscale 1 2
timestamp 1604502729
<< locali >>
rect 85 252 161 386
rect 195 252 257 386
rect 1252 364 1318 414
rect 1114 236 1223 310
rect 1257 226 1291 364
rect 1645 364 1715 596
rect 1257 154 1323 226
rect 1681 210 1715 364
rect 1641 176 1715 210
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 17 454 89 596
rect 129 488 163 649
rect 485 564 551 649
rect 602 581 833 615
rect 197 530 393 564
rect 197 454 231 530
rect 359 496 566 530
rect 17 420 231 454
rect 265 462 325 496
rect 265 428 495 462
rect 265 420 325 428
rect 17 218 51 420
rect 291 218 325 420
rect 17 108 89 218
rect 125 17 191 218
rect 225 70 325 218
rect 359 344 427 394
rect 359 192 393 344
rect 461 310 495 428
rect 427 260 495 310
rect 532 360 566 496
rect 602 428 636 581
rect 670 481 733 547
rect 602 394 665 428
rect 532 294 597 360
rect 631 290 665 394
rect 699 376 733 481
rect 767 410 833 581
rect 905 530 1028 649
rect 1062 482 1128 596
rect 1162 516 1228 649
rect 1342 516 1408 649
rect 1062 470 1391 482
rect 875 448 1391 470
rect 875 410 1128 448
rect 699 342 1012 376
rect 631 260 706 290
rect 427 226 706 260
rect 631 224 706 226
rect 743 245 826 308
rect 359 190 425 192
rect 743 190 777 245
rect 860 211 894 342
rect 947 270 1012 342
rect 1046 364 1128 410
rect 1046 226 1080 364
rect 359 156 777 190
rect 811 177 894 211
rect 359 70 425 156
rect 811 122 845 177
rect 459 17 567 120
rect 665 72 845 122
rect 879 17 929 143
rect 975 70 1080 226
rect 1357 330 1391 448
rect 1325 264 1391 330
rect 1443 310 1509 572
rect 1555 364 1605 649
rect 1751 364 1801 649
rect 1443 244 1646 310
rect 1139 17 1205 202
rect 1357 17 1409 210
rect 1443 70 1509 244
rect 1555 17 1607 210
rect 1749 17 1801 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
<< metal1 >>
rect 0 683 1824 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 0 617 1824 649
rect 0 17 1824 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
rect 0 -49 1824 -17
<< labels >>
rlabel locali s 85 252 161 386 6 D
port 1 nsew signal input
rlabel locali s 1257 226 1291 364 6 Q
port 2 nsew signal output
rlabel locali s 1257 154 1323 226 6 Q
port 2 nsew signal output
rlabel locali s 1252 364 1318 414 6 Q
port 2 nsew signal output
rlabel locali s 1681 210 1715 364 6 Q_N
port 3 nsew signal output
rlabel locali s 1645 364 1715 596 6 Q_N
port 3 nsew signal output
rlabel locali s 1641 176 1715 210 6 Q_N
port 3 nsew signal output
rlabel locali s 1114 236 1223 310 6 RESET_B
port 4 nsew signal input
rlabel locali s 195 252 257 386 6 GATE_N
port 5 nsew clock input
rlabel metal1 s 0 -49 1824 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 1824 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1824 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3115144
string GDS_START 3101144
<< end >>
