magic
tech sky130A
magscale 1 2
timestamp 1604502741
<< locali >>
rect 182 236 257 334
rect 982 236 1048 310
rect 1362 290 1414 356
rect 1737 364 1825 596
rect 1791 294 1825 364
rect 1933 310 1999 596
rect 1933 294 1988 310
rect 1791 260 1988 294
rect 1791 217 1832 260
rect 1766 70 1832 217
rect 1938 70 1988 260
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 17 436 73 596
rect 113 436 179 649
rect 213 581 765 615
rect 17 250 51 436
rect 213 402 279 581
rect 731 551 765 581
rect 320 513 697 547
rect 320 436 386 513
rect 85 368 325 402
rect 85 294 140 368
rect 17 150 89 250
rect 291 184 325 368
rect 427 318 477 479
rect 511 375 629 479
rect 359 284 561 318
rect 359 150 393 284
rect 17 116 393 150
rect 427 124 477 250
rect 511 158 561 284
rect 595 124 629 375
rect 17 114 89 116
rect 427 90 629 124
rect 663 85 697 513
rect 731 381 865 551
rect 731 287 797 347
rect 731 153 765 287
rect 831 253 865 381
rect 799 187 865 253
rect 907 226 941 596
rect 981 364 1047 649
rect 1193 581 1500 615
rect 1081 384 1159 560
rect 1087 258 1121 384
rect 1193 350 1227 581
rect 1261 384 1328 547
rect 1367 424 1417 547
rect 1466 542 1500 581
rect 1466 458 1550 542
rect 1367 390 1482 424
rect 1155 292 1227 350
rect 907 153 948 226
rect 1087 224 1260 258
rect 731 119 948 153
rect 982 156 1192 190
rect 982 85 1016 156
rect 125 17 207 82
rect 663 51 1016 85
rect 1050 17 1100 122
rect 1142 85 1192 156
rect 1226 153 1260 224
rect 1294 187 1328 384
rect 1364 153 1414 255
rect 1226 119 1414 153
rect 1448 85 1482 390
rect 1142 51 1482 85
rect 1516 149 1550 458
rect 1589 466 1700 649
rect 1589 364 1623 466
rect 1657 317 1703 430
rect 1859 364 1893 649
rect 1584 251 1757 317
rect 2039 364 2089 649
rect 1516 83 1630 149
rect 1666 17 1732 217
rect 1868 17 1902 226
rect 2024 17 2090 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
<< metal1 >>
rect 0 683 2112 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 0 617 2112 649
rect 0 17 2112 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
rect 0 -49 2112 -17
<< obsm1 >>
rect 499 421 557 430
rect 1075 421 1133 430
rect 499 393 1133 421
rect 499 384 557 393
rect 1075 384 1133 393
rect 1267 421 1325 430
rect 1651 421 1709 430
rect 1267 393 1709 421
rect 1267 384 1325 393
rect 1651 384 1709 393
<< labels >>
rlabel locali s 182 236 257 334 6 A
port 1 nsew signal input
rlabel locali s 982 236 1048 310 6 B
port 2 nsew signal input
rlabel locali s 1362 290 1414 356 6 C
port 3 nsew signal input
rlabel locali s 1938 70 1988 260 6 X
port 4 nsew signal output
rlabel locali s 1933 310 1999 596 6 X
port 4 nsew signal output
rlabel locali s 1933 294 1988 310 6 X
port 4 nsew signal output
rlabel locali s 1791 294 1825 364 6 X
port 4 nsew signal output
rlabel locali s 1791 260 1988 294 6 X
port 4 nsew signal output
rlabel locali s 1791 217 1832 260 6 X
port 4 nsew signal output
rlabel locali s 1766 70 1832 217 6 X
port 4 nsew signal output
rlabel locali s 1737 364 1825 596 6 X
port 4 nsew signal output
rlabel metal1 s 0 -49 2112 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 617 2112 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2112 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 602122
string GDS_START 586892
<< end >>
