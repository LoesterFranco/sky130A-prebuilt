magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 17 370 87 596
rect 17 236 51 370
rect 199 298 265 360
rect 307 298 373 360
rect 409 298 481 360
rect 17 96 90 236
rect 313 51 563 128
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 121 394 213 649
rect 247 428 313 596
rect 347 462 429 649
rect 463 428 529 596
rect 247 394 529 428
rect 85 270 165 336
rect 124 264 165 270
rect 569 264 619 596
rect 124 230 619 264
rect 124 17 240 196
rect 456 162 522 230
rect 558 162 631 196
rect 597 17 631 162
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel locali s 409 298 481 360 6 A1
port 1 nsew signal input
rlabel locali s 307 298 373 360 6 A2
port 2 nsew signal input
rlabel locali s 199 298 265 360 6 A3
port 3 nsew signal input
rlabel locali s 313 51 563 128 6 B1
port 4 nsew signal input
rlabel locali s 17 370 87 596 6 X
port 5 nsew signal output
rlabel locali s 17 236 51 370 6 X
port 5 nsew signal output
rlabel locali s 17 96 90 236 6 X
port 5 nsew signal output
rlabel metal1 s 0 -49 672 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 672 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3816918
string GDS_START 3809900
<< end >>
