magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 644 561
rect 103 357 173 417
rect 311 427 361 527
rect 17 199 69 265
rect 103 161 137 357
rect 171 285 251 323
rect 471 299 539 527
rect 171 199 205 285
rect 246 215 319 251
rect 103 127 233 161
rect 19 17 85 93
rect 183 59 233 127
rect 281 153 319 215
rect 361 199 433 265
rect 467 203 550 265
rect 281 69 341 153
rect 393 83 433 199
rect 471 17 539 161
rect 0 -17 644 17
<< obsli1 >>
rect 17 451 269 493
rect 17 367 69 451
rect 219 391 269 451
rect 403 391 437 493
rect 219 357 437 391
rect 403 349 437 357
<< metal1 >>
rect 0 496 644 592
rect 0 -48 644 48
<< labels >>
rlabel locali s 281 153 319 215 6 A1
port 1 nsew signal input
rlabel locali s 281 69 341 153 6 A1
port 1 nsew signal input
rlabel locali s 246 215 319 251 6 A1
port 1 nsew signal input
rlabel locali s 393 83 433 199 6 A2
port 2 nsew signal input
rlabel locali s 361 199 433 265 6 A2
port 2 nsew signal input
rlabel locali s 467 203 550 265 6 A3
port 3 nsew signal input
rlabel locali s 171 285 251 323 6 B1
port 4 nsew signal input
rlabel locali s 171 199 205 285 6 B1
port 4 nsew signal input
rlabel locali s 17 199 69 265 6 B2
port 5 nsew signal input
rlabel locali s 183 59 233 127 6 Y
port 6 nsew signal output
rlabel locali s 103 357 173 417 6 Y
port 6 nsew signal output
rlabel locali s 103 161 137 357 6 Y
port 6 nsew signal output
rlabel locali s 103 127 233 161 6 Y
port 6 nsew signal output
rlabel locali s 471 17 539 161 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 19 17 85 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 644 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 644 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 471 299 539 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 311 427 361 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 644 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 644 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3647352
string GDS_START 3641386
<< end >>
