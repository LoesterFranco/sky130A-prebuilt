magic
tech sky130A
magscale 1 2
timestamp 1601050039
<< nwell >>
rect -38 261 1694 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 80 47 110 177
rect 164 47 194 177
rect 264 47 294 131
rect 359 47 389 131
rect 443 47 473 131
rect 527 47 557 131
rect 611 47 641 131
rect 799 47 829 131
rect 883 47 913 131
rect 967 47 997 131
rect 1056 47 1086 131
rect 1164 47 1194 131
rect 1236 47 1266 131
rect 1332 47 1362 131
rect 1431 47 1461 177
rect 1539 47 1569 177
<< pmoshvt >>
rect 80 297 110 497
rect 164 297 194 497
rect 259 371 289 497
rect 348 371 378 497
rect 443 371 473 497
rect 527 371 557 497
rect 611 371 641 497
rect 799 369 829 497
rect 883 369 913 497
rect 967 369 997 497
rect 1056 369 1086 497
rect 1141 369 1171 497
rect 1236 371 1266 497
rect 1344 371 1374 497
rect 1439 297 1469 497
rect 1523 297 1553 497
<< ndiff >>
rect 28 97 80 177
rect 28 63 36 97
rect 70 63 80 97
rect 28 47 80 63
rect 110 97 164 177
rect 110 63 120 97
rect 154 63 164 97
rect 110 47 164 63
rect 194 131 246 177
rect 1379 131 1431 177
rect 194 93 264 131
rect 194 59 220 93
rect 254 59 264 93
rect 194 47 264 59
rect 294 47 359 131
rect 389 106 443 131
rect 389 72 399 106
rect 433 72 443 106
rect 389 47 443 72
rect 473 106 527 131
rect 473 72 483 106
rect 517 72 527 106
rect 473 47 527 72
rect 557 89 611 131
rect 557 55 567 89
rect 601 55 611 89
rect 557 47 611 55
rect 641 106 693 131
rect 641 72 651 106
rect 685 72 693 106
rect 641 47 693 72
rect 747 98 799 131
rect 747 64 755 98
rect 789 64 799 98
rect 747 47 799 64
rect 829 106 883 131
rect 829 72 839 106
rect 873 72 883 106
rect 829 47 883 72
rect 913 89 967 131
rect 913 55 923 89
rect 957 55 967 89
rect 913 47 967 55
rect 997 106 1056 131
rect 997 72 1007 106
rect 1041 72 1056 106
rect 997 47 1056 72
rect 1086 101 1164 131
rect 1086 67 1108 101
rect 1142 67 1164 101
rect 1086 47 1164 67
rect 1194 47 1236 131
rect 1266 47 1332 131
rect 1362 89 1431 131
rect 1362 55 1372 89
rect 1406 55 1431 89
rect 1362 47 1431 55
rect 1461 165 1539 177
rect 1461 131 1495 165
rect 1529 131 1539 165
rect 1461 97 1539 131
rect 1461 63 1495 97
rect 1529 63 1539 97
rect 1461 47 1539 63
rect 1569 97 1621 177
rect 1569 63 1579 97
rect 1613 63 1621 97
rect 1569 47 1621 63
<< pdiff >>
rect 28 477 80 497
rect 28 443 36 477
rect 70 443 80 477
rect 28 409 80 443
rect 28 375 36 409
rect 70 375 80 409
rect 28 297 80 375
rect 110 477 164 497
rect 110 443 120 477
rect 154 443 164 477
rect 110 409 164 443
rect 110 375 120 409
rect 154 375 164 409
rect 110 297 164 375
rect 194 489 259 497
rect 194 455 212 489
rect 246 455 259 489
rect 194 371 259 455
rect 289 371 348 497
rect 378 484 443 497
rect 378 450 399 484
rect 433 450 443 484
rect 378 416 443 450
rect 378 382 399 416
rect 433 382 443 416
rect 378 371 443 382
rect 473 456 527 497
rect 473 422 483 456
rect 517 422 527 456
rect 473 371 527 422
rect 557 489 611 497
rect 557 455 567 489
rect 601 455 611 489
rect 557 371 611 455
rect 641 456 693 497
rect 641 422 651 456
rect 685 422 693 456
rect 641 371 693 422
rect 747 485 799 497
rect 747 451 755 485
rect 789 451 799 485
rect 747 417 799 451
rect 747 383 755 417
rect 789 383 799 417
rect 194 297 244 371
rect 747 369 799 383
rect 829 472 883 497
rect 829 438 839 472
rect 873 438 883 472
rect 829 369 883 438
rect 913 489 967 497
rect 913 455 923 489
rect 957 455 967 489
rect 913 369 967 455
rect 997 472 1056 497
rect 997 438 1007 472
rect 1041 438 1056 472
rect 997 369 1056 438
rect 1086 477 1141 497
rect 1086 443 1097 477
rect 1131 443 1141 477
rect 1086 369 1141 443
rect 1171 371 1236 497
rect 1266 371 1344 497
rect 1374 489 1439 497
rect 1374 455 1394 489
rect 1428 455 1439 489
rect 1374 371 1439 455
rect 1171 369 1221 371
rect 1389 297 1439 371
rect 1469 477 1523 497
rect 1469 443 1479 477
rect 1513 443 1523 477
rect 1469 409 1523 443
rect 1469 375 1479 409
rect 1513 375 1523 409
rect 1469 297 1523 375
rect 1553 477 1605 497
rect 1553 443 1563 477
rect 1597 443 1605 477
rect 1553 409 1605 443
rect 1553 375 1563 409
rect 1597 375 1605 409
rect 1553 297 1605 375
<< ndiffc >>
rect 36 63 70 97
rect 120 63 154 97
rect 220 59 254 93
rect 399 72 433 106
rect 483 72 517 106
rect 567 55 601 89
rect 651 72 685 106
rect 755 64 789 98
rect 839 72 873 106
rect 923 55 957 89
rect 1007 72 1041 106
rect 1108 67 1142 101
rect 1372 55 1406 89
rect 1495 131 1529 165
rect 1495 63 1529 97
rect 1579 63 1613 97
<< pdiffc >>
rect 36 443 70 477
rect 36 375 70 409
rect 120 443 154 477
rect 120 375 154 409
rect 212 455 246 489
rect 399 450 433 484
rect 399 382 433 416
rect 483 422 517 456
rect 567 455 601 489
rect 651 422 685 456
rect 755 451 789 485
rect 755 383 789 417
rect 839 438 873 472
rect 923 455 957 489
rect 1007 438 1041 472
rect 1097 443 1131 477
rect 1394 455 1428 489
rect 1479 443 1513 477
rect 1479 375 1513 409
rect 1563 443 1597 477
rect 1563 375 1597 409
<< poly >>
rect 80 497 110 523
rect 164 497 194 523
rect 259 497 289 523
rect 348 497 378 523
rect 443 497 473 523
rect 527 497 557 523
rect 611 497 641 523
rect 799 497 829 523
rect 883 497 913 523
rect 967 497 997 523
rect 1056 497 1086 523
rect 1141 497 1171 523
rect 1236 497 1266 523
rect 1344 497 1374 523
rect 1439 497 1469 523
rect 1523 497 1553 523
rect 80 265 110 297
rect 164 265 194 297
rect 259 265 289 371
rect 348 339 378 371
rect 335 323 389 339
rect 335 289 345 323
rect 379 289 389 323
rect 335 273 389 289
rect 80 249 194 265
rect 80 215 124 249
rect 158 215 194 249
rect 80 199 194 215
rect 239 249 293 265
rect 239 215 249 249
rect 283 229 293 249
rect 283 215 294 229
rect 239 199 294 215
rect 80 177 110 199
rect 164 177 194 199
rect 264 131 294 199
rect 359 131 389 273
rect 443 271 473 371
rect 527 272 557 371
rect 611 354 641 371
rect 799 354 829 369
rect 611 324 829 354
rect 883 337 913 369
rect 754 321 829 324
rect 754 287 764 321
rect 798 287 829 321
rect 431 255 485 271
rect 431 221 441 255
rect 475 221 485 255
rect 431 205 485 221
rect 527 256 581 272
rect 754 271 829 287
rect 871 321 925 337
rect 871 287 881 321
rect 915 287 925 321
rect 871 271 925 287
rect 527 222 537 256
rect 571 222 581 256
rect 527 206 581 222
rect 443 131 473 205
rect 527 131 557 206
rect 799 176 829 271
rect 884 176 914 271
rect 967 241 997 369
rect 1056 241 1086 369
rect 1141 337 1171 369
rect 1236 339 1266 371
rect 1140 321 1194 337
rect 1140 287 1150 321
rect 1184 287 1194 321
rect 1140 271 1194 287
rect 611 146 829 176
rect 611 131 641 146
rect 799 131 829 146
rect 883 146 914 176
rect 956 225 1010 241
rect 956 191 966 225
rect 1000 191 1010 225
rect 956 175 1010 191
rect 1056 225 1110 241
rect 1056 191 1066 225
rect 1100 191 1110 225
rect 1056 175 1110 191
rect 883 131 913 146
rect 967 131 997 175
rect 1056 131 1086 175
rect 1164 131 1194 271
rect 1236 323 1290 339
rect 1236 289 1246 323
rect 1280 289 1290 323
rect 1236 273 1290 289
rect 1236 131 1266 273
rect 1344 265 1374 371
rect 1439 265 1469 297
rect 1523 265 1553 297
rect 1332 249 1386 265
rect 1332 215 1342 249
rect 1376 215 1386 249
rect 1332 199 1386 215
rect 1431 249 1569 265
rect 1431 215 1442 249
rect 1476 215 1510 249
rect 1544 215 1569 249
rect 1431 199 1569 215
rect 1332 131 1362 199
rect 1431 177 1461 199
rect 1539 177 1569 199
rect 80 21 110 47
rect 164 21 194 47
rect 264 21 294 47
rect 359 21 389 47
rect 443 21 473 47
rect 527 21 557 47
rect 611 21 641 47
rect 799 21 829 47
rect 883 21 913 47
rect 967 21 997 47
rect 1056 21 1086 47
rect 1164 21 1194 47
rect 1236 21 1266 47
rect 1332 21 1362 47
rect 1431 21 1461 47
rect 1539 21 1569 47
<< polycont >>
rect 345 289 379 323
rect 124 215 158 249
rect 249 215 283 249
rect 764 287 798 321
rect 441 221 475 255
rect 881 287 915 321
rect 537 222 571 256
rect 1150 287 1184 321
rect 966 191 1000 225
rect 1066 191 1100 225
rect 1246 289 1280 323
rect 1342 215 1376 249
rect 1442 215 1476 249
rect 1510 215 1544 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 36 477 70 527
rect 36 409 70 443
rect 120 477 162 493
rect 154 443 162 477
rect 196 489 262 527
rect 196 455 212 489
rect 246 455 262 489
rect 380 484 449 493
rect 120 409 162 443
rect 380 450 399 484
rect 433 450 449 484
rect 380 416 449 450
rect 36 359 70 375
rect 113 375 120 390
rect 154 375 162 409
rect 113 356 162 375
rect 261 382 399 416
rect 433 382 449 416
rect 483 456 517 493
rect 551 489 617 527
rect 551 455 567 489
rect 601 455 617 489
rect 651 456 698 493
rect 483 421 517 422
rect 685 422 698 456
rect 651 421 698 422
rect 483 387 698 421
rect 739 485 805 527
rect 739 451 755 485
rect 789 451 805 485
rect 739 417 805 451
rect 739 383 755 417
rect 789 383 805 417
rect 839 472 873 493
rect 907 489 973 527
rect 907 455 923 489
rect 957 455 973 489
rect 1007 472 1041 493
rect 839 421 873 438
rect 1007 421 1041 438
rect 1097 477 1337 493
rect 1131 443 1337 477
rect 1378 489 1444 527
rect 1378 455 1394 489
rect 1428 455 1444 489
rect 1479 477 1513 493
rect 1097 425 1337 443
rect 839 387 1041 421
rect 1303 421 1337 425
rect 113 317 147 356
rect 261 333 295 382
rect 188 320 295 333
rect 17 283 147 317
rect 181 299 295 320
rect 329 323 431 338
rect 181 286 222 299
rect 329 289 345 323
rect 379 289 397 323
rect 465 314 683 348
rect 17 181 74 283
rect 181 249 215 286
rect 108 215 124 249
rect 158 215 215 249
rect 17 147 138 181
rect 36 97 70 113
rect 104 97 138 147
rect 181 165 215 215
rect 249 255 301 265
rect 465 255 499 314
rect 249 249 305 255
rect 283 221 305 249
rect 339 221 351 255
rect 425 221 441 255
rect 475 221 499 255
rect 537 256 615 272
rect 571 255 615 256
rect 571 222 581 255
rect 537 221 581 222
rect 283 215 351 221
rect 249 199 351 215
rect 537 206 615 221
rect 649 250 683 314
rect 731 323 814 349
rect 1134 337 1184 391
rect 1303 387 1436 421
rect 731 321 769 323
rect 731 287 764 321
rect 803 289 814 323
rect 798 287 814 289
rect 859 321 1184 337
rect 859 287 881 321
rect 915 303 1150 321
rect 915 287 931 303
rect 1134 287 1150 303
rect 1230 323 1367 347
rect 1230 289 1246 323
rect 1280 289 1321 323
rect 1355 289 1367 323
rect 1402 328 1436 387
rect 1479 409 1513 443
rect 1563 477 1597 527
rect 1563 409 1597 443
rect 1513 375 1529 393
rect 1479 359 1529 375
rect 1563 359 1597 375
rect 1402 294 1460 328
rect 859 250 893 287
rect 1134 271 1184 287
rect 649 193 893 250
rect 944 221 953 255
rect 987 225 1016 255
rect 944 191 966 221
rect 1000 191 1016 225
rect 1050 191 1066 225
rect 1100 191 1187 225
rect 1221 221 1229 255
rect 1263 249 1392 255
rect 1263 221 1342 249
rect 1221 215 1342 221
rect 1376 215 1392 249
rect 1221 199 1392 215
rect 1426 249 1460 294
rect 1495 317 1529 359
rect 1495 283 1639 317
rect 1426 215 1442 249
rect 1476 215 1510 249
rect 1544 215 1560 249
rect 1084 187 1187 191
rect 385 165 397 187
rect 181 153 397 165
rect 431 153 433 187
rect 181 131 433 153
rect 307 106 433 131
rect 104 63 120 97
rect 154 63 170 97
rect 36 17 70 63
rect 204 59 220 93
rect 254 59 270 93
rect 204 17 270 59
rect 307 72 399 106
rect 307 51 433 72
rect 483 123 685 157
rect 483 106 517 123
rect 651 106 685 123
rect 483 51 517 72
rect 551 55 567 89
rect 601 55 617 89
rect 551 17 617 55
rect 839 123 1041 157
rect 1084 153 1137 187
rect 1171 153 1187 187
rect 1426 165 1460 215
rect 1594 181 1639 283
rect 839 106 873 123
rect 651 51 685 72
rect 739 64 755 98
rect 789 64 805 98
rect 739 17 805 64
rect 1007 106 1041 123
rect 1276 131 1460 165
rect 1495 165 1639 181
rect 1529 147 1639 165
rect 1529 131 1545 147
rect 839 51 873 72
rect 907 55 923 89
rect 957 55 973 89
rect 907 17 973 55
rect 1007 51 1041 72
rect 1108 101 1142 119
rect 1276 101 1310 131
rect 1142 67 1310 101
rect 1495 97 1545 131
rect 1108 51 1310 67
rect 1356 55 1372 89
rect 1406 55 1422 89
rect 1356 17 1422 55
rect 1479 63 1495 97
rect 1529 63 1545 97
rect 1479 51 1545 63
rect 1579 97 1613 113
rect 1579 17 1613 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 397 289 431 323
rect 305 221 339 255
rect 581 221 615 255
rect 769 321 803 323
rect 769 289 798 321
rect 798 289 803 321
rect 1321 289 1355 323
rect 953 225 987 255
rect 953 221 966 225
rect 966 221 987 225
rect 1229 221 1263 255
rect 397 153 431 187
rect 1137 153 1171 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
<< metal1 >>
rect 0 561 1656 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 0 496 1656 527
rect 385 323 443 329
rect 385 289 397 323
rect 431 320 443 323
rect 757 323 815 329
rect 757 320 769 323
rect 431 292 769 320
rect 431 289 443 292
rect 385 283 443 289
rect 757 289 769 292
rect 803 320 815 323
rect 1309 323 1367 329
rect 1309 320 1321 323
rect 803 292 1321 320
rect 803 289 815 292
rect 757 283 815 289
rect 1309 289 1321 292
rect 1355 289 1367 323
rect 1309 283 1367 289
rect 293 255 351 261
rect 293 221 305 255
rect 339 252 351 255
rect 569 255 627 261
rect 569 252 581 255
rect 339 224 581 252
rect 339 221 351 224
rect 293 215 351 221
rect 569 221 581 224
rect 615 252 627 255
rect 941 255 999 261
rect 941 252 953 255
rect 615 224 953 252
rect 615 221 627 224
rect 569 215 627 221
rect 941 221 953 224
rect 987 252 999 255
rect 1217 255 1275 261
rect 1217 252 1229 255
rect 987 224 1229 252
rect 987 221 999 224
rect 941 215 999 221
rect 1217 221 1229 224
rect 1263 221 1275 255
rect 1217 215 1275 221
rect 385 187 443 193
rect 385 153 397 187
rect 431 184 443 187
rect 1125 187 1183 193
rect 1125 184 1137 187
rect 431 156 1137 184
rect 431 153 443 156
rect 385 147 443 153
rect 1125 153 1137 156
rect 1171 153 1183 187
rect 1125 147 1183 153
rect 0 17 1656 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
rect 0 -48 1656 -17
<< labels >>
flabel corelocali s 121 425 155 459 0 FreeSans 200 0 0 0 COUT
port 8 nsew
flabel corelocali s 121 357 155 391 0 FreeSans 200 0 0 0 COUT
port 8 nsew
flabel corelocali s 1597 221 1631 255 0 FreeSans 200 0 0 0 SUM
port 9 nsew
flabel corelocali s 305 221 339 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 397 289 431 323 0 FreeSans 200 0 0 0 B
port 2 nsew
flabel corelocali s 1137 357 1171 391 0 FreeSans 200 0 0 0 CIN
port 3 nsew
flabel corelocali s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel corelocali s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
rlabel comment s 0 0 0 0 4 fa_2
<< properties >>
string FIXED_BBOX 0 0 1656 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2032722
string GDS_START 2019124
string path 11.000 9.975 6.950 9.975 6.950 7.475 
<< end >>
