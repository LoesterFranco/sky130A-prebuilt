magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 1766 704
<< pwell >>
rect 0 0 1728 49
<< scnmos >>
rect 84 74 114 222
rect 184 74 214 222
rect 284 74 314 222
rect 424 74 454 222
rect 524 74 554 222
rect 610 74 640 222
rect 696 74 726 222
rect 782 74 812 222
rect 980 74 1010 222
rect 1066 74 1096 222
rect 1152 74 1182 222
rect 1238 74 1268 222
rect 1324 74 1354 222
rect 1410 74 1440 222
rect 1496 74 1526 222
rect 1614 74 1644 222
<< pmoshvt >>
rect 337 368 367 592
rect 437 368 467 592
rect 527 368 557 592
rect 693 368 723 592
rect 897 368 927 592
rect 1063 368 1093 592
rect 1425 368 1455 592
rect 1611 368 1641 592
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 152 184 222
rect 114 118 139 152
rect 173 118 184 152
rect 114 74 184 118
rect 214 210 284 222
rect 214 176 239 210
rect 273 176 284 210
rect 214 120 284 176
rect 214 86 239 120
rect 273 86 284 120
rect 214 74 284 86
rect 314 152 424 222
rect 314 118 339 152
rect 373 118 424 152
rect 314 74 424 118
rect 454 210 524 222
rect 454 176 465 210
rect 499 176 524 210
rect 454 120 524 176
rect 454 86 465 120
rect 499 86 524 120
rect 454 74 524 86
rect 554 207 610 222
rect 554 173 565 207
rect 599 173 610 207
rect 554 74 610 173
rect 640 120 696 222
rect 640 86 651 120
rect 685 86 696 120
rect 640 74 696 86
rect 726 207 782 222
rect 726 173 737 207
rect 771 173 782 207
rect 726 74 782 173
rect 812 132 862 222
rect 930 142 980 222
rect 812 120 869 132
rect 812 86 823 120
rect 857 86 869 120
rect 812 74 869 86
rect 923 126 980 142
rect 923 92 935 126
rect 969 92 980 126
rect 923 74 980 92
rect 1010 210 1066 222
rect 1010 176 1021 210
rect 1055 176 1066 210
rect 1010 74 1066 176
rect 1096 126 1152 222
rect 1096 92 1107 126
rect 1141 92 1152 126
rect 1096 74 1152 92
rect 1182 210 1238 222
rect 1182 176 1193 210
rect 1227 176 1238 210
rect 1182 74 1238 176
rect 1268 126 1324 222
rect 1268 92 1279 126
rect 1313 92 1324 126
rect 1268 74 1324 92
rect 1354 210 1410 222
rect 1354 176 1365 210
rect 1399 176 1410 210
rect 1354 74 1410 176
rect 1440 126 1496 222
rect 1440 92 1451 126
rect 1485 92 1496 126
rect 1440 74 1496 92
rect 1526 210 1614 222
rect 1526 176 1553 210
rect 1587 176 1614 210
rect 1526 74 1614 176
rect 1644 138 1694 222
rect 1644 126 1701 138
rect 1644 92 1655 126
rect 1689 92 1701 126
rect 1644 74 1701 92
<< pdiff >>
rect 27 580 337 592
rect 27 546 48 580
rect 82 546 128 580
rect 162 546 209 580
rect 243 546 289 580
rect 323 546 337 580
rect 27 508 337 546
rect 27 474 48 508
rect 82 474 128 508
rect 162 474 209 508
rect 243 474 289 508
rect 323 474 337 508
rect 27 440 337 474
rect 27 406 48 440
rect 82 406 128 440
rect 162 406 209 440
rect 243 406 289 440
rect 323 406 337 440
rect 27 368 337 406
rect 367 580 437 592
rect 367 546 380 580
rect 414 546 437 580
rect 367 500 437 546
rect 367 466 380 500
rect 414 466 437 500
rect 367 424 437 466
rect 367 390 380 424
rect 414 390 437 424
rect 367 368 437 390
rect 467 580 527 592
rect 467 546 480 580
rect 514 546 527 580
rect 467 508 527 546
rect 467 474 480 508
rect 514 474 527 508
rect 467 368 527 474
rect 557 580 693 592
rect 557 546 570 580
rect 604 546 646 580
rect 680 546 693 580
rect 557 500 693 546
rect 557 466 570 500
rect 604 466 646 500
rect 680 466 693 500
rect 557 424 693 466
rect 557 390 570 424
rect 604 390 646 424
rect 680 390 693 424
rect 557 368 693 390
rect 723 580 897 592
rect 723 546 736 580
rect 770 546 850 580
rect 884 546 897 580
rect 723 500 897 546
rect 723 466 736 500
rect 770 466 850 500
rect 884 466 897 500
rect 723 368 897 466
rect 927 580 1063 592
rect 927 546 940 580
rect 974 546 1016 580
rect 1050 546 1063 580
rect 927 500 1063 546
rect 927 466 940 500
rect 974 466 1016 500
rect 1050 466 1063 500
rect 927 424 1063 466
rect 927 390 940 424
rect 974 390 1016 424
rect 1050 390 1063 424
rect 927 368 1063 390
rect 1093 580 1425 592
rect 1093 546 1106 580
rect 1140 546 1174 580
rect 1208 546 1242 580
rect 1276 546 1310 580
rect 1344 546 1378 580
rect 1412 546 1425 580
rect 1093 500 1425 546
rect 1093 466 1106 500
rect 1140 466 1174 500
rect 1208 466 1242 500
rect 1276 466 1310 500
rect 1344 466 1378 500
rect 1412 466 1425 500
rect 1093 368 1425 466
rect 1455 580 1611 592
rect 1455 546 1468 580
rect 1502 546 1564 580
rect 1598 546 1611 580
rect 1455 500 1611 546
rect 1455 466 1468 500
rect 1502 466 1564 500
rect 1598 466 1611 500
rect 1455 424 1611 466
rect 1455 390 1468 424
rect 1502 390 1564 424
rect 1598 390 1611 424
rect 1455 368 1611 390
rect 1641 580 1700 592
rect 1641 546 1654 580
rect 1688 546 1700 580
rect 1641 500 1700 546
rect 1641 466 1654 500
rect 1688 466 1700 500
rect 1641 368 1700 466
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 139 118 173 152
rect 239 176 273 210
rect 239 86 273 120
rect 339 118 373 152
rect 465 176 499 210
rect 465 86 499 120
rect 565 173 599 207
rect 651 86 685 120
rect 737 173 771 207
rect 823 86 857 120
rect 935 92 969 126
rect 1021 176 1055 210
rect 1107 92 1141 126
rect 1193 176 1227 210
rect 1279 92 1313 126
rect 1365 176 1399 210
rect 1451 92 1485 126
rect 1553 176 1587 210
rect 1655 92 1689 126
<< pdiffc >>
rect 48 546 82 580
rect 128 546 162 580
rect 209 546 243 580
rect 289 546 323 580
rect 48 474 82 508
rect 128 474 162 508
rect 209 474 243 508
rect 289 474 323 508
rect 48 406 82 440
rect 128 406 162 440
rect 209 406 243 440
rect 289 406 323 440
rect 380 546 414 580
rect 380 466 414 500
rect 380 390 414 424
rect 480 546 514 580
rect 480 474 514 508
rect 570 546 604 580
rect 646 546 680 580
rect 570 466 604 500
rect 646 466 680 500
rect 570 390 604 424
rect 646 390 680 424
rect 736 546 770 580
rect 850 546 884 580
rect 736 466 770 500
rect 850 466 884 500
rect 940 546 974 580
rect 1016 546 1050 580
rect 940 466 974 500
rect 1016 466 1050 500
rect 940 390 974 424
rect 1016 390 1050 424
rect 1106 546 1140 580
rect 1174 546 1208 580
rect 1242 546 1276 580
rect 1310 546 1344 580
rect 1378 546 1412 580
rect 1106 466 1140 500
rect 1174 466 1208 500
rect 1242 466 1276 500
rect 1310 466 1344 500
rect 1378 466 1412 500
rect 1468 546 1502 580
rect 1564 546 1598 580
rect 1468 466 1502 500
rect 1564 466 1598 500
rect 1468 390 1502 424
rect 1564 390 1598 424
rect 1654 546 1688 580
rect 1654 466 1688 500
<< poly >>
rect 337 592 367 618
rect 437 592 467 618
rect 527 592 557 618
rect 693 592 723 618
rect 897 592 927 618
rect 1063 592 1093 618
rect 1425 592 1455 618
rect 1611 592 1641 618
rect 337 353 367 368
rect 437 353 467 368
rect 527 353 557 368
rect 693 353 723 368
rect 897 353 927 368
rect 1063 353 1093 368
rect 1425 353 1455 368
rect 1611 353 1641 368
rect 334 336 370 353
rect 434 336 470 353
rect 84 320 470 336
rect 84 286 132 320
rect 166 286 200 320
rect 234 286 268 320
rect 302 286 336 320
rect 370 286 404 320
rect 438 286 470 320
rect 84 270 470 286
rect 524 336 560 353
rect 690 336 726 353
rect 894 336 930 353
rect 1060 336 1096 353
rect 1422 336 1458 353
rect 1608 336 1644 353
rect 524 320 812 336
rect 524 286 540 320
rect 574 286 608 320
rect 642 286 676 320
rect 710 286 744 320
rect 778 286 812 320
rect 524 270 812 286
rect 894 320 1268 336
rect 894 286 910 320
rect 944 286 978 320
rect 1012 286 1046 320
rect 1080 286 1114 320
rect 1148 286 1182 320
rect 1216 286 1268 320
rect 894 270 1268 286
rect 84 222 114 270
rect 184 222 214 270
rect 284 222 314 270
rect 424 222 454 270
rect 524 222 554 270
rect 610 222 640 270
rect 696 222 726 270
rect 782 222 812 270
rect 980 222 1010 270
rect 1066 222 1096 270
rect 1152 222 1182 270
rect 1238 222 1268 270
rect 1324 320 1644 336
rect 1324 286 1363 320
rect 1397 286 1431 320
rect 1465 286 1499 320
rect 1533 286 1567 320
rect 1601 286 1644 320
rect 1324 270 1644 286
rect 1324 222 1354 270
rect 1410 222 1440 270
rect 1496 222 1526 270
rect 1614 222 1644 270
rect 84 48 114 74
rect 184 48 214 74
rect 284 48 314 74
rect 424 48 454 74
rect 524 48 554 74
rect 610 48 640 74
rect 696 48 726 74
rect 782 48 812 74
rect 980 48 1010 74
rect 1066 48 1096 74
rect 1152 48 1182 74
rect 1238 48 1268 74
rect 1324 48 1354 74
rect 1410 48 1440 74
rect 1496 48 1526 74
rect 1614 48 1644 74
<< polycont >>
rect 132 286 166 320
rect 200 286 234 320
rect 268 286 302 320
rect 336 286 370 320
rect 404 286 438 320
rect 540 286 574 320
rect 608 286 642 320
rect 676 286 710 320
rect 744 286 778 320
rect 910 286 944 320
rect 978 286 1012 320
rect 1046 286 1080 320
rect 1114 286 1148 320
rect 1182 286 1216 320
rect 1363 286 1397 320
rect 1431 286 1465 320
rect 1499 286 1533 320
rect 1567 286 1601 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 23 580 330 649
rect 23 546 48 580
rect 82 546 128 580
rect 162 546 209 580
rect 243 546 289 580
rect 323 546 330 580
rect 23 508 330 546
rect 23 474 48 508
rect 82 474 128 508
rect 162 474 209 508
rect 243 474 289 508
rect 323 474 330 508
rect 23 440 330 474
rect 23 406 48 440
rect 82 406 128 440
rect 162 406 209 440
rect 243 406 289 440
rect 323 406 330 440
rect 23 390 330 406
rect 364 580 430 596
rect 364 546 380 580
rect 414 546 430 580
rect 364 500 430 546
rect 364 466 380 500
rect 414 466 430 500
rect 364 424 430 466
rect 464 580 530 649
rect 464 546 480 580
rect 514 546 530 580
rect 464 508 530 546
rect 464 474 480 508
rect 514 474 530 508
rect 464 458 530 474
rect 564 580 686 596
rect 564 546 570 580
rect 604 546 646 580
rect 680 546 686 580
rect 564 500 686 546
rect 564 466 570 500
rect 604 466 646 500
rect 680 466 686 500
rect 564 424 686 466
rect 720 580 900 649
rect 720 546 736 580
rect 770 546 850 580
rect 884 546 900 580
rect 720 500 900 546
rect 720 466 736 500
rect 770 466 850 500
rect 884 466 900 500
rect 720 458 900 466
rect 934 580 1056 596
rect 934 546 940 580
rect 974 546 1016 580
rect 1050 546 1056 580
rect 934 500 1056 546
rect 934 466 940 500
rect 974 466 1016 500
rect 1050 466 1056 500
rect 934 424 1056 466
rect 1090 580 1428 649
rect 1090 546 1106 580
rect 1140 546 1174 580
rect 1208 546 1242 580
rect 1276 546 1310 580
rect 1344 546 1378 580
rect 1412 546 1428 580
rect 1090 500 1428 546
rect 1090 466 1106 500
rect 1140 466 1174 500
rect 1208 466 1242 500
rect 1276 466 1310 500
rect 1344 466 1378 500
rect 1412 466 1428 500
rect 1090 458 1428 466
rect 1464 580 1602 596
rect 1464 546 1468 580
rect 1502 546 1564 580
rect 1598 546 1602 580
rect 1464 500 1602 546
rect 1464 466 1468 500
rect 1502 466 1564 500
rect 1598 466 1602 500
rect 1464 424 1602 466
rect 1638 580 1704 649
rect 1638 546 1654 580
rect 1688 546 1704 580
rect 1638 500 1704 546
rect 1638 466 1654 500
rect 1688 466 1704 500
rect 1638 458 1704 466
rect 364 390 380 424
rect 414 390 570 424
rect 604 390 646 424
rect 680 390 940 424
rect 974 390 1016 424
rect 1050 390 1468 424
rect 1502 390 1564 424
rect 1598 390 1703 424
rect 25 320 455 356
rect 25 286 132 320
rect 166 286 200 320
rect 234 286 268 320
rect 302 286 336 320
rect 370 286 404 320
rect 438 286 455 320
rect 25 270 455 286
rect 505 320 839 356
rect 505 286 540 320
rect 574 286 608 320
rect 642 286 676 320
rect 710 286 744 320
rect 778 286 839 320
rect 505 270 839 286
rect 889 320 1232 356
rect 889 286 910 320
rect 944 286 978 320
rect 1012 286 1046 320
rect 1080 286 1114 320
rect 1148 286 1182 320
rect 1216 286 1232 320
rect 889 270 1232 286
rect 1347 320 1617 356
rect 1347 286 1363 320
rect 1397 286 1431 320
rect 1465 286 1499 320
rect 1533 286 1567 320
rect 1601 286 1617 320
rect 1347 270 1617 286
rect 23 210 515 236
rect 1657 226 1703 390
rect 23 176 39 210
rect 73 202 239 210
rect 73 176 89 202
rect 23 120 89 176
rect 223 176 239 202
rect 273 202 465 210
rect 273 176 289 202
rect 23 86 39 120
rect 73 86 89 120
rect 23 70 89 86
rect 123 152 189 168
rect 123 118 139 152
rect 173 118 189 152
rect 123 17 189 118
rect 223 120 289 176
rect 449 176 465 202
rect 499 176 515 210
rect 223 86 239 120
rect 273 86 289 120
rect 223 70 289 86
rect 323 152 389 168
rect 323 118 339 152
rect 373 118 389 152
rect 323 17 389 118
rect 449 136 515 176
rect 549 210 1243 226
rect 549 207 1021 210
rect 549 173 565 207
rect 599 173 737 207
rect 771 176 1021 207
rect 1055 176 1193 210
rect 1227 176 1243 210
rect 1349 210 1703 226
rect 1349 176 1365 210
rect 1399 176 1553 210
rect 1587 176 1703 210
rect 771 173 787 176
rect 549 170 787 173
rect 1019 160 1057 176
rect 1191 160 1229 176
rect 1363 160 1401 176
rect 1551 160 1589 176
rect 449 120 873 136
rect 449 86 465 120
rect 499 86 651 120
rect 685 86 823 120
rect 857 86 873 120
rect 449 70 873 86
rect 919 126 985 142
rect 919 92 935 126
rect 969 104 985 126
rect 1091 126 1157 142
rect 1091 104 1107 126
rect 969 92 1107 104
rect 1141 104 1157 126
rect 1263 126 1329 142
rect 1263 104 1279 126
rect 1141 92 1279 104
rect 1313 104 1329 126
rect 1435 126 1501 142
rect 1435 104 1451 126
rect 1313 92 1451 104
rect 1485 104 1501 126
rect 1639 126 1705 142
rect 1639 104 1655 126
rect 1485 92 1655 104
rect 1689 92 1705 126
rect 919 70 1705 92
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
<< metal1 >>
rect 0 683 1728 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 0 617 1728 649
rect 0 17 1728 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
rect 0 -49 1728 -17
<< labels >>
rlabel comment s 0 0 0 0 4 nand4_4
flabel pwell s 0 0 1728 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 1728 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 1728 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 1728 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 D
port 4 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 4 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 D
port 4 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 D
port 4 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 D
port 4 nsew
flabel corelocali s 1375 316 1409 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 1471 316 1505 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 1567 316 1601 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 1663 242 1697 276 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 1663 316 1697 350 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 1087 316 1121 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 1183 316 1217 350 0 FreeSans 340 0 0 0 B
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 1728 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1762834
string GDS_START 1748584
<< end >>
