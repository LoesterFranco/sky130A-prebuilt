magic
tech sky130A
magscale 1 2
timestamp 1599588232
<< locali >>
rect 167 424 233 596
rect 143 390 233 424
rect 21 236 87 310
rect 143 304 177 390
rect 121 270 177 304
rect 211 270 277 356
rect 313 336 359 578
rect 409 384 459 578
rect 425 336 459 384
rect 313 270 391 336
rect 425 270 505 336
rect 562 270 647 356
rect 121 202 155 270
rect 25 70 155 202
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 23 530 133 649
rect 23 364 109 530
rect 599 390 649 649
rect 191 202 644 236
rect 191 70 241 202
rect 275 17 341 168
rect 378 70 444 202
rect 478 17 544 168
rect 578 70 644 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel locali s 562 270 647 356 6 A1
port 1 nsew signal input
rlabel locali s 425 336 459 384 6 A2
port 2 nsew signal input
rlabel locali s 425 270 505 336 6 A2
port 2 nsew signal input
rlabel locali s 409 384 459 578 6 A2
port 2 nsew signal input
rlabel locali s 313 336 359 578 6 A3
port 3 nsew signal input
rlabel locali s 313 270 391 336 6 A3
port 3 nsew signal input
rlabel locali s 211 270 277 356 6 A4
port 4 nsew signal input
rlabel locali s 21 236 87 310 6 B1
port 5 nsew signal input
rlabel locali s 167 424 233 596 6 Y
port 6 nsew signal output
rlabel locali s 143 390 233 424 6 Y
port 6 nsew signal output
rlabel locali s 143 304 177 390 6 Y
port 6 nsew signal output
rlabel locali s 121 270 177 304 6 Y
port 6 nsew signal output
rlabel locali s 121 202 155 270 6 Y
port 6 nsew signal output
rlabel locali s 25 70 155 202 6 Y
port 6 nsew signal output
rlabel metal1 s 0 -49 672 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 8 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 9 nsew power bidirectional
rlabel metal1 s 0 617 672 715 6 VPWR
port 10 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 745928
string GDS_START 739168
<< end >>
