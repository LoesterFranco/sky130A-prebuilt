magic
tech sky130A
magscale 1 2
timestamp 1604502705
<< nwell >>
rect -38 332 806 704
<< pwell >>
rect 0 0 768 49
<< scnmos >>
rect 132 100 162 248
rect 234 120 264 248
rect 329 123 359 251
rect 423 123 453 251
rect 509 123 539 251
rect 624 123 654 251
<< pmoshvt >>
rect 92 368 122 592
rect 228 392 258 592
rect 318 392 348 592
rect 426 392 456 592
rect 516 392 546 592
rect 594 392 624 592
<< ndiff >>
rect 279 248 329 251
rect 79 220 132 248
rect 79 186 87 220
rect 121 186 132 220
rect 79 146 132 186
rect 79 112 87 146
rect 121 112 132 146
rect 79 100 132 112
rect 162 172 234 248
rect 162 138 173 172
rect 207 138 234 172
rect 162 120 234 138
rect 264 123 329 248
rect 359 123 423 251
rect 453 218 509 251
rect 453 184 464 218
rect 498 184 509 218
rect 453 123 509 184
rect 539 221 624 251
rect 539 187 566 221
rect 600 187 624 221
rect 539 123 624 187
rect 654 238 707 251
rect 654 204 665 238
rect 699 204 707 238
rect 654 123 707 204
rect 264 120 314 123
rect 162 100 215 120
<< pdiff >>
rect 37 580 92 592
rect 37 546 45 580
rect 79 546 92 580
rect 37 500 92 546
rect 37 466 45 500
rect 79 466 92 500
rect 37 420 92 466
rect 37 386 45 420
rect 79 386 92 420
rect 37 368 92 386
rect 122 580 228 592
rect 122 546 158 580
rect 192 546 228 580
rect 122 510 228 546
rect 122 476 158 510
rect 192 476 228 510
rect 122 440 228 476
rect 122 406 158 440
rect 192 406 228 440
rect 122 392 228 406
rect 258 580 318 592
rect 258 546 271 580
rect 305 546 318 580
rect 258 510 318 546
rect 258 476 271 510
rect 305 476 318 510
rect 258 440 318 476
rect 258 406 271 440
rect 305 406 318 440
rect 258 392 318 406
rect 348 580 426 592
rect 348 546 365 580
rect 399 546 426 580
rect 348 508 426 546
rect 348 474 365 508
rect 399 474 426 508
rect 348 392 426 474
rect 456 580 516 592
rect 456 546 469 580
rect 503 546 516 580
rect 456 509 516 546
rect 456 475 469 509
rect 503 475 516 509
rect 456 438 516 475
rect 456 404 469 438
rect 503 404 516 438
rect 456 392 516 404
rect 546 392 594 592
rect 624 580 679 592
rect 624 546 637 580
rect 671 546 679 580
rect 624 509 679 546
rect 624 475 637 509
rect 671 475 679 509
rect 624 438 679 475
rect 624 404 637 438
rect 671 404 679 438
rect 624 392 679 404
rect 122 368 175 392
<< ndiffc >>
rect 87 186 121 220
rect 87 112 121 146
rect 173 138 207 172
rect 464 184 498 218
rect 566 187 600 221
rect 665 204 699 238
<< pdiffc >>
rect 45 546 79 580
rect 45 466 79 500
rect 45 386 79 420
rect 158 546 192 580
rect 158 476 192 510
rect 158 406 192 440
rect 271 546 305 580
rect 271 476 305 510
rect 271 406 305 440
rect 365 546 399 580
rect 365 474 399 508
rect 469 546 503 580
rect 469 475 503 509
rect 469 404 503 438
rect 637 546 671 580
rect 637 475 671 509
rect 637 404 671 438
<< poly >>
rect 92 592 122 618
rect 228 592 258 618
rect 318 592 348 618
rect 426 592 456 618
rect 516 592 546 618
rect 594 592 624 618
rect 228 377 258 392
rect 318 377 348 392
rect 426 377 456 392
rect 516 377 546 392
rect 594 377 624 392
rect 92 353 122 368
rect 225 356 261 377
rect 315 356 351 377
rect 89 336 125 353
rect 207 340 273 356
rect 89 320 162 336
rect 89 286 112 320
rect 146 286 162 320
rect 207 306 223 340
rect 257 306 273 340
rect 207 290 273 306
rect 315 340 381 356
rect 315 306 331 340
rect 365 306 381 340
rect 315 290 381 306
rect 89 270 162 286
rect 132 248 162 270
rect 234 248 264 290
rect 329 251 359 290
rect 423 266 459 377
rect 513 296 549 377
rect 509 266 549 296
rect 591 296 627 377
rect 591 266 654 296
rect 423 251 453 266
rect 509 251 539 266
rect 624 251 654 266
rect 132 74 162 100
rect 234 94 264 120
rect 329 97 359 123
rect 423 101 453 123
rect 509 101 539 123
rect 624 101 654 123
rect 401 85 467 101
rect 401 51 417 85
rect 451 51 467 85
rect 401 35 467 51
rect 509 85 575 101
rect 509 51 525 85
rect 559 51 575 85
rect 509 35 575 51
rect 624 85 743 101
rect 624 51 693 85
rect 727 51 743 85
rect 624 35 743 51
<< polycont >>
rect 112 286 146 320
rect 223 306 257 340
rect 331 306 365 340
rect 417 51 451 85
rect 525 51 559 85
rect 693 51 727 85
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 25 580 95 596
rect 25 546 45 580
rect 79 546 95 580
rect 25 500 95 546
rect 25 466 45 500
rect 79 466 95 500
rect 25 420 95 466
rect 25 386 45 420
rect 79 386 95 420
rect 129 580 221 649
rect 129 546 158 580
rect 192 546 221 580
rect 129 510 221 546
rect 129 476 158 510
rect 192 476 221 510
rect 129 440 221 476
rect 129 406 158 440
rect 192 406 221 440
rect 129 390 221 406
rect 255 580 321 596
rect 255 546 271 580
rect 305 546 321 580
rect 255 510 321 546
rect 255 476 271 510
rect 305 476 321 510
rect 255 440 321 476
rect 361 580 419 649
rect 361 546 365 580
rect 399 546 419 580
rect 361 508 419 546
rect 361 474 365 508
rect 399 474 419 508
rect 361 458 419 474
rect 453 580 519 596
rect 453 546 469 580
rect 503 546 519 580
rect 453 509 519 546
rect 453 475 469 509
rect 503 475 519 509
rect 255 406 271 440
rect 305 424 321 440
rect 453 438 519 475
rect 453 424 469 438
rect 305 406 469 424
rect 255 404 469 406
rect 503 404 519 438
rect 255 390 519 404
rect 453 388 519 390
rect 621 580 715 596
rect 621 546 637 580
rect 671 546 715 580
rect 621 509 715 546
rect 621 475 637 509
rect 671 475 715 509
rect 621 438 715 475
rect 621 404 637 438
rect 671 404 715 438
rect 621 388 715 404
rect 25 370 95 386
rect 25 236 59 370
rect 223 340 273 356
rect 96 320 189 336
rect 96 286 112 320
rect 146 286 189 320
rect 257 306 273 340
rect 223 290 273 306
rect 313 340 381 356
rect 313 306 331 340
rect 365 306 381 340
rect 649 323 715 388
rect 313 290 381 306
rect 96 270 189 286
rect 155 256 189 270
rect 448 289 715 323
rect 448 256 514 289
rect 25 220 121 236
rect 155 222 514 256
rect 649 238 715 289
rect 25 202 87 220
rect 71 186 87 202
rect 448 218 514 222
rect 71 146 121 186
rect 71 112 87 146
rect 71 96 121 112
rect 157 172 223 188
rect 157 138 173 172
rect 207 138 223 172
rect 448 184 464 218
rect 498 184 514 218
rect 448 168 514 184
rect 550 221 615 237
rect 550 187 566 221
rect 600 187 615 221
rect 649 204 665 238
rect 699 204 715 238
rect 649 203 715 204
rect 550 171 615 187
rect 579 169 615 171
rect 157 17 223 138
rect 579 135 643 169
rect 313 88 467 134
rect 401 85 467 88
rect 401 51 417 85
rect 451 51 467 85
rect 505 101 545 134
rect 505 85 575 101
rect 505 51 525 85
rect 559 51 575 85
rect 609 17 643 135
rect 677 85 743 134
rect 677 51 693 85
rect 727 51 743 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a311o_1
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 10 nsew
flabel corelocali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 10 nsew
flabel corelocali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 10 nsew
flabel corelocali s 703 94 737 128 0 FreeSans 340 0 0 0 C1
port 5 nsew
flabel corelocali s 511 94 545 128 0 FreeSans 340 0 0 0 B1
port 4 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 319 94 353 128 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 415 94 449 128 0 FreeSans 340 0 0 0 A1
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 768 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3609368
string GDS_START 3601836
<< end >>
