magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 644 561
rect 108 455 174 527
rect 295 439 329 527
rect 29 299 386 335
rect 29 207 129 299
rect 163 199 285 265
rect 321 249 386 299
rect 321 215 387 249
rect 20 17 79 173
rect 463 157 523 423
rect 560 199 615 325
rect 191 123 523 157
rect 191 51 260 123
rect 352 17 418 89
rect 459 51 523 123
rect 559 17 625 165
rect 0 -17 644 17
<< obsli1 >>
rect 22 421 74 493
rect 210 421 244 493
rect 363 457 618 493
rect 22 405 244 421
rect 363 405 429 457
rect 22 371 429 405
rect 557 359 618 457
<< metal1 >>
rect 0 496 644 592
rect 0 -48 644 48
<< labels >>
rlabel locali s 163 199 285 265 6 A1
port 1 nsew signal input
rlabel locali s 321 249 386 299 6 A2
port 2 nsew signal input
rlabel locali s 321 215 387 249 6 A2
port 2 nsew signal input
rlabel locali s 29 299 386 335 6 A2
port 2 nsew signal input
rlabel locali s 29 207 129 299 6 A2
port 2 nsew signal input
rlabel locali s 560 199 615 325 6 B1
port 3 nsew signal input
rlabel locali s 463 157 523 423 6 Y
port 4 nsew signal output
rlabel locali s 459 51 523 123 6 Y
port 4 nsew signal output
rlabel locali s 191 123 523 157 6 Y
port 4 nsew signal output
rlabel locali s 191 51 260 123 6 Y
port 4 nsew signal output
rlabel locali s 559 17 625 165 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 352 17 418 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 20 17 79 173 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 644 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 644 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 295 439 329 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 108 455 174 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 644 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 644 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 4064022
string GDS_START 4058158
<< end >>
