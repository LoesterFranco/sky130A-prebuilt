magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1564 561
rect 17 297 85 527
rect 119 345 153 493
rect 187 379 253 527
rect 287 345 321 493
rect 355 379 489 527
rect 591 379 657 527
rect 771 379 809 527
rect 119 297 321 345
rect 1391 379 1457 527
rect 119 263 153 297
rect 17 211 153 263
rect 423 211 616 263
rect 650 211 895 263
rect 931 211 1170 263
rect 1204 211 1354 263
rect 1390 211 1547 263
rect 119 177 153 211
rect 17 17 85 177
rect 119 143 321 177
rect 119 51 153 143
rect 187 17 253 109
rect 287 51 321 143
rect 355 17 405 109
rect 985 17 1121 101
rect 1223 17 1289 101
rect 1391 17 1457 101
rect 0 -17 1564 17
<< obsli1 >>
rect 523 345 557 493
rect 691 345 725 493
rect 867 459 1289 493
rect 867 379 933 459
rect 967 345 1001 425
rect 355 297 1001 345
rect 1051 297 1105 459
rect 1139 345 1189 425
rect 1223 379 1289 459
rect 1323 345 1357 425
rect 1491 345 1547 493
rect 1139 297 1547 345
rect 355 263 389 297
rect 187 211 389 263
rect 355 177 389 211
rect 355 143 609 177
rect 439 135 609 143
rect 643 101 677 177
rect 711 135 1547 177
rect 439 51 861 101
rect 897 51 951 135
rect 1155 51 1189 135
rect 1323 51 1357 135
rect 1491 51 1547 135
<< metal1 >>
rect 0 496 1564 592
rect 0 -48 1564 48
<< labels >>
rlabel locali s 1390 211 1547 263 6 A1
port 1 nsew signal input
rlabel locali s 1204 211 1354 263 6 A2
port 2 nsew signal input
rlabel locali s 931 211 1170 263 6 A3
port 3 nsew signal input
rlabel locali s 650 211 895 263 6 B1
port 4 nsew signal input
rlabel locali s 423 211 616 263 6 C1
port 5 nsew signal input
rlabel locali s 287 345 321 493 6 X
port 6 nsew signal output
rlabel locali s 287 51 321 143 6 X
port 6 nsew signal output
rlabel locali s 119 345 153 493 6 X
port 6 nsew signal output
rlabel locali s 119 297 321 345 6 X
port 6 nsew signal output
rlabel locali s 119 263 153 297 6 X
port 6 nsew signal output
rlabel locali s 119 177 153 211 6 X
port 6 nsew signal output
rlabel locali s 119 143 321 177 6 X
port 6 nsew signal output
rlabel locali s 119 51 153 143 6 X
port 6 nsew signal output
rlabel locali s 17 211 153 263 6 X
port 6 nsew signal output
rlabel locali s 1391 17 1457 101 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1223 17 1289 101 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 985 17 1121 101 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 355 17 405 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 187 17 253 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 17 17 85 177 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 1564 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1564 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1391 379 1457 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 771 379 809 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 591 379 657 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 355 379 489 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 187 379 253 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 17 297 85 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 1564 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 1564 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1564 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 768168
string GDS_START 755876
<< end >>
