magic
tech sky130A
magscale 1 2
timestamp 1601050082
<< locali >>
rect 25 260 101 356
rect 345 410 411 476
rect 377 296 411 410
rect 377 230 455 296
rect 1549 406 1621 596
rect 1587 226 1621 406
rect 1553 70 1621 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 23 424 89 596
rect 129 458 163 649
rect 203 559 269 596
rect 315 593 387 649
rect 742 593 820 649
rect 421 559 708 585
rect 964 581 1175 615
rect 964 559 998 581
rect 203 551 998 559
rect 203 525 455 551
rect 674 525 998 551
rect 23 390 169 424
rect 135 310 169 390
rect 203 344 295 525
rect 135 226 227 310
rect 23 192 227 226
rect 23 70 73 192
rect 109 17 159 158
rect 193 85 227 192
rect 261 270 343 344
rect 445 364 511 491
rect 551 485 591 517
rect 551 451 827 485
rect 551 425 591 451
rect 445 330 523 364
rect 261 119 295 270
rect 489 264 523 330
rect 557 332 591 425
rect 628 366 708 417
rect 557 298 640 332
rect 489 230 572 264
rect 329 162 504 196
rect 329 85 363 162
rect 193 51 363 85
rect 397 17 436 128
rect 470 85 504 162
rect 538 119 572 230
rect 606 189 640 298
rect 674 291 708 366
rect 793 391 827 451
rect 861 425 930 491
rect 793 325 862 391
rect 674 257 751 291
rect 896 283 930 425
rect 606 123 683 189
rect 717 172 751 257
rect 785 240 930 283
rect 964 308 998 525
rect 1032 376 1066 547
rect 1109 410 1175 581
rect 1247 504 1313 649
rect 1032 342 1151 376
rect 964 274 1083 308
rect 785 206 983 240
rect 1017 230 1083 274
rect 1117 280 1151 342
rect 1217 372 1283 448
rect 1358 372 1408 572
rect 1448 406 1514 649
rect 1217 338 1553 372
rect 1217 314 1283 338
rect 1382 280 1448 304
rect 1117 246 1448 280
rect 949 189 983 206
rect 1117 189 1151 246
rect 1382 238 1448 246
rect 1485 270 1553 338
rect 717 138 915 172
rect 717 85 751 138
rect 470 51 751 85
rect 797 17 847 104
rect 881 85 915 138
rect 949 119 1015 189
rect 1049 139 1151 189
rect 1112 85 1178 102
rect 881 51 1178 85
rect 1245 17 1311 212
rect 1485 204 1519 270
rect 1655 364 1705 649
rect 1357 170 1519 204
rect 1357 70 1423 170
rect 1460 17 1519 136
rect 1655 17 1705 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
<< metal1 >>
rect 0 683 1728 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 0 617 1728 649
rect 0 17 1728 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
rect 0 -49 1728 -17
<< labels >>
rlabel locali s 377 296 411 410 6 D
port 1 nsew signal input
rlabel locali s 377 230 455 296 6 D
port 1 nsew signal input
rlabel locali s 345 410 411 476 6 D
port 1 nsew signal input
rlabel locali s 1587 226 1621 406 6 Q
port 2 nsew signal output
rlabel locali s 1553 70 1621 226 6 Q
port 2 nsew signal output
rlabel locali s 1549 406 1621 596 6 Q
port 2 nsew signal output
rlabel locali s 25 260 101 356 6 CLK
port 3 nsew clock input
rlabel metal1 s 0 -49 1728 49 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1728 715 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1728 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2652250
string GDS_START 2638882
<< end >>
