magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 806 704
<< pwell >>
rect 0 0 768 49
<< scnmos >>
rect 113 74 143 222
rect 191 74 221 222
rect 305 74 335 222
rect 419 74 449 222
rect 533 74 563 222
rect 619 74 649 222
<< pmoshvt >>
rect 104 392 134 592
rect 194 392 224 592
rect 326 392 356 592
rect 416 392 446 592
rect 540 368 570 592
rect 630 368 660 592
<< ndiff >>
rect 56 210 113 222
rect 56 176 68 210
rect 102 176 113 210
rect 56 120 113 176
rect 56 86 68 120
rect 102 86 113 120
rect 56 74 113 86
rect 143 74 191 222
rect 221 74 305 222
rect 335 74 419 222
rect 449 202 533 222
rect 449 168 469 202
rect 503 168 533 202
rect 449 116 533 168
rect 449 82 469 116
rect 503 82 533 116
rect 449 74 533 82
rect 563 199 619 222
rect 563 165 574 199
rect 608 165 619 199
rect 563 74 619 165
rect 649 200 723 222
rect 649 166 681 200
rect 715 166 723 200
rect 649 120 723 166
rect 649 86 660 120
rect 694 86 723 120
rect 649 74 723 86
<< pdiff >>
rect 27 580 104 592
rect 27 546 39 580
rect 73 546 104 580
rect 27 510 104 546
rect 27 476 39 510
rect 73 476 104 510
rect 27 440 104 476
rect 27 406 39 440
rect 73 406 104 440
rect 27 392 104 406
rect 134 580 194 592
rect 134 546 147 580
rect 181 546 194 580
rect 134 509 194 546
rect 134 475 147 509
rect 181 475 194 509
rect 134 438 194 475
rect 134 404 147 438
rect 181 404 194 438
rect 134 392 194 404
rect 224 580 326 592
rect 224 546 259 580
rect 293 546 326 580
rect 224 456 326 546
rect 224 422 259 456
rect 293 422 326 456
rect 224 392 326 422
rect 356 580 416 592
rect 356 546 369 580
rect 403 546 416 580
rect 356 509 416 546
rect 356 475 369 509
rect 403 475 416 509
rect 356 438 416 475
rect 356 404 369 438
rect 403 404 416 438
rect 356 392 416 404
rect 446 576 540 592
rect 446 542 476 576
rect 510 542 540 576
rect 446 392 540 542
rect 487 368 540 392
rect 570 414 630 592
rect 570 380 583 414
rect 617 380 630 414
rect 570 368 630 380
rect 660 576 741 592
rect 660 542 692 576
rect 726 542 741 576
rect 660 368 741 542
<< ndiffc >>
rect 68 176 102 210
rect 68 86 102 120
rect 469 168 503 202
rect 469 82 503 116
rect 574 165 608 199
rect 681 166 715 200
rect 660 86 694 120
<< pdiffc >>
rect 39 546 73 580
rect 39 476 73 510
rect 39 406 73 440
rect 147 546 181 580
rect 147 475 181 509
rect 147 404 181 438
rect 259 546 293 580
rect 259 422 293 456
rect 369 546 403 580
rect 369 475 403 509
rect 369 404 403 438
rect 476 542 510 576
rect 583 380 617 414
rect 692 542 726 576
<< poly >>
rect 104 592 134 618
rect 194 592 224 618
rect 326 592 356 618
rect 416 592 446 618
rect 540 592 570 618
rect 630 592 660 618
rect 104 377 134 392
rect 194 377 224 392
rect 326 377 356 392
rect 416 377 446 392
rect 101 326 137 377
rect 23 310 137 326
rect 23 276 39 310
rect 73 290 137 310
rect 191 310 227 377
rect 323 310 359 377
rect 416 358 449 377
rect 419 310 449 358
rect 540 353 570 368
rect 630 353 660 368
rect 537 320 573 353
rect 627 326 663 353
rect 627 320 747 326
rect 533 310 747 320
rect 191 294 257 310
rect 73 276 143 290
rect 23 260 143 276
rect 113 222 143 260
rect 191 260 207 294
rect 241 260 257 294
rect 191 244 257 260
rect 305 294 371 310
rect 305 260 321 294
rect 355 260 371 294
rect 305 244 371 260
rect 419 294 485 310
rect 419 260 435 294
rect 469 260 485 294
rect 419 244 485 260
rect 533 276 697 310
rect 731 276 747 310
rect 533 260 747 276
rect 191 222 221 244
rect 305 222 335 244
rect 419 222 449 244
rect 533 222 563 260
rect 619 222 649 260
rect 113 48 143 74
rect 191 48 221 74
rect 305 48 335 74
rect 419 48 449 74
rect 533 48 563 74
rect 619 48 649 74
<< polycont >>
rect 39 276 73 310
rect 207 260 241 294
rect 321 260 355 294
rect 435 260 469 294
rect 697 276 731 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 23 580 89 649
rect 23 546 39 580
rect 73 546 89 580
rect 23 510 89 546
rect 23 476 39 510
rect 73 476 89 510
rect 23 440 89 476
rect 23 406 39 440
rect 73 406 89 440
rect 23 390 89 406
rect 123 580 197 596
rect 123 546 147 580
rect 181 546 197 580
rect 123 509 197 546
rect 123 475 147 509
rect 181 475 197 509
rect 123 438 197 475
rect 123 404 147 438
rect 181 404 197 438
rect 243 580 309 649
rect 243 546 259 580
rect 293 546 309 580
rect 243 456 309 546
rect 243 422 259 456
rect 293 422 309 456
rect 243 412 309 422
rect 353 580 419 596
rect 353 546 369 580
rect 403 546 419 580
rect 353 509 419 546
rect 460 576 526 649
rect 460 542 476 576
rect 510 542 526 576
rect 460 532 526 542
rect 674 576 745 649
rect 674 542 692 576
rect 726 542 745 576
rect 674 532 745 542
rect 353 475 369 509
rect 403 498 419 509
rect 403 475 747 498
rect 353 464 747 475
rect 353 438 419 464
rect 123 378 197 404
rect 353 404 369 438
rect 403 404 419 438
rect 353 378 419 404
rect 23 310 89 356
rect 23 276 39 310
rect 73 276 89 310
rect 23 260 89 276
rect 123 344 419 378
rect 567 414 647 430
rect 567 380 583 414
rect 617 380 647 414
rect 123 226 157 344
rect 52 210 157 226
rect 52 176 68 210
rect 102 192 157 210
rect 191 294 263 310
rect 191 260 207 294
rect 241 260 263 294
rect 102 176 118 192
rect 52 120 118 176
rect 52 86 68 120
rect 102 86 118 120
rect 191 88 263 260
rect 305 294 371 310
rect 305 260 321 294
rect 355 260 371 294
rect 305 88 371 260
rect 409 294 485 310
rect 409 260 435 294
rect 469 260 485 294
rect 409 236 485 260
rect 567 226 647 380
rect 681 310 747 464
rect 681 276 697 310
rect 731 276 747 310
rect 681 260 747 276
rect 453 168 469 202
rect 503 168 519 202
rect 453 116 519 168
rect 558 199 647 226
rect 558 165 574 199
rect 608 165 647 199
rect 558 154 647 165
rect 681 200 731 216
rect 715 166 731 200
rect 681 120 731 166
rect 52 70 118 86
rect 453 82 469 116
rect 503 82 519 116
rect 453 17 519 82
rect 644 86 660 120
rect 694 86 731 120
rect 644 17 731 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel comment s 0 0 0 0 4 and4_2
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 415 242 449 276 0 FreeSans 340 0 0 0 D
port 4 nsew
flabel corelocali s 319 94 353 128 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 319 168 353 202 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 319 242 353 276 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 223 94 257 128 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 223 168 257 202 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 223 242 257 276 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 607 168 641 202 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 607 242 641 276 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 607 390 641 424 0 FreeSans 340 0 0 0 X
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 768 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3220954
string GDS_START 3213750
<< end >>
