magic
tech sky130A
magscale 1 2
timestamp 1604502729
<< locali >>
rect 25 260 91 356
rect 211 364 288 440
rect 211 226 245 364
rect 393 270 459 356
rect 501 270 567 356
rect 601 270 681 356
rect 211 70 277 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 130 542 196 649
rect 329 542 395 649
rect 548 542 614 649
rect 770 542 841 649
rect 23 508 89 540
rect 23 474 797 508
rect 23 390 159 474
rect 125 226 159 390
rect 23 192 159 226
rect 322 390 729 440
rect 322 326 356 390
rect 279 260 356 326
rect 763 336 797 474
rect 723 270 797 336
rect 322 226 356 260
rect 23 108 89 192
rect 125 17 175 158
rect 322 192 814 226
rect 311 17 433 158
rect 748 70 814 192
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel locali s 25 260 91 356 6 A_N
port 1 nsew signal input
rlabel locali s 601 270 681 356 6 B
port 2 nsew signal input
rlabel locali s 501 270 567 356 6 C
port 3 nsew signal input
rlabel locali s 393 270 459 356 6 D
port 4 nsew signal input
rlabel locali s 211 364 288 440 6 X
port 5 nsew signal output
rlabel locali s 211 226 245 364 6 X
port 5 nsew signal output
rlabel locali s 211 70 277 226 6 X
port 5 nsew signal output
rlabel metal1 s 0 -49 864 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 864 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3352610
string GDS_START 3346012
<< end >>
