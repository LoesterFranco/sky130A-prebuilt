magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 1195 323 1245 425
rect 1383 323 1433 425
rect 1571 323 1621 425
rect 1759 323 1809 425
rect 1195 289 1913 323
rect 17 213 101 257
rect 1158 215 1776 255
rect 17 51 63 213
rect 1810 181 1913 289
rect 425 145 1913 181
rect 425 51 501 145
rect 613 51 689 145
rect 801 51 877 145
rect 989 51 1065 145
rect 1177 51 1253 145
rect 1365 51 1441 145
rect 1553 51 1629 145
rect 1741 51 1817 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 25 291 69 527
rect 103 291 189 493
rect 233 291 292 527
rect 335 333 399 493
rect 443 367 493 527
rect 537 333 587 493
rect 631 367 681 527
rect 725 333 775 493
rect 819 367 869 527
rect 913 333 963 493
rect 1007 367 1057 527
rect 1101 459 1903 493
rect 1101 333 1151 459
rect 335 291 1151 333
rect 1289 357 1339 459
rect 1477 357 1527 459
rect 1665 357 1715 459
rect 1853 357 1903 459
rect 145 257 189 291
rect 145 215 1104 257
rect 145 213 247 215
rect 97 17 141 179
rect 175 51 247 213
rect 289 17 391 181
rect 545 17 579 111
rect 733 17 767 111
rect 921 17 955 111
rect 1109 17 1143 111
rect 1297 17 1331 111
rect 1485 17 1519 111
rect 1673 17 1707 111
rect 1861 17 1915 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< labels >>
rlabel locali s 17 213 101 257 6 A
port 1 nsew signal input
rlabel locali s 17 51 63 213 6 A
port 1 nsew signal input
rlabel locali s 1158 215 1776 255 6 SLEEP
port 2 nsew signal input
rlabel locali s 1810 181 1913 289 6 X
port 3 nsew signal output
rlabel locali s 1759 323 1809 425 6 X
port 3 nsew signal output
rlabel locali s 1741 51 1817 145 6 X
port 3 nsew signal output
rlabel locali s 1571 323 1621 425 6 X
port 3 nsew signal output
rlabel locali s 1553 51 1629 145 6 X
port 3 nsew signal output
rlabel locali s 1383 323 1433 425 6 X
port 3 nsew signal output
rlabel locali s 1365 51 1441 145 6 X
port 3 nsew signal output
rlabel locali s 1195 323 1245 425 6 X
port 3 nsew signal output
rlabel locali s 1195 289 1913 323 6 X
port 3 nsew signal output
rlabel locali s 1177 51 1253 145 6 X
port 3 nsew signal output
rlabel locali s 989 51 1065 145 6 X
port 3 nsew signal output
rlabel locali s 801 51 877 145 6 X
port 3 nsew signal output
rlabel locali s 613 51 689 145 6 X
port 3 nsew signal output
rlabel locali s 425 145 1913 181 6 X
port 3 nsew signal output
rlabel locali s 425 51 501 145 6 X
port 3 nsew signal output
rlabel metal1 s 0 -48 1932 48 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 496 1932 592 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1932 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2644196
string GDS_START 2630010
<< end >>
