magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 736 561
rect 17 315 80 527
rect 206 426 329 527
rect 29 149 82 265
rect 291 391 329 426
rect 363 425 458 493
rect 291 353 357 391
rect 492 358 535 527
rect 575 359 632 493
rect 17 17 71 115
rect 402 153 484 249
rect 598 289 632 359
rect 666 325 719 527
rect 598 185 719 289
rect 402 61 444 153
rect 598 143 632 185
rect 482 17 548 116
rect 583 51 632 143
rect 666 17 719 149
rect 0 -17 736 17
<< obsli1 >>
rect 116 249 171 381
rect 210 319 257 392
rect 402 319 440 378
rect 210 285 564 319
rect 116 203 283 249
rect 116 61 171 203
rect 317 114 368 285
rect 211 61 368 114
rect 518 199 564 285
<< metal1 >>
rect 0 496 736 592
rect 0 -48 736 48
<< labels >>
rlabel locali s 29 149 82 265 6 A_N
port 1 nsew signal input
rlabel locali s 363 425 458 493 6 B
port 2 nsew signal input
rlabel locali s 402 153 484 249 6 C
port 3 nsew signal input
rlabel locali s 402 61 444 153 6 C
port 3 nsew signal input
rlabel locali s 598 289 632 359 6 X
port 4 nsew signal output
rlabel locali s 598 185 719 289 6 X
port 4 nsew signal output
rlabel locali s 598 143 632 185 6 X
port 4 nsew signal output
rlabel locali s 583 51 632 143 6 X
port 4 nsew signal output
rlabel locali s 575 359 632 493 6 X
port 4 nsew signal output
rlabel locali s 666 17 719 149 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 482 17 548 116 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 17 17 71 115 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 736 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 736 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 666 325 719 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 492 358 535 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 291 391 329 426 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 291 353 357 391 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 206 426 329 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 17 315 80 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 736 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 736 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3794272
string GDS_START 3787724
<< end >>
