magic
tech sky130A
magscale 1 2
timestamp 1604502741
<< locali >>
rect 20 238 146 372
rect 665 363 748 612
rect 690 224 748 363
rect 665 71 748 224
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 19 441 80 545
rect 115 476 181 649
rect 283 479 344 545
rect 19 406 261 441
rect 195 204 261 406
rect 19 164 261 204
rect 295 322 344 479
rect 397 399 469 438
rect 565 433 631 649
rect 397 365 631 399
rect 582 325 631 365
rect 295 276 548 322
rect 19 61 82 164
rect 117 17 183 130
rect 295 127 344 276
rect 582 259 656 325
rect 582 242 631 259
rect 397 208 631 242
rect 397 142 469 208
rect 283 61 344 127
rect 565 17 631 174
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel locali s 20 238 146 372 6 A
port 1 nsew signal input
rlabel locali s 690 224 748 363 6 X
port 2 nsew signal output
rlabel locali s 665 363 748 612 6 X
port 2 nsew signal output
rlabel locali s 665 71 748 224 6 X
port 2 nsew signal output
rlabel metal1 s 0 -49 768 49 8 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 617 768 715 6 VPWR
port 4 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 2239424
string GDS_START 2232990
<< end >>
