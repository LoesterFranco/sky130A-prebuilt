magic
tech sky130A
magscale 1 2
timestamp 1604502710
<< nwell >>
rect -38 332 902 704
<< pwell >>
rect 0 0 864 49
<< scpmos >>
rect 83 392 119 592
rect 183 392 219 592
rect 425 392 461 592
rect 525 392 561 592
rect 625 392 661 592
rect 745 392 781 592
<< nmoslvt >>
rect 89 74 119 202
rect 167 74 197 202
rect 431 74 461 202
rect 509 74 539 202
rect 667 74 697 202
rect 745 74 775 202
<< ndiff >>
rect 32 188 89 202
rect 32 154 44 188
rect 78 154 89 188
rect 32 120 89 154
rect 32 86 44 120
rect 78 86 89 120
rect 32 74 89 86
rect 119 74 167 202
rect 197 120 431 202
rect 197 86 208 120
rect 242 86 297 120
rect 331 86 386 120
rect 420 86 431 120
rect 197 74 431 86
rect 461 74 509 202
rect 539 190 667 202
rect 539 156 550 190
rect 584 156 622 190
rect 656 156 667 190
rect 539 116 667 156
rect 539 82 550 116
rect 584 82 622 116
rect 656 82 667 116
rect 539 74 667 82
rect 697 74 745 202
rect 775 188 832 202
rect 775 154 786 188
rect 820 154 832 188
rect 775 120 832 154
rect 775 86 786 120
rect 820 86 832 120
rect 775 74 832 86
<< pdiff >>
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 511 83 546
rect 27 477 39 511
rect 73 477 83 511
rect 27 442 83 477
rect 27 408 39 442
rect 73 408 83 442
rect 27 392 83 408
rect 119 580 183 592
rect 119 546 139 580
rect 173 546 183 580
rect 119 510 183 546
rect 119 476 139 510
rect 173 476 183 510
rect 119 392 183 476
rect 219 531 285 592
rect 219 497 239 531
rect 273 497 285 531
rect 219 442 285 497
rect 219 408 239 442
rect 273 408 285 442
rect 219 392 285 408
rect 369 531 425 592
rect 369 497 381 531
rect 415 497 425 531
rect 369 442 425 497
rect 369 408 381 442
rect 415 408 425 442
rect 369 392 425 408
rect 461 580 525 592
rect 461 546 481 580
rect 515 546 525 580
rect 461 510 525 546
rect 461 476 481 510
rect 515 476 525 510
rect 461 392 525 476
rect 561 580 625 592
rect 561 546 581 580
rect 615 546 625 580
rect 561 511 625 546
rect 561 477 581 511
rect 615 477 625 511
rect 561 442 625 477
rect 561 408 581 442
rect 615 408 625 442
rect 561 392 625 408
rect 661 580 745 592
rect 661 546 681 580
rect 715 546 745 580
rect 661 510 745 546
rect 661 476 681 510
rect 715 476 745 510
rect 661 392 745 476
rect 781 580 837 592
rect 781 546 791 580
rect 825 546 837 580
rect 781 511 837 546
rect 781 477 791 511
rect 825 477 837 511
rect 781 442 837 477
rect 781 408 791 442
rect 825 408 837 442
rect 781 392 837 408
<< ndiffc >>
rect 44 154 78 188
rect 44 86 78 120
rect 208 86 242 120
rect 297 86 331 120
rect 386 86 420 120
rect 550 156 584 190
rect 622 156 656 190
rect 550 82 584 116
rect 622 82 656 116
rect 786 154 820 188
rect 786 86 820 120
<< pdiffc >>
rect 39 546 73 580
rect 39 477 73 511
rect 39 408 73 442
rect 139 546 173 580
rect 139 476 173 510
rect 239 497 273 531
rect 239 408 273 442
rect 381 497 415 531
rect 381 408 415 442
rect 481 546 515 580
rect 481 476 515 510
rect 581 546 615 580
rect 581 477 615 511
rect 581 408 615 442
rect 681 546 715 580
rect 681 476 715 510
rect 791 546 825 580
rect 791 477 825 511
rect 791 408 825 442
<< poly >>
rect 83 592 119 618
rect 183 592 219 618
rect 425 592 461 618
rect 525 592 561 618
rect 625 592 661 618
rect 745 592 781 618
rect 83 290 119 392
rect 183 358 219 392
rect 425 358 461 392
rect 525 358 561 392
rect 625 358 661 392
rect 53 274 119 290
rect 53 240 69 274
rect 103 240 119 274
rect 53 224 119 240
rect 89 202 119 224
rect 167 342 263 358
rect 167 308 213 342
rect 247 308 263 342
rect 167 274 263 308
rect 167 240 213 274
rect 247 240 263 274
rect 167 224 263 240
rect 395 342 461 358
rect 395 308 411 342
rect 445 308 461 342
rect 395 274 461 308
rect 395 240 411 274
rect 445 240 461 274
rect 395 224 461 240
rect 167 202 197 224
rect 431 202 461 224
rect 509 342 575 358
rect 509 308 525 342
rect 559 308 575 342
rect 509 274 575 308
rect 509 240 525 274
rect 559 240 575 274
rect 509 224 575 240
rect 625 342 697 358
rect 625 308 647 342
rect 681 308 697 342
rect 625 274 697 308
rect 625 240 647 274
rect 681 240 697 274
rect 625 224 697 240
rect 509 202 539 224
rect 667 202 697 224
rect 745 302 781 392
rect 745 286 843 302
rect 745 252 793 286
rect 827 252 843 286
rect 745 236 843 252
rect 745 202 775 236
rect 89 48 119 74
rect 167 48 197 74
rect 431 48 461 74
rect 509 48 539 74
rect 667 48 697 74
rect 745 48 775 74
<< polycont >>
rect 69 240 103 274
rect 213 308 247 342
rect 213 240 247 274
rect 411 308 445 342
rect 411 240 445 274
rect 525 308 559 342
rect 525 240 559 274
rect 647 308 681 342
rect 647 240 681 274
rect 793 252 827 286
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 23 580 89 596
rect 23 546 39 580
rect 73 546 89 580
rect 23 511 89 546
rect 23 477 39 511
rect 73 477 89 511
rect 23 442 89 477
rect 123 581 531 615
rect 123 580 189 581
rect 123 546 139 580
rect 173 546 189 580
rect 465 580 531 581
rect 123 510 189 546
rect 123 476 139 510
rect 173 476 189 510
rect 123 460 189 476
rect 223 531 331 547
rect 223 497 239 531
rect 273 497 331 531
rect 23 408 39 442
rect 73 426 89 442
rect 223 442 331 497
rect 223 426 239 442
rect 73 408 239 426
rect 273 408 331 442
rect 23 392 331 408
rect 365 531 431 547
rect 365 497 381 531
rect 415 497 431 531
rect 365 442 431 497
rect 465 546 481 580
rect 515 546 531 580
rect 465 510 531 546
rect 465 476 481 510
rect 515 476 531 510
rect 465 460 531 476
rect 565 580 631 596
rect 565 546 581 580
rect 615 546 631 580
rect 565 511 631 546
rect 565 477 581 511
rect 615 477 631 511
rect 365 408 381 442
rect 415 426 431 442
rect 565 442 631 477
rect 665 580 731 649
rect 665 546 681 580
rect 715 546 731 580
rect 665 510 731 546
rect 665 476 681 510
rect 715 476 731 510
rect 665 460 731 476
rect 775 580 841 596
rect 775 546 791 580
rect 825 546 841 580
rect 775 511 841 546
rect 775 477 791 511
rect 825 477 841 511
rect 565 426 581 442
rect 415 408 581 426
rect 615 426 631 442
rect 775 442 841 477
rect 775 426 791 442
rect 615 408 791 426
rect 825 408 841 442
rect 365 392 841 408
rect 25 274 119 358
rect 25 240 69 274
rect 103 240 119 274
rect 25 224 119 240
rect 197 342 263 358
rect 197 308 213 342
rect 247 308 263 342
rect 197 274 263 308
rect 197 240 213 274
rect 247 240 263 274
rect 197 224 263 240
rect 297 356 331 392
rect 297 190 359 356
rect 395 342 461 358
rect 395 308 411 342
rect 445 308 461 342
rect 395 274 461 308
rect 395 240 411 274
rect 445 240 461 274
rect 395 224 461 240
rect 505 342 575 358
rect 505 308 525 342
rect 559 308 575 342
rect 505 274 575 308
rect 505 240 525 274
rect 559 240 575 274
rect 505 224 575 240
rect 631 342 743 358
rect 631 308 647 342
rect 681 308 743 342
rect 631 274 743 308
rect 631 240 647 274
rect 681 240 743 274
rect 631 224 743 240
rect 777 286 843 356
rect 777 252 793 286
rect 827 252 843 286
rect 777 236 843 252
rect 28 188 550 190
rect 28 154 44 188
rect 78 156 550 188
rect 584 156 622 190
rect 656 156 672 190
rect 78 154 94 156
rect 28 120 94 154
rect 28 86 44 120
rect 78 86 94 120
rect 28 70 94 86
rect 192 86 208 120
rect 242 86 297 120
rect 331 86 386 120
rect 420 86 436 120
rect 192 17 436 86
rect 505 116 672 156
rect 505 82 550 116
rect 584 82 622 116
rect 656 82 672 116
rect 505 66 672 82
rect 770 188 836 190
rect 770 154 786 188
rect 820 154 836 188
rect 770 120 836 154
rect 770 86 786 120
rect 820 86 836 120
rect 770 17 836 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 8 nsew
flabel nbase s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 9 nsew
rlabel comment s 0 0 0 0 4 a222oi_1
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 10 nsew
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 7 nsew
flabel corelocali s 223 242 257 276 0 FreeSans 340 0 0 0 C2
port 6 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 C2
port 6 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 C1
port 5 nsew
flabel corelocali s 511 242 545 276 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 799 242 833 276 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 703 242 737 276 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 319 168 353 202 0 FreeSans 340 0 0 0 Y
port 11 nsew
flabel corelocali s 319 242 353 276 0 FreeSans 340 0 0 0 Y
port 11 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 Y
port 11 nsew
flabel corelocali s 415 242 449 276 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 B2
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 864 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3567888
string GDS_START 3559246
<< end >>
