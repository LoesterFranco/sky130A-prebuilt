magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 828 561
rect 19 299 85 527
rect 19 17 85 161
rect 119 151 157 493
rect 203 367 253 527
rect 467 435 517 527
rect 667 435 717 527
rect 280 215 346 259
rect 400 199 467 325
rect 537 287 618 325
rect 537 199 571 287
rect 667 249 710 325
rect 617 215 710 249
rect 119 59 153 151
rect 667 149 710 215
rect 757 146 801 325
rect 187 17 253 93
rect 375 17 441 93
rect 0 -17 828 17
<< obsli1 >>
rect 291 333 357 485
rect 391 393 425 493
rect 559 393 593 493
rect 759 393 793 493
rect 391 359 793 393
rect 196 299 357 333
rect 196 161 230 299
rect 196 127 509 161
rect 299 51 341 127
rect 475 93 509 127
rect 475 59 809 93
<< metal1 >>
rect 0 496 828 592
rect 0 -48 828 48
<< labels >>
rlabel locali s 757 146 801 325 6 A1
port 1 nsew signal input
rlabel locali s 667 249 710 325 6 A2
port 2 nsew signal input
rlabel locali s 667 149 710 215 6 A2
port 2 nsew signal input
rlabel locali s 617 215 710 249 6 A2
port 2 nsew signal input
rlabel locali s 537 287 618 325 6 A3
port 3 nsew signal input
rlabel locali s 537 199 571 287 6 A3
port 3 nsew signal input
rlabel locali s 400 199 467 325 6 A4
port 4 nsew signal input
rlabel locali s 280 215 346 259 6 B1
port 5 nsew signal input
rlabel locali s 119 151 157 493 6 X
port 6 nsew signal output
rlabel locali s 119 59 153 151 6 X
port 6 nsew signal output
rlabel locali s 375 17 441 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 187 17 253 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 19 17 85 161 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 828 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 828 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 667 435 717 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 467 435 517 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 203 367 253 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 19 299 85 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 828 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 828 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3691120
string GDS_START 3682866
<< end >>
