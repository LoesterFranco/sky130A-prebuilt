magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 2630 704
rect 705 316 918 332
<< pwell >>
rect 0 0 2592 49
<< scnmos >>
rect 101 74 131 158
rect 179 74 209 158
rect 375 87 405 171
rect 461 87 491 171
rect 533 87 563 171
rect 733 74 763 222
rect 928 74 958 222
rect 1126 90 1156 174
rect 1319 90 1349 174
rect 1409 90 1439 174
rect 1545 90 1575 218
rect 1767 74 1797 222
rect 1865 74 1895 222
rect 1967 74 1997 158
rect 2045 74 2075 158
rect 2266 74 2296 158
rect 2464 74 2494 222
<< pmoshvt >>
rect 84 508 114 592
rect 162 508 192 592
rect 388 436 418 564
rect 524 436 554 520
rect 602 436 632 520
rect 797 352 827 576
rect 1067 368 1097 592
rect 1262 508 1292 592
rect 1352 508 1382 592
rect 1453 508 1483 592
rect 1562 405 1592 573
rect 1764 392 1794 592
rect 1951 392 1981 592
rect 2058 502 2088 586
rect 2142 502 2172 586
rect 2284 458 2314 586
rect 2478 368 2508 592
<< ndiff >>
rect 676 186 733 222
rect 44 132 101 158
rect 44 98 56 132
rect 90 98 101 132
rect 44 74 101 98
rect 131 74 179 158
rect 209 120 265 158
rect 209 86 220 120
rect 254 86 265 120
rect 319 146 375 171
rect 319 112 330 146
rect 364 112 375 146
rect 319 87 375 112
rect 405 146 461 171
rect 405 112 416 146
rect 450 112 461 146
rect 405 87 461 112
rect 491 87 533 171
rect 563 146 620 171
rect 563 112 574 146
rect 608 112 620 146
rect 563 87 620 112
rect 676 152 688 186
rect 722 152 733 186
rect 676 118 733 152
rect 209 74 265 86
rect 676 84 688 118
rect 722 84 733 118
rect 676 74 733 84
rect 763 202 818 222
rect 763 168 774 202
rect 808 168 818 202
rect 763 120 818 168
rect 763 86 774 120
rect 808 86 818 120
rect 763 74 818 86
rect 872 210 928 222
rect 872 176 883 210
rect 917 176 928 210
rect 872 120 928 176
rect 872 86 883 120
rect 917 86 928 120
rect 872 74 928 86
rect 958 210 1015 222
rect 958 176 969 210
rect 1003 176 1015 210
rect 958 120 1015 176
rect 1495 174 1545 218
rect 958 86 969 120
rect 1003 86 1015 120
rect 1069 157 1126 174
rect 1069 123 1081 157
rect 1115 123 1126 157
rect 1069 90 1126 123
rect 1156 153 1319 174
rect 1156 119 1261 153
rect 1295 119 1319 153
rect 1156 90 1319 119
rect 1349 90 1409 174
rect 1439 136 1545 174
rect 1439 102 1450 136
rect 1484 102 1545 136
rect 1439 90 1545 102
rect 1575 187 1632 218
rect 1575 153 1586 187
rect 1620 153 1632 187
rect 1575 90 1632 153
rect 1710 128 1767 222
rect 1710 94 1722 128
rect 1756 94 1767 128
rect 958 74 1015 86
rect 1710 74 1767 94
rect 1797 74 1865 222
rect 1895 200 1952 222
rect 1895 166 1906 200
rect 1940 166 1952 200
rect 1895 158 1952 166
rect 2407 210 2464 222
rect 2407 176 2419 210
rect 2453 176 2464 210
rect 1895 120 1967 158
rect 1895 86 1906 120
rect 1940 86 1967 120
rect 1895 74 1967 86
rect 1997 74 2045 158
rect 2075 117 2266 158
rect 2075 83 2086 117
rect 2120 83 2221 117
rect 2255 83 2266 117
rect 2075 74 2266 83
rect 2296 131 2353 158
rect 2296 97 2307 131
rect 2341 97 2353 131
rect 2296 74 2353 97
rect 2407 120 2464 176
rect 2407 86 2419 120
rect 2453 86 2464 120
rect 2407 74 2464 86
rect 2494 210 2565 222
rect 2494 176 2519 210
rect 2553 176 2565 210
rect 2494 120 2565 176
rect 2494 86 2519 120
rect 2553 86 2565 120
rect 2494 74 2565 86
<< pdiff >>
rect 27 567 84 592
rect 27 533 37 567
rect 71 533 84 567
rect 27 508 84 533
rect 114 508 162 592
rect 192 567 251 592
rect 192 533 205 567
rect 239 533 251 567
rect 1012 580 1067 592
rect 741 564 797 576
rect 192 508 251 533
rect 329 516 388 564
rect 329 482 341 516
rect 375 482 388 516
rect 329 436 388 482
rect 418 520 471 564
rect 741 530 750 564
rect 784 530 797 564
rect 418 508 524 520
rect 418 474 477 508
rect 511 474 524 508
rect 418 436 524 474
rect 554 436 602 520
rect 632 495 687 520
rect 632 461 645 495
rect 679 461 687 495
rect 632 436 687 461
rect 741 352 797 530
rect 827 405 882 576
rect 1012 546 1020 580
rect 1054 546 1067 580
rect 827 371 840 405
rect 874 371 882 405
rect 827 352 882 371
rect 1012 368 1067 546
rect 1097 421 1152 592
rect 1206 567 1262 592
rect 1206 533 1215 567
rect 1249 533 1262 567
rect 1206 508 1262 533
rect 1292 567 1352 592
rect 1292 533 1305 567
rect 1339 533 1352 567
rect 1292 508 1352 533
rect 1382 508 1453 592
rect 1483 584 1544 592
rect 1483 550 1498 584
rect 1532 573 1544 584
rect 1705 584 1764 592
rect 1532 550 1562 573
rect 1483 508 1562 550
rect 1097 387 1110 421
rect 1144 387 1152 421
rect 1097 368 1152 387
rect 1509 405 1562 508
rect 1592 448 1651 573
rect 1592 414 1605 448
rect 1639 414 1651 448
rect 1592 405 1651 414
rect 1705 550 1717 584
rect 1751 550 1764 584
rect 1705 392 1764 550
rect 1794 392 1951 592
rect 1981 586 2040 592
rect 1981 584 2058 586
rect 1981 550 1994 584
rect 2028 550 2058 584
rect 1981 511 2058 550
rect 1981 477 1994 511
rect 2028 502 2058 511
rect 2088 502 2142 586
rect 2172 555 2284 586
rect 2172 521 2211 555
rect 2245 521 2284 555
rect 2172 502 2284 521
rect 2028 477 2040 502
rect 1981 438 2040 477
rect 1981 404 1994 438
rect 2028 404 2040 438
rect 1981 392 2040 404
rect 2231 458 2284 502
rect 2314 574 2369 586
rect 2314 540 2327 574
rect 2361 540 2369 574
rect 2314 504 2369 540
rect 2314 470 2327 504
rect 2361 470 2369 504
rect 2314 458 2369 470
rect 2423 580 2478 592
rect 2423 546 2431 580
rect 2465 546 2478 580
rect 2423 497 2478 546
rect 2423 463 2431 497
rect 2465 463 2478 497
rect 2423 414 2478 463
rect 2423 380 2431 414
rect 2465 380 2478 414
rect 2423 368 2478 380
rect 2508 580 2565 592
rect 2508 546 2521 580
rect 2555 546 2565 580
rect 2508 497 2565 546
rect 2508 463 2521 497
rect 2555 463 2565 497
rect 2508 414 2565 463
rect 2508 380 2521 414
rect 2555 380 2565 414
rect 2508 368 2565 380
<< ndiffc >>
rect 56 98 90 132
rect 220 86 254 120
rect 330 112 364 146
rect 416 112 450 146
rect 574 112 608 146
rect 688 152 722 186
rect 688 84 722 118
rect 774 168 808 202
rect 774 86 808 120
rect 883 176 917 210
rect 883 86 917 120
rect 969 176 1003 210
rect 969 86 1003 120
rect 1081 123 1115 157
rect 1261 119 1295 153
rect 1450 102 1484 136
rect 1586 153 1620 187
rect 1722 94 1756 128
rect 1906 166 1940 200
rect 2419 176 2453 210
rect 1906 86 1940 120
rect 2086 83 2120 117
rect 2221 83 2255 117
rect 2307 97 2341 131
rect 2419 86 2453 120
rect 2519 176 2553 210
rect 2519 86 2553 120
<< pdiffc >>
rect 37 533 71 567
rect 205 533 239 567
rect 341 482 375 516
rect 750 530 784 564
rect 477 474 511 508
rect 645 461 679 495
rect 1020 546 1054 580
rect 840 371 874 405
rect 1215 533 1249 567
rect 1305 533 1339 567
rect 1498 550 1532 584
rect 1110 387 1144 421
rect 1605 414 1639 448
rect 1717 550 1751 584
rect 1994 550 2028 584
rect 1994 477 2028 511
rect 2211 521 2245 555
rect 1994 404 2028 438
rect 2327 540 2361 574
rect 2327 470 2361 504
rect 2431 546 2465 580
rect 2431 463 2465 497
rect 2431 380 2465 414
rect 2521 546 2555 580
rect 2521 463 2555 497
rect 2521 380 2555 414
<< poly >>
rect 84 592 114 618
rect 162 592 192 618
rect 388 564 418 590
rect 797 576 827 602
rect 1067 592 1097 618
rect 1262 592 1292 618
rect 1352 592 1382 618
rect 1453 592 1483 618
rect 84 493 114 508
rect 162 493 192 508
rect 81 398 117 493
rect 159 476 195 493
rect 159 446 225 476
rect 195 402 225 446
rect 524 520 554 546
rect 602 520 632 546
rect 388 421 418 436
rect 524 421 554 436
rect 602 421 632 436
rect 71 382 137 398
rect 71 348 87 382
rect 121 348 137 382
rect 71 314 137 348
rect 71 280 87 314
rect 121 280 137 314
rect 71 246 137 280
rect 195 386 261 402
rect 195 352 211 386
rect 245 352 261 386
rect 195 318 261 352
rect 195 284 211 318
rect 245 284 261 318
rect 333 391 557 421
rect 333 288 363 391
rect 599 343 635 421
rect 914 412 980 428
rect 914 378 930 412
rect 964 378 980 412
rect 411 327 491 343
rect 411 293 427 327
rect 461 293 491 327
rect 195 268 261 284
rect 303 272 369 288
rect 411 277 491 293
rect 71 212 87 246
rect 121 212 137 246
rect 303 238 319 272
rect 353 238 369 272
rect 303 220 369 238
rect 71 196 137 212
rect 101 158 131 196
rect 179 190 405 220
rect 179 158 209 190
rect 375 171 405 190
rect 461 171 491 277
rect 533 327 635 343
rect 797 337 827 352
rect 914 346 980 378
rect 1562 573 1592 599
rect 1764 592 1794 618
rect 1951 592 1981 618
rect 1262 493 1292 508
rect 1352 493 1382 508
rect 1453 493 1483 508
rect 1259 460 1295 493
rect 1349 466 1385 493
rect 1184 444 1295 460
rect 1184 410 1200 444
rect 1234 430 1295 444
rect 1337 450 1408 466
rect 1234 410 1250 430
rect 1184 394 1250 410
rect 1337 416 1358 450
rect 1392 416 1408 450
rect 1337 400 1408 416
rect 1067 353 1097 368
rect 1064 346 1100 353
rect 1337 346 1367 400
rect 914 344 1367 346
rect 533 293 549 327
rect 583 293 635 327
rect 794 310 830 337
rect 533 259 635 293
rect 533 225 549 259
rect 583 225 635 259
rect 690 294 830 310
rect 914 310 930 344
rect 964 316 1367 344
rect 964 310 980 316
rect 914 294 980 310
rect 690 260 706 294
rect 740 280 830 294
rect 740 260 763 280
rect 690 244 763 260
rect 533 209 635 225
rect 733 222 763 244
rect 928 222 958 294
rect 533 171 563 209
rect 101 48 131 74
rect 179 48 209 74
rect 375 61 405 87
rect 461 61 491 87
rect 533 61 563 87
rect 1126 174 1156 316
rect 1450 306 1486 493
rect 1562 390 1592 405
rect 2058 586 2088 612
rect 2142 586 2172 612
rect 2284 586 2314 612
rect 2478 592 2508 618
rect 2058 487 2088 502
rect 2142 487 2172 502
rect 1559 373 1595 390
rect 1764 377 1794 392
rect 1951 377 1981 392
rect 1540 357 1606 373
rect 1540 323 1556 357
rect 1590 323 1606 357
rect 1540 307 1606 323
rect 1761 321 1797 377
rect 1948 360 1984 377
rect 1409 290 1492 306
rect 1301 246 1367 262
rect 1301 212 1317 246
rect 1351 212 1367 246
rect 1301 196 1367 212
rect 1409 256 1442 290
rect 1476 256 1492 290
rect 1409 240 1492 256
rect 1319 174 1349 196
rect 1409 174 1439 240
rect 1545 218 1575 307
rect 1654 305 1797 321
rect 1947 344 2013 360
rect 1947 310 1963 344
rect 1997 310 2013 344
rect 1654 271 1670 305
rect 1704 271 1738 305
rect 1772 271 1797 305
rect 1654 255 1797 271
rect 1767 222 1797 255
rect 1839 294 1905 310
rect 1947 294 2013 310
rect 2055 317 2091 487
rect 2139 470 2175 487
rect 2133 454 2199 470
rect 2133 420 2149 454
rect 2183 420 2199 454
rect 2284 443 2314 458
rect 2133 404 2199 420
rect 2055 301 2121 317
rect 1839 260 1855 294
rect 1889 260 1905 294
rect 1839 244 1905 260
rect 1865 222 1895 244
rect 733 48 763 74
rect 928 48 958 74
rect 1126 64 1156 90
rect 1319 64 1349 90
rect 1409 64 1439 90
rect 1545 64 1575 90
rect 1967 158 1997 294
rect 2055 267 2071 301
rect 2105 267 2121 301
rect 2055 251 2121 267
rect 2163 203 2193 404
rect 2281 267 2317 443
rect 2478 353 2508 368
rect 2475 267 2511 353
rect 2045 173 2193 203
rect 2235 251 2511 267
rect 2235 217 2251 251
rect 2285 237 2511 251
rect 2285 217 2317 237
rect 2464 222 2494 237
rect 2235 201 2317 217
rect 2045 158 2075 173
rect 2266 158 2296 201
rect 1767 48 1797 74
rect 1865 48 1895 74
rect 1967 48 1997 74
rect 2045 48 2075 74
rect 2266 48 2296 74
rect 2464 48 2494 74
<< polycont >>
rect 87 348 121 382
rect 87 280 121 314
rect 211 352 245 386
rect 211 284 245 318
rect 930 378 964 412
rect 427 293 461 327
rect 87 212 121 246
rect 319 238 353 272
rect 1200 410 1234 444
rect 1358 416 1392 450
rect 549 293 583 327
rect 549 225 583 259
rect 930 310 964 344
rect 706 260 740 294
rect 1556 323 1590 357
rect 1317 212 1351 246
rect 1442 256 1476 290
rect 1963 310 1997 344
rect 1670 271 1704 305
rect 1738 271 1772 305
rect 2149 420 2183 454
rect 1855 260 1889 294
rect 2071 267 2105 301
rect 2251 217 2285 251
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2592 683
rect 17 567 87 596
rect 17 533 37 567
rect 71 533 87 567
rect 17 470 87 533
rect 189 567 239 649
rect 189 533 205 567
rect 189 504 239 533
rect 273 581 443 615
rect 273 470 307 581
rect 17 436 307 470
rect 341 516 375 547
rect 17 162 51 436
rect 85 382 161 398
rect 85 348 87 382
rect 121 348 161 382
rect 85 314 161 348
rect 85 280 87 314
rect 121 280 161 314
rect 85 246 161 280
rect 85 212 87 246
rect 121 212 161 246
rect 85 196 161 212
rect 195 386 261 402
rect 195 352 211 386
rect 245 356 261 386
rect 341 356 375 482
rect 409 424 443 581
rect 477 508 527 649
rect 734 564 800 649
rect 734 530 750 564
rect 784 530 800 564
rect 1004 580 1054 649
rect 1004 546 1020 580
rect 1004 530 1054 546
rect 1199 567 1249 596
rect 1199 538 1215 567
rect 1088 533 1215 538
rect 511 474 527 508
rect 477 458 527 474
rect 620 496 695 524
rect 1088 504 1249 533
rect 1283 567 1355 596
rect 1283 533 1305 567
rect 1339 533 1355 567
rect 1482 584 1548 649
rect 1482 550 1498 584
rect 1532 550 1548 584
rect 1701 584 1767 649
rect 1701 550 1717 584
rect 1751 550 1767 584
rect 1994 584 2044 600
rect 2028 550 2044 584
rect 1283 504 1355 533
rect 1088 496 1122 504
rect 620 495 1122 496
rect 620 461 645 495
rect 679 462 1122 495
rect 679 461 695 462
rect 620 424 695 461
rect 409 390 654 424
rect 245 352 477 356
rect 195 327 477 352
rect 195 322 427 327
rect 195 318 261 322
rect 195 284 211 318
rect 245 284 261 318
rect 411 293 427 322
rect 461 293 477 327
rect 195 188 261 284
rect 303 272 369 288
rect 411 277 477 293
rect 511 350 586 356
rect 545 327 586 350
rect 545 316 549 327
rect 511 293 549 316
rect 583 293 586 327
rect 303 238 319 272
rect 353 238 369 272
rect 303 222 369 238
rect 511 259 586 293
rect 511 225 549 259
rect 583 225 586 259
rect 511 209 586 225
rect 17 132 106 162
rect 195 154 364 188
rect 620 175 654 390
rect 790 412 980 428
rect 790 405 930 412
rect 790 371 840 405
rect 874 378 930 405
rect 964 378 980 412
rect 874 371 980 378
rect 790 344 980 371
rect 790 310 930 344
rect 964 310 980 344
rect 690 294 756 310
rect 690 260 706 294
rect 740 260 756 294
rect 690 236 756 260
rect 790 294 980 310
rect 1026 330 1060 462
rect 1165 444 1249 460
rect 1165 428 1200 444
rect 1094 421 1200 428
rect 1094 387 1110 421
rect 1144 410 1200 421
rect 1234 410 1249 444
rect 1144 394 1249 410
rect 1144 387 1199 394
rect 1094 364 1199 387
rect 1026 296 1131 330
rect 790 202 824 294
rect 17 98 56 132
rect 90 98 106 132
rect 314 146 364 154
rect 17 68 106 98
rect 204 86 220 120
rect 254 86 270 120
rect 204 17 270 86
rect 314 112 330 146
rect 314 83 364 112
rect 400 146 466 175
rect 400 112 416 146
rect 450 112 466 146
rect 400 17 466 112
rect 558 146 654 175
rect 558 112 574 146
rect 608 112 654 146
rect 558 83 654 112
rect 688 186 722 202
rect 688 118 722 152
rect 688 17 722 84
rect 758 168 774 202
rect 808 168 824 202
rect 758 120 824 168
rect 758 86 774 120
rect 808 86 824 120
rect 758 70 824 86
rect 867 210 917 226
rect 867 176 883 210
rect 867 120 917 176
rect 867 86 883 120
rect 867 17 917 86
rect 953 210 1019 226
rect 953 176 969 210
rect 1003 176 1019 210
rect 953 120 1019 176
rect 953 86 969 120
rect 1003 86 1019 120
rect 1065 157 1131 296
rect 1065 123 1081 157
rect 1115 123 1131 157
rect 1065 119 1131 123
rect 953 85 1019 86
rect 1165 85 1199 364
rect 1283 360 1317 504
rect 1389 482 1960 516
rect 1389 466 1423 482
rect 1351 450 1423 466
rect 1351 416 1358 450
rect 1392 416 1423 450
rect 1351 400 1423 416
rect 1589 414 1605 448
rect 1639 414 1688 448
rect 1540 360 1606 366
rect 1233 357 1606 360
rect 1233 326 1556 357
rect 1233 153 1267 326
rect 1540 323 1556 326
rect 1590 323 1606 357
rect 1654 321 1688 414
rect 1926 345 1960 482
rect 1994 511 2044 550
rect 2028 477 2044 511
rect 2169 555 2277 649
rect 2169 521 2211 555
rect 2245 521 2277 555
rect 2169 505 2277 521
rect 2311 574 2377 590
rect 2311 540 2327 574
rect 2361 540 2377 574
rect 1994 438 2044 477
rect 2311 504 2377 540
rect 2311 470 2327 504
rect 2361 470 2377 504
rect 2311 464 2377 470
rect 2028 419 2044 438
rect 2133 454 2377 464
rect 2133 420 2149 454
rect 2183 420 2377 454
rect 2133 419 2377 420
rect 2028 404 2081 419
rect 1994 385 2081 404
rect 2047 351 2189 385
rect 1926 344 2013 345
rect 1654 305 1788 321
rect 1926 310 1963 344
rect 1997 310 2013 344
rect 1426 290 1492 292
rect 1301 246 1392 262
rect 1426 256 1442 290
rect 1476 289 1492 290
rect 1654 289 1670 305
rect 1476 271 1670 289
rect 1704 271 1738 305
rect 1772 271 1788 305
rect 1476 256 1788 271
rect 1426 255 1788 256
rect 1822 294 1892 310
rect 1926 309 2013 310
rect 1822 260 1855 294
rect 1889 275 1892 294
rect 2055 301 2121 317
rect 2055 275 2071 301
rect 1889 267 2071 275
rect 2105 267 2121 301
rect 1889 260 2121 267
rect 1301 212 1317 246
rect 1351 221 1392 246
rect 1351 212 1552 221
rect 1301 187 1552 212
rect 1233 119 1261 153
rect 1295 119 1324 153
rect 1358 85 1392 187
rect 953 51 1392 85
rect 1434 136 1484 153
rect 1434 102 1450 136
rect 1434 17 1484 102
rect 1518 85 1552 187
rect 1586 187 1620 255
rect 1822 241 2121 260
rect 2155 267 2189 351
rect 2329 350 2377 419
rect 2329 316 2335 350
rect 2369 316 2377 350
rect 2329 310 2377 316
rect 2415 580 2481 596
rect 2415 546 2431 580
rect 2465 546 2481 580
rect 2415 497 2481 546
rect 2415 463 2431 497
rect 2465 463 2481 497
rect 2415 414 2481 463
rect 2415 380 2431 414
rect 2465 380 2481 414
rect 2415 310 2481 380
rect 2521 580 2571 649
rect 2555 546 2571 580
rect 2521 497 2571 546
rect 2555 463 2571 497
rect 2521 414 2571 463
rect 2555 380 2571 414
rect 2521 364 2571 380
rect 2155 251 2301 267
rect 1822 221 1856 241
rect 1586 119 1620 153
rect 1654 187 1856 221
rect 2155 217 2251 251
rect 2285 217 2301 251
rect 2155 201 2301 217
rect 1890 200 2189 201
rect 1654 85 1688 187
rect 1890 166 1906 200
rect 1940 167 2189 200
rect 1940 166 1956 167
rect 1518 51 1688 85
rect 1722 128 1772 153
rect 1756 94 1772 128
rect 1722 17 1772 94
rect 1890 120 1956 166
rect 2335 162 2369 310
rect 2415 226 2469 310
rect 1890 86 1906 120
rect 1940 86 1956 120
rect 1890 70 1956 86
rect 2070 117 2262 133
rect 2070 83 2086 117
rect 2120 83 2221 117
rect 2255 83 2262 117
rect 2070 17 2262 83
rect 2298 131 2369 162
rect 2298 97 2307 131
rect 2341 97 2369 131
rect 2298 67 2369 97
rect 2403 210 2469 226
rect 2403 176 2419 210
rect 2453 176 2469 210
rect 2403 120 2469 176
rect 2403 86 2419 120
rect 2453 86 2469 120
rect 2403 70 2469 86
rect 2503 210 2569 226
rect 2503 176 2519 210
rect 2553 176 2569 210
rect 2503 120 2569 176
rect 2503 86 2519 120
rect 2553 86 2569 120
rect 2503 17 2569 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2592 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 511 316 545 350
rect 2335 316 2369 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
<< metal1 >>
rect 0 683 2592 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2592 683
rect 0 617 2592 649
rect 499 350 557 356
rect 499 316 511 350
rect 545 347 557 350
rect 2323 350 2381 356
rect 2323 347 2335 350
rect 545 319 2335 347
rect 545 316 557 319
rect 499 310 557 316
rect 2323 316 2335 319
rect 2369 316 2381 350
rect 2323 310 2381 316
rect 0 17 2592 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2592 17
rect 0 -49 2592 -17
<< labels >>
rlabel comment s 0 0 0 0 4 edfxtp_1
flabel comment s 1135 336 1135 336 0 FreeSans 200 0 0 0 no_jumper_check
flabel pwell s 0 0 2592 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 0 617 2592 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 2592 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 2592 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 319 242 353 276 0 FreeSans 340 0 0 0 DE
port 3 nsew
flabel corelocali s 127 242 161 276 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 703 242 737 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 2431 316 2465 350 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 2431 390 2465 424 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 2431 464 2465 498 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 2431 538 2465 572 0 FreeSans 340 0 0 0 Q
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 2592 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2149800
string GDS_START 2131308
<< end >>
