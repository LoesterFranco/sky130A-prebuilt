magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1196 561
rect 17 299 69 527
rect 103 333 169 493
rect 203 367 253 527
rect 375 333 441 425
rect 103 301 441 333
rect 122 289 441 301
rect 991 357 1057 527
rect 21 215 88 255
rect 122 177 169 289
rect 300 215 465 255
rect 519 215 716 255
rect 756 215 908 255
rect 944 215 1179 255
rect 103 127 169 177
rect 291 17 341 109
rect 475 17 509 109
rect 643 17 690 109
rect 839 17 873 109
rect 1007 17 1041 109
rect 0 -17 1196 17
<< obsli1 >>
rect 291 459 509 493
rect 291 367 341 459
rect 475 323 509 459
rect 543 459 889 493
rect 543 367 609 459
rect 643 323 693 425
rect 475 289 693 323
rect 739 323 789 425
rect 823 367 889 459
rect 923 323 957 493
rect 1091 323 1141 493
rect 739 289 1141 323
rect 17 93 69 181
rect 203 147 1141 181
rect 203 93 253 147
rect 17 51 253 93
rect 375 51 441 147
rect 543 51 609 147
rect 739 51 805 147
rect 907 51 973 147
rect 1075 51 1141 147
<< metal1 >>
rect 0 496 1196 592
rect 0 -48 1196 48
<< labels >>
rlabel locali s 944 215 1179 255 6 A1
port 1 nsew signal input
rlabel locali s 756 215 908 255 6 A2
port 2 nsew signal input
rlabel locali s 519 215 716 255 6 A3
port 3 nsew signal input
rlabel locali s 300 215 465 255 6 A4
port 4 nsew signal input
rlabel locali s 21 215 88 255 6 B1
port 5 nsew signal input
rlabel locali s 375 333 441 425 6 Y
port 6 nsew signal output
rlabel locali s 122 289 441 301 6 Y
port 6 nsew signal output
rlabel locali s 122 177 169 289 6 Y
port 6 nsew signal output
rlabel locali s 103 333 169 493 6 Y
port 6 nsew signal output
rlabel locali s 103 301 441 333 6 Y
port 6 nsew signal output
rlabel locali s 103 127 169 177 6 Y
port 6 nsew signal output
rlabel locali s 1007 17 1041 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 839 17 873 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 643 17 690 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 475 17 509 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 291 17 341 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 1196 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1196 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 991 357 1057 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 203 367 253 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 17 299 69 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 1196 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 1196 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 972736
string GDS_START 961692
<< end >>
