magic
tech sky130A
magscale 1 2
timestamp 1599588209
<< nwell >>
rect -38 332 2534 704
<< pwell >>
rect 0 0 2496 49
<< scpmos >>
rect 108 464 138 592
rect 208 464 238 592
rect 292 464 322 592
rect 382 464 412 592
rect 490 464 520 592
rect 638 368 668 592
rect 892 368 922 592
rect 1094 506 1124 590
rect 1184 506 1214 590
rect 1292 506 1322 590
rect 1416 423 1446 591
rect 1626 423 1656 591
rect 1734 476 1764 560
rect 1818 476 1848 560
rect 1919 392 1949 560
rect 2009 392 2039 560
rect 2110 368 2140 592
rect 2200 368 2230 592
rect 2290 368 2320 592
rect 2380 368 2410 592
<< nmoslvt >>
rect 93 74 123 158
rect 193 74 223 158
rect 271 74 301 158
rect 422 74 452 158
rect 500 74 530 158
rect 600 74 630 222
rect 798 74 828 222
rect 996 100 1026 184
rect 1132 100 1162 184
rect 1257 100 1287 184
rect 1441 74 1471 184
rect 1557 74 1587 184
rect 1736 74 1766 158
rect 1814 74 1844 158
rect 2012 74 2042 222
rect 2107 74 2137 222
rect 2210 74 2240 222
rect 2296 74 2326 222
rect 2382 74 2412 222
<< ndiff >>
rect 550 158 600 222
rect 36 130 93 158
rect 36 96 48 130
rect 82 96 93 130
rect 36 74 93 96
rect 123 130 193 158
rect 123 96 148 130
rect 182 96 193 130
rect 123 74 193 96
rect 223 74 271 158
rect 301 128 422 158
rect 301 94 344 128
rect 378 94 422 128
rect 301 74 422 94
rect 452 74 500 158
rect 530 133 600 158
rect 530 99 541 133
rect 575 99 600 133
rect 530 74 600 99
rect 630 202 687 222
rect 630 168 641 202
rect 675 168 687 202
rect 630 120 687 168
rect 630 86 641 120
rect 675 86 687 120
rect 630 74 687 86
rect 741 127 798 222
rect 741 93 753 127
rect 787 93 798 127
rect 741 74 798 93
rect 828 210 885 222
rect 828 176 839 210
rect 873 176 885 210
rect 828 120 885 176
rect 828 86 839 120
rect 873 86 885 120
rect 939 170 996 184
rect 939 136 951 170
rect 985 136 996 170
rect 939 100 996 136
rect 1026 170 1132 184
rect 1026 136 1087 170
rect 1121 136 1132 170
rect 1026 100 1132 136
rect 1162 100 1257 184
rect 1287 120 1441 184
rect 1287 100 1314 120
rect 828 74 885 86
rect 1302 86 1314 100
rect 1348 86 1441 120
rect 1302 74 1441 86
rect 1471 161 1557 184
rect 1471 127 1494 161
rect 1528 127 1557 161
rect 1471 74 1557 127
rect 1587 158 1721 184
rect 1955 210 2012 222
rect 1955 176 1967 210
rect 2001 176 2012 210
rect 1587 140 1736 158
rect 1587 106 1675 140
rect 1709 106 1736 140
rect 1587 74 1736 106
rect 1766 74 1814 158
rect 1844 125 1901 158
rect 1844 91 1855 125
rect 1889 91 1901 125
rect 1844 74 1901 91
rect 1955 120 2012 176
rect 1955 86 1967 120
rect 2001 86 2012 120
rect 1955 74 2012 86
rect 2042 192 2107 222
rect 2042 158 2053 192
rect 2087 158 2107 192
rect 2042 116 2107 158
rect 2042 82 2053 116
rect 2087 82 2107 116
rect 2042 74 2107 82
rect 2137 210 2210 222
rect 2137 176 2165 210
rect 2199 176 2210 210
rect 2137 120 2210 176
rect 2137 86 2165 120
rect 2199 86 2210 120
rect 2137 74 2210 86
rect 2240 123 2296 222
rect 2240 89 2251 123
rect 2285 89 2296 123
rect 2240 74 2296 89
rect 2326 210 2382 222
rect 2326 176 2337 210
rect 2371 176 2382 210
rect 2326 120 2382 176
rect 2326 86 2337 120
rect 2371 86 2382 120
rect 2326 74 2382 86
rect 2412 131 2469 222
rect 2412 97 2423 131
rect 2457 97 2469 131
rect 2412 74 2469 97
<< pdiff >>
rect 1340 621 1398 633
rect 49 580 108 592
rect 49 546 61 580
rect 95 546 108 580
rect 49 510 108 546
rect 49 476 61 510
rect 95 476 108 510
rect 49 464 108 476
rect 138 580 208 592
rect 138 546 161 580
rect 195 546 208 580
rect 138 510 208 546
rect 138 476 161 510
rect 195 476 208 510
rect 138 464 208 476
rect 238 464 292 592
rect 322 580 382 592
rect 322 546 335 580
rect 369 546 382 580
rect 322 512 382 546
rect 322 478 335 512
rect 369 478 382 512
rect 322 464 382 478
rect 412 464 490 592
rect 520 580 638 592
rect 520 546 562 580
rect 596 546 638 580
rect 520 464 638 546
rect 585 368 638 464
rect 668 421 727 592
rect 668 387 681 421
rect 715 387 727 421
rect 668 368 727 387
rect 781 580 892 592
rect 781 546 819 580
rect 853 546 892 580
rect 781 368 892 546
rect 922 421 981 592
rect 1340 590 1352 621
rect 1035 568 1094 590
rect 1035 534 1047 568
rect 1081 534 1094 568
rect 1035 506 1094 534
rect 1124 565 1184 590
rect 1124 531 1137 565
rect 1171 531 1184 565
rect 1124 506 1184 531
rect 1214 506 1292 590
rect 1322 587 1352 590
rect 1386 591 1398 621
rect 1386 587 1416 591
rect 1322 506 1416 587
rect 922 387 935 421
rect 969 387 981 421
rect 922 368 981 387
rect 1363 423 1416 506
rect 1446 469 1626 591
rect 1446 435 1480 469
rect 1514 435 1626 469
rect 1446 423 1626 435
rect 1656 560 1716 591
rect 2057 560 2110 592
rect 1656 548 1734 560
rect 1656 514 1670 548
rect 1704 514 1734 548
rect 1656 476 1734 514
rect 1764 476 1818 560
rect 1848 535 1919 560
rect 1848 501 1861 535
rect 1895 501 1919 535
rect 1848 476 1919 501
rect 1656 469 1716 476
rect 1656 435 1670 469
rect 1704 435 1716 469
rect 1656 423 1716 435
rect 1866 392 1919 476
rect 1949 548 2009 560
rect 1949 514 1962 548
rect 1996 514 2009 548
rect 1949 444 2009 514
rect 1949 410 1962 444
rect 1996 410 2009 444
rect 1949 392 2009 410
rect 2039 548 2110 560
rect 2039 514 2061 548
rect 2095 514 2110 548
rect 2039 438 2110 514
rect 2039 404 2061 438
rect 2095 404 2110 438
rect 2039 392 2110 404
rect 2057 368 2110 392
rect 2140 580 2200 592
rect 2140 546 2153 580
rect 2187 546 2200 580
rect 2140 497 2200 546
rect 2140 463 2153 497
rect 2187 463 2200 497
rect 2140 414 2200 463
rect 2140 380 2153 414
rect 2187 380 2200 414
rect 2140 368 2200 380
rect 2230 580 2290 592
rect 2230 546 2243 580
rect 2277 546 2290 580
rect 2230 478 2290 546
rect 2230 444 2243 478
rect 2277 444 2290 478
rect 2230 368 2290 444
rect 2320 580 2380 592
rect 2320 546 2333 580
rect 2367 546 2380 580
rect 2320 497 2380 546
rect 2320 463 2333 497
rect 2367 463 2380 497
rect 2320 414 2380 463
rect 2320 380 2333 414
rect 2367 380 2380 414
rect 2320 368 2380 380
rect 2410 580 2469 592
rect 2410 546 2423 580
rect 2457 546 2469 580
rect 2410 471 2469 546
rect 2410 437 2423 471
rect 2457 437 2469 471
rect 2410 368 2469 437
<< ndiffc >>
rect 48 96 82 130
rect 148 96 182 130
rect 344 94 378 128
rect 541 99 575 133
rect 641 168 675 202
rect 641 86 675 120
rect 753 93 787 127
rect 839 176 873 210
rect 839 86 873 120
rect 951 136 985 170
rect 1087 136 1121 170
rect 1314 86 1348 120
rect 1494 127 1528 161
rect 1967 176 2001 210
rect 1675 106 1709 140
rect 1855 91 1889 125
rect 1967 86 2001 120
rect 2053 158 2087 192
rect 2053 82 2087 116
rect 2165 176 2199 210
rect 2165 86 2199 120
rect 2251 89 2285 123
rect 2337 176 2371 210
rect 2337 86 2371 120
rect 2423 97 2457 131
<< pdiffc >>
rect 61 546 95 580
rect 61 476 95 510
rect 161 546 195 580
rect 161 476 195 510
rect 335 546 369 580
rect 335 478 369 512
rect 562 546 596 580
rect 681 387 715 421
rect 819 546 853 580
rect 1047 534 1081 568
rect 1137 531 1171 565
rect 1352 587 1386 621
rect 935 387 969 421
rect 1480 435 1514 469
rect 1670 514 1704 548
rect 1861 501 1895 535
rect 1670 435 1704 469
rect 1962 514 1996 548
rect 1962 410 1996 444
rect 2061 514 2095 548
rect 2061 404 2095 438
rect 2153 546 2187 580
rect 2153 463 2187 497
rect 2153 380 2187 414
rect 2243 546 2277 580
rect 2243 444 2277 478
rect 2333 546 2367 580
rect 2333 463 2367 497
rect 2333 380 2367 414
rect 2423 546 2457 580
rect 2423 437 2457 471
<< poly >>
rect 108 592 138 618
rect 208 592 238 618
rect 292 592 322 618
rect 382 592 412 618
rect 490 592 520 618
rect 638 592 668 618
rect 892 592 922 618
rect 108 449 138 464
rect 208 449 238 464
rect 292 449 322 464
rect 382 449 412 464
rect 490 449 520 464
rect 39 419 241 449
rect 39 257 69 419
rect 117 355 223 371
rect 289 357 325 449
rect 379 428 415 449
rect 373 412 439 428
rect 373 378 389 412
rect 423 378 439 412
rect 117 321 133 355
rect 167 321 223 355
rect 117 305 223 321
rect 39 241 151 257
rect 39 227 101 241
rect 85 207 101 227
rect 135 207 151 241
rect 85 191 151 207
rect 93 158 123 191
rect 193 158 223 305
rect 265 341 331 357
rect 265 307 281 341
rect 315 307 331 341
rect 265 291 331 307
rect 373 344 439 378
rect 373 310 389 344
rect 423 310 439 344
rect 487 388 523 449
rect 487 372 553 388
rect 487 338 503 372
rect 537 338 553 372
rect 1094 590 1124 616
rect 1184 590 1214 616
rect 1292 590 1322 616
rect 1416 591 1446 617
rect 1626 591 1656 617
rect 2110 592 2140 618
rect 2200 592 2230 618
rect 2290 592 2320 618
rect 2380 592 2410 618
rect 1094 491 1124 506
rect 1184 491 1214 506
rect 1292 491 1322 506
rect 1091 474 1127 491
rect 1015 458 1127 474
rect 1015 424 1031 458
rect 1065 444 1127 458
rect 1181 456 1217 491
rect 1065 424 1081 444
rect 1015 408 1081 424
rect 1181 440 1247 456
rect 1181 406 1197 440
rect 1231 406 1247 440
rect 638 353 668 368
rect 892 353 922 368
rect 1181 366 1247 406
rect 487 322 553 338
rect 373 294 439 310
rect 271 158 301 291
rect 373 230 452 246
rect 373 196 389 230
rect 423 196 452 230
rect 373 180 452 196
rect 422 158 452 180
rect 500 158 530 322
rect 635 310 671 353
rect 889 326 925 353
rect 996 336 1247 366
rect 996 326 1026 336
rect 769 310 1026 326
rect 635 294 721 310
rect 635 274 671 294
rect 600 260 671 274
rect 705 260 721 294
rect 769 276 785 310
rect 819 296 1026 310
rect 819 276 835 296
rect 769 260 835 276
rect 600 244 721 260
rect 600 222 630 244
rect 798 222 828 260
rect 996 184 1026 296
rect 1289 288 1325 491
rect 1734 560 1764 586
rect 1818 560 1848 586
rect 1919 560 1949 586
rect 2009 560 2039 586
rect 1734 461 1764 476
rect 1818 461 1848 476
rect 1416 408 1446 423
rect 1626 408 1656 423
rect 1413 388 1449 408
rect 1623 391 1659 408
rect 1367 372 1471 388
rect 1367 338 1383 372
rect 1417 338 1471 372
rect 1367 322 1471 338
rect 1554 375 1659 391
rect 1554 341 1570 375
rect 1604 355 1659 375
rect 1604 341 1665 355
rect 1731 343 1767 461
rect 1554 325 1665 341
rect 1257 272 1325 288
rect 1132 256 1215 272
rect 1132 222 1165 256
rect 1199 222 1215 256
rect 1132 206 1215 222
rect 1257 238 1275 272
rect 1309 238 1325 272
rect 1257 222 1325 238
rect 1132 184 1162 206
rect 1257 184 1287 222
rect 1441 184 1471 322
rect 1527 261 1593 277
rect 1527 227 1543 261
rect 1577 227 1593 261
rect 1527 211 1593 227
rect 1635 229 1665 325
rect 1707 327 1773 343
rect 1707 293 1723 327
rect 1757 293 1773 327
rect 1707 277 1773 293
rect 1815 277 1851 461
rect 1919 377 1949 392
rect 2009 377 2039 392
rect 1916 360 1952 377
rect 1893 344 1959 360
rect 1893 310 1909 344
rect 1943 324 1959 344
rect 2006 324 2042 377
rect 2110 353 2140 368
rect 2200 353 2230 368
rect 2290 353 2320 368
rect 2380 353 2410 368
rect 1943 310 2042 324
rect 1893 294 2042 310
rect 1821 246 1851 277
rect 1821 230 1933 246
rect 1557 184 1587 211
rect 1635 199 1766 229
rect 1821 210 1883 230
rect 996 74 1026 100
rect 1132 74 1162 100
rect 1257 74 1287 100
rect 1736 158 1766 199
rect 1814 196 1883 210
rect 1917 196 1933 230
rect 2012 222 2042 294
rect 2107 326 2143 353
rect 2197 326 2233 353
rect 2287 326 2323 353
rect 2377 326 2413 353
rect 2107 310 2413 326
rect 2107 276 2123 310
rect 2157 276 2191 310
rect 2225 276 2259 310
rect 2293 276 2413 310
rect 2107 260 2413 276
rect 2107 222 2137 260
rect 2210 222 2240 260
rect 2296 222 2326 260
rect 2382 222 2412 260
rect 1814 180 1933 196
rect 1814 158 1844 180
rect 93 48 123 74
rect 193 48 223 74
rect 271 48 301 74
rect 422 48 452 74
rect 500 48 530 74
rect 600 48 630 74
rect 798 48 828 74
rect 1441 48 1471 74
rect 1557 48 1587 74
rect 1736 48 1766 74
rect 1814 48 1844 74
rect 2012 48 2042 74
rect 2107 48 2137 74
rect 2210 48 2240 74
rect 2296 48 2326 74
rect 2382 48 2412 74
<< polycont >>
rect 389 378 423 412
rect 133 321 167 355
rect 101 207 135 241
rect 281 307 315 341
rect 389 310 423 344
rect 503 338 537 372
rect 1031 424 1065 458
rect 1197 406 1231 440
rect 389 196 423 230
rect 671 260 705 294
rect 785 276 819 310
rect 1383 338 1417 372
rect 1570 341 1604 375
rect 1165 222 1199 256
rect 1275 238 1309 272
rect 1543 227 1577 261
rect 1723 293 1757 327
rect 1909 310 1943 344
rect 1883 196 1917 230
rect 2123 276 2157 310
rect 2191 276 2225 310
rect 2259 276 2293 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2496 683
rect 17 580 111 596
rect 17 546 61 580
rect 95 546 111 580
rect 17 510 111 546
rect 17 476 61 510
rect 95 476 111 510
rect 17 425 111 476
rect 145 580 211 649
rect 145 546 161 580
rect 195 546 211 580
rect 145 510 211 546
rect 145 476 161 510
rect 195 476 211 510
rect 145 460 211 476
rect 319 580 385 596
rect 319 546 335 580
rect 369 546 385 580
rect 517 580 641 649
rect 517 546 562 580
rect 596 546 641 580
rect 777 580 895 649
rect 1336 621 1402 649
rect 777 546 819 580
rect 853 546 895 580
rect 1031 568 1081 594
rect 319 512 385 546
rect 1031 542 1047 568
rect 929 534 1047 542
rect 929 512 1081 534
rect 319 478 335 512
rect 369 508 1081 512
rect 1115 565 1187 594
rect 1336 587 1352 621
rect 1386 587 1402 621
rect 1336 571 1402 587
rect 1115 531 1137 565
rect 1171 531 1187 565
rect 1654 548 1720 564
rect 369 478 963 508
rect 1115 502 1187 531
rect 1221 503 1620 537
rect 319 462 385 478
rect 373 425 439 428
rect 17 412 439 425
rect 17 391 389 412
rect 17 355 183 391
rect 373 378 389 391
rect 423 378 439 412
rect 17 321 133 355
rect 167 321 183 355
rect 17 305 183 321
rect 217 341 331 357
rect 217 307 281 341
rect 315 307 331 341
rect 17 157 51 305
rect 217 291 331 307
rect 373 344 439 378
rect 373 310 389 344
rect 423 310 439 344
rect 487 372 553 430
rect 487 338 503 372
rect 537 338 553 372
rect 487 310 553 338
rect 373 294 439 310
rect 587 270 621 478
rect 665 421 731 444
rect 665 387 681 421
rect 715 398 731 421
rect 715 387 833 398
rect 665 364 833 387
rect 771 310 833 364
rect 85 241 439 257
rect 85 207 101 241
rect 135 230 439 241
rect 135 207 389 230
rect 85 196 389 207
rect 423 196 439 230
rect 85 191 439 196
rect 313 162 439 191
rect 473 236 621 270
rect 655 294 737 310
rect 655 260 671 294
rect 705 260 737 294
rect 655 236 737 260
rect 771 276 785 310
rect 819 276 833 310
rect 867 330 901 478
rect 1015 458 1081 474
rect 1015 444 1031 458
rect 935 424 1031 444
rect 1065 424 1081 458
rect 935 421 1081 424
rect 969 408 1081 421
rect 969 387 985 408
rect 935 364 985 387
rect 867 296 985 330
rect 771 260 833 276
rect 17 130 98 157
rect 17 96 48 130
rect 82 96 98 130
rect 17 70 98 96
rect 132 130 198 157
rect 132 96 148 130
rect 182 96 198 130
rect 473 128 507 236
rect 771 202 805 260
rect 625 168 641 202
rect 675 168 805 202
rect 839 210 889 226
rect 873 176 889 210
rect 132 17 198 96
rect 296 94 344 128
rect 378 94 507 128
rect 296 78 507 94
rect 541 133 591 162
rect 575 99 591 133
rect 541 17 591 99
rect 625 120 691 168
rect 625 86 641 120
rect 675 86 691 120
rect 625 70 691 86
rect 737 127 803 134
rect 737 93 753 127
rect 787 93 803 127
rect 737 17 803 93
rect 839 120 889 176
rect 873 86 889 120
rect 935 170 985 296
rect 935 136 951 170
rect 935 119 985 136
rect 839 85 889 86
rect 1019 85 1053 408
rect 1115 356 1149 502
rect 1221 456 1255 503
rect 1183 440 1255 456
rect 1183 406 1197 440
rect 1231 406 1255 440
rect 1443 435 1480 469
rect 1514 435 1552 469
rect 1183 390 1255 406
rect 1367 372 1432 388
rect 1367 356 1383 372
rect 1087 338 1383 356
rect 1417 338 1432 372
rect 1087 322 1432 338
rect 1087 170 1121 322
rect 1466 288 1500 435
rect 1586 391 1620 503
rect 1654 514 1670 548
rect 1704 514 1720 548
rect 1654 469 1720 514
rect 1845 535 1911 649
rect 1845 501 1861 535
rect 1895 501 1911 535
rect 1845 472 1911 501
rect 1946 548 2027 564
rect 1946 514 1962 548
rect 1996 514 2027 548
rect 1654 435 1670 469
rect 1704 438 1720 469
rect 1946 444 2027 514
rect 1704 435 1837 438
rect 1654 404 1837 435
rect 1554 375 1620 391
rect 1554 341 1570 375
rect 1604 341 1620 375
rect 1803 360 1837 404
rect 1946 410 1962 444
rect 1996 410 2027 444
rect 1946 394 2027 410
rect 1803 344 1959 360
rect 1554 325 1620 341
rect 1707 327 1769 343
rect 1259 272 1500 288
rect 1707 293 1723 327
rect 1757 293 1769 327
rect 1707 282 1769 293
rect 1087 119 1121 136
rect 1155 256 1215 272
rect 1155 222 1165 256
rect 1199 222 1215 256
rect 1259 238 1275 272
rect 1309 238 1500 272
rect 1259 222 1500 238
rect 1155 188 1215 222
rect 1155 154 1432 188
rect 1155 85 1189 154
rect 839 51 1189 85
rect 1298 86 1314 120
rect 1348 86 1364 120
rect 1298 17 1364 86
rect 1398 93 1432 154
rect 1466 177 1500 222
rect 1534 261 1769 282
rect 1534 227 1543 261
rect 1577 248 1769 261
rect 1803 310 1909 344
rect 1943 310 1959 344
rect 1803 294 1959 310
rect 1993 326 2027 394
rect 2061 548 2095 649
rect 2061 438 2095 514
rect 2061 388 2095 404
rect 2137 580 2203 596
rect 2137 546 2153 580
rect 2187 546 2203 580
rect 2137 497 2203 546
rect 2137 463 2153 497
rect 2187 463 2203 497
rect 2137 414 2203 463
rect 2243 580 2293 649
rect 2277 546 2293 580
rect 2243 478 2293 546
rect 2277 444 2293 478
rect 2243 428 2293 444
rect 2333 580 2371 596
rect 2367 546 2371 580
rect 2333 497 2371 546
rect 2367 463 2371 497
rect 2137 380 2153 414
rect 2187 394 2203 414
rect 2333 414 2371 463
rect 2407 580 2473 649
rect 2407 546 2423 580
rect 2457 546 2473 580
rect 2407 471 2473 546
rect 2407 437 2423 471
rect 2457 437 2473 471
rect 2187 380 2333 394
rect 2367 403 2371 414
rect 2367 380 2471 403
rect 2137 360 2471 380
rect 1993 310 2309 326
rect 1577 227 1625 248
rect 1534 211 1625 227
rect 1803 214 1837 294
rect 1993 276 2123 310
rect 2157 276 2191 310
rect 2225 276 2259 310
rect 2293 276 2309 310
rect 1993 260 2309 276
rect 1466 161 1557 177
rect 1466 127 1494 161
rect 1528 127 1557 161
rect 1591 93 1625 211
rect 1398 59 1625 93
rect 1659 180 1837 214
rect 1871 230 2027 260
rect 1871 196 1883 230
rect 1917 226 2027 230
rect 2352 226 2471 360
rect 1917 196 1933 226
rect 1871 180 1933 196
rect 1967 210 2001 226
rect 1659 140 1725 180
rect 2149 210 2471 226
rect 1659 106 1675 140
rect 1709 106 1725 140
rect 1659 70 1725 106
rect 1839 125 1905 146
rect 1839 91 1855 125
rect 1889 91 1905 125
rect 1839 17 1905 91
rect 1967 120 2001 176
rect 1967 70 2001 86
rect 2037 158 2053 192
rect 2087 158 2103 192
rect 2037 116 2103 158
rect 2037 82 2053 116
rect 2087 82 2103 116
rect 2037 17 2103 82
rect 2149 176 2165 210
rect 2199 176 2337 210
rect 2371 176 2471 210
rect 2149 120 2199 176
rect 2149 86 2165 120
rect 2149 70 2199 86
rect 2235 123 2301 142
rect 2235 89 2251 123
rect 2285 89 2301 123
rect 2235 17 2301 89
rect 2335 120 2373 176
rect 2335 86 2337 120
rect 2371 86 2373 120
rect 2335 70 2373 86
rect 2407 131 2473 142
rect 2407 97 2423 131
rect 2457 97 2473 131
rect 2407 17 2473 97
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2496 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
<< metal1 >>
rect 0 683 2496 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2496 683
rect 0 617 2496 649
rect 0 17 2496 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2496 17
rect 0 -49 2496 -17
<< labels >>
rlabel comment s 0 0 0 0 4 sdfxtp_4
flabel comment s 1000 314 1000 314 0 FreeSans 200 0 0 0 no_jumper_check
flabel pwell s 0 0 2496 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nwell s 0 617 2496 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 2496 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 2496 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 319 168 353 202 0 FreeSans 340 0 0 0 SCE
port 4 nsew
flabel corelocali s 703 242 737 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 SCD
port 3 nsew
flabel corelocali s 511 390 545 424 0 FreeSans 340 0 0 0 SCD
port 3 nsew
flabel corelocali s 2431 242 2465 276 0 FreeSans 340 0 0 0 Q
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 2496 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 331718
string GDS_START 314256
<< end >>
