magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 736 561
rect 122 265 156 492
rect 191 343 241 527
rect 511 369 577 527
rect 651 432 719 493
rect 122 199 225 265
rect 300 199 381 323
rect 653 299 719 432
rect 483 153 551 265
rect 674 165 719 299
rect 175 17 241 97
rect 509 17 576 94
rect 651 51 719 165
rect 0 -17 736 17
<< obsli1 >>
rect 27 165 79 425
rect 331 363 449 416
rect 415 333 449 363
rect 415 299 619 333
rect 415 165 449 299
rect 585 265 619 299
rect 27 131 449 165
rect 585 199 640 265
rect 27 51 79 131
rect 331 128 449 131
rect 331 51 397 128
<< metal1 >>
rect 0 496 736 592
rect 0 -48 736 48
<< labels >>
rlabel locali s 122 265 156 492 6 A
port 1 nsew signal input
rlabel locali s 122 199 225 265 6 A
port 1 nsew signal input
rlabel locali s 300 199 381 323 6 B
port 2 nsew signal input
rlabel locali s 483 153 551 265 6 C
port 3 nsew signal input
rlabel locali s 674 165 719 299 6 X
port 4 nsew signal output
rlabel locali s 653 299 719 432 6 X
port 4 nsew signal output
rlabel locali s 651 432 719 493 6 X
port 4 nsew signal output
rlabel locali s 651 51 719 165 6 X
port 4 nsew signal output
rlabel locali s 509 17 576 94 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 175 17 241 97 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 736 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 736 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 511 369 577 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 191 343 241 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 736 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 736 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1622170
string GDS_START 1616046
<< end >>
