magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 2392 561
rect 35 289 69 527
rect 307 357 341 527
rect 475 357 509 527
rect 643 367 677 527
rect 811 367 845 527
rect 979 367 1013 527
rect 1047 323 1113 493
rect 1147 367 1181 527
rect 1215 323 1281 493
rect 1315 367 1349 527
rect 1383 323 1449 493
rect 1483 367 1517 527
rect 1551 323 1617 493
rect 1651 367 1685 527
rect 1719 323 1785 493
rect 1819 367 1853 527
rect 1887 323 1953 493
rect 1987 367 2021 527
rect 2055 323 2121 493
rect 2155 367 2189 527
rect 2223 323 2289 493
rect 2323 367 2357 527
rect 1047 289 2375 323
rect 22 215 88 255
rect 2324 181 2375 289
rect 35 17 69 181
rect 1047 147 2375 181
rect 307 17 341 113
rect 475 17 509 113
rect 643 17 677 113
rect 811 17 845 113
rect 979 17 1013 113
rect 1047 52 1113 147
rect 1047 51 1097 52
rect 1147 17 1181 113
rect 1215 52 1281 147
rect 1231 51 1265 52
rect 1315 17 1349 113
rect 1383 52 1449 147
rect 1399 51 1433 52
rect 1483 17 1517 113
rect 1551 52 1617 147
rect 1651 17 1685 113
rect 1719 52 1785 147
rect 1819 17 1853 113
rect 1887 52 1953 147
rect 1987 17 2021 113
rect 2055 52 2121 147
rect 2155 17 2189 113
rect 2223 52 2289 147
rect 2323 17 2357 113
rect 0 -17 2392 17
<< obsli1 >>
rect 103 289 169 493
rect 207 323 273 493
rect 375 323 441 493
rect 543 323 609 493
rect 711 323 777 493
rect 879 323 945 493
rect 207 289 509 323
rect 543 289 1013 323
rect 122 255 169 289
rect 475 255 509 289
rect 978 255 1013 289
rect 122 215 441 255
rect 475 215 937 255
rect 978 215 2290 255
rect 122 181 169 215
rect 475 181 509 215
rect 978 181 1013 215
rect 103 52 169 181
rect 207 147 509 181
rect 543 147 1013 181
rect 207 52 273 147
rect 375 52 441 147
rect 543 52 609 147
rect 711 52 777 147
rect 879 52 945 147
<< metal1 >>
rect 0 496 2392 592
rect 0 -48 2392 48
<< labels >>
rlabel locali s 22 215 88 255 6 A
port 1 nsew signal input
rlabel locali s 2324 181 2375 289 6 X
port 2 nsew signal output
rlabel locali s 2223 323 2289 493 6 X
port 2 nsew signal output
rlabel locali s 2223 52 2289 147 6 X
port 2 nsew signal output
rlabel locali s 2055 323 2121 493 6 X
port 2 nsew signal output
rlabel locali s 2055 52 2121 147 6 X
port 2 nsew signal output
rlabel locali s 1887 323 1953 493 6 X
port 2 nsew signal output
rlabel locali s 1887 52 1953 147 6 X
port 2 nsew signal output
rlabel locali s 1719 323 1785 493 6 X
port 2 nsew signal output
rlabel locali s 1719 52 1785 147 6 X
port 2 nsew signal output
rlabel locali s 1551 323 1617 493 6 X
port 2 nsew signal output
rlabel locali s 1551 52 1617 147 6 X
port 2 nsew signal output
rlabel locali s 1399 51 1433 52 6 X
port 2 nsew signal output
rlabel locali s 1383 323 1449 493 6 X
port 2 nsew signal output
rlabel locali s 1383 52 1449 147 6 X
port 2 nsew signal output
rlabel locali s 1231 51 1265 52 6 X
port 2 nsew signal output
rlabel locali s 1215 323 1281 493 6 X
port 2 nsew signal output
rlabel locali s 1215 52 1281 147 6 X
port 2 nsew signal output
rlabel locali s 1047 323 1113 493 6 X
port 2 nsew signal output
rlabel locali s 1047 289 2375 323 6 X
port 2 nsew signal output
rlabel locali s 1047 147 2375 181 6 X
port 2 nsew signal output
rlabel locali s 1047 52 1113 147 6 X
port 2 nsew signal output
rlabel locali s 1047 51 1097 52 6 X
port 2 nsew signal output
rlabel locali s 2323 17 2357 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 2155 17 2189 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1987 17 2021 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1819 17 1853 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1651 17 1685 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1483 17 1517 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1315 17 1349 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1147 17 1181 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 979 17 1013 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 811 17 845 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 643 17 677 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 475 17 509 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 307 17 341 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 35 17 69 181 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 0 -17 2392 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 2392 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 2323 367 2357 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 2155 367 2189 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1987 367 2021 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1819 367 1853 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1651 367 1685 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1483 367 1517 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1315 367 1349 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1147 367 1181 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 979 367 1013 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 811 367 845 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 643 367 677 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 475 357 509 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 307 357 341 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 35 289 69 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 0 527 2392 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 496 2392 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2392 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3075520
string GDS_START 3057318
<< end >>
