magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1932 561
rect 17 357 89 527
rect 194 373 261 527
rect 17 199 86 323
rect 17 17 89 165
rect 194 265 261 339
rect 483 447 549 527
rect 651 447 717 527
rect 819 447 885 527
rect 987 447 1053 527
rect 194 199 286 265
rect 399 289 1915 345
rect 194 124 261 199
rect 1865 171 1915 289
rect 194 17 261 89
rect 531 17 597 97
rect 699 17 765 97
rect 867 17 933 97
rect 1035 17 1101 97
rect 1255 123 1915 171
rect 0 -17 1932 17
<< obsli1 >>
rect 123 323 160 493
rect 120 255 160 323
rect 120 221 121 255
rect 155 221 160 255
rect 120 199 160 221
rect 123 56 160 199
rect 295 299 365 493
rect 399 413 449 493
rect 583 413 617 493
rect 751 413 785 493
rect 919 413 953 493
rect 1087 413 1915 493
rect 399 379 1915 413
rect 320 255 365 299
rect 320 205 1185 255
rect 1235 221 1316 255
rect 1350 221 1831 255
rect 1235 205 1831 221
rect 320 165 397 205
rect 295 51 397 165
rect 431 131 1221 171
rect 431 51 497 131
rect 631 55 665 131
rect 799 51 833 131
rect 967 55 1001 131
rect 1135 89 1221 131
rect 1135 51 1915 89
<< obsli1c >>
rect 121 221 155 255
rect 1316 221 1350 255
<< metal1 >>
rect 0 496 1932 592
rect 0 -48 1932 48
<< obsm1 >>
rect 109 255 167 261
rect 109 221 121 255
rect 155 252 167 255
rect 1304 255 1362 261
rect 1304 252 1316 255
rect 155 224 1316 252
rect 155 221 167 224
rect 109 215 167 221
rect 1304 221 1316 224
rect 1350 221 1362 255
rect 1304 215 1362 221
<< labels >>
rlabel locali s 17 199 86 323 6 A
port 1 nsew signal input
rlabel locali s 194 265 261 339 6 TE_B
port 2 nsew signal input
rlabel locali s 194 199 286 265 6 TE_B
port 2 nsew signal input
rlabel locali s 194 124 261 199 6 TE_B
port 2 nsew signal input
rlabel locali s 1865 171 1915 289 6 Z
port 3 nsew signal output
rlabel locali s 1255 123 1915 171 6 Z
port 3 nsew signal output
rlabel locali s 399 289 1915 345 6 Z
port 3 nsew signal output
rlabel locali s 1035 17 1101 97 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 867 17 933 97 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 699 17 765 97 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 531 17 597 97 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 194 17 261 89 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 17 17 89 165 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 1932 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1932 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 987 447 1053 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 819 447 885 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 651 447 717 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 483 447 549 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 194 373 261 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 17 357 89 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 1932 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 1932 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1932 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2884376
string GDS_START 2870464
<< end >>
