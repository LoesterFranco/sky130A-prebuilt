magic
tech sky130A
magscale 1 2
timestamp 1599588232
<< locali >>
rect 25 270 286 356
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2400 683
rect 24 424 90 596
rect 130 458 164 649
rect 204 424 270 596
rect 310 458 344 649
rect 24 390 354 424
rect 320 326 354 390
rect 388 394 454 596
rect 494 428 528 649
rect 568 394 634 596
rect 674 428 708 649
rect 748 394 814 596
rect 388 360 814 394
rect 854 384 888 649
rect 928 424 994 596
rect 928 404 946 424
rect 923 390 946 404
rect 980 390 994 424
rect 923 384 994 390
rect 1034 384 1068 649
rect 1108 424 1174 596
rect 1108 404 1124 424
rect 1102 390 1124 404
rect 1158 390 1174 424
rect 1102 384 1174 390
rect 1214 384 1248 649
rect 1288 424 1354 596
rect 1288 404 1304 424
rect 1284 390 1304 404
rect 1338 390 1354 424
rect 1284 384 1354 390
rect 1394 384 1428 649
rect 1468 424 1534 596
rect 1468 390 1484 424
rect 1518 390 1534 424
rect 1468 384 1534 390
rect 1574 384 1608 649
rect 1648 424 1714 596
rect 1648 404 1664 424
rect 1653 390 1664 404
rect 1698 390 1714 424
rect 1653 384 1714 390
rect 1754 384 1799 649
rect 1838 424 1904 596
rect 1838 404 1854 424
rect 1839 390 1854 404
rect 1888 390 1904 424
rect 1839 384 1904 390
rect 1944 384 1991 649
rect 2028 424 2094 596
rect 2028 404 2044 424
rect 2025 390 2044 404
rect 2078 390 2094 424
rect 2025 384 2094 390
rect 2134 384 2177 649
rect 2218 424 2284 596
rect 2218 404 2234 424
rect 2211 390 2234 404
rect 2268 390 2284 424
rect 748 350 814 360
rect 320 260 692 326
rect 748 316 845 350
rect 879 316 887 350
rect 748 260 887 316
rect 320 236 354 260
rect 23 202 354 236
rect 737 226 787 260
rect 23 70 73 202
rect 109 17 175 168
rect 223 70 257 202
rect 395 192 787 226
rect 293 17 359 168
rect 395 70 429 192
rect 465 17 515 158
rect 551 70 601 192
rect 637 17 703 158
rect 737 70 787 192
rect 823 17 889 226
rect 923 70 973 384
rect 1007 316 1018 350
rect 1052 316 1061 350
rect 1007 260 1061 316
rect 1009 17 1059 221
rect 1102 70 1145 384
rect 1180 316 1196 350
rect 1230 316 1246 350
rect 1180 260 1246 316
rect 1181 17 1247 221
rect 1284 70 1331 384
rect 1368 316 1384 350
rect 1418 316 1434 350
rect 1368 260 1434 316
rect 1367 17 1433 221
rect 1468 70 1517 384
rect 1552 316 1567 350
rect 1601 316 1618 350
rect 1552 260 1618 316
rect 1553 17 1619 221
rect 1653 70 1703 384
rect 1737 316 1753 350
rect 1787 316 1803 350
rect 1737 260 1803 316
rect 1739 17 1805 221
rect 1839 70 1889 384
rect 1923 316 1938 350
rect 1972 316 1989 350
rect 1923 260 1989 316
rect 1925 17 1991 221
rect 2025 70 2075 384
rect 2211 358 2284 390
rect 2324 364 2374 649
rect 2109 316 2125 350
rect 2159 316 2175 350
rect 2109 260 2175 316
rect 2111 17 2177 221
rect 2211 70 2277 358
rect 2311 17 2377 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2400 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 946 390 980 424
rect 1124 390 1158 424
rect 1304 390 1338 424
rect 1484 390 1518 424
rect 1664 390 1698 424
rect 1854 390 1888 424
rect 2044 390 2078 424
rect 2234 390 2268 424
rect 845 316 879 350
rect 1018 316 1052 350
rect 1196 316 1230 350
rect 1384 316 1418 350
rect 1567 316 1601 350
rect 1753 316 1787 350
rect 1938 316 1972 350
rect 2125 316 2159 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
<< metal1 >>
rect 0 683 2400 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2400 683
rect 0 617 2400 649
rect 0 616 50 617
rect 932 424 2280 430
rect 932 390 946 424
rect 980 390 1124 424
rect 1158 390 1304 424
rect 1338 390 1484 424
rect 1518 390 1664 424
rect 1698 390 1854 424
rect 1888 390 2044 424
rect 2078 390 2234 424
rect 2268 390 2280 424
rect 932 384 2280 390
rect 0 49 50 50
rect 0 17 2400 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2400 17
rect 0 -49 2400 -17
<< obsm1 >>
rect 831 350 2171 356
rect 831 316 845 350
rect 879 316 1018 350
rect 1052 316 1196 350
rect 1230 316 1384 350
rect 1418 316 1567 350
rect 1601 316 1753 350
rect 1787 316 1938 350
rect 1972 316 2125 350
rect 2159 316 2171 350
rect 831 310 2171 316
<< labels >>
rlabel locali s 25 270 286 356 6 A
port 1 nsew signal input
rlabel metal1 s 932 384 2280 430 6 Y
port 2 nsew signal output
rlabel metal1 s 0 -49 2400 49 8 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 4 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 617 2400 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2400 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3469900
string GDS_START 3449780
<< end >>
