magic
tech sky130A
magscale 1 2
timestamp 1604502741
<< locali >>
rect 87 252 167 386
rect 201 338 267 430
rect 1153 364 1226 596
rect 1192 220 1226 364
rect 1158 70 1226 220
rect 1543 70 1610 596
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 19 420 109 596
rect 147 464 213 649
rect 247 512 313 596
rect 476 546 542 649
rect 247 478 829 512
rect 247 464 335 478
rect 19 218 53 420
rect 301 304 335 464
rect 369 376 582 444
rect 652 410 761 444
rect 415 342 668 376
rect 227 252 381 304
rect 19 150 89 218
rect 227 184 293 252
rect 415 218 449 342
rect 339 184 449 218
rect 507 150 573 302
rect 19 116 573 150
rect 607 294 668 342
rect 607 101 641 294
rect 702 260 736 410
rect 795 360 829 478
rect 896 412 1004 649
rect 1044 378 1112 580
rect 770 294 829 360
rect 863 344 1112 378
rect 1260 420 1310 649
rect 863 294 929 344
rect 1078 320 1112 344
rect 978 260 1044 310
rect 702 226 1044 260
rect 1078 254 1158 320
rect 702 211 827 226
rect 675 145 827 211
rect 1078 192 1112 254
rect 1344 326 1413 596
rect 1453 364 1503 649
rect 1344 260 1500 326
rect 125 17 191 82
rect 468 17 535 82
rect 607 51 852 101
rect 941 17 1007 192
rect 1041 70 1112 192
rect 1260 17 1310 226
rect 1344 108 1412 260
rect 1458 17 1508 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
rlabel locali s 87 252 167 386 6 D
port 1 nsew signal input
rlabel locali s 1192 220 1226 364 6 Q
port 2 nsew signal output
rlabel locali s 1158 70 1226 220 6 Q
port 2 nsew signal output
rlabel locali s 1153 364 1226 596 6 Q
port 2 nsew signal output
rlabel locali s 1543 70 1610 596 6 Q_N
port 3 nsew signal output
rlabel locali s 201 338 267 430 6 GATE_N
port 4 nsew clock input
rlabel metal1 s 0 -49 1632 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 617 1632 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 2143298
string GDS_START 2130664
<< end >>
