magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 18 425 379 483
rect 18 151 88 265
rect 132 199 271 323
rect 561 299 615 493
rect 305 199 419 265
rect 581 152 615 299
rect 561 83 615 152
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 18 357 366 391
rect 423 367 479 527
rect 18 299 82 357
rect 332 333 366 357
rect 332 299 487 333
rect 453 265 487 299
rect 453 199 511 265
rect 453 165 487 199
rect 135 131 487 165
rect 19 17 85 117
rect 135 61 169 131
rect 209 17 285 97
rect 329 61 363 131
rect 397 17 483 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 305 199 419 265 6 A
port 1 nsew signal input
rlabel locali s 18 425 379 483 6 B
port 2 nsew signal input
rlabel locali s 132 199 271 323 6 C
port 3 nsew signal input
rlabel locali s 18 151 88 265 6 D
port 4 nsew signal input
rlabel locali s 581 152 615 299 6 X
port 5 nsew signal output
rlabel locali s 561 299 615 493 6 X
port 5 nsew signal output
rlabel locali s 561 83 615 152 6 X
port 5 nsew signal output
rlabel metal1 s 0 -48 644 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 498236
string GDS_START 491974
<< end >>
