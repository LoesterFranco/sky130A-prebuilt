magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 552 561
rect 17 206 73 493
rect 107 372 249 527
rect 17 51 85 206
rect 213 215 307 261
rect 388 255 431 478
rect 467 383 533 527
rect 489 255 535 323
rect 341 219 431 255
rect 341 215 407 219
rect 469 215 535 255
rect 119 17 153 109
rect 399 17 433 109
rect 0 -17 552 17
<< obsli1 >>
rect 283 338 349 493
rect 119 295 349 338
rect 119 181 176 295
rect 119 143 261 181
rect 201 115 261 143
rect 299 143 535 181
rect 299 127 365 143
rect 201 113 264 115
rect 201 111 266 113
rect 201 110 268 111
rect 201 108 269 110
rect 201 107 270 108
rect 201 105 271 107
rect 201 104 272 105
rect 201 51 273 104
rect 467 51 535 143
<< metal1 >>
rect 0 496 552 592
rect 0 -48 552 48
<< labels >>
rlabel locali s 489 255 535 323 6 A1
port 1 nsew signal input
rlabel locali s 469 215 535 255 6 A1
port 1 nsew signal input
rlabel locali s 388 255 431 478 6 A2
port 2 nsew signal input
rlabel locali s 341 219 431 255 6 A2
port 2 nsew signal input
rlabel locali s 341 215 407 219 6 A2
port 2 nsew signal input
rlabel locali s 213 215 307 261 6 B1
port 3 nsew signal input
rlabel locali s 17 206 73 493 6 X
port 4 nsew signal output
rlabel locali s 17 51 85 206 6 X
port 4 nsew signal output
rlabel locali s 399 17 433 109 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 119 17 153 109 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 552 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 552 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 467 383 533 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 107 372 249 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 552 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 552 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 552 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1297996
string GDS_START 1292424
<< end >>
