magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 667 323 743 493
rect 855 323 931 493
rect 1043 323 1119 493
rect 1231 323 1307 493
rect 1419 323 1495 493
rect 1607 323 1683 493
rect 1795 323 1871 493
rect 1983 323 2059 493
rect 2172 323 2227 472
rect 667 289 2227 323
rect 17 215 547 255
rect 2127 181 2227 289
rect 667 147 2227 181
rect 667 52 743 147
rect 667 51 727 52
rect 855 52 931 147
rect 881 51 915 52
rect 1043 52 1119 147
rect 1069 51 1103 52
rect 1231 52 1307 147
rect 1419 52 1495 147
rect 1607 52 1683 147
rect 1795 52 1871 147
rect 1983 52 2059 147
rect 2172 73 2227 147
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2300 561
rect 35 289 69 527
rect 103 323 179 493
rect 223 367 257 527
rect 291 323 367 493
rect 411 367 445 527
rect 479 323 555 493
rect 599 367 633 527
rect 787 367 821 527
rect 975 367 1009 527
rect 1163 367 1197 527
rect 1351 367 1385 527
rect 1539 367 1573 527
rect 1727 367 1761 527
rect 1915 367 1949 527
rect 2103 367 2137 527
rect 103 289 633 323
rect 598 255 633 289
rect 598 215 2035 255
rect 598 181 633 215
rect 35 17 69 181
rect 103 147 633 181
rect 103 52 179 147
rect 223 17 257 113
rect 291 52 367 147
rect 411 17 445 113
rect 479 52 555 147
rect 599 17 633 113
rect 787 17 821 113
rect 975 17 1009 113
rect 1163 17 1197 113
rect 1351 17 1385 113
rect 1539 17 1573 113
rect 1727 17 1761 113
rect 1915 17 1949 113
rect 2103 17 2137 113
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2300 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
<< metal1 >>
rect 0 561 2300 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2300 561
rect 0 496 2300 527
rect 0 17 2300 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2300 17
rect 0 -48 2300 -17
<< labels >>
rlabel locali s 17 215 547 255 6 A
port 1 nsew signal input
rlabel locali s 2172 323 2227 472 6 X
port 2 nsew signal output
rlabel locali s 2172 73 2227 147 6 X
port 2 nsew signal output
rlabel locali s 2127 181 2227 289 6 X
port 2 nsew signal output
rlabel locali s 1983 323 2059 493 6 X
port 2 nsew signal output
rlabel locali s 1983 52 2059 147 6 X
port 2 nsew signal output
rlabel locali s 1795 323 1871 493 6 X
port 2 nsew signal output
rlabel locali s 1795 52 1871 147 6 X
port 2 nsew signal output
rlabel locali s 1607 323 1683 493 6 X
port 2 nsew signal output
rlabel locali s 1607 52 1683 147 6 X
port 2 nsew signal output
rlabel locali s 1419 323 1495 493 6 X
port 2 nsew signal output
rlabel locali s 1419 52 1495 147 6 X
port 2 nsew signal output
rlabel locali s 1231 323 1307 493 6 X
port 2 nsew signal output
rlabel locali s 1231 52 1307 147 6 X
port 2 nsew signal output
rlabel locali s 1069 51 1103 52 6 X
port 2 nsew signal output
rlabel locali s 1043 323 1119 493 6 X
port 2 nsew signal output
rlabel locali s 1043 52 1119 147 6 X
port 2 nsew signal output
rlabel locali s 881 51 915 52 6 X
port 2 nsew signal output
rlabel locali s 855 323 931 493 6 X
port 2 nsew signal output
rlabel locali s 855 52 931 147 6 X
port 2 nsew signal output
rlabel locali s 667 323 743 493 6 X
port 2 nsew signal output
rlabel locali s 667 289 2227 323 6 X
port 2 nsew signal output
rlabel locali s 667 147 2227 181 6 X
port 2 nsew signal output
rlabel locali s 667 52 743 147 6 X
port 2 nsew signal output
rlabel locali s 667 51 727 52 6 X
port 2 nsew signal output
rlabel metal1 s 0 -48 2300 48 8 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 496 2300 592 6 VPWR
port 4 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2300 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1656102
string GDS_START 1639570
<< end >>
