magic
tech sky130A
magscale 1 2
timestamp 1604502710
<< nwell >>
rect -38 332 902 704
<< pwell >>
rect 0 0 864 49
<< scpmos >>
rect 122 368 158 592
rect 225 392 261 592
rect 303 392 339 592
rect 497 392 533 592
rect 587 392 623 592
rect 683 392 719 592
<< nmoslvt >>
rect 129 88 159 236
rect 227 126 257 236
rect 313 126 343 236
rect 489 126 519 254
rect 575 126 605 254
rect 683 126 713 254
<< ndiff >>
rect 439 236 489 254
rect 76 214 129 236
rect 76 180 84 214
rect 118 180 129 214
rect 76 134 129 180
rect 76 100 84 134
rect 118 100 129 134
rect 76 88 129 100
rect 159 202 227 236
rect 159 168 170 202
rect 204 168 227 202
rect 159 134 227 168
rect 159 100 170 134
rect 204 126 227 134
rect 257 186 313 236
rect 257 152 268 186
rect 302 152 313 186
rect 257 126 313 152
rect 343 172 489 236
rect 343 138 368 172
rect 402 138 444 172
rect 478 138 489 172
rect 343 126 489 138
rect 519 241 575 254
rect 519 207 530 241
rect 564 207 575 241
rect 519 126 575 207
rect 605 126 683 254
rect 713 230 766 254
rect 713 196 724 230
rect 758 196 766 230
rect 713 126 766 196
rect 204 100 212 126
rect 159 88 212 100
<< pdiff >>
rect 70 580 122 592
rect 70 546 78 580
rect 112 546 122 580
rect 70 497 122 546
rect 70 463 78 497
rect 112 463 122 497
rect 70 414 122 463
rect 70 380 78 414
rect 112 380 122 414
rect 70 368 122 380
rect 158 580 225 592
rect 158 546 168 580
rect 202 546 225 580
rect 158 470 225 546
rect 158 436 168 470
rect 202 436 225 470
rect 158 392 225 436
rect 261 392 303 592
rect 339 547 391 592
rect 339 513 349 547
rect 383 513 391 547
rect 339 460 391 513
rect 339 426 349 460
rect 383 426 391 460
rect 339 392 391 426
rect 445 544 497 592
rect 445 510 453 544
rect 487 510 497 544
rect 445 392 497 510
rect 533 580 587 592
rect 533 546 543 580
rect 577 546 587 580
rect 533 510 587 546
rect 533 476 543 510
rect 577 476 587 510
rect 533 440 587 476
rect 533 406 543 440
rect 577 406 587 440
rect 533 392 587 406
rect 623 580 683 592
rect 623 546 636 580
rect 670 546 683 580
rect 623 508 683 546
rect 623 474 636 508
rect 670 474 683 508
rect 623 392 683 474
rect 719 580 771 592
rect 719 546 729 580
rect 763 546 771 580
rect 719 509 771 546
rect 719 475 729 509
rect 763 475 771 509
rect 719 438 771 475
rect 719 404 729 438
rect 763 404 771 438
rect 719 392 771 404
rect 158 368 210 392
<< ndiffc >>
rect 84 180 118 214
rect 84 100 118 134
rect 170 168 204 202
rect 170 100 204 134
rect 268 152 302 186
rect 368 138 402 172
rect 444 138 478 172
rect 530 207 564 241
rect 724 196 758 230
<< pdiffc >>
rect 78 546 112 580
rect 78 463 112 497
rect 78 380 112 414
rect 168 546 202 580
rect 168 436 202 470
rect 349 513 383 547
rect 349 426 383 460
rect 453 510 487 544
rect 543 546 577 580
rect 543 476 577 510
rect 543 406 577 440
rect 636 546 670 580
rect 636 474 670 508
rect 729 546 763 580
rect 729 475 763 509
rect 729 404 763 438
<< poly >>
rect 122 592 158 618
rect 225 592 261 618
rect 303 592 339 618
rect 497 592 533 618
rect 587 592 623 618
rect 683 592 719 618
rect 122 330 158 368
rect 93 314 159 330
rect 225 324 261 392
rect 303 346 339 392
rect 497 356 533 392
rect 587 356 623 392
rect 309 324 339 346
rect 467 340 533 356
rect 93 280 109 314
rect 143 280 159 314
rect 93 264 159 280
rect 129 236 159 264
rect 201 308 267 324
rect 201 274 217 308
rect 251 274 267 308
rect 201 258 267 274
rect 309 308 375 324
rect 309 274 325 308
rect 359 274 375 308
rect 467 306 483 340
rect 517 306 533 340
rect 467 290 533 306
rect 575 340 641 356
rect 575 306 591 340
rect 625 306 641 340
rect 575 290 641 306
rect 309 258 375 274
rect 227 236 257 258
rect 313 236 343 258
rect 489 254 519 290
rect 575 254 605 290
rect 683 269 719 392
rect 683 254 713 269
rect 227 100 257 126
rect 313 100 343 126
rect 489 104 519 126
rect 453 88 519 104
rect 575 100 605 126
rect 683 104 713 126
rect 129 62 159 88
rect 453 54 469 88
rect 503 54 519 88
rect 453 38 519 54
rect 683 88 763 104
rect 683 54 713 88
rect 747 54 763 88
rect 683 38 763 54
<< polycont >>
rect 109 280 143 314
rect 217 274 251 308
rect 325 274 359 308
rect 483 306 517 340
rect 591 306 625 340
rect 469 54 503 88
rect 713 54 747 88
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 25 580 112 596
rect 25 546 78 580
rect 25 497 112 546
rect 25 463 78 497
rect 25 414 112 463
rect 152 580 218 649
rect 152 546 168 580
rect 202 546 218 580
rect 152 470 218 546
rect 152 436 168 470
rect 202 436 218 470
rect 152 426 218 436
rect 265 581 503 615
rect 25 380 78 414
rect 265 392 299 581
rect 333 513 349 547
rect 383 513 399 547
rect 333 460 399 513
rect 437 544 503 581
rect 437 510 453 544
rect 487 510 503 544
rect 437 494 503 510
rect 543 580 577 596
rect 543 510 577 546
rect 333 426 349 460
rect 383 426 506 460
rect 25 364 112 380
rect 25 230 59 364
rect 146 358 438 392
rect 146 330 180 358
rect 93 314 180 330
rect 93 280 109 314
rect 143 280 180 314
rect 93 264 180 280
rect 214 308 267 324
rect 214 274 217 308
rect 251 274 267 308
rect 214 236 267 274
rect 309 308 370 324
rect 309 274 325 308
rect 359 274 370 308
rect 309 236 370 274
rect 404 242 438 358
rect 472 356 506 426
rect 543 440 577 476
rect 617 580 689 649
rect 617 546 636 580
rect 670 546 689 580
rect 617 508 689 546
rect 617 474 636 508
rect 670 474 689 508
rect 617 458 689 474
rect 729 580 779 596
rect 763 546 779 580
rect 729 509 779 546
rect 763 475 779 509
rect 729 438 779 475
rect 577 406 729 424
rect 543 404 729 406
rect 763 404 779 438
rect 543 390 779 404
rect 729 388 779 390
rect 472 340 533 356
rect 472 306 483 340
rect 517 306 533 340
rect 472 290 533 306
rect 575 340 647 356
rect 575 306 591 340
rect 625 306 647 340
rect 575 290 647 306
rect 404 241 580 242
rect 25 214 118 230
rect 25 180 84 214
rect 404 207 530 241
rect 564 207 580 241
rect 404 206 580 207
rect 708 230 774 258
rect 708 202 724 230
rect 25 134 118 180
rect 25 100 84 134
rect 25 84 118 100
rect 154 168 170 202
rect 204 168 220 202
rect 154 134 220 168
rect 154 100 170 134
rect 204 100 220 134
rect 154 17 220 100
rect 257 186 318 202
rect 257 152 268 186
rect 302 152 318 186
rect 629 196 724 202
rect 758 196 774 230
rect 257 104 318 152
rect 352 138 368 172
rect 402 138 444 172
rect 478 138 587 172
rect 257 88 519 104
rect 257 54 469 88
rect 503 54 519 88
rect 257 51 519 54
rect 553 17 587 138
rect 629 168 774 196
rect 629 17 663 168
rect 697 88 839 134
rect 697 54 713 88
rect 747 54 839 88
rect 697 51 839 54
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
rlabel comment s 0 0 0 0 4 a2bb2o_1
flabel comment s 501 280 501 280 0 FreeSans 200 0 0 0 no_jumper_check
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 223 242 257 276 0 FreeSans 340 0 0 0 A1_N
port 1 nsew
flabel corelocali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 703 94 737 128 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 799 94 833 128 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 319 242 353 276 0 FreeSans 340 0 0 0 A2_N
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 864 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3494330
string GDS_START 3486380
<< end >>
