magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 17 195 69 265
rect 187 215 266 255
rect 304 215 381 341
rect 447 215 523 341
rect 709 409 769 493
rect 709 375 898 409
rect 567 215 665 257
rect 836 181 898 375
rect 709 147 898 181
rect 709 53 785 147
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 50 334 116 493
rect 160 370 202 527
rect 340 409 491 493
rect 236 375 593 409
rect 236 334 270 375
rect 50 299 270 334
rect 109 289 270 299
rect 109 161 153 289
rect 559 325 593 375
rect 629 359 675 527
rect 803 443 881 527
rect 559 291 743 325
rect 699 257 743 291
rect 699 215 775 257
rect 34 127 153 161
rect 227 147 597 181
rect 227 129 314 147
rect 34 51 100 127
rect 134 59 401 93
rect 453 17 487 111
rect 521 54 597 147
rect 641 17 675 181
rect 829 17 863 113
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
rlabel locali s 567 215 665 257 6 A1
port 1 nsew signal input
rlabel locali s 447 215 523 341 6 A2
port 2 nsew signal input
rlabel locali s 187 215 266 255 6 B1
port 3 nsew signal input
rlabel locali s 304 215 381 341 6 B2
port 4 nsew signal input
rlabel locali s 17 195 69 265 6 C1
port 5 nsew signal input
rlabel locali s 836 181 898 375 6 X
port 6 nsew signal output
rlabel locali s 709 409 769 493 6 X
port 6 nsew signal output
rlabel locali s 709 375 898 409 6 X
port 6 nsew signal output
rlabel locali s 709 147 898 181 6 X
port 6 nsew signal output
rlabel locali s 709 53 785 147 6 X
port 6 nsew signal output
rlabel metal1 s 0 -48 920 48 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 496 920 592 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 920 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 855110
string GDS_START 847288
<< end >>
