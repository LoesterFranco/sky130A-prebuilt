magic
tech sky130A
magscale 1 2
timestamp 1601050088
<< locali >>
rect 123 424 189 547
rect 313 424 379 547
rect 123 390 379 424
rect 25 270 286 356
rect 323 236 379 390
rect 123 202 389 236
rect 123 132 189 202
rect 323 132 389 202
rect 996 260 1130 326
rect 1081 236 1130 260
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 23 581 479 615
rect 23 390 89 581
rect 223 458 273 581
rect 413 362 479 581
rect 513 396 563 649
rect 603 362 653 596
rect 693 396 745 649
rect 879 596 957 598
rect 785 362 835 596
rect 413 328 835 362
rect 879 364 1039 596
rect 1079 364 1129 649
rect 879 328 957 364
rect 423 260 889 294
rect 23 85 89 226
rect 223 85 289 160
rect 423 85 489 260
rect 23 51 489 85
rect 523 17 589 226
rect 623 70 689 260
rect 723 17 789 226
rect 823 70 889 260
rect 923 226 957 328
rect 923 70 1001 226
rect 1035 17 1101 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
rlabel locali s 25 270 286 356 6 A
port 1 nsew signal input
rlabel locali s 1081 236 1130 260 6 TE
port 2 nsew signal input
rlabel locali s 996 260 1130 326 6 TE
port 2 nsew signal input
rlabel locali s 323 236 379 390 6 Z
port 3 nsew signal output
rlabel locali s 323 132 389 202 6 Z
port 3 nsew signal output
rlabel locali s 313 424 379 547 6 Z
port 3 nsew signal output
rlabel locali s 123 424 189 547 6 Z
port 3 nsew signal output
rlabel locali s 123 390 379 424 6 Z
port 3 nsew signal output
rlabel locali s 123 202 389 236 6 Z
port 3 nsew signal output
rlabel locali s 123 132 189 202 6 Z
port 3 nsew signal output
rlabel metal1 s 0 -49 1152 49 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 617 1152 715 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 2388520
string GDS_START 2379252
<< end >>
