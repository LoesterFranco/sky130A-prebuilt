magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 335 2342 704
rect -38 332 288 335
rect 620 332 2342 335
rect 620 324 1412 332
rect 1108 311 1412 324
<< pwell >>
rect 0 0 2304 49
<< scnmos >>
rect 95 78 125 162
rect 173 78 203 162
rect 379 119 409 267
rect 495 119 525 267
rect 702 119 732 203
rect 802 119 832 203
rect 880 119 910 203
rect 958 119 988 203
rect 1076 74 1106 202
rect 1194 74 1224 202
rect 1404 74 1434 158
rect 1482 74 1512 158
rect 1594 74 1624 158
rect 1672 74 1702 158
rect 1873 74 1903 222
rect 2088 74 2118 184
rect 2188 74 2218 222
<< pmoshvt >>
rect 86 508 116 592
rect 176 508 206 592
rect 378 392 408 592
rect 470 392 500 592
rect 675 463 705 547
rect 766 463 796 547
rect 844 463 874 547
rect 971 463 1001 547
rect 1203 347 1233 547
rect 1293 347 1323 547
rect 1435 471 1465 555
rect 1519 471 1549 555
rect 1621 471 1651 555
rect 1711 471 1741 555
rect 1814 368 1844 592
rect 2085 424 2115 592
rect 2188 368 2218 592
<< ndiff >>
rect 322 200 379 267
rect 322 166 334 200
rect 368 166 379 200
rect 38 137 95 162
rect 38 103 50 137
rect 84 103 95 137
rect 38 78 95 103
rect 125 78 173 162
rect 203 137 268 162
rect 203 103 222 137
rect 256 103 268 137
rect 322 119 379 166
rect 409 160 495 267
rect 409 126 434 160
rect 468 126 495 160
rect 409 119 495 126
rect 525 225 575 267
rect 525 161 584 225
rect 525 127 538 161
rect 572 127 584 161
rect 525 119 584 127
rect 643 179 702 203
rect 643 145 657 179
rect 691 145 702 179
rect 643 119 702 145
rect 732 179 802 203
rect 732 145 757 179
rect 791 145 802 179
rect 732 119 802 145
rect 832 119 880 203
rect 910 119 958 203
rect 988 202 1042 203
rect 1121 218 1179 230
rect 1121 202 1133 218
rect 988 119 1076 202
rect 203 78 268 103
rect 424 96 474 119
rect 1003 82 1076 119
rect 1003 48 1015 82
rect 1049 74 1076 82
rect 1106 184 1133 202
rect 1167 202 1179 218
rect 1167 184 1194 202
rect 1106 74 1194 184
rect 1224 158 1274 202
rect 1816 210 1873 222
rect 1816 176 1828 210
rect 1862 176 1873 210
rect 1224 130 1404 158
rect 1224 96 1322 130
rect 1356 96 1404 130
rect 1224 74 1404 96
rect 1434 74 1482 158
rect 1512 128 1594 158
rect 1512 94 1536 128
rect 1570 94 1594 128
rect 1512 74 1594 94
rect 1624 74 1672 158
rect 1702 133 1759 158
rect 1702 99 1713 133
rect 1747 99 1759 133
rect 1702 74 1759 99
rect 1816 120 1873 176
rect 1816 86 1828 120
rect 1862 86 1873 120
rect 1816 74 1873 86
rect 1903 210 1974 222
rect 1903 176 1928 210
rect 1962 176 1974 210
rect 2133 210 2188 222
rect 2133 184 2141 210
rect 1903 120 1974 176
rect 1903 86 1928 120
rect 1962 86 1974 120
rect 1903 74 1974 86
rect 2031 145 2088 184
rect 2031 111 2043 145
rect 2077 111 2088 145
rect 2031 74 2088 111
rect 2118 176 2141 184
rect 2175 176 2188 210
rect 2118 120 2188 176
rect 2118 86 2141 120
rect 2175 86 2188 120
rect 2118 74 2188 86
rect 2218 210 2275 222
rect 2218 176 2229 210
rect 2263 176 2275 210
rect 2218 120 2275 176
rect 2218 86 2229 120
rect 2263 86 2275 120
rect 2218 74 2275 86
rect 1049 48 1061 74
rect 1003 36 1061 48
<< pdiff >>
rect 27 567 86 592
rect 27 533 39 567
rect 73 533 86 567
rect 27 508 86 533
rect 116 567 176 592
rect 116 533 129 567
rect 163 533 176 567
rect 116 508 176 533
rect 206 584 265 592
rect 206 550 219 584
rect 253 550 265 584
rect 206 508 265 550
rect 319 434 378 592
rect 319 400 331 434
rect 365 400 378 434
rect 319 392 378 400
rect 408 584 470 592
rect 408 550 421 584
rect 455 550 470 584
rect 408 392 470 550
rect 500 448 557 592
rect 500 414 511 448
rect 545 414 557 448
rect 500 392 557 414
rect 892 567 953 579
rect 892 547 905 567
rect 617 522 675 547
rect 617 488 629 522
rect 663 488 675 522
rect 617 463 675 488
rect 705 539 766 547
rect 705 505 719 539
rect 753 505 766 539
rect 705 463 766 505
rect 796 463 844 547
rect 874 533 905 547
rect 939 547 953 567
rect 1759 567 1814 592
rect 1759 555 1767 567
rect 1382 547 1435 555
rect 939 533 971 547
rect 874 463 971 533
rect 1001 520 1057 547
rect 1001 486 1015 520
rect 1049 486 1057 520
rect 1001 463 1057 486
rect 1144 535 1203 547
rect 1144 501 1156 535
rect 1190 501 1203 535
rect 1144 466 1203 501
rect 1144 432 1156 466
rect 1190 432 1203 466
rect 1144 398 1203 432
rect 1144 364 1156 398
rect 1190 364 1203 398
rect 1144 347 1203 364
rect 1233 535 1293 547
rect 1233 501 1246 535
rect 1280 501 1293 535
rect 1233 464 1293 501
rect 1233 430 1246 464
rect 1280 430 1293 464
rect 1233 393 1293 430
rect 1233 359 1246 393
rect 1280 359 1293 393
rect 1233 347 1293 359
rect 1323 523 1435 547
rect 1323 489 1361 523
rect 1395 489 1435 523
rect 1323 471 1435 489
rect 1465 471 1519 555
rect 1549 530 1621 555
rect 1549 496 1567 530
rect 1601 496 1621 530
rect 1549 471 1621 496
rect 1651 530 1711 555
rect 1651 496 1664 530
rect 1698 496 1711 530
rect 1651 471 1711 496
rect 1741 533 1767 555
rect 1801 533 1814 567
rect 1741 471 1814 533
rect 1323 347 1376 471
rect 1759 437 1767 471
rect 1801 437 1814 471
rect 1759 368 1814 437
rect 1844 580 1967 592
rect 1844 546 1857 580
rect 1891 546 1925 580
rect 1959 546 1967 580
rect 1844 497 1967 546
rect 1844 463 1857 497
rect 1891 463 1925 497
rect 1959 463 1967 497
rect 1844 414 1967 463
rect 2026 579 2085 592
rect 2026 545 2038 579
rect 2072 545 2085 579
rect 2026 471 2085 545
rect 2026 437 2038 471
rect 2072 437 2085 471
rect 2026 424 2085 437
rect 2115 580 2188 592
rect 2115 546 2135 580
rect 2169 546 2188 580
rect 2115 497 2188 546
rect 2115 463 2135 497
rect 2169 463 2188 497
rect 2115 424 2188 463
rect 1844 380 1857 414
rect 1891 380 1925 414
rect 1959 380 1967 414
rect 2133 414 2188 424
rect 1844 368 1967 380
rect 2133 380 2141 414
rect 2175 380 2188 414
rect 2133 368 2188 380
rect 2218 580 2277 592
rect 2218 546 2231 580
rect 2265 546 2277 580
rect 2218 497 2277 546
rect 2218 463 2231 497
rect 2265 463 2277 497
rect 2218 414 2277 463
rect 2218 380 2231 414
rect 2265 380 2277 414
rect 2218 368 2277 380
<< ndiffc >>
rect 334 166 368 200
rect 50 103 84 137
rect 222 103 256 137
rect 434 126 468 160
rect 538 127 572 161
rect 657 145 691 179
rect 757 145 791 179
rect 1015 48 1049 82
rect 1133 184 1167 218
rect 1828 176 1862 210
rect 1322 96 1356 130
rect 1536 94 1570 128
rect 1713 99 1747 133
rect 1828 86 1862 120
rect 1928 176 1962 210
rect 1928 86 1962 120
rect 2043 111 2077 145
rect 2141 176 2175 210
rect 2141 86 2175 120
rect 2229 176 2263 210
rect 2229 86 2263 120
<< pdiffc >>
rect 39 533 73 567
rect 129 533 163 567
rect 219 550 253 584
rect 331 400 365 434
rect 421 550 455 584
rect 511 414 545 448
rect 629 488 663 522
rect 719 505 753 539
rect 905 533 939 567
rect 1015 486 1049 520
rect 1156 501 1190 535
rect 1156 432 1190 466
rect 1156 364 1190 398
rect 1246 501 1280 535
rect 1246 430 1280 464
rect 1246 359 1280 393
rect 1361 489 1395 523
rect 1567 496 1601 530
rect 1664 496 1698 530
rect 1767 533 1801 567
rect 1767 437 1801 471
rect 1857 546 1891 580
rect 1925 546 1959 580
rect 1857 463 1891 497
rect 1925 463 1959 497
rect 2038 545 2072 579
rect 2038 437 2072 471
rect 2135 546 2169 580
rect 2135 463 2169 497
rect 1857 380 1891 414
rect 1925 380 1959 414
rect 2141 380 2175 414
rect 2231 546 2265 580
rect 2231 463 2265 497
rect 2231 380 2265 414
<< poly >>
rect 86 592 116 618
rect 176 592 206 618
rect 378 592 408 618
rect 470 592 500 618
rect 572 615 1326 645
rect 86 493 116 508
rect 176 493 206 508
rect 83 470 119 493
rect 44 386 125 470
rect 44 352 60 386
rect 94 352 125 386
rect 44 318 125 352
rect 44 284 60 318
rect 94 284 125 318
rect 44 250 125 284
rect 44 216 60 250
rect 94 216 125 250
rect 44 200 125 216
rect 95 162 125 200
rect 173 428 209 493
rect 173 412 266 428
rect 173 378 216 412
rect 250 378 266 412
rect 173 344 266 378
rect 378 355 408 392
rect 470 355 500 392
rect 572 355 602 615
rect 675 547 705 573
rect 763 562 799 615
rect 766 547 796 562
rect 844 547 874 573
rect 971 547 1001 573
rect 1203 547 1233 573
rect 1290 562 1326 615
rect 1814 592 1844 618
rect 2085 592 2115 618
rect 2188 592 2218 618
rect 1293 547 1323 562
rect 1435 555 1465 581
rect 1519 555 1549 581
rect 1621 555 1651 581
rect 1711 555 1741 581
rect 675 442 705 463
rect 675 397 710 442
rect 766 437 796 463
rect 844 448 874 463
rect 971 448 1001 463
rect 841 431 877 448
rect 968 431 1004 448
rect 841 415 926 431
rect 841 401 876 415
rect 173 310 216 344
rect 250 310 266 344
rect 173 276 266 310
rect 357 339 428 355
rect 357 305 378 339
rect 412 305 428 339
rect 357 282 428 305
rect 470 339 602 355
rect 644 381 710 397
rect 644 347 660 381
rect 694 347 710 381
rect 644 342 710 347
rect 860 381 876 401
rect 910 381 926 415
rect 860 347 926 381
rect 644 339 818 342
rect 470 305 511 339
rect 545 314 602 339
rect 646 335 818 339
rect 648 333 818 335
rect 652 331 818 333
rect 659 324 818 331
rect 545 310 606 314
rect 667 312 818 324
rect 545 306 611 310
rect 545 305 613 306
rect 470 304 613 305
rect 470 302 617 304
rect 470 300 619 302
rect 470 297 621 300
rect 470 294 624 297
rect 470 282 629 294
rect 173 242 216 276
rect 250 242 266 276
rect 379 267 409 282
rect 495 267 525 282
rect 592 280 629 282
rect 595 278 629 280
rect 597 276 629 278
rect 599 270 629 276
rect 173 226 266 242
rect 173 162 203 226
rect 599 240 732 270
rect 702 203 732 240
rect 788 248 818 312
rect 860 313 876 347
rect 910 313 926 347
rect 860 297 926 313
rect 968 415 1112 431
rect 968 381 1062 415
rect 1096 381 1112 415
rect 968 365 1112 381
rect 788 218 832 248
rect 802 203 832 218
rect 880 203 910 297
rect 968 248 998 365
rect 1435 456 1465 471
rect 1519 456 1549 471
rect 1621 456 1651 471
rect 1711 456 1741 471
rect 1432 439 1468 456
rect 1408 423 1474 439
rect 1408 389 1424 423
rect 1458 389 1474 423
rect 1408 373 1474 389
rect 1203 332 1233 347
rect 1293 332 1323 347
rect 1200 323 1236 332
rect 1046 307 1236 323
rect 1046 273 1062 307
rect 1096 293 1236 307
rect 1290 325 1326 332
rect 1290 295 1434 325
rect 1096 273 1112 293
rect 1046 257 1112 273
rect 958 218 998 248
rect 958 203 988 218
rect 1076 202 1106 257
rect 1194 230 1362 247
rect 379 93 409 119
rect 495 93 525 119
rect 702 93 732 119
rect 802 93 832 119
rect 880 93 910 119
rect 95 52 125 78
rect 173 51 203 78
rect 958 51 988 119
rect 173 21 988 51
rect 1194 217 1312 230
rect 1194 202 1224 217
rect 1296 196 1312 217
rect 1346 196 1362 230
rect 1296 180 1362 196
rect 1404 158 1434 295
rect 1516 246 1552 456
rect 1618 433 1654 456
rect 1482 230 1552 246
rect 1482 196 1502 230
rect 1536 196 1552 230
rect 1482 180 1552 196
rect 1594 417 1660 433
rect 1594 383 1610 417
rect 1644 383 1660 417
rect 1594 367 1660 383
rect 1482 158 1512 180
rect 1594 158 1624 367
rect 1708 319 1744 456
rect 2085 409 2115 424
rect 1814 353 1844 368
rect 1811 319 1847 353
rect 2082 319 2118 409
rect 2188 353 2218 368
rect 2185 326 2221 353
rect 1666 303 2118 319
rect 1666 269 1682 303
rect 1716 269 2118 303
rect 1666 253 2118 269
rect 2160 310 2226 326
rect 2160 276 2176 310
rect 2210 276 2226 310
rect 2160 260 2226 276
rect 1672 158 1702 253
rect 1873 222 1903 253
rect 2088 184 2118 253
rect 2188 222 2218 260
rect 1076 48 1106 74
rect 1194 48 1224 74
rect 1404 48 1434 74
rect 1482 48 1512 74
rect 1594 48 1624 74
rect 1672 48 1702 74
rect 1873 48 1903 74
rect 2088 48 2118 74
rect 2188 48 2218 74
<< polycont >>
rect 60 352 94 386
rect 60 284 94 318
rect 60 216 94 250
rect 216 378 250 412
rect 216 310 250 344
rect 378 305 412 339
rect 660 347 694 381
rect 876 381 910 415
rect 511 305 545 339
rect 216 242 250 276
rect 876 313 910 347
rect 1062 381 1096 415
rect 1424 389 1458 423
rect 1062 273 1096 307
rect 1312 196 1346 230
rect 1502 196 1536 230
rect 1610 383 1644 417
rect 1682 269 1716 303
rect 2176 276 2210 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2304 683
rect 23 567 73 649
rect 23 533 39 567
rect 23 504 73 533
rect 113 567 169 596
rect 113 533 129 567
rect 163 533 169 567
rect 203 584 269 649
rect 203 550 219 584
rect 253 550 269 584
rect 405 584 471 649
rect 405 550 421 584
rect 455 550 471 584
rect 888 567 957 649
rect 113 526 169 533
rect 113 516 178 526
rect 613 522 669 538
rect 281 516 393 518
rect 613 516 629 522
rect 113 504 629 516
rect 138 488 629 504
rect 663 488 669 522
rect 703 505 719 539
rect 753 505 854 539
rect 888 533 905 567
rect 939 533 957 567
rect 998 520 1065 536
rect 998 508 1015 520
rect 138 484 669 488
rect 138 482 306 484
rect 378 482 669 484
rect 138 462 285 482
rect 629 471 669 482
rect 802 499 854 505
rect 989 499 1015 508
rect 802 486 1015 499
rect 1049 486 1065 520
rect 25 386 104 439
rect 25 352 60 386
rect 94 352 104 386
rect 25 318 104 352
rect 25 284 60 318
rect 94 284 104 318
rect 25 250 104 284
rect 25 216 60 250
rect 94 216 104 250
rect 25 200 104 216
rect 138 166 172 462
rect 319 434 365 450
rect 319 428 331 434
rect 206 424 260 428
rect 206 412 223 424
rect 206 378 216 412
rect 257 390 260 424
rect 250 378 260 390
rect 206 344 260 378
rect 206 310 216 344
rect 250 310 260 344
rect 206 276 260 310
rect 206 242 216 276
rect 250 242 260 276
rect 206 226 260 242
rect 294 400 331 428
rect 294 373 365 400
rect 495 414 511 448
rect 545 416 595 448
rect 629 437 768 471
rect 545 414 600 416
rect 495 413 600 414
rect 495 412 604 413
rect 495 408 605 412
rect 495 403 610 408
rect 495 381 700 403
rect 495 373 660 381
rect 294 228 328 373
rect 583 365 660 373
rect 589 359 660 365
rect 409 339 455 356
rect 595 347 660 359
rect 694 347 700 381
rect 362 305 378 339
rect 412 305 455 339
rect 495 310 511 339
rect 362 262 455 305
rect 489 305 511 310
rect 545 305 561 339
rect 489 298 561 305
rect 595 315 700 347
rect 489 228 555 298
rect 595 278 632 315
rect 294 200 555 228
rect 294 166 334 200
rect 368 195 555 200
rect 589 241 632 278
rect 734 274 768 437
rect 368 194 512 195
rect 368 166 384 194
rect 34 137 172 166
rect 34 103 50 137
rect 84 132 172 137
rect 206 137 256 166
rect 84 103 100 132
rect 34 74 100 103
rect 206 103 222 137
rect 294 119 384 166
rect 589 161 623 241
rect 666 240 768 274
rect 802 465 1065 486
rect 1156 535 1206 649
rect 1190 501 1206 535
rect 1156 466 1206 501
rect 666 207 707 240
rect 418 126 434 160
rect 468 126 484 160
rect 206 17 256 103
rect 418 17 484 126
rect 522 127 538 161
rect 572 127 623 161
rect 522 85 623 127
rect 657 179 707 207
rect 802 206 836 465
rect 978 456 1021 465
rect 691 145 707 179
rect 657 119 707 145
rect 741 179 836 206
rect 870 415 926 431
rect 870 381 876 415
rect 910 381 926 415
rect 870 347 926 381
rect 870 313 876 347
rect 910 313 926 347
rect 870 218 926 313
rect 978 323 1012 456
rect 1190 432 1206 466
rect 1046 424 1122 431
rect 1046 415 1087 424
rect 1046 381 1062 415
rect 1121 390 1122 424
rect 1096 381 1122 390
rect 1046 365 1122 381
rect 1156 398 1206 432
rect 1190 364 1206 398
rect 1156 348 1206 364
rect 1246 535 1296 551
rect 1280 501 1296 535
rect 1246 464 1296 501
rect 1340 523 1533 539
rect 1340 489 1361 523
rect 1395 489 1533 523
rect 1340 473 1533 489
rect 1280 430 1296 464
rect 1246 393 1296 430
rect 1280 359 1296 393
rect 978 307 1112 323
rect 1246 314 1296 359
rect 978 289 1062 307
rect 1046 273 1062 289
rect 1096 273 1112 307
rect 1046 257 1112 273
rect 1149 280 1296 314
rect 1330 423 1465 439
rect 1330 389 1424 423
rect 1458 389 1465 423
rect 1330 373 1465 389
rect 1149 218 1183 280
rect 1330 246 1364 373
rect 1499 319 1533 473
rect 1567 530 1612 649
rect 1762 567 1805 649
rect 1601 496 1612 530
rect 1567 467 1612 496
rect 1652 530 1728 546
rect 1652 496 1664 530
rect 1698 496 1728 530
rect 1652 467 1728 496
rect 1567 424 1660 433
rect 1601 417 1660 424
rect 1601 390 1610 417
rect 1567 383 1610 390
rect 1644 383 1660 417
rect 1567 367 1660 383
rect 1694 387 1728 467
rect 1762 533 1767 567
rect 1801 533 1805 567
rect 1762 471 1805 533
rect 1762 437 1767 471
rect 1801 437 1805 471
rect 1762 421 1805 437
rect 1852 580 1990 597
rect 1852 546 1857 580
rect 1891 546 1925 580
rect 1959 546 1990 580
rect 1852 497 1990 546
rect 1852 463 1857 497
rect 1891 463 1925 497
rect 1959 463 1990 497
rect 1852 414 1990 463
rect 1694 353 1794 387
rect 1852 380 1857 414
rect 1891 380 1925 414
rect 1959 380 1990 414
rect 1852 362 1990 380
rect 870 184 1133 218
rect 1167 184 1183 218
rect 1217 230 1364 246
rect 1217 196 1312 230
rect 1346 196 1364 230
rect 741 145 757 179
rect 791 145 836 179
rect 1217 180 1364 196
rect 1398 303 1726 319
rect 1398 285 1682 303
rect 1217 150 1251 180
rect 741 119 836 145
rect 870 116 1251 150
rect 1398 146 1432 285
rect 1666 269 1682 285
rect 1716 269 1726 303
rect 1666 253 1726 269
rect 1486 230 1552 246
rect 1486 196 1502 230
rect 1536 214 1552 230
rect 1760 214 1794 353
rect 1536 196 1794 214
rect 1486 180 1794 196
rect 1285 130 1432 146
rect 870 85 904 116
rect 522 51 904 85
rect 1285 96 1322 130
rect 1356 96 1432 130
rect 999 48 1015 82
rect 1049 48 1065 82
rect 1285 80 1432 96
rect 1507 128 1599 136
rect 1507 94 1536 128
rect 1570 94 1599 128
rect 999 17 1065 48
rect 1507 17 1599 94
rect 1697 133 1794 180
rect 1697 99 1713 133
rect 1747 99 1794 133
rect 1697 70 1794 99
rect 1828 210 1878 226
rect 1862 176 1878 210
rect 1828 120 1878 176
rect 1862 86 1878 120
rect 1828 17 1878 86
rect 1912 210 1990 362
rect 1912 176 1928 210
rect 1962 176 1990 210
rect 1912 120 1990 176
rect 1912 86 1928 120
rect 1962 86 1990 120
rect 1912 70 1990 86
rect 2038 579 2088 595
rect 2072 545 2088 579
rect 2038 471 2088 545
rect 2072 437 2088 471
rect 2038 326 2088 437
rect 2122 580 2181 649
rect 2122 546 2135 580
rect 2169 546 2181 580
rect 2122 497 2181 546
rect 2122 463 2135 497
rect 2169 463 2181 497
rect 2122 414 2181 463
rect 2122 380 2141 414
rect 2175 380 2181 414
rect 2122 364 2181 380
rect 2215 580 2287 596
rect 2215 546 2231 580
rect 2265 546 2287 580
rect 2215 497 2287 546
rect 2215 463 2231 497
rect 2265 463 2287 497
rect 2215 414 2287 463
rect 2215 380 2231 414
rect 2265 380 2287 414
rect 2215 364 2287 380
rect 2038 310 2219 326
rect 2038 276 2176 310
rect 2210 276 2219 310
rect 2038 260 2219 276
rect 2038 145 2088 260
rect 2253 226 2287 364
rect 2038 111 2043 145
rect 2077 111 2088 145
rect 2038 70 2088 111
rect 2129 210 2179 226
rect 2129 176 2141 210
rect 2175 176 2179 210
rect 2129 120 2179 176
rect 2129 86 2141 120
rect 2175 86 2179 120
rect 2129 17 2179 86
rect 2213 210 2287 226
rect 2213 176 2229 210
rect 2263 176 2287 210
rect 2213 120 2287 176
rect 2213 86 2229 120
rect 2263 86 2287 120
rect 2213 70 2287 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2304 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 223 412 257 424
rect 223 390 250 412
rect 250 390 257 412
rect 1087 415 1121 424
rect 1087 390 1096 415
rect 1096 390 1121 415
rect 1567 390 1601 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
<< metal1 >>
rect 0 683 2304 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2304 683
rect 0 617 2304 649
rect 211 424 269 430
rect 211 390 223 424
rect 257 421 269 424
rect 1075 424 1133 430
rect 1075 421 1087 424
rect 257 393 1087 421
rect 257 390 269 393
rect 211 384 269 390
rect 1075 390 1087 393
rect 1121 421 1133 424
rect 1555 424 1613 430
rect 1555 421 1567 424
rect 1121 393 1567 421
rect 1121 390 1133 393
rect 1075 384 1133 390
rect 1555 390 1567 393
rect 1601 390 1613 424
rect 1555 384 1613 390
rect 0 17 2304 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2304 17
rect 0 -49 2304 -17
<< labels >>
flabel comment s 602 36 602 36 0 FreeSans 300 0 0 0 no_jumper_check
flabel comment s 940 630 940 630 0 FreeSans 300 0 0 0 no_jumper_check
rlabel comment s 0 0 0 0 4 dfrbp_1
flabel pwell s 0 0 2304 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 0 617 2304 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 223 390 257 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew
flabel metal1 s 0 617 2304 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 2304 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 2239 94 2273 128 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 2239 168 2273 202 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 2239 390 2273 424 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 31 390 65 424 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 1951 390 1985 424 0 FreeSans 340 0 0 0 Q_N
port 9 nsew
flabel corelocali s 1951 464 1985 498 0 FreeSans 340 0 0 0 Q_N
port 9 nsew
flabel corelocali s 1951 538 1985 572 0 FreeSans 340 0 0 0 Q_N
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 2304 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2549030
string GDS_START 2530424
<< end >>
