magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 2246 582
<< pwell >>
rect 27 -17 61 17
<< scnmos >>
rect 83 47 113 177
rect 177 47 207 177
rect 271 47 301 177
rect 375 47 405 177
rect 459 47 489 177
rect 553 47 583 177
rect 647 47 677 177
rect 751 47 781 177
rect 939 47 969 177
rect 1033 47 1063 177
rect 1127 47 1157 177
rect 1231 47 1261 177
rect 1413 47 1443 177
rect 1507 47 1537 177
rect 1601 47 1631 177
rect 1705 47 1735 177
rect 1789 47 1819 177
rect 1883 47 1913 177
rect 1977 47 2007 177
rect 2081 47 2111 177
<< pmoshvt >>
rect 85 297 121 497
rect 179 297 215 497
rect 273 297 309 497
rect 367 297 403 497
rect 461 297 497 497
rect 555 297 591 497
rect 649 297 685 497
rect 743 297 779 497
rect 935 297 971 497
rect 1029 297 1065 497
rect 1123 297 1159 497
rect 1217 297 1253 497
rect 1415 297 1451 497
rect 1509 297 1545 497
rect 1603 297 1639 497
rect 1697 297 1733 497
rect 1791 297 1827 497
rect 1885 297 1921 497
rect 1979 297 2015 497
rect 2073 297 2109 497
<< ndiff >>
rect 27 95 83 177
rect 27 61 39 95
rect 73 61 83 95
rect 27 47 83 61
rect 113 163 177 177
rect 113 129 133 163
rect 167 129 177 163
rect 113 47 177 129
rect 207 95 271 177
rect 207 61 227 95
rect 261 61 271 95
rect 207 47 271 61
rect 301 163 375 177
rect 301 129 321 163
rect 355 129 375 163
rect 301 47 375 129
rect 405 163 459 177
rect 405 129 415 163
rect 449 129 459 163
rect 405 95 459 129
rect 405 61 415 95
rect 449 61 459 95
rect 405 47 459 61
rect 489 95 553 177
rect 489 61 509 95
rect 543 61 553 95
rect 489 47 553 61
rect 583 163 647 177
rect 583 129 603 163
rect 637 129 647 163
rect 583 95 647 129
rect 583 61 603 95
rect 637 61 647 95
rect 583 47 647 61
rect 677 95 751 177
rect 677 61 697 95
rect 731 61 751 95
rect 677 47 751 61
rect 781 163 833 177
rect 781 129 791 163
rect 825 129 833 163
rect 781 95 833 129
rect 781 61 791 95
rect 825 61 833 95
rect 781 47 833 61
rect 887 133 939 177
rect 887 99 895 133
rect 929 99 939 133
rect 887 47 939 99
rect 969 163 1033 177
rect 969 129 989 163
rect 1023 129 1033 163
rect 969 47 1033 129
rect 1063 95 1127 177
rect 1063 61 1083 95
rect 1117 61 1127 95
rect 1063 47 1127 61
rect 1157 163 1231 177
rect 1157 129 1177 163
rect 1211 129 1231 163
rect 1157 47 1231 129
rect 1261 95 1413 177
rect 1261 61 1271 95
rect 1305 61 1369 95
rect 1403 61 1413 95
rect 1261 47 1413 61
rect 1443 95 1507 177
rect 1443 61 1463 95
rect 1497 61 1507 95
rect 1443 47 1507 61
rect 1537 163 1601 177
rect 1537 129 1557 163
rect 1591 129 1601 163
rect 1537 95 1601 129
rect 1537 61 1557 95
rect 1591 61 1601 95
rect 1537 47 1601 61
rect 1631 95 1705 177
rect 1631 61 1651 95
rect 1685 61 1705 95
rect 1631 47 1705 61
rect 1735 163 1789 177
rect 1735 129 1745 163
rect 1779 129 1789 163
rect 1735 95 1789 129
rect 1735 61 1745 95
rect 1779 61 1789 95
rect 1735 47 1789 61
rect 1819 95 1883 177
rect 1819 61 1839 95
rect 1873 61 1883 95
rect 1819 47 1883 61
rect 1913 163 1977 177
rect 1913 129 1933 163
rect 1967 129 1977 163
rect 1913 95 1977 129
rect 1913 61 1933 95
rect 1967 61 1977 95
rect 1913 47 1977 61
rect 2007 95 2081 177
rect 2007 61 2027 95
rect 2061 61 2081 95
rect 2007 47 2081 61
rect 2111 163 2163 177
rect 2111 129 2121 163
rect 2155 129 2163 163
rect 2111 95 2163 129
rect 2111 61 2121 95
rect 2155 61 2163 95
rect 2111 47 2163 61
<< pdiff >>
rect 27 477 85 497
rect 27 443 39 477
rect 73 443 85 477
rect 27 409 85 443
rect 27 375 39 409
rect 73 375 85 409
rect 27 297 85 375
rect 121 477 179 497
rect 121 443 133 477
rect 167 443 179 477
rect 121 409 179 443
rect 121 375 133 409
rect 167 375 179 409
rect 121 341 179 375
rect 121 307 133 341
rect 167 307 179 341
rect 121 297 179 307
rect 215 477 273 497
rect 215 443 227 477
rect 261 443 273 477
rect 215 409 273 443
rect 215 375 227 409
rect 261 375 273 409
rect 215 297 273 375
rect 309 477 367 497
rect 309 443 321 477
rect 355 443 367 477
rect 309 409 367 443
rect 309 375 321 409
rect 355 375 367 409
rect 309 341 367 375
rect 309 307 321 341
rect 355 307 367 341
rect 309 297 367 307
rect 403 477 461 497
rect 403 443 415 477
rect 449 443 461 477
rect 403 409 461 443
rect 403 375 415 409
rect 449 375 461 409
rect 403 297 461 375
rect 497 477 555 497
rect 497 443 509 477
rect 543 443 555 477
rect 497 409 555 443
rect 497 375 509 409
rect 543 375 555 409
rect 497 341 555 375
rect 497 307 509 341
rect 543 307 555 341
rect 497 297 555 307
rect 591 477 649 497
rect 591 443 603 477
rect 637 443 649 477
rect 591 409 649 443
rect 591 375 603 409
rect 637 375 649 409
rect 591 297 649 375
rect 685 477 743 497
rect 685 443 697 477
rect 731 443 743 477
rect 685 409 743 443
rect 685 375 697 409
rect 731 375 743 409
rect 685 341 743 375
rect 685 307 697 341
rect 731 307 743 341
rect 685 297 743 307
rect 779 477 935 497
rect 779 443 791 477
rect 825 443 889 477
rect 923 443 935 477
rect 779 409 935 443
rect 779 375 791 409
rect 825 375 889 409
rect 923 375 935 409
rect 779 297 935 375
rect 971 477 1029 497
rect 971 443 983 477
rect 1017 443 1029 477
rect 971 409 1029 443
rect 971 375 983 409
rect 1017 375 1029 409
rect 971 341 1029 375
rect 971 307 983 341
rect 1017 307 1029 341
rect 971 297 1029 307
rect 1065 477 1123 497
rect 1065 443 1077 477
rect 1111 443 1123 477
rect 1065 409 1123 443
rect 1065 375 1077 409
rect 1111 375 1123 409
rect 1065 297 1123 375
rect 1159 477 1217 497
rect 1159 443 1171 477
rect 1205 443 1217 477
rect 1159 409 1217 443
rect 1159 375 1171 409
rect 1205 375 1217 409
rect 1159 341 1217 375
rect 1159 307 1171 341
rect 1205 307 1217 341
rect 1159 297 1217 307
rect 1253 477 1307 497
rect 1253 443 1265 477
rect 1299 443 1307 477
rect 1253 409 1307 443
rect 1253 375 1265 409
rect 1299 375 1307 409
rect 1253 297 1307 375
rect 1361 477 1415 497
rect 1361 443 1369 477
rect 1403 443 1415 477
rect 1361 409 1415 443
rect 1361 375 1369 409
rect 1403 375 1415 409
rect 1361 297 1415 375
rect 1451 409 1509 497
rect 1451 375 1463 409
rect 1497 375 1509 409
rect 1451 341 1509 375
rect 1451 307 1463 341
rect 1497 307 1509 341
rect 1451 297 1509 307
rect 1545 477 1603 497
rect 1545 443 1557 477
rect 1591 443 1603 477
rect 1545 409 1603 443
rect 1545 375 1557 409
rect 1591 375 1603 409
rect 1545 297 1603 375
rect 1639 409 1697 497
rect 1639 375 1651 409
rect 1685 375 1697 409
rect 1639 341 1697 375
rect 1639 307 1651 341
rect 1685 307 1697 341
rect 1639 297 1697 307
rect 1733 477 1791 497
rect 1733 443 1745 477
rect 1779 443 1791 477
rect 1733 409 1791 443
rect 1733 375 1745 409
rect 1779 375 1791 409
rect 1733 341 1791 375
rect 1733 307 1745 341
rect 1779 307 1791 341
rect 1733 297 1791 307
rect 1827 477 1885 497
rect 1827 443 1839 477
rect 1873 443 1885 477
rect 1827 409 1885 443
rect 1827 375 1839 409
rect 1873 375 1885 409
rect 1827 297 1885 375
rect 1921 477 1979 497
rect 1921 443 1933 477
rect 1967 443 1979 477
rect 1921 409 1979 443
rect 1921 375 1933 409
rect 1967 375 1979 409
rect 1921 341 1979 375
rect 1921 307 1933 341
rect 1967 307 1979 341
rect 1921 297 1979 307
rect 2015 477 2073 497
rect 2015 443 2027 477
rect 2061 443 2073 477
rect 2015 409 2073 443
rect 2015 375 2027 409
rect 2061 375 2073 409
rect 2015 297 2073 375
rect 2109 477 2167 497
rect 2109 443 2121 477
rect 2155 443 2167 477
rect 2109 409 2167 443
rect 2109 375 2121 409
rect 2155 375 2167 409
rect 2109 341 2167 375
rect 2109 307 2121 341
rect 2155 307 2167 341
rect 2109 297 2167 307
<< ndiffc >>
rect 39 61 73 95
rect 133 129 167 163
rect 227 61 261 95
rect 321 129 355 163
rect 415 129 449 163
rect 415 61 449 95
rect 509 61 543 95
rect 603 129 637 163
rect 603 61 637 95
rect 697 61 731 95
rect 791 129 825 163
rect 791 61 825 95
rect 895 99 929 133
rect 989 129 1023 163
rect 1083 61 1117 95
rect 1177 129 1211 163
rect 1271 61 1305 95
rect 1369 61 1403 95
rect 1463 61 1497 95
rect 1557 129 1591 163
rect 1557 61 1591 95
rect 1651 61 1685 95
rect 1745 129 1779 163
rect 1745 61 1779 95
rect 1839 61 1873 95
rect 1933 129 1967 163
rect 1933 61 1967 95
rect 2027 61 2061 95
rect 2121 129 2155 163
rect 2121 61 2155 95
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 133 443 167 477
rect 133 375 167 409
rect 133 307 167 341
rect 227 443 261 477
rect 227 375 261 409
rect 321 443 355 477
rect 321 375 355 409
rect 321 307 355 341
rect 415 443 449 477
rect 415 375 449 409
rect 509 443 543 477
rect 509 375 543 409
rect 509 307 543 341
rect 603 443 637 477
rect 603 375 637 409
rect 697 443 731 477
rect 697 375 731 409
rect 697 307 731 341
rect 791 443 825 477
rect 889 443 923 477
rect 791 375 825 409
rect 889 375 923 409
rect 983 443 1017 477
rect 983 375 1017 409
rect 983 307 1017 341
rect 1077 443 1111 477
rect 1077 375 1111 409
rect 1171 443 1205 477
rect 1171 375 1205 409
rect 1171 307 1205 341
rect 1265 443 1299 477
rect 1265 375 1299 409
rect 1369 443 1403 477
rect 1369 375 1403 409
rect 1463 375 1497 409
rect 1463 307 1497 341
rect 1557 443 1591 477
rect 1557 375 1591 409
rect 1651 375 1685 409
rect 1651 307 1685 341
rect 1745 443 1779 477
rect 1745 375 1779 409
rect 1745 307 1779 341
rect 1839 443 1873 477
rect 1839 375 1873 409
rect 1933 443 1967 477
rect 1933 375 1967 409
rect 1933 307 1967 341
rect 2027 443 2061 477
rect 2027 375 2061 409
rect 2121 443 2155 477
rect 2121 375 2155 409
rect 2121 307 2155 341
<< poly >>
rect 85 497 121 523
rect 179 497 215 523
rect 273 497 309 523
rect 367 497 403 523
rect 461 497 497 523
rect 555 497 591 523
rect 649 497 685 523
rect 743 497 779 523
rect 935 497 971 523
rect 1029 497 1065 523
rect 1123 497 1159 523
rect 1217 497 1253 523
rect 1415 497 1451 523
rect 1509 497 1545 523
rect 1603 497 1639 523
rect 1697 497 1733 523
rect 1791 497 1827 523
rect 1885 497 1921 523
rect 1979 497 2015 523
rect 2073 497 2109 523
rect 85 282 121 297
rect 179 282 215 297
rect 273 282 309 297
rect 367 282 403 297
rect 461 282 497 297
rect 555 282 591 297
rect 649 282 685 297
rect 743 282 779 297
rect 935 282 971 297
rect 1029 282 1065 297
rect 1123 282 1159 297
rect 1217 282 1253 297
rect 1415 282 1451 297
rect 1509 282 1545 297
rect 1603 282 1639 297
rect 1697 282 1733 297
rect 1791 282 1827 297
rect 1885 282 1921 297
rect 1979 282 2015 297
rect 2073 282 2109 297
rect 83 265 123 282
rect 177 265 217 282
rect 271 265 311 282
rect 365 265 405 282
rect 83 249 405 265
rect 83 215 101 249
rect 135 215 179 249
rect 213 215 257 249
rect 291 215 335 249
rect 369 215 405 249
rect 83 199 405 215
rect 83 177 113 199
rect 177 177 207 199
rect 271 177 301 199
rect 375 177 405 199
rect 459 265 499 282
rect 553 265 593 282
rect 647 265 687 282
rect 741 265 781 282
rect 459 249 781 265
rect 459 215 475 249
rect 509 215 553 249
rect 587 215 631 249
rect 665 215 709 249
rect 743 215 781 249
rect 459 199 781 215
rect 933 265 973 282
rect 1027 265 1067 282
rect 1121 265 1161 282
rect 1215 265 1255 282
rect 1413 265 1453 282
rect 1507 265 1547 282
rect 1601 265 1641 282
rect 1695 265 1735 282
rect 933 249 1261 265
rect 933 215 955 249
rect 989 215 1033 249
rect 1067 215 1111 249
rect 1145 215 1189 249
rect 1223 215 1261 249
rect 933 199 1261 215
rect 459 177 489 199
rect 553 177 583 199
rect 647 177 677 199
rect 751 177 781 199
rect 939 177 969 199
rect 1033 177 1063 199
rect 1127 177 1157 199
rect 1231 177 1261 199
rect 1413 249 1735 265
rect 1413 215 1429 249
rect 1463 215 1507 249
rect 1541 215 1585 249
rect 1619 215 1663 249
rect 1697 215 1735 249
rect 1413 199 1735 215
rect 1413 177 1443 199
rect 1507 177 1537 199
rect 1601 177 1631 199
rect 1705 177 1735 199
rect 1789 265 1829 282
rect 1883 265 1923 282
rect 1977 265 2017 282
rect 2071 265 2111 282
rect 1789 249 2111 265
rect 1789 215 1799 249
rect 1833 215 1877 249
rect 1911 215 1955 249
rect 1989 215 2033 249
rect 2067 215 2111 249
rect 1789 199 2111 215
rect 1789 177 1819 199
rect 1883 177 1913 199
rect 1977 177 2007 199
rect 2081 177 2111 199
rect 83 21 113 47
rect 177 21 207 47
rect 271 21 301 47
rect 375 21 405 47
rect 459 21 489 47
rect 553 21 583 47
rect 647 21 677 47
rect 751 21 781 47
rect 939 21 969 47
rect 1033 21 1063 47
rect 1127 21 1157 47
rect 1231 21 1261 47
rect 1413 21 1443 47
rect 1507 21 1537 47
rect 1601 21 1631 47
rect 1705 21 1735 47
rect 1789 21 1819 47
rect 1883 21 1913 47
rect 1977 21 2007 47
rect 2081 21 2111 47
<< polycont >>
rect 101 215 135 249
rect 179 215 213 249
rect 257 215 291 249
rect 335 215 369 249
rect 475 215 509 249
rect 553 215 587 249
rect 631 215 665 249
rect 709 215 743 249
rect 955 215 989 249
rect 1033 215 1067 249
rect 1111 215 1145 249
rect 1189 215 1223 249
rect 1429 215 1463 249
rect 1507 215 1541 249
rect 1585 215 1619 249
rect 1663 215 1697 249
rect 1799 215 1833 249
rect 1877 215 1911 249
rect 1955 215 1989 249
rect 2033 215 2067 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 31 477 81 527
rect 31 443 39 477
rect 73 443 81 477
rect 31 409 81 443
rect 31 375 39 409
rect 73 375 81 409
rect 31 359 81 375
rect 125 477 175 493
rect 125 443 133 477
rect 167 443 175 477
rect 125 409 175 443
rect 125 375 133 409
rect 167 375 175 409
rect 125 341 175 375
rect 219 477 269 527
rect 219 443 227 477
rect 261 443 269 477
rect 219 409 269 443
rect 219 375 227 409
rect 261 375 269 409
rect 219 359 269 375
rect 313 477 363 493
rect 313 443 321 477
rect 355 443 363 477
rect 313 409 363 443
rect 313 375 321 409
rect 355 375 363 409
rect 125 325 133 341
rect 17 307 133 325
rect 167 325 175 341
rect 313 341 363 375
rect 407 477 457 527
rect 407 443 415 477
rect 449 443 457 477
rect 407 409 457 443
rect 407 375 415 409
rect 449 375 457 409
rect 407 359 457 375
rect 501 477 551 493
rect 501 443 509 477
rect 543 443 551 477
rect 501 409 551 443
rect 501 375 509 409
rect 543 375 551 409
rect 313 325 321 341
rect 167 307 321 325
rect 355 325 363 341
rect 501 341 551 375
rect 595 477 645 527
rect 595 443 603 477
rect 637 443 645 477
rect 595 409 645 443
rect 595 375 603 409
rect 637 375 645 409
rect 595 359 645 375
rect 689 477 739 493
rect 689 443 697 477
rect 731 443 739 477
rect 689 409 739 443
rect 689 375 697 409
rect 731 375 739 409
rect 501 325 509 341
rect 355 307 509 325
rect 543 325 551 341
rect 689 341 739 375
rect 783 477 931 527
rect 783 443 791 477
rect 825 443 889 477
rect 923 443 931 477
rect 783 409 931 443
rect 783 375 791 409
rect 825 375 889 409
rect 923 375 931 409
rect 783 359 931 375
rect 975 477 1025 493
rect 975 443 983 477
rect 1017 443 1025 477
rect 975 409 1025 443
rect 975 375 983 409
rect 1017 375 1025 409
rect 689 325 697 341
rect 543 307 697 325
rect 731 325 739 341
rect 975 341 1025 375
rect 1069 477 1119 527
rect 1069 443 1077 477
rect 1111 443 1119 477
rect 1069 409 1119 443
rect 1069 375 1077 409
rect 1111 375 1119 409
rect 1069 359 1119 375
rect 1163 477 1213 493
rect 1163 443 1171 477
rect 1205 443 1213 477
rect 1163 409 1213 443
rect 1163 375 1171 409
rect 1205 375 1213 409
rect 731 307 863 325
rect 17 291 863 307
rect 975 307 983 341
rect 1017 325 1025 341
rect 1163 341 1213 375
rect 1257 477 1307 527
rect 1257 443 1265 477
rect 1299 443 1307 477
rect 1257 409 1307 443
rect 1257 375 1265 409
rect 1299 375 1307 409
rect 1257 359 1307 375
rect 1355 477 1787 493
rect 1355 443 1369 477
rect 1403 459 1557 477
rect 1403 443 1411 459
rect 1355 409 1411 443
rect 1549 443 1557 459
rect 1591 459 1745 477
rect 1591 443 1599 459
rect 1355 375 1369 409
rect 1403 375 1411 409
rect 1355 359 1411 375
rect 1455 409 1505 425
rect 1455 375 1463 409
rect 1497 375 1505 409
rect 1163 325 1171 341
rect 1017 307 1171 325
rect 1205 325 1213 341
rect 1455 341 1505 375
rect 1549 409 1599 443
rect 1737 443 1745 459
rect 1779 443 1787 477
rect 1549 375 1557 409
rect 1591 375 1599 409
rect 1549 359 1599 375
rect 1643 409 1693 425
rect 1643 375 1651 409
rect 1685 375 1693 409
rect 1455 325 1463 341
rect 1205 307 1463 325
rect 1497 325 1505 341
rect 1643 341 1693 375
rect 1643 325 1651 341
rect 1497 307 1651 325
rect 1685 307 1693 341
rect 975 291 1693 307
rect 1737 409 1787 443
rect 1737 375 1745 409
rect 1779 375 1787 409
rect 1737 341 1787 375
rect 1831 477 1881 527
rect 1831 443 1839 477
rect 1873 443 1881 477
rect 1831 409 1881 443
rect 1831 375 1839 409
rect 1873 375 1881 409
rect 1831 359 1881 375
rect 1925 477 1975 493
rect 1925 443 1933 477
rect 1967 443 1975 477
rect 1925 409 1975 443
rect 1925 375 1933 409
rect 1967 375 1975 409
rect 1737 307 1745 341
rect 1779 325 1787 341
rect 1925 341 1975 375
rect 2019 477 2069 527
rect 2019 443 2027 477
rect 2061 443 2069 477
rect 2019 409 2069 443
rect 2019 375 2027 409
rect 2061 375 2069 409
rect 2019 359 2069 375
rect 2113 477 2175 493
rect 2113 443 2121 477
rect 2155 443 2175 477
rect 2113 409 2175 443
rect 2113 375 2121 409
rect 2155 375 2175 409
rect 1925 325 1933 341
rect 1779 307 1933 325
rect 1967 325 1975 341
rect 2113 341 2175 375
rect 2113 325 2121 341
rect 1967 307 2121 325
rect 2155 307 2175 341
rect 1737 291 2175 307
rect 17 181 51 291
rect 829 257 863 291
rect 85 249 405 257
rect 85 215 101 249
rect 135 215 179 249
rect 213 215 257 249
rect 291 215 335 249
rect 369 215 405 249
rect 459 249 781 257
rect 459 215 475 249
rect 509 215 553 249
rect 587 215 631 249
rect 665 215 709 249
rect 743 215 781 249
rect 829 249 1261 257
rect 829 215 955 249
rect 989 215 1033 249
rect 1067 215 1111 249
rect 1145 215 1189 249
rect 1223 215 1261 249
rect 1295 181 1361 291
rect 1413 249 1735 257
rect 1413 215 1429 249
rect 1463 215 1507 249
rect 1541 215 1585 249
rect 1619 215 1663 249
rect 1697 215 1735 249
rect 1769 249 2188 257
rect 1769 215 1799 249
rect 1833 215 1877 249
rect 1911 215 1955 249
rect 1989 215 2033 249
rect 2067 215 2188 249
rect 17 163 371 181
rect 17 129 133 163
rect 167 129 321 163
rect 355 129 371 163
rect 415 163 841 181
rect 449 145 603 163
rect 449 129 465 145
rect 415 95 465 129
rect 577 129 603 145
rect 637 145 791 163
rect 637 129 653 145
rect 20 61 39 95
rect 73 61 227 95
rect 261 61 415 95
rect 449 61 465 95
rect 20 51 465 61
rect 509 95 543 111
rect 509 17 543 61
rect 577 95 653 129
rect 765 129 791 145
rect 825 129 841 163
rect 577 61 603 95
rect 637 61 653 95
rect 577 51 653 61
rect 697 95 731 111
rect 697 17 731 61
rect 765 95 841 129
rect 765 61 791 95
rect 825 61 841 95
rect 765 51 841 61
rect 892 133 929 167
rect 892 99 895 133
rect 973 163 1361 181
rect 973 129 989 163
rect 1023 129 1177 163
rect 1211 129 1361 163
rect 1395 163 2171 181
rect 1395 147 1557 163
rect 892 95 929 99
rect 1395 95 1429 147
rect 1531 129 1557 147
rect 1591 145 1745 163
rect 1591 129 1607 145
rect 892 61 1083 95
rect 1117 61 1271 95
rect 1305 61 1369 95
rect 1403 61 1429 95
rect 892 51 1429 61
rect 1463 95 1497 111
rect 1463 17 1497 61
rect 1531 95 1607 129
rect 1719 129 1745 145
rect 1779 145 1933 163
rect 1779 129 1795 145
rect 1531 61 1557 95
rect 1591 61 1607 95
rect 1531 51 1607 61
rect 1651 95 1685 111
rect 1651 17 1685 61
rect 1719 95 1795 129
rect 1907 129 1933 145
rect 1967 145 2121 163
rect 1967 129 1983 145
rect 1719 61 1745 95
rect 1779 61 1795 95
rect 1719 51 1795 61
rect 1839 95 1873 111
rect 1839 17 1873 61
rect 1907 95 1983 129
rect 2095 129 2121 145
rect 2155 129 2171 163
rect 1907 61 1933 95
rect 1967 61 1983 95
rect 1907 51 1983 61
rect 2027 95 2061 111
rect 2027 17 2061 61
rect 2095 95 2171 129
rect 2095 61 2121 95
rect 2155 61 2171 95
rect 2095 51 2171 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
<< metal1 >>
rect 0 561 2208 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 0 496 2208 527
rect 0 17 2208 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
rect 0 -48 2208 -17
<< labels >>
flabel corelocali s 596 238 596 238 0 FreeSans 400 0 0 0 A1_N
port 1 nsew
flabel corelocali s 1960 221 1994 255 0 FreeSans 400 0 0 0 B1
port 3 nsew
flabel corelocali s 1549 221 1583 255 0 FreeSans 400 0 0 0 B2
port 4 nsew
flabel corelocali s 228 238 228 238 0 FreeSans 400 0 0 0 A2_N
port 2 nsew
flabel corelocali s 1317 289 1351 323 0 FreeSans 400 0 0 0 Y
port 9 nsew
flabel nbase s 27 527 61 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel pwell s 27 -17 61 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel metal1 s 27 -17 61 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel metal1 s 27 527 61 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
rlabel comment s 0 0 0 0 4 o2bb2ai_4
<< properties >>
string FIXED_BBOX 0 0 2208 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 686526
string GDS_START 670836
<< end >>
