magic
tech sky130A
magscale 1 2
timestamp 1599588232
<< locali >>
rect 85 196 167 398
rect 313 290 381 356
rect 743 236 877 310
rect 2585 364 2668 596
rect 2798 364 2863 596
rect 2585 200 2619 364
rect 2553 124 2619 200
rect 2829 230 2863 364
rect 2791 74 2863 230
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2880 683
rect 17 492 89 596
rect 191 526 241 649
rect 275 581 445 615
rect 275 492 309 581
rect 17 458 309 492
rect 17 150 51 458
rect 343 424 377 547
rect 411 492 445 581
rect 479 526 529 649
rect 631 496 709 592
rect 743 530 809 649
rect 1021 530 1087 649
rect 1121 578 1289 612
rect 1121 496 1155 578
rect 1330 544 1396 596
rect 1539 577 1605 649
rect 631 492 1155 496
rect 411 462 1155 492
rect 1310 510 1396 544
rect 1639 551 1881 585
rect 1639 543 1673 551
rect 411 458 709 462
rect 201 390 533 424
rect 201 256 267 390
rect 201 222 400 256
rect 17 84 120 150
rect 218 17 284 162
rect 330 96 400 222
rect 467 196 533 390
rect 575 350 641 398
rect 575 316 607 350
rect 575 196 641 316
rect 675 162 709 458
rect 833 362 993 428
rect 911 202 945 362
rect 1043 294 1077 462
rect 1191 428 1271 476
rect 1111 394 1271 428
rect 1111 362 1225 394
rect 1043 260 1157 294
rect 434 17 500 162
rect 600 70 709 162
rect 743 17 777 202
rect 813 168 945 202
rect 813 70 879 168
rect 917 17 983 134
rect 1019 85 1069 226
rect 1107 119 1157 260
rect 1191 85 1225 362
rect 1310 382 1344 510
rect 1430 509 1673 543
rect 1430 476 1464 509
rect 1378 416 1464 476
rect 1740 475 1806 517
rect 1646 425 1806 475
rect 1586 382 1652 391
rect 1310 348 1652 382
rect 1310 337 1344 348
rect 1259 303 1344 337
rect 1586 329 1652 348
rect 1259 119 1293 303
rect 1441 295 1507 314
rect 1740 295 1806 425
rect 1847 358 1881 551
rect 1915 392 1981 649
rect 2089 431 2155 596
rect 2299 465 2456 649
rect 2089 397 2289 431
rect 2490 424 2540 569
rect 1847 324 2125 358
rect 1327 227 1377 269
rect 1441 261 1806 295
rect 2059 292 2125 324
rect 1327 193 1562 227
rect 1327 85 1377 193
rect 1019 51 1377 85
rect 1444 17 1494 159
rect 1528 85 1562 193
rect 1596 119 1630 261
rect 1840 258 2017 290
rect 2167 258 2221 360
rect 1840 227 2221 258
rect 1664 224 2221 227
rect 2255 297 2289 397
rect 2323 361 2540 424
rect 2708 364 2758 649
rect 2323 350 2497 361
rect 2323 345 2431 350
rect 2465 316 2497 350
rect 2255 231 2397 297
rect 1664 193 1874 224
rect 1664 85 1698 193
rect 2255 190 2289 231
rect 1528 51 1698 85
rect 1732 17 1782 154
rect 1908 124 2289 190
rect 2331 17 2397 197
rect 2431 85 2497 316
rect 2653 264 2795 330
rect 2653 85 2687 264
rect 2431 51 2687 85
rect 2721 17 2755 230
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2880 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 607 316 641 350
rect 2431 316 2465 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
<< metal1 >>
rect 0 683 2880 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2880 683
rect 0 617 2880 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 2880 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2880 17
rect 0 -49 2880 -17
<< obsm1 >>
rect 595 350 653 356
rect 595 316 607 350
rect 641 347 653 350
rect 2419 350 2477 356
rect 2419 347 2431 350
rect 641 319 2431 347
rect 641 316 653 319
rect 595 310 653 316
rect 2419 316 2431 319
rect 2465 316 2477 350
rect 2419 310 2477 316
<< labels >>
rlabel locali s 85 196 167 398 6 D
port 1 nsew signal input
rlabel locali s 313 290 381 356 6 DE
port 2 nsew signal input
rlabel locali s 2585 364 2668 596 6 Q
port 3 nsew signal output
rlabel locali s 2585 200 2619 364 6 Q
port 3 nsew signal output
rlabel locali s 2553 124 2619 200 6 Q
port 3 nsew signal output
rlabel locali s 2829 230 2863 364 6 Q_N
port 4 nsew signal output
rlabel locali s 2798 364 2863 596 6 Q_N
port 4 nsew signal output
rlabel locali s 2791 74 2863 230 6 Q_N
port 4 nsew signal output
rlabel locali s 743 236 877 310 6 CLK
port 5 nsew clock input
rlabel metal1 s 0 -49 2880 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 7 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 617 2880 715 6 VPWR
port 9 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2880 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 2393690
string GDS_START 2373356
<< end >>
