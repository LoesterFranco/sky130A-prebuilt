magic
tech sky130A
magscale 1 2
timestamp 1601050088
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 23 364 73 649
rect 113 424 177 599
rect 113 390 129 424
rect 163 390 177 424
rect 113 266 177 390
rect 211 388 269 649
rect 303 424 369 596
rect 303 390 319 424
rect 353 390 369 424
rect 303 388 369 390
rect 409 388 459 649
rect 493 424 559 596
rect 493 390 509 424
rect 543 390 559 424
rect 493 388 559 390
rect 599 388 649 649
rect 683 424 742 596
rect 683 390 699 424
rect 733 390 742 424
rect 214 350 276 354
rect 214 316 229 350
rect 263 316 276 350
rect 214 270 276 316
rect 123 226 177 266
rect 37 17 89 226
rect 123 70 189 226
rect 223 17 275 226
rect 311 70 369 388
rect 404 350 462 354
rect 404 316 417 350
rect 451 316 462 350
rect 404 270 462 316
rect 405 17 461 226
rect 497 70 559 388
rect 594 350 649 354
rect 594 316 605 350
rect 639 316 649 350
rect 594 270 649 316
rect 595 17 649 226
rect 683 70 742 390
rect 783 388 830 649
rect 868 424 926 596
rect 868 390 879 424
rect 913 390 926 424
rect 868 388 926 390
rect 962 388 1019 649
rect 1053 424 1116 596
rect 1053 390 1069 424
rect 1103 390 1116 424
rect 777 350 833 354
rect 777 316 788 350
rect 822 316 833 350
rect 777 270 833 316
rect 778 17 830 226
rect 868 70 919 388
rect 954 350 1017 354
rect 954 316 970 350
rect 1004 316 1017 350
rect 954 270 1017 316
rect 1053 257 1116 390
rect 1153 388 1219 649
rect 1253 424 1319 596
rect 1253 390 1269 424
rect 1303 390 1319 424
rect 1151 350 1218 354
rect 1151 316 1169 350
rect 1203 316 1218 350
rect 1151 270 1218 316
rect 1253 257 1319 390
rect 1353 388 1419 649
rect 1453 424 1509 596
rect 1453 390 1469 424
rect 1503 390 1509 424
rect 1354 350 1418 354
rect 1354 316 1368 350
rect 1402 316 1418 350
rect 1354 270 1418 316
rect 1053 236 1105 257
rect 1253 236 1305 257
rect 953 17 1005 226
rect 1043 70 1105 236
rect 1141 17 1205 226
rect 1239 70 1305 236
rect 1453 226 1509 390
rect 1547 364 1609 649
rect 1341 17 1409 226
rect 1443 70 1509 226
rect 1543 17 1609 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 129 390 163 424
rect 319 390 353 424
rect 509 390 543 424
rect 699 390 733 424
rect 229 316 263 350
rect 417 316 451 350
rect 605 316 639 350
rect 879 390 913 424
rect 1069 390 1103 424
rect 788 316 822 350
rect 970 316 1004 350
rect 1269 390 1303 424
rect 1169 316 1203 350
rect 1469 390 1503 424
rect 1368 316 1402 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 117 424 1515 430
rect 117 390 129 424
rect 163 390 319 424
rect 353 390 509 424
rect 543 390 699 424
rect 733 390 879 424
rect 913 390 1069 424
rect 1103 390 1269 424
rect 1303 390 1469 424
rect 1503 390 1515 424
rect 117 384 1515 390
rect 217 350 1414 356
rect 217 316 229 350
rect 263 316 417 350
rect 451 316 605 350
rect 639 316 788 350
rect 822 316 970 350
rect 1004 316 1169 350
rect 1203 316 1368 350
rect 1402 316 1414 350
rect 217 310 1414 316
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
rlabel metal1 s 217 310 1414 356 6 A
port 1 nsew signal input
rlabel metal1 s 117 384 1515 430 6 Y
port 2 nsew signal output
rlabel metal1 s 0 -49 1632 49 8 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 617 1632 715 6 VPWR
port 4 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1803336
string GDS_START 1789728
<< end >>
