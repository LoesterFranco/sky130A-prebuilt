magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 655 357 707 493
rect 17 215 125 255
rect 163 215 257 257
rect 213 135 257 215
rect 305 213 417 257
rect 305 135 349 213
rect 455 196 525 257
rect 673 117 707 357
rect 655 51 707 117
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 18 449 85 493
rect 308 451 379 527
rect 18 343 69 449
rect 413 417 479 493
rect 113 377 479 417
rect 517 387 583 527
rect 18 299 607 343
rect 18 17 119 170
rect 573 157 607 299
rect 422 123 607 157
rect 422 93 456 123
rect 174 51 456 93
rect 517 17 583 89
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel locali s 305 213 417 257 6 A1
port 1 nsew signal input
rlabel locali s 305 135 349 213 6 A1
port 1 nsew signal input
rlabel locali s 455 196 525 257 6 A2
port 2 nsew signal input
rlabel locali s 213 135 257 215 6 B1
port 3 nsew signal input
rlabel locali s 163 215 257 257 6 B1
port 3 nsew signal input
rlabel locali s 17 215 125 255 6 B2
port 4 nsew signal input
rlabel locali s 673 117 707 357 6 X
port 5 nsew signal output
rlabel locali s 655 357 707 493 6 X
port 5 nsew signal output
rlabel locali s 655 51 707 117 6 X
port 5 nsew signal output
rlabel metal1 s 0 -48 736 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 736 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1259064
string GDS_START 1252572
<< end >>
