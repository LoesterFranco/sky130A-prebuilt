magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 806 704
<< pwell >>
rect 0 0 768 49
<< scnmos >>
rect 158 85 358 169
rect 413 85 613 169
<< pmoshvt >>
rect 160 392 360 592
rect 415 392 615 592
<< ndiff >>
rect 42 145 158 169
rect 42 111 113 145
rect 147 111 158 145
rect 42 85 158 111
rect 358 145 413 169
rect 358 111 369 145
rect 403 111 413 145
rect 358 85 413 111
rect 613 145 741 169
rect 613 111 624 145
rect 658 111 741 145
rect 613 85 741 111
<< pdiff >>
rect 27 580 160 592
rect 27 546 113 580
rect 147 546 160 580
rect 27 509 160 546
rect 27 475 113 509
rect 147 475 160 509
rect 27 392 160 475
rect 360 580 415 592
rect 360 546 371 580
rect 405 546 415 580
rect 360 509 415 546
rect 360 475 371 509
rect 405 475 415 509
rect 360 438 415 475
rect 360 404 371 438
rect 405 404 415 438
rect 360 392 415 404
rect 615 580 741 592
rect 615 546 626 580
rect 660 546 741 580
rect 615 509 741 546
rect 615 475 626 509
rect 660 475 741 509
rect 615 392 741 475
<< ndiffc >>
rect 113 111 147 145
rect 369 111 403 145
rect 624 111 658 145
<< pdiffc >>
rect 113 546 147 580
rect 113 475 147 509
rect 371 546 405 580
rect 371 475 405 509
rect 371 404 405 438
rect 626 546 660 580
rect 626 475 660 509
<< poly >>
rect 160 592 360 618
rect 415 592 615 618
rect 160 366 360 392
rect 415 366 615 392
rect 160 301 226 366
rect 160 267 176 301
rect 210 267 226 301
rect 160 251 226 267
rect 292 300 479 316
rect 292 266 308 300
rect 342 266 429 300
rect 463 266 479 300
rect 292 238 479 266
rect 549 301 615 366
rect 549 267 565 301
rect 599 267 615 301
rect 549 251 615 267
rect 292 209 358 238
rect 158 169 358 209
rect 413 209 479 238
rect 413 169 613 209
rect 158 47 358 85
rect 413 47 613 85
<< polycont >>
rect 176 267 210 301
rect 308 266 342 300
rect 429 266 463 300
rect 565 267 599 301
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 113 580 163 649
rect 147 546 163 580
rect 113 509 163 546
rect 147 475 163 509
rect 113 457 163 475
rect 292 580 479 649
rect 292 546 371 580
rect 405 546 479 580
rect 292 509 479 546
rect 292 475 371 509
rect 405 475 479 509
rect 292 438 479 475
rect 610 580 660 649
rect 610 546 626 580
rect 610 509 660 546
rect 610 475 626 509
rect 610 459 660 475
rect 292 404 371 438
rect 405 404 479 438
rect 160 301 226 317
rect 160 267 176 301
rect 210 267 226 301
rect 160 162 226 267
rect 292 300 479 404
rect 292 266 308 300
rect 342 266 429 300
rect 463 266 479 300
rect 292 250 479 266
rect 534 301 615 317
rect 534 267 565 301
rect 599 267 615 301
rect 113 145 226 162
rect 534 162 615 267
rect 147 111 226 145
rect 113 17 226 111
rect 353 145 419 161
rect 353 111 369 145
rect 403 111 419 145
rect 353 17 419 111
rect 534 145 658 162
rect 534 111 624 145
rect 534 17 658 111
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel comment s 0 0 0 0 4 decap_8
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 2 nsew
flabel nbase s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 3 nsew
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 1 nsew
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 768 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3437810
string GDS_START 3433956
<< end >>
