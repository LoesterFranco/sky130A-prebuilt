magic
tech sky130A
magscale 1 2
timestamp 1604502741
<< locali >>
rect 18 378 78 613
rect 18 53 78 288
<< obsli1 >>
rect 0 649 31 683
rect 65 649 96 683
rect 0 -17 31 17
rect 65 -17 96 17
<< obsli1c >>
rect 31 649 65 683
rect 31 -17 65 17
<< metal1 >>
rect 0 683 96 715
rect 0 649 31 683
rect 65 649 96 683
rect 0 617 96 649
rect 0 17 96 49
rect 0 -17 31 17
rect 65 -17 96 17
rect 0 -49 96 -17
<< labels >>
rlabel metal1 s 0 -49 96 49 8 VGND
port 1 nsew ground bidirectional
rlabel locali s 18 53 78 288 6 VNB
port 2 nsew ground bidirectional
rlabel locali s 18 378 78 613 6 VPB
port 3 nsew power bidirectional
rlabel metal1 s 0 617 96 715 6 VPWR
port 4 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE WELLTAP
string FIXED_BBOX 0 0 96 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 469724
string GDS_START 467024
<< end >>
