magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 460 561
rect 108 447 174 527
rect 17 191 102 345
rect 208 357 443 493
rect 324 119 360 357
rect 394 153 443 323
rect 108 17 288 89
rect 324 51 443 119
rect 0 -17 460 17
<< obsli1 >>
rect 17 413 74 493
rect 17 379 174 413
rect 137 323 174 379
rect 137 157 290 323
rect 17 123 290 157
rect 17 51 74 123
<< metal1 >>
rect 0 496 460 592
rect 0 -48 460 48
<< labels >>
rlabel locali s 394 153 443 323 6 A
port 1 nsew signal input
rlabel locali s 17 191 102 345 6 TE_B
port 2 nsew signal input
rlabel locali s 324 119 360 357 6 Z
port 3 nsew signal output
rlabel locali s 324 51 443 119 6 Z
port 3 nsew signal output
rlabel locali s 208 357 443 493 6 Z
port 3 nsew signal output
rlabel locali s 108 17 288 89 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 460 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 460 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 108 447 174 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 460 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 460 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 460 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2893796
string GDS_START 2888730
<< end >>
