magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 111 364 183 596
rect 111 226 145 364
rect 293 236 359 310
rect 111 70 179 226
rect 461 249 595 356
rect 643 326 743 356
rect 643 260 907 326
rect 643 249 743 260
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 27 364 77 649
rect 217 424 356 649
rect 393 424 557 551
rect 697 458 763 649
rect 871 424 937 572
rect 393 390 937 424
rect 217 356 427 390
rect 871 364 937 390
rect 217 330 251 356
rect 179 264 251 330
rect 27 17 77 226
rect 393 215 427 356
rect 866 215 932 226
rect 215 17 359 202
rect 393 181 932 215
rect 393 70 552 181
rect 668 17 768 136
rect 866 70 932 181
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
rlabel locali s 293 236 359 310 6 A
port 1 nsew signal input
rlabel locali s 461 249 595 356 6 B
port 2 nsew signal input
rlabel locali s 643 326 743 356 6 C
port 3 nsew signal input
rlabel locali s 643 260 907 326 6 C
port 3 nsew signal input
rlabel locali s 643 249 743 260 6 C
port 3 nsew signal input
rlabel locali s 111 364 183 596 6 X
port 4 nsew signal output
rlabel locali s 111 226 145 364 6 X
port 4 nsew signal output
rlabel locali s 111 70 179 226 6 X
port 4 nsew signal output
rlabel metal1 s 0 -49 960 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 617 960 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1883740
string GDS_START 1875916
<< end >>
