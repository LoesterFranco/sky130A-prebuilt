magic
tech sky130A
magscale 1 2
timestamp 1599588244
<< locali >>
rect 217 492 313 596
rect 217 458 451 492
rect 21 260 167 356
rect 203 270 269 356
rect 417 226 451 458
rect 371 70 451 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 23 424 89 540
rect 130 458 183 649
rect 347 530 414 649
rect 23 390 337 424
rect 303 326 337 390
rect 303 260 383 326
rect 303 226 337 260
rect 23 192 337 226
rect 23 108 76 192
rect 110 17 244 158
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< metal1 >>
rect 0 683 480 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 0 617 480 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 480 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
rect 0 -49 480 -17
<< labels >>
rlabel locali s 21 260 167 356 6 A_N
port 1 nsew signal input
rlabel locali s 203 270 269 356 6 B
port 2 nsew signal input
rlabel locali s 417 226 451 458 6 Y
port 3 nsew signal output
rlabel locali s 371 70 451 226 6 Y
port 3 nsew signal output
rlabel locali s 217 492 313 596 6 Y
port 3 nsew signal output
rlabel locali s 217 458 451 492 6 Y
port 3 nsew signal output
rlabel metal1 s 0 -49 480 49 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 5 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 617 480 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 480 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 2008040
string GDS_START 2003424
<< end >>
