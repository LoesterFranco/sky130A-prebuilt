magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 17 215 85 328
rect 202 283 484 340
rect 202 181 254 283
rect 202 147 448 181
rect 202 57 286 147
rect 401 51 448 147
rect 560 199 622 340
rect 666 199 714 340
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 17 408 69 444
rect 120 442 192 527
rect 304 442 380 527
rect 491 442 569 527
rect 774 442 891 485
rect 17 374 806 408
rect 17 362 163 374
rect 129 181 163 362
rect 17 147 163 181
rect 288 215 523 249
rect 17 58 69 147
rect 134 17 168 113
rect 330 17 364 113
rect 489 165 523 215
rect 772 199 806 374
rect 850 165 891 442
rect 489 131 891 165
rect 492 17 568 97
rect 680 17 768 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
rlabel locali s 560 199 622 340 6 A
port 1 nsew signal input
rlabel locali s 666 199 714 340 6 B
port 2 nsew signal input
rlabel locali s 17 215 85 328 6 C_N
port 3 nsew signal input
rlabel locali s 401 51 448 147 6 X
port 4 nsew signal output
rlabel locali s 202 283 484 340 6 X
port 4 nsew signal output
rlabel locali s 202 181 254 283 6 X
port 4 nsew signal output
rlabel locali s 202 147 448 181 6 X
port 4 nsew signal output
rlabel locali s 202 57 286 147 6 X
port 4 nsew signal output
rlabel metal1 s 0 -48 920 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 920 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 920 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 491918
string GDS_START 485228
<< end >>
