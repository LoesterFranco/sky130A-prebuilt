magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 998 704
<< pwell >>
rect 0 0 960 49
<< scnmos >>
rect 91 74 121 222
rect 177 74 207 222
rect 263 74 293 222
rect 357 74 387 222
rect 553 74 583 222
rect 727 74 757 222
<< pmoshvt >>
rect 84 368 114 592
rect 174 368 204 592
rect 264 368 294 592
rect 354 368 384 592
rect 556 368 586 592
rect 646 368 676 592
rect 736 368 766 592
rect 826 368 856 592
<< ndiff >>
rect 38 202 91 222
rect 38 168 46 202
rect 80 168 91 202
rect 38 124 91 168
rect 38 90 46 124
rect 80 90 91 124
rect 38 74 91 90
rect 121 177 177 222
rect 121 143 132 177
rect 166 143 177 177
rect 121 74 177 143
rect 207 184 263 222
rect 207 150 218 184
rect 252 150 263 184
rect 207 116 263 150
rect 207 82 218 116
rect 252 82 263 116
rect 207 74 263 82
rect 293 116 357 222
rect 293 82 308 116
rect 342 82 357 116
rect 293 74 357 82
rect 387 184 446 222
rect 387 150 398 184
rect 432 150 446 184
rect 387 116 446 150
rect 387 82 398 116
rect 432 82 446 116
rect 387 74 446 82
rect 500 127 553 222
rect 500 93 508 127
rect 542 93 553 127
rect 500 74 553 93
rect 583 202 727 222
rect 583 168 594 202
rect 628 168 668 202
rect 702 168 727 202
rect 583 116 727 168
rect 583 82 594 116
rect 628 82 668 116
rect 702 82 727 116
rect 583 74 727 82
rect 757 194 814 222
rect 757 160 768 194
rect 802 160 814 194
rect 757 120 814 160
rect 757 86 768 120
rect 802 86 814 120
rect 757 74 814 86
<< pdiff >>
rect 29 580 84 592
rect 29 546 37 580
rect 71 546 84 580
rect 29 497 84 546
rect 29 463 37 497
rect 71 463 84 497
rect 29 414 84 463
rect 29 380 37 414
rect 71 380 84 414
rect 29 368 84 380
rect 114 580 174 592
rect 114 546 127 580
rect 161 546 174 580
rect 114 497 174 546
rect 114 463 127 497
rect 161 463 174 497
rect 114 414 174 463
rect 114 380 127 414
rect 161 380 174 414
rect 114 368 174 380
rect 204 580 264 592
rect 204 546 217 580
rect 251 546 264 580
rect 204 492 264 546
rect 204 458 217 492
rect 251 458 264 492
rect 204 368 264 458
rect 294 580 354 592
rect 294 546 307 580
rect 341 546 354 580
rect 294 505 354 546
rect 294 471 307 505
rect 341 471 354 505
rect 294 424 354 471
rect 294 390 307 424
rect 341 390 354 424
rect 294 368 354 390
rect 384 582 443 592
rect 384 548 397 582
rect 431 548 443 582
rect 384 514 443 548
rect 384 480 397 514
rect 431 480 443 514
rect 384 368 443 480
rect 497 582 556 592
rect 497 548 509 582
rect 543 548 556 582
rect 497 514 556 548
rect 497 480 509 514
rect 543 480 556 514
rect 497 368 556 480
rect 586 531 646 592
rect 586 497 599 531
rect 633 497 646 531
rect 586 446 646 497
rect 586 412 599 446
rect 633 412 646 446
rect 586 368 646 412
rect 676 580 736 592
rect 676 546 689 580
rect 723 546 736 580
rect 676 462 736 546
rect 676 428 689 462
rect 723 428 736 462
rect 676 368 736 428
rect 766 547 826 592
rect 766 513 779 547
rect 813 513 826 547
rect 766 479 826 513
rect 766 445 779 479
rect 813 445 826 479
rect 766 411 826 445
rect 766 377 779 411
rect 813 377 826 411
rect 766 368 826 377
rect 856 580 911 592
rect 856 546 869 580
rect 903 546 911 580
rect 856 497 911 546
rect 856 463 869 497
rect 903 463 911 497
rect 856 414 911 463
rect 856 380 869 414
rect 903 380 911 414
rect 856 368 911 380
<< ndiffc >>
rect 46 168 80 202
rect 46 90 80 124
rect 132 143 166 177
rect 218 150 252 184
rect 218 82 252 116
rect 308 82 342 116
rect 398 150 432 184
rect 398 82 432 116
rect 508 93 542 127
rect 594 168 628 202
rect 668 168 702 202
rect 594 82 628 116
rect 668 82 702 116
rect 768 160 802 194
rect 768 86 802 120
<< pdiffc >>
rect 37 546 71 580
rect 37 463 71 497
rect 37 380 71 414
rect 127 546 161 580
rect 127 463 161 497
rect 127 380 161 414
rect 217 546 251 580
rect 217 458 251 492
rect 307 546 341 580
rect 307 471 341 505
rect 307 390 341 424
rect 397 548 431 582
rect 397 480 431 514
rect 509 548 543 582
rect 509 480 543 514
rect 599 497 633 531
rect 599 412 633 446
rect 689 546 723 580
rect 689 428 723 462
rect 779 513 813 547
rect 779 445 813 479
rect 779 377 813 411
rect 869 546 903 580
rect 869 463 903 497
rect 869 380 903 414
<< poly >>
rect 84 592 114 618
rect 174 592 204 618
rect 264 592 294 618
rect 354 592 384 618
rect 556 592 586 618
rect 646 592 676 618
rect 736 592 766 618
rect 826 592 856 618
rect 84 353 114 368
rect 174 353 204 368
rect 264 353 294 368
rect 354 353 384 368
rect 556 353 586 368
rect 646 353 676 368
rect 736 353 766 368
rect 826 353 856 368
rect 81 310 117 353
rect 171 310 207 353
rect 261 336 297 353
rect 351 336 387 353
rect 32 294 207 310
rect 32 260 48 294
rect 82 260 207 294
rect 249 320 387 336
rect 249 286 265 320
rect 299 286 337 320
rect 371 286 387 320
rect 249 270 387 286
rect 32 244 207 260
rect 91 222 121 244
rect 177 222 207 244
rect 263 222 293 270
rect 357 222 387 270
rect 553 310 589 353
rect 643 310 679 353
rect 733 310 769 353
rect 823 310 859 353
rect 553 294 685 310
rect 553 260 635 294
rect 669 260 685 294
rect 553 244 685 260
rect 727 294 859 310
rect 727 260 809 294
rect 843 260 859 294
rect 727 244 859 260
rect 553 222 583 244
rect 727 222 757 244
rect 91 48 121 74
rect 177 48 207 74
rect 263 48 293 74
rect 357 48 387 74
rect 553 48 583 74
rect 727 48 757 74
<< polycont >>
rect 48 260 82 294
rect 265 286 299 320
rect 337 286 371 320
rect 635 260 669 294
rect 809 260 843 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 21 580 71 649
rect 21 546 37 580
rect 21 497 71 546
rect 21 463 37 497
rect 21 414 71 463
rect 21 380 37 414
rect 21 364 71 380
rect 111 580 161 596
rect 111 546 127 580
rect 111 497 161 546
rect 111 463 127 497
rect 111 424 161 463
rect 201 580 267 649
rect 201 546 217 580
rect 251 546 267 580
rect 201 492 267 546
rect 201 458 217 492
rect 251 458 267 492
rect 307 580 341 596
rect 307 505 341 546
rect 381 582 447 649
rect 381 548 397 582
rect 431 548 447 582
rect 381 514 447 548
rect 381 480 397 514
rect 431 480 447 514
rect 493 582 919 615
rect 493 548 509 582
rect 543 581 919 582
rect 543 548 559 581
rect 493 514 559 548
rect 689 580 723 581
rect 493 480 509 514
rect 543 480 559 514
rect 593 531 649 547
rect 593 497 599 531
rect 633 497 649 531
rect 307 446 341 471
rect 593 446 649 497
rect 307 424 599 446
rect 111 414 307 424
rect 111 380 127 414
rect 161 390 307 414
rect 341 412 599 424
rect 633 412 649 446
rect 869 580 919 581
rect 689 462 723 546
rect 689 412 723 428
rect 763 513 779 547
rect 813 513 829 547
rect 763 479 829 513
rect 763 445 779 479
rect 813 445 829 479
rect 341 390 471 412
rect 763 411 829 445
rect 111 364 161 380
rect 763 378 779 411
rect 505 377 779 378
rect 813 377 829 411
rect 217 320 455 356
rect 25 294 96 310
rect 25 260 48 294
rect 82 260 96 294
rect 217 286 265 320
rect 299 286 337 320
rect 371 286 455 320
rect 505 344 829 377
rect 903 546 919 580
rect 869 497 919 546
rect 903 463 919 497
rect 869 414 919 463
rect 903 380 919 414
rect 869 364 919 380
rect 25 236 96 260
rect 505 252 551 344
rect 130 218 551 252
rect 601 294 743 310
rect 601 260 635 294
rect 669 260 743 294
rect 601 236 743 260
rect 793 294 935 310
rect 793 260 809 294
rect 843 260 935 294
rect 793 236 935 260
rect 30 168 46 202
rect 80 168 96 202
rect 30 124 96 168
rect 130 177 166 218
rect 517 202 551 218
rect 130 143 132 177
rect 130 127 166 143
rect 202 150 218 184
rect 252 150 398 184
rect 432 150 448 184
rect 517 168 594 202
rect 628 168 668 202
rect 702 168 718 202
rect 30 90 46 124
rect 80 90 96 124
rect 30 85 96 90
rect 202 116 252 150
rect 398 116 448 150
rect 202 85 218 116
rect 30 82 218 85
rect 30 51 252 82
rect 288 82 308 116
rect 342 82 362 116
rect 288 66 362 82
rect 432 82 448 116
rect 398 66 448 82
rect 492 127 558 134
rect 492 93 508 127
rect 542 93 558 127
rect 288 17 322 66
rect 492 17 558 93
rect 592 116 718 168
rect 592 82 594 116
rect 628 82 668 116
rect 702 82 718 116
rect 592 66 718 82
rect 752 194 818 202
rect 752 160 768 194
rect 802 160 818 194
rect 752 120 818 160
rect 752 86 768 120
rect 802 86 818 120
rect 752 17 818 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a211oi_2
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 511 242 545 276 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 799 242 833 276 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 895 242 929 276 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 607 242 641 276 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 703 242 737 276 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 A1
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 960 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3965440
string GDS_START 3956502
<< end >>
