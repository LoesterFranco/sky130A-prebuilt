magic
tech sky130A
magscale 1 2
timestamp 1601050047
<< nwell >>
rect -38 332 710 704
<< pwell >>
rect 0 0 672 49
<< scpmos >>
rect 86 368 116 536
rect 193 368 223 592
rect 326 368 356 592
rect 440 368 470 568
rect 524 368 554 568
<< nmoslvt >>
rect 85 112 115 222
rect 187 74 217 222
rect 274 74 304 222
rect 443 74 473 202
rect 542 74 572 202
<< ndiff >>
rect 28 184 85 222
rect 28 150 40 184
rect 74 150 85 184
rect 28 112 85 150
rect 115 152 187 222
rect 115 118 142 152
rect 176 118 187 152
rect 115 112 187 118
rect 130 74 187 112
rect 217 210 274 222
rect 217 176 228 210
rect 262 176 274 210
rect 217 120 274 176
rect 217 86 228 120
rect 262 86 274 120
rect 217 74 274 86
rect 304 202 354 222
rect 304 146 443 202
rect 304 112 315 146
rect 349 112 397 146
rect 431 112 443 146
rect 304 74 443 112
rect 473 190 542 202
rect 473 156 497 190
rect 531 156 542 190
rect 473 120 542 156
rect 473 86 497 120
rect 531 86 542 120
rect 473 74 542 86
rect 572 146 645 202
rect 572 112 583 146
rect 617 112 645 146
rect 572 74 645 112
<< pdiff >>
rect 134 573 193 592
rect 134 539 146 573
rect 180 539 193 573
rect 134 536 193 539
rect 27 524 86 536
rect 27 490 39 524
rect 73 490 86 524
rect 27 440 86 490
rect 27 406 39 440
rect 73 406 86 440
rect 27 368 86 406
rect 116 368 193 536
rect 223 414 326 592
rect 223 380 257 414
rect 291 380 326 414
rect 223 368 326 380
rect 356 573 415 592
rect 356 539 369 573
rect 403 568 415 573
rect 403 539 440 568
rect 356 368 440 539
rect 470 368 524 568
rect 554 556 637 568
rect 554 522 591 556
rect 625 522 637 556
rect 554 485 637 522
rect 554 451 591 485
rect 625 451 637 485
rect 554 414 637 451
rect 554 380 591 414
rect 625 380 637 414
rect 554 368 637 380
<< ndiffc >>
rect 40 150 74 184
rect 142 118 176 152
rect 228 176 262 210
rect 228 86 262 120
rect 315 112 349 146
rect 397 112 431 146
rect 497 156 531 190
rect 497 86 531 120
rect 583 112 617 146
<< pdiffc >>
rect 146 539 180 573
rect 39 490 73 524
rect 39 406 73 440
rect 257 380 291 414
rect 369 539 403 573
rect 591 522 625 556
rect 591 451 625 485
rect 591 380 625 414
<< poly >>
rect 193 592 223 618
rect 326 592 356 618
rect 86 536 116 562
rect 440 568 470 594
rect 524 568 554 594
rect 86 353 116 368
rect 193 353 223 368
rect 326 353 356 368
rect 440 353 470 368
rect 524 353 554 368
rect 83 336 119 353
rect 44 320 119 336
rect 44 286 60 320
rect 94 286 119 320
rect 190 326 226 353
rect 323 326 359 353
rect 437 336 473 353
rect 190 310 359 326
rect 190 290 309 310
rect 44 270 119 286
rect 187 276 309 290
rect 343 276 359 310
rect 85 222 115 270
rect 187 260 359 276
rect 407 320 473 336
rect 407 286 423 320
rect 457 286 473 320
rect 407 270 473 286
rect 187 222 217 260
rect 274 222 304 260
rect 85 86 115 112
rect 443 202 473 270
rect 521 330 557 353
rect 521 314 587 330
rect 521 280 537 314
rect 571 280 587 314
rect 521 264 587 280
rect 542 202 572 264
rect 187 48 217 74
rect 274 48 304 74
rect 443 48 473 74
rect 542 48 572 74
<< polycont >>
rect 60 286 94 320
rect 309 276 343 310
rect 423 286 457 320
rect 537 280 571 314
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 130 573 196 649
rect 23 524 89 540
rect 23 490 39 524
rect 73 490 89 524
rect 130 539 146 573
rect 180 539 196 573
rect 130 516 196 539
rect 353 573 419 649
rect 353 539 369 573
rect 403 539 419 573
rect 353 516 419 539
rect 575 556 655 572
rect 575 522 591 556
rect 625 522 655 556
rect 23 482 89 490
rect 575 485 655 522
rect 23 448 541 482
rect 23 440 178 448
rect 23 406 39 440
rect 73 406 178 440
rect 23 390 178 406
rect 25 320 110 356
rect 25 286 60 320
rect 94 286 110 320
rect 25 270 110 286
rect 144 236 178 390
rect 24 202 178 236
rect 212 380 257 414
rect 291 380 329 414
rect 212 364 329 380
rect 212 226 246 364
rect 293 310 359 326
rect 293 276 309 310
rect 343 276 359 310
rect 293 260 359 276
rect 407 320 473 356
rect 407 286 423 320
rect 457 286 473 320
rect 407 270 473 286
rect 507 330 541 448
rect 575 451 591 485
rect 625 451 655 485
rect 575 414 655 451
rect 575 380 591 414
rect 625 380 655 414
rect 575 364 655 380
rect 507 314 587 330
rect 507 280 537 314
rect 571 280 587 314
rect 507 264 587 280
rect 325 230 359 260
rect 621 230 655 364
rect 212 210 278 226
rect 24 184 90 202
rect 24 150 40 184
rect 74 150 90 184
rect 212 176 228 210
rect 262 176 278 210
rect 325 196 655 230
rect 24 108 90 150
rect 126 152 176 168
rect 126 118 142 152
rect 126 17 176 118
rect 212 120 278 176
rect 481 190 547 196
rect 212 86 228 120
rect 262 86 278 120
rect 212 70 278 86
rect 312 146 447 162
rect 312 112 315 146
rect 349 112 397 146
rect 431 112 447 146
rect 312 17 447 112
rect 481 156 497 190
rect 531 156 547 190
rect 481 120 547 156
rect 481 86 497 120
rect 531 86 547 120
rect 481 70 547 86
rect 583 146 649 162
rect 617 112 649 146
rect 583 17 649 112
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel comment s 0 0 0 0 4 or2b_2
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 223 94 257 128 0 FreeSans 340 0 0 0 X
port 7 nsew
flabel corelocali s 223 168 257 202 0 FreeSans 340 0 0 0 X
port 7 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 B_N
port 2 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 672 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 785978
string GDS_START 780324
<< end >>
