magic
tech sky130A
magscale 1 2
timestamp 1601050082
<< locali >>
rect 555 424 621 596
rect 133 390 621 424
rect 25 236 99 356
rect 133 236 167 390
rect 201 270 267 356
rect 309 270 375 356
rect 409 270 551 356
rect 585 270 651 356
rect 133 202 616 236
rect 217 70 408 202
rect 550 70 616 202
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 63 458 113 649
rect 153 492 219 596
rect 253 526 335 649
rect 369 492 435 596
rect 153 458 435 492
rect 68 17 134 168
rect 442 17 516 168
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel locali s 309 270 375 356 6 A1
port 1 nsew signal input
rlabel locali s 201 270 267 356 6 A2
port 2 nsew signal input
rlabel locali s 25 236 99 356 6 A3
port 3 nsew signal input
rlabel locali s 409 270 551 356 6 B1
port 4 nsew signal input
rlabel locali s 585 270 651 356 6 C1
port 5 nsew signal input
rlabel locali s 555 424 621 596 6 Y
port 6 nsew signal output
rlabel locali s 550 70 616 202 6 Y
port 6 nsew signal output
rlabel locali s 217 70 408 202 6 Y
port 6 nsew signal output
rlabel locali s 133 390 621 424 6 Y
port 6 nsew signal output
rlabel locali s 133 236 167 390 6 Y
port 6 nsew signal output
rlabel locali s 133 202 616 236 6 Y
port 6 nsew signal output
rlabel metal1 s 0 -49 672 49 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 617 672 715 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3582166
string GDS_START 3575678
<< end >>
