magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 19 459 275 493
rect 19 323 85 459
rect 207 439 275 459
rect 19 289 627 323
rect 25 153 125 255
rect 163 215 263 255
rect 213 135 263 215
rect 305 211 417 255
rect 305 135 347 211
rect 453 199 525 255
rect 559 165 627 289
rect 419 131 627 165
rect 419 101 455 131
rect 174 51 455 101
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 311 451 382 527
rect 129 396 163 423
rect 421 396 455 433
rect 129 357 455 396
rect 512 371 565 527
rect 19 17 119 119
rect 501 17 567 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 305 211 417 255 6 A1
port 1 nsew signal input
rlabel locali s 305 135 347 211 6 A1
port 1 nsew signal input
rlabel locali s 453 199 525 255 6 A2
port 2 nsew signal input
rlabel locali s 213 135 263 215 6 B1
port 3 nsew signal input
rlabel locali s 163 215 263 255 6 B1
port 3 nsew signal input
rlabel locali s 25 153 125 255 6 B2
port 4 nsew signal input
rlabel locali s 559 165 627 289 6 Y
port 5 nsew signal output
rlabel locali s 419 131 627 165 6 Y
port 5 nsew signal output
rlabel locali s 419 101 455 131 6 Y
port 5 nsew signal output
rlabel locali s 207 439 275 459 6 Y
port 5 nsew signal output
rlabel locali s 174 51 455 101 6 Y
port 5 nsew signal output
rlabel locali s 19 459 275 493 6 Y
port 5 nsew signal output
rlabel locali s 19 323 85 459 6 Y
port 5 nsew signal output
rlabel locali s 19 289 627 323 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -48 644 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1282794
string GDS_START 1276988
<< end >>
