magic
tech sky130A
magscale 1 2
timestamp 1601050056
<< nwell >>
rect -38 332 1670 704
rect 768 312 1178 332
<< pwell >>
rect 0 0 1632 49
<< scpmos >>
rect 81 424 117 592
rect 159 424 195 592
rect 372 368 408 536
rect 570 379 606 547
rect 675 451 711 535
rect 753 451 789 535
rect 858 356 894 580
rect 1056 348 1092 516
rect 1162 374 1198 574
rect 1295 374 1331 574
rect 1412 368 1448 592
rect 1502 368 1538 592
<< nmoslvt >>
rect 84 112 114 222
rect 170 112 200 222
rect 288 74 318 222
rect 550 74 580 184
rect 655 81 685 165
rect 733 81 763 165
rect 869 81 899 229
rect 1067 74 1097 222
rect 1168 74 1198 222
rect 1240 74 1270 222
rect 1434 74 1464 222
rect 1520 74 1550 222
<< ndiff >>
rect 27 183 84 222
rect 27 149 39 183
rect 73 149 84 183
rect 27 112 84 149
rect 114 183 170 222
rect 114 149 125 183
rect 159 149 170 183
rect 114 112 170 149
rect 200 112 288 222
rect 215 74 288 112
rect 318 210 375 222
rect 318 176 329 210
rect 363 176 375 210
rect 318 74 375 176
rect 429 123 550 184
rect 429 89 441 123
rect 475 89 550 123
rect 429 74 550 89
rect 580 165 640 184
rect 819 165 869 229
rect 580 153 655 165
rect 580 119 593 153
rect 627 119 655 153
rect 580 81 655 119
rect 685 81 733 165
rect 763 129 869 165
rect 763 95 774 129
rect 808 95 869 129
rect 763 81 869 95
rect 899 184 956 229
rect 899 150 910 184
rect 944 150 956 184
rect 899 81 956 150
rect 1010 202 1067 222
rect 1010 168 1022 202
rect 1056 168 1067 202
rect 1010 120 1067 168
rect 1010 86 1022 120
rect 1056 86 1067 120
rect 580 74 630 81
rect 215 40 227 74
rect 261 40 273 74
rect 1010 74 1067 86
rect 1097 202 1168 222
rect 1097 168 1122 202
rect 1156 168 1168 202
rect 1097 120 1168 168
rect 1097 86 1122 120
rect 1156 86 1168 120
rect 1097 74 1168 86
rect 1198 74 1240 222
rect 1270 210 1325 222
rect 1270 176 1281 210
rect 1315 176 1325 210
rect 1270 120 1325 176
rect 1270 86 1281 120
rect 1315 86 1325 120
rect 1270 74 1325 86
rect 1379 131 1434 222
rect 1379 97 1389 131
rect 1423 97 1434 131
rect 1379 74 1434 97
rect 1464 210 1520 222
rect 1464 176 1475 210
rect 1509 176 1520 210
rect 1464 120 1520 176
rect 1464 86 1475 120
rect 1509 86 1520 120
rect 1464 74 1520 86
rect 1550 210 1605 222
rect 1550 176 1561 210
rect 1595 176 1605 210
rect 1550 120 1605 176
rect 1550 86 1561 120
rect 1595 86 1605 120
rect 1550 74 1605 86
rect 215 28 273 40
<< pdiff >>
rect 27 580 81 592
rect 27 546 37 580
rect 71 546 81 580
rect 27 476 81 546
rect 27 442 37 476
rect 71 442 81 476
rect 27 424 81 442
rect 117 424 159 592
rect 195 580 249 592
rect 195 546 205 580
rect 239 546 249 580
rect 195 498 249 546
rect 195 464 205 498
rect 239 464 249 498
rect 195 424 249 464
rect 303 582 357 594
rect 303 548 313 582
rect 347 548 357 582
rect 303 536 357 548
rect 303 368 372 536
rect 408 414 462 536
rect 408 380 418 414
rect 452 380 462 414
rect 408 368 462 380
rect 516 535 570 547
rect 516 501 526 535
rect 560 501 570 535
rect 516 427 570 501
rect 516 393 526 427
rect 560 393 570 427
rect 516 379 570 393
rect 606 535 660 547
rect 804 568 858 580
rect 804 535 814 568
rect 606 510 675 535
rect 606 476 616 510
rect 650 476 675 510
rect 606 451 675 476
rect 711 451 753 535
rect 789 534 814 535
rect 848 534 858 568
rect 789 469 858 534
rect 789 451 814 469
rect 606 379 660 451
rect 804 435 814 451
rect 848 435 858 469
rect 804 356 858 435
rect 894 568 948 580
rect 1346 580 1412 592
rect 1346 574 1358 580
rect 894 534 904 568
rect 938 534 948 568
rect 1107 562 1162 574
rect 894 485 948 534
rect 1107 528 1118 562
rect 1152 528 1162 562
rect 1107 516 1162 528
rect 894 451 904 485
rect 938 451 948 485
rect 894 402 948 451
rect 894 368 904 402
rect 938 368 948 402
rect 894 356 948 368
rect 1002 394 1056 516
rect 1002 360 1012 394
rect 1046 360 1056 394
rect 1002 348 1056 360
rect 1092 374 1162 516
rect 1198 562 1295 574
rect 1198 528 1251 562
rect 1285 528 1295 562
rect 1198 491 1295 528
rect 1198 457 1251 491
rect 1285 457 1295 491
rect 1198 420 1295 457
rect 1198 386 1251 420
rect 1285 386 1295 420
rect 1198 374 1295 386
rect 1331 546 1358 574
rect 1392 546 1412 580
rect 1331 478 1412 546
rect 1331 444 1358 478
rect 1392 444 1412 478
rect 1331 374 1412 444
rect 1092 348 1142 374
rect 1362 368 1412 374
rect 1448 580 1502 592
rect 1448 546 1458 580
rect 1492 546 1502 580
rect 1448 497 1502 546
rect 1448 463 1458 497
rect 1492 463 1502 497
rect 1448 414 1502 463
rect 1448 380 1458 414
rect 1492 380 1502 414
rect 1448 368 1502 380
rect 1538 580 1594 592
rect 1538 546 1548 580
rect 1582 546 1594 580
rect 1538 497 1594 546
rect 1538 463 1548 497
rect 1582 463 1594 497
rect 1538 414 1594 463
rect 1538 380 1548 414
rect 1582 380 1594 414
rect 1538 368 1594 380
<< ndiffc >>
rect 39 149 73 183
rect 125 149 159 183
rect 329 176 363 210
rect 441 89 475 123
rect 593 119 627 153
rect 774 95 808 129
rect 910 150 944 184
rect 1022 168 1056 202
rect 1022 86 1056 120
rect 227 40 261 74
rect 1122 168 1156 202
rect 1122 86 1156 120
rect 1281 176 1315 210
rect 1281 86 1315 120
rect 1389 97 1423 131
rect 1475 176 1509 210
rect 1475 86 1509 120
rect 1561 176 1595 210
rect 1561 86 1595 120
<< pdiffc >>
rect 37 546 71 580
rect 37 442 71 476
rect 205 546 239 580
rect 205 464 239 498
rect 313 548 347 582
rect 418 380 452 414
rect 526 501 560 535
rect 526 393 560 427
rect 616 476 650 510
rect 814 534 848 568
rect 814 435 848 469
rect 904 534 938 568
rect 1118 528 1152 562
rect 904 451 938 485
rect 904 368 938 402
rect 1012 360 1046 394
rect 1251 528 1285 562
rect 1251 457 1285 491
rect 1251 386 1285 420
rect 1358 546 1392 580
rect 1358 444 1392 478
rect 1458 546 1492 580
rect 1458 463 1492 497
rect 1458 380 1492 414
rect 1548 546 1582 580
rect 1548 463 1582 497
rect 1548 380 1582 414
<< poly >>
rect 81 592 117 618
rect 159 592 195 618
rect 372 615 711 645
rect 372 536 408 615
rect 570 547 606 573
rect 81 392 117 424
rect 44 376 117 392
rect 44 342 60 376
rect 94 342 117 376
rect 44 308 117 342
rect 159 392 195 424
rect 159 376 225 392
rect 159 342 175 376
rect 209 342 225 376
rect 675 535 711 615
rect 858 580 894 606
rect 753 535 789 561
rect 675 425 711 451
rect 753 383 789 451
rect 159 326 225 342
rect 44 274 60 308
rect 94 274 117 308
rect 44 258 117 274
rect 84 222 114 258
rect 170 222 200 326
rect 372 272 408 368
rect 570 343 606 379
rect 706 367 789 383
rect 538 327 658 343
rect 538 293 554 327
rect 588 293 658 327
rect 706 333 722 367
rect 756 333 789 367
rect 1162 574 1198 600
rect 1295 574 1331 600
rect 1412 592 1448 618
rect 1502 592 1538 618
rect 1056 516 1092 542
rect 706 317 789 333
rect 858 317 894 356
rect 538 277 658 293
rect 288 256 496 272
rect 288 242 446 256
rect 288 222 318 242
rect 430 222 446 242
rect 480 229 496 256
rect 628 269 658 277
rect 628 239 685 269
rect 480 222 580 229
rect 84 86 114 112
rect 170 86 200 112
rect 430 199 580 222
rect 550 184 580 199
rect 655 165 685 239
rect 733 165 763 317
rect 831 301 899 317
rect 831 267 847 301
rect 881 267 899 301
rect 831 251 899 267
rect 869 229 899 251
rect 1056 310 1092 348
rect 1162 310 1198 374
rect 1295 326 1331 374
rect 1412 326 1448 368
rect 1502 326 1538 368
rect 1056 294 1198 310
rect 1056 260 1083 294
rect 1117 260 1198 294
rect 1056 244 1198 260
rect 1067 222 1097 244
rect 1168 222 1198 244
rect 1240 310 1331 326
rect 1240 276 1256 310
rect 1290 276 1331 310
rect 1240 260 1331 276
rect 1379 310 1538 326
rect 1379 276 1395 310
rect 1429 290 1538 310
rect 1429 276 1550 290
rect 1379 260 1550 276
rect 1240 222 1270 260
rect 1434 222 1464 260
rect 1520 222 1550 260
rect 288 48 318 74
rect 550 48 580 74
rect 655 55 685 81
rect 733 55 763 81
rect 869 55 899 81
rect 1067 48 1097 74
rect 1168 48 1198 74
rect 1240 48 1270 74
rect 1434 48 1464 74
rect 1520 48 1550 74
<< polycont >>
rect 60 342 94 376
rect 175 342 209 376
rect 60 274 94 308
rect 554 293 588 327
rect 722 333 756 367
rect 446 222 480 256
rect 847 267 881 301
rect 1083 260 1117 294
rect 1256 276 1290 310
rect 1395 276 1429 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 21 580 87 649
rect 21 546 37 580
rect 71 546 87 580
rect 21 476 87 546
rect 21 442 37 476
rect 71 442 87 476
rect 189 580 255 596
rect 189 546 205 580
rect 239 546 255 580
rect 189 498 255 546
rect 297 582 363 649
rect 297 548 313 582
rect 347 548 363 582
rect 798 568 848 649
rect 297 532 363 548
rect 510 535 560 551
rect 510 501 526 535
rect 510 498 560 501
rect 189 464 205 498
rect 239 464 560 498
rect 21 426 87 442
rect 25 376 110 392
rect 25 342 60 376
rect 94 342 110 376
rect 25 308 110 342
rect 159 376 260 430
rect 159 342 175 376
rect 209 342 260 376
rect 159 326 260 342
rect 25 274 60 308
rect 94 274 110 308
rect 294 278 328 464
rect 25 258 110 274
rect 144 244 328 278
rect 362 414 468 430
rect 362 380 418 414
rect 452 380 468 414
rect 362 343 468 380
rect 510 427 560 464
rect 600 510 672 539
rect 600 476 616 510
rect 650 476 672 510
rect 600 447 672 476
rect 510 393 526 427
rect 510 377 560 393
rect 362 327 604 343
rect 362 309 554 327
rect 144 224 178 244
rect 23 183 73 224
rect 23 149 39 183
rect 23 17 73 149
rect 109 183 178 224
rect 362 210 396 309
rect 538 293 554 309
rect 588 293 604 327
rect 538 277 604 293
rect 638 283 672 447
rect 798 534 814 568
rect 798 469 848 534
rect 798 435 814 469
rect 798 419 848 435
rect 888 568 965 584
rect 888 534 904 568
rect 938 534 965 568
rect 888 485 965 534
rect 1102 562 1168 649
rect 1342 580 1408 649
rect 1102 528 1118 562
rect 1152 528 1168 562
rect 1102 512 1168 528
rect 1235 562 1301 578
rect 1235 528 1251 562
rect 1285 528 1301 562
rect 888 451 904 485
rect 938 478 965 485
rect 1235 491 1301 528
rect 938 451 1201 478
rect 888 444 1201 451
rect 888 402 965 444
rect 888 385 904 402
rect 706 368 904 385
rect 938 368 965 402
rect 706 367 965 368
rect 706 333 722 367
rect 756 351 965 367
rect 756 333 772 351
rect 706 317 772 333
rect 831 301 897 317
rect 831 283 847 301
rect 109 149 125 183
rect 159 149 178 183
rect 313 176 329 210
rect 363 176 396 210
rect 430 256 496 272
rect 430 222 446 256
rect 480 240 496 256
rect 638 267 847 283
rect 881 267 897 301
rect 638 249 897 267
rect 480 222 543 240
rect 430 206 543 222
rect 109 142 178 149
rect 109 123 475 142
rect 109 108 441 123
rect 425 89 441 108
rect 211 40 227 74
rect 261 40 277 74
rect 425 70 475 89
rect 509 85 543 206
rect 638 169 672 249
rect 931 215 965 351
rect 577 153 672 169
rect 577 119 593 153
rect 627 119 672 153
rect 706 181 876 215
rect 706 85 740 181
rect 509 51 740 85
rect 774 129 808 147
rect 211 17 277 40
rect 774 17 808 95
rect 842 85 876 181
rect 910 184 965 215
rect 944 150 965 184
rect 910 119 965 150
rect 999 394 1062 410
rect 999 360 1012 394
rect 1046 360 1062 394
rect 999 344 1062 360
rect 999 202 1033 344
rect 1167 326 1201 444
rect 1235 457 1251 491
rect 1285 457 1301 491
rect 1235 420 1301 457
rect 1342 546 1358 580
rect 1392 546 1408 580
rect 1342 478 1408 546
rect 1342 444 1358 478
rect 1392 444 1408 478
rect 1342 428 1408 444
rect 1442 580 1513 596
rect 1442 546 1458 580
rect 1492 546 1513 580
rect 1442 497 1513 546
rect 1442 463 1458 497
rect 1492 463 1513 497
rect 1235 386 1251 420
rect 1285 394 1301 420
rect 1442 414 1513 463
rect 1285 386 1408 394
rect 1235 360 1408 386
rect 1442 380 1458 414
rect 1492 380 1513 414
rect 1442 364 1513 380
rect 1548 580 1598 649
rect 1582 546 1598 580
rect 1548 497 1598 546
rect 1582 463 1598 497
rect 1548 414 1598 463
rect 1582 380 1598 414
rect 1548 364 1598 380
rect 1374 326 1408 360
rect 1167 310 1306 326
rect 1067 294 1133 310
rect 1067 260 1083 294
rect 1117 260 1133 294
rect 1167 276 1256 310
rect 1290 276 1306 310
rect 1167 260 1306 276
rect 1374 310 1445 326
rect 1374 276 1395 310
rect 1429 276 1445 310
rect 1374 260 1445 276
rect 1067 236 1133 260
rect 1374 226 1408 260
rect 1479 226 1513 364
rect 1265 210 1408 226
rect 999 168 1022 202
rect 1056 168 1072 202
rect 999 120 1072 168
rect 999 86 1022 120
rect 1056 86 1072 120
rect 999 85 1072 86
rect 842 51 1072 85
rect 1106 168 1122 202
rect 1156 168 1172 202
rect 1106 120 1172 168
rect 1106 86 1122 120
rect 1156 86 1172 120
rect 1106 17 1172 86
rect 1265 176 1281 210
rect 1315 192 1408 210
rect 1459 210 1525 226
rect 1315 176 1331 192
rect 1265 120 1331 176
rect 1459 176 1475 210
rect 1509 176 1525 210
rect 1265 86 1281 120
rect 1315 86 1331 120
rect 1265 70 1331 86
rect 1373 131 1423 158
rect 1373 97 1389 131
rect 1373 17 1423 97
rect 1459 120 1525 176
rect 1459 86 1475 120
rect 1509 86 1525 120
rect 1459 70 1525 86
rect 1561 210 1611 226
rect 1595 176 1611 210
rect 1561 120 1611 176
rect 1595 86 1611 120
rect 1561 17 1611 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
rlabel comment s 0 0 0 0 4 sdlclkp_2
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 1471 390 1505 424 0 FreeSans 340 0 0 0 GCLK
port 8 nsew
flabel corelocali s 1471 464 1505 498 0 FreeSans 340 0 0 0 GCLK
port 8 nsew
flabel corelocali s 1471 538 1505 572 0 FreeSans 340 0 0 0 GCLK
port 8 nsew
flabel corelocali s 1087 242 1121 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 223 390 257 424 0 FreeSans 340 0 0 0 GATE
port 2 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 SCE
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 1632 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 276222
string GDS_START 264174
<< end >>
