magic
tech sky130A
magscale 1 2
timestamp 1601050047
<< nwell >>
rect -38 332 1382 704
<< pwell >>
rect 0 0 1344 49
<< scpmos >>
rect 86 392 116 592
rect 176 392 206 592
rect 276 392 306 592
rect 376 392 406 592
rect 486 392 516 592
rect 576 392 606 592
rect 676 392 706 592
rect 776 392 806 592
rect 886 368 916 592
rect 983 368 1013 592
rect 1128 368 1158 592
rect 1218 368 1248 592
<< nmoslvt >>
rect 84 136 114 264
rect 184 136 214 264
rect 270 136 300 264
rect 378 136 408 264
rect 483 136 513 264
rect 570 136 600 264
rect 671 136 701 264
rect 757 136 787 264
rect 971 74 1001 222
rect 1057 74 1087 222
rect 1143 74 1173 222
rect 1229 74 1259 222
<< ndiff >>
rect 27 252 84 264
rect 27 218 39 252
rect 73 218 84 252
rect 27 182 84 218
rect 27 148 39 182
rect 73 148 84 182
rect 27 136 84 148
rect 114 185 184 264
rect 114 151 139 185
rect 173 151 184 185
rect 114 136 184 151
rect 214 211 270 264
rect 214 177 225 211
rect 259 177 270 211
rect 214 136 270 177
rect 300 185 378 264
rect 300 151 325 185
rect 359 151 378 185
rect 300 136 378 151
rect 408 229 483 264
rect 408 195 425 229
rect 459 195 483 229
rect 408 136 483 195
rect 513 183 570 264
rect 513 149 525 183
rect 559 149 570 183
rect 513 136 570 149
rect 600 252 671 264
rect 600 218 618 252
rect 652 218 671 252
rect 600 136 671 218
rect 701 183 757 264
rect 701 149 712 183
rect 746 149 757 183
rect 701 136 757 149
rect 787 252 844 264
rect 787 218 798 252
rect 832 218 844 252
rect 787 136 844 218
rect 898 100 971 222
rect 898 66 910 100
rect 944 74 971 100
rect 1001 210 1057 222
rect 1001 176 1012 210
rect 1046 176 1057 210
rect 1001 120 1057 176
rect 1001 86 1012 120
rect 1046 86 1057 120
rect 1001 74 1057 86
rect 1087 142 1143 222
rect 1087 108 1098 142
rect 1132 108 1143 142
rect 1087 74 1143 108
rect 1173 210 1229 222
rect 1173 176 1184 210
rect 1218 176 1229 210
rect 1173 120 1229 176
rect 1173 86 1184 120
rect 1218 86 1229 120
rect 1173 74 1229 86
rect 1259 202 1317 222
rect 1259 168 1271 202
rect 1305 168 1317 202
rect 1259 120 1317 168
rect 1259 86 1271 120
rect 1305 86 1317 120
rect 1259 74 1317 86
rect 944 66 956 74
rect 898 54 956 66
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 509 86 546
rect 27 475 39 509
rect 73 475 86 509
rect 27 438 86 475
rect 27 404 39 438
rect 73 404 86 438
rect 27 392 86 404
rect 116 580 176 592
rect 116 546 129 580
rect 163 546 176 580
rect 116 510 176 546
rect 116 476 129 510
rect 163 476 176 510
rect 116 440 176 476
rect 116 406 129 440
rect 163 406 176 440
rect 116 392 176 406
rect 206 531 276 592
rect 206 497 229 531
rect 263 497 276 531
rect 206 440 276 497
rect 206 406 229 440
rect 263 406 276 440
rect 206 392 276 406
rect 306 580 376 592
rect 306 546 329 580
rect 363 546 376 580
rect 306 508 376 546
rect 306 474 329 508
rect 363 474 376 508
rect 306 392 376 474
rect 406 580 486 592
rect 406 546 429 580
rect 463 546 486 580
rect 406 508 486 546
rect 406 474 429 508
rect 463 474 486 508
rect 406 392 486 474
rect 516 580 576 592
rect 516 546 529 580
rect 563 546 576 580
rect 516 508 576 546
rect 516 474 529 508
rect 563 474 576 508
rect 516 392 576 474
rect 606 531 676 592
rect 606 497 629 531
rect 663 497 676 531
rect 606 440 676 497
rect 606 406 629 440
rect 663 406 676 440
rect 606 392 676 406
rect 706 580 776 592
rect 706 546 729 580
rect 763 546 776 580
rect 706 508 776 546
rect 706 474 729 508
rect 763 474 776 508
rect 706 392 776 474
rect 806 580 886 592
rect 806 546 836 580
rect 870 546 886 580
rect 806 500 886 546
rect 806 466 836 500
rect 870 466 886 500
rect 806 420 886 466
rect 806 392 836 420
rect 824 386 836 392
rect 870 386 886 420
rect 824 368 886 386
rect 916 580 983 592
rect 916 546 936 580
rect 970 546 983 580
rect 916 500 983 546
rect 916 466 936 500
rect 970 466 983 500
rect 916 420 983 466
rect 916 386 936 420
rect 970 386 983 420
rect 916 368 983 386
rect 1013 580 1128 592
rect 1013 546 1056 580
rect 1090 546 1128 580
rect 1013 488 1128 546
rect 1013 454 1056 488
rect 1090 454 1128 488
rect 1013 368 1128 454
rect 1158 580 1218 592
rect 1158 546 1171 580
rect 1205 546 1218 580
rect 1158 500 1218 546
rect 1158 466 1171 500
rect 1205 466 1218 500
rect 1158 420 1218 466
rect 1158 386 1171 420
rect 1205 386 1218 420
rect 1158 368 1218 386
rect 1248 580 1317 592
rect 1248 546 1271 580
rect 1305 546 1317 580
rect 1248 497 1317 546
rect 1248 463 1271 497
rect 1305 463 1317 497
rect 1248 414 1317 463
rect 1248 380 1271 414
rect 1305 380 1317 414
rect 1248 368 1317 380
<< ndiffc >>
rect 39 218 73 252
rect 39 148 73 182
rect 139 151 173 185
rect 225 177 259 211
rect 325 151 359 185
rect 425 195 459 229
rect 525 149 559 183
rect 618 218 652 252
rect 712 149 746 183
rect 798 218 832 252
rect 910 66 944 100
rect 1012 176 1046 210
rect 1012 86 1046 120
rect 1098 108 1132 142
rect 1184 176 1218 210
rect 1184 86 1218 120
rect 1271 168 1305 202
rect 1271 86 1305 120
<< pdiffc >>
rect 39 546 73 580
rect 39 475 73 509
rect 39 404 73 438
rect 129 546 163 580
rect 129 476 163 510
rect 129 406 163 440
rect 229 497 263 531
rect 229 406 263 440
rect 329 546 363 580
rect 329 474 363 508
rect 429 546 463 580
rect 429 474 463 508
rect 529 546 563 580
rect 529 474 563 508
rect 629 497 663 531
rect 629 406 663 440
rect 729 546 763 580
rect 729 474 763 508
rect 836 546 870 580
rect 836 466 870 500
rect 836 386 870 420
rect 936 546 970 580
rect 936 466 970 500
rect 936 386 970 420
rect 1056 546 1090 580
rect 1056 454 1090 488
rect 1171 546 1205 580
rect 1171 466 1205 500
rect 1171 386 1205 420
rect 1271 546 1305 580
rect 1271 463 1305 497
rect 1271 380 1305 414
<< poly >>
rect 86 592 116 618
rect 176 592 206 618
rect 276 592 306 618
rect 376 592 406 618
rect 486 592 516 618
rect 576 592 606 618
rect 676 592 706 618
rect 776 592 806 618
rect 886 592 916 618
rect 983 592 1013 618
rect 1128 592 1158 618
rect 1218 592 1248 618
rect 86 377 116 392
rect 176 377 206 392
rect 276 377 306 392
rect 376 377 406 392
rect 486 377 516 392
rect 576 377 606 392
rect 676 377 706 392
rect 776 377 806 392
rect 83 309 119 377
rect 173 356 209 377
rect 273 356 309 377
rect 373 356 409 377
rect 169 340 309 356
rect 83 279 114 309
rect 169 306 185 340
rect 219 306 253 340
rect 287 320 309 340
rect 369 340 435 356
rect 287 306 303 320
rect 169 290 303 306
rect 369 306 385 340
rect 419 306 435 340
rect 369 290 435 306
rect 84 264 114 279
rect 184 264 214 290
rect 270 279 303 290
rect 270 264 300 279
rect 378 264 408 290
rect 483 279 519 377
rect 573 356 609 377
rect 673 356 709 377
rect 567 340 709 356
rect 567 306 583 340
rect 617 306 651 340
rect 685 306 709 340
rect 773 309 809 377
rect 886 353 916 368
rect 983 353 1013 368
rect 1128 353 1158 368
rect 1218 353 1248 368
rect 567 290 709 306
rect 483 264 513 279
rect 570 264 600 290
rect 671 279 709 290
rect 757 279 809 309
rect 883 336 919 353
rect 980 336 1016 353
rect 1125 336 1161 353
rect 1215 336 1251 353
rect 883 320 1251 336
rect 883 286 899 320
rect 933 286 967 320
rect 1001 286 1035 320
rect 1069 286 1103 320
rect 1137 300 1251 320
rect 1137 286 1259 300
rect 671 264 701 279
rect 757 264 787 279
rect 883 270 1259 286
rect 971 222 1001 270
rect 1057 222 1087 270
rect 1143 222 1173 270
rect 1229 222 1259 270
rect 84 62 114 136
rect 184 110 214 136
rect 270 110 300 136
rect 378 62 408 136
rect 483 114 513 136
rect 84 32 408 62
rect 456 98 522 114
rect 570 110 600 136
rect 671 110 701 136
rect 456 64 472 98
rect 506 64 522 98
rect 456 62 522 64
rect 757 62 787 136
rect 456 32 787 62
rect 971 48 1001 74
rect 1057 48 1087 74
rect 1143 48 1173 74
rect 1229 48 1259 74
<< polycont >>
rect 185 306 219 340
rect 253 306 287 340
rect 385 306 419 340
rect 583 306 617 340
rect 651 306 685 340
rect 899 286 933 320
rect 967 286 1001 320
rect 1035 286 1069 320
rect 1103 286 1137 320
rect 472 64 506 98
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 23 580 73 649
rect 23 546 39 580
rect 23 509 73 546
rect 23 475 39 509
rect 23 438 73 475
rect 23 404 39 438
rect 23 388 73 404
rect 113 581 379 615
rect 113 580 179 581
rect 113 546 129 580
rect 163 546 179 580
rect 313 580 379 581
rect 113 510 179 546
rect 113 476 129 510
rect 163 476 179 510
rect 113 440 179 476
rect 113 406 129 440
rect 163 406 179 440
rect 113 390 179 406
rect 213 531 279 547
rect 213 497 229 531
rect 263 497 279 531
rect 213 440 279 497
rect 313 546 329 580
rect 363 546 379 580
rect 313 508 379 546
rect 313 474 329 508
rect 363 474 379 508
rect 313 458 379 474
rect 413 580 479 649
rect 413 546 429 580
rect 463 546 479 580
rect 413 508 479 546
rect 413 474 429 508
rect 463 474 479 508
rect 413 458 479 474
rect 513 581 779 615
rect 513 580 579 581
rect 513 546 529 580
rect 563 546 579 580
rect 713 580 779 581
rect 513 508 579 546
rect 513 474 529 508
rect 563 474 579 508
rect 513 458 579 474
rect 613 531 679 547
rect 613 497 629 531
rect 663 497 679 531
rect 213 406 229 440
rect 263 424 279 440
rect 613 440 679 497
rect 713 546 729 580
rect 763 546 779 580
rect 713 508 779 546
rect 713 474 729 508
rect 763 474 779 508
rect 713 458 779 474
rect 820 580 886 649
rect 820 546 836 580
rect 870 546 886 580
rect 820 500 886 546
rect 820 466 836 500
rect 870 466 886 500
rect 613 424 629 440
rect 263 406 629 424
rect 663 424 679 440
rect 663 406 769 424
rect 213 390 769 406
rect 169 340 303 356
rect 169 306 185 340
rect 219 306 253 340
rect 287 306 303 340
rect 169 290 303 306
rect 369 340 455 356
rect 369 306 385 340
rect 419 306 455 340
rect 369 290 455 306
rect 505 340 701 356
rect 505 306 583 340
rect 617 306 651 340
rect 685 306 701 340
rect 505 290 701 306
rect 735 336 769 390
rect 820 420 886 466
rect 820 386 836 420
rect 870 386 886 420
rect 820 370 886 386
rect 920 580 986 596
rect 920 546 936 580
rect 970 546 986 580
rect 920 500 986 546
rect 920 466 936 500
rect 970 466 986 500
rect 920 420 986 466
rect 1040 580 1106 649
rect 1040 546 1056 580
rect 1090 546 1106 580
rect 1040 488 1106 546
rect 1040 454 1056 488
rect 1090 454 1106 488
rect 1040 438 1106 454
rect 1155 580 1221 596
rect 1155 546 1171 580
rect 1205 546 1221 580
rect 1155 500 1221 546
rect 1155 466 1171 500
rect 1205 466 1221 500
rect 920 386 936 420
rect 970 404 986 420
rect 1155 420 1221 466
rect 1155 404 1171 420
rect 970 386 1171 404
rect 1205 386 1221 420
rect 920 370 1221 386
rect 735 320 1153 336
rect 735 302 899 320
rect 883 286 899 302
rect 933 286 967 320
rect 1001 286 1035 320
rect 1069 286 1103 320
rect 1137 286 1153 320
rect 883 270 1153 286
rect 1187 282 1221 370
rect 1255 580 1321 649
rect 1255 546 1271 580
rect 1305 546 1321 580
rect 1255 497 1321 546
rect 1255 463 1271 497
rect 1305 463 1321 497
rect 1255 414 1321 463
rect 1255 380 1271 414
rect 1305 380 1321 414
rect 1255 364 1321 380
rect 23 256 89 268
rect 782 256 848 268
rect 23 252 848 256
rect 23 218 39 252
rect 73 229 618 252
rect 73 222 425 229
rect 73 218 89 222
rect 23 182 89 218
rect 225 211 275 222
rect 23 148 39 182
rect 73 148 89 182
rect 23 132 89 148
rect 123 185 189 188
rect 123 151 139 185
rect 173 151 189 185
rect 123 17 189 151
rect 259 177 275 211
rect 409 195 425 222
rect 459 218 618 229
rect 652 218 798 252
rect 832 218 848 252
rect 459 195 475 218
rect 225 132 275 177
rect 309 185 375 188
rect 309 151 325 185
rect 359 151 375 185
rect 409 168 475 195
rect 883 184 917 270
rect 1187 236 1319 282
rect 509 183 917 184
rect 309 17 375 151
rect 509 149 525 183
rect 559 149 712 183
rect 746 150 917 183
rect 996 210 1221 236
rect 996 176 1012 210
rect 1046 202 1184 210
rect 746 149 762 150
rect 509 148 762 149
rect 409 114 455 134
rect 696 132 762 148
rect 996 120 1046 176
rect 1218 176 1221 210
rect 409 98 522 114
rect 409 64 472 98
rect 506 64 522 98
rect 409 51 522 64
rect 894 100 960 116
rect 894 66 910 100
rect 944 66 960 100
rect 996 86 1012 120
rect 996 70 1046 86
rect 1082 142 1148 158
rect 1082 108 1098 142
rect 1132 108 1148 142
rect 894 17 960 66
rect 1082 17 1148 108
rect 1184 120 1221 176
rect 1218 86 1221 120
rect 1184 70 1221 86
rect 1255 168 1271 202
rect 1305 168 1321 202
rect 1255 120 1321 168
rect 1255 86 1271 120
rect 1305 86 1321 120
rect 1255 17 1321 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
<< metal1 >>
rect 0 683 1344 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 0 617 1344 649
rect 0 17 1344 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
rect 0 -49 1344 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o22a_4
flabel pwell s 0 0 1344 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 1344 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 1344 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 1344 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 415 94 449 128 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 1279 242 1313 276 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 B2
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 1344 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1309014
string GDS_START 1298006
<< end >>
