magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 644 561
rect 286 451 357 527
rect 491 371 541 527
rect 575 357 627 493
rect 17 215 115 255
rect 153 215 248 257
rect 18 17 109 170
rect 204 135 248 215
rect 297 215 363 257
rect 297 135 339 215
rect 397 208 479 269
rect 593 117 627 357
rect 475 17 541 89
rect 575 51 627 117
rect 0 -17 644 17
<< obsli1 >>
rect 18 449 85 493
rect 18 325 69 449
rect 119 417 165 425
rect 391 417 441 493
rect 119 377 441 417
rect 119 359 156 377
rect 274 375 441 377
rect 187 337 253 343
rect 187 325 547 337
rect 18 303 559 325
rect 18 291 253 303
rect 519 296 559 303
rect 525 181 559 296
rect 505 157 559 181
rect 390 148 559 157
rect 390 123 541 148
rect 390 93 424 123
rect 164 51 424 93
<< metal1 >>
rect 0 496 644 592
rect 0 -48 644 48
<< labels >>
rlabel locali s 297 215 363 257 6 A1
port 1 nsew signal input
rlabel locali s 297 135 339 215 6 A1
port 1 nsew signal input
rlabel locali s 397 208 479 269 6 A2
port 2 nsew signal input
rlabel locali s 204 135 248 215 6 B1
port 3 nsew signal input
rlabel locali s 153 215 248 257 6 B1
port 3 nsew signal input
rlabel locali s 17 215 115 255 6 B2
port 4 nsew signal input
rlabel locali s 593 117 627 357 6 X
port 5 nsew signal output
rlabel locali s 575 357 627 493 6 X
port 5 nsew signal output
rlabel locali s 575 51 627 117 6 X
port 5 nsew signal output
rlabel locali s 475 17 541 89 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 18 17 109 170 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 644 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 644 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 491 371 541 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 286 451 357 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 644 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 644 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 4134734
string GDS_START 4128146
<< end >>
