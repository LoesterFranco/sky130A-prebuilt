magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 644 561
rect 18 299 72 527
rect 106 357 309 493
rect 18 199 72 265
rect 18 137 69 199
rect 106 165 140 357
rect 174 199 248 323
rect 282 199 340 323
rect 386 199 445 493
rect 539 299 627 527
rect 515 199 627 265
rect 103 131 169 165
rect 303 17 437 97
rect 539 17 627 165
rect 0 -17 644 17
<< obsli1 >>
rect 203 131 505 165
rect 203 97 269 131
rect 18 51 269 97
rect 471 75 505 131
<< metal1 >>
rect 0 496 644 592
rect 0 -48 644 48
<< labels >>
rlabel locali s 515 199 627 265 6 A1
port 1 nsew signal input
rlabel locali s 386 199 445 493 6 A2
port 2 nsew signal input
rlabel locali s 282 199 340 323 6 A3
port 3 nsew signal input
rlabel locali s 18 199 72 265 6 B1
port 4 nsew signal input
rlabel locali s 18 137 69 199 6 B1
port 4 nsew signal input
rlabel locali s 174 199 248 323 6 B2
port 5 nsew signal input
rlabel locali s 106 357 309 493 6 Y
port 6 nsew signal output
rlabel locali s 106 165 140 357 6 Y
port 6 nsew signal output
rlabel locali s 103 131 169 165 6 Y
port 6 nsew signal output
rlabel locali s 539 17 627 165 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 303 17 437 97 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 644 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 644 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 539 299 627 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 18 299 72 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 644 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 644 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 912600
string GDS_START 905924
<< end >>
