magic
tech sky130A
magscale 1 2
timestamp 1601050047
<< nwell >>
rect -38 332 2054 704
<< pwell >>
rect 0 0 2016 49
<< scpmos >>
rect 86 368 116 592
rect 176 368 206 592
rect 266 368 296 592
rect 356 368 386 592
rect 448 368 478 592
rect 546 368 576 592
rect 646 368 676 592
rect 746 368 776 592
rect 1033 368 1063 592
rect 1123 368 1153 592
rect 1213 368 1243 592
rect 1319 368 1349 592
rect 1419 368 1449 592
rect 1509 368 1539 592
rect 1619 368 1649 592
rect 1709 368 1739 592
rect 1810 368 1840 536
rect 1900 368 1930 536
<< nmoslvt >>
rect 84 85 114 233
rect 170 85 200 233
rect 256 85 286 233
rect 359 85 389 233
rect 445 85 475 233
rect 545 85 575 233
rect 640 85 670 233
rect 726 85 756 233
rect 1048 98 1078 246
rect 1134 98 1164 246
rect 1252 82 1282 230
rect 1338 82 1368 230
rect 1456 82 1486 230
rect 1542 82 1572 230
rect 1674 82 1704 230
rect 1760 82 1790 230
rect 1860 82 1890 230
<< ndiff >>
rect 27 221 84 233
rect 27 187 39 221
rect 73 187 84 221
rect 27 131 84 187
rect 27 97 39 131
rect 73 97 84 131
rect 27 85 84 97
rect 114 152 170 233
rect 114 118 125 152
rect 159 118 170 152
rect 114 85 170 118
rect 200 181 256 233
rect 200 147 211 181
rect 245 147 256 181
rect 200 85 256 147
rect 286 152 359 233
rect 286 118 297 152
rect 331 118 359 152
rect 286 85 359 118
rect 389 225 445 233
rect 389 191 400 225
rect 434 191 445 225
rect 389 153 445 191
rect 389 119 400 153
rect 434 119 445 153
rect 389 85 445 119
rect 475 153 545 233
rect 475 119 500 153
rect 534 119 545 153
rect 475 85 545 119
rect 575 221 640 233
rect 575 187 590 221
rect 624 187 640 221
rect 575 85 640 187
rect 670 153 726 233
rect 670 119 681 153
rect 715 119 726 153
rect 670 85 726 119
rect 756 221 813 233
rect 756 187 767 221
rect 801 187 813 221
rect 756 85 813 187
rect 975 98 1048 246
rect 1078 234 1134 246
rect 1078 200 1089 234
rect 1123 200 1134 234
rect 1078 98 1134 200
rect 1164 230 1214 246
rect 1164 98 1252 230
rect 975 82 1033 98
rect 975 48 987 82
rect 1021 48 1033 82
rect 1179 82 1252 98
rect 1282 218 1338 230
rect 1282 184 1293 218
rect 1327 184 1338 218
rect 1282 82 1338 184
rect 1368 82 1456 230
rect 1486 202 1542 230
rect 1486 168 1497 202
rect 1531 168 1542 202
rect 1486 128 1542 168
rect 1486 94 1497 128
rect 1531 94 1542 128
rect 1486 82 1542 94
rect 1572 128 1674 230
rect 1572 94 1606 128
rect 1640 94 1674 128
rect 1572 82 1674 94
rect 1704 202 1760 230
rect 1704 168 1715 202
rect 1749 168 1760 202
rect 1704 128 1760 168
rect 1704 94 1715 128
rect 1749 94 1760 128
rect 1704 82 1760 94
rect 1790 202 1860 230
rect 1790 168 1815 202
rect 1849 168 1860 202
rect 1790 128 1860 168
rect 1790 94 1815 128
rect 1849 94 1860 128
rect 1790 82 1860 94
rect 1890 202 1961 230
rect 1890 168 1915 202
rect 1949 168 1961 202
rect 1890 128 1961 168
rect 1890 94 1915 128
rect 1949 94 1961 128
rect 1890 82 1961 94
rect 975 36 1033 48
rect 1179 48 1191 82
rect 1225 48 1237 82
rect 1179 36 1237 48
rect 1383 48 1395 82
rect 1429 48 1441 82
rect 1383 36 1441 48
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 497 86 546
rect 27 463 39 497
rect 73 463 86 497
rect 27 414 86 463
rect 27 380 39 414
rect 73 380 86 414
rect 27 368 86 380
rect 116 580 176 592
rect 116 546 129 580
rect 163 546 176 580
rect 116 500 176 546
rect 116 466 129 500
rect 163 466 176 500
rect 116 368 176 466
rect 206 531 266 592
rect 206 497 219 531
rect 253 497 266 531
rect 206 424 266 497
rect 206 390 219 424
rect 253 390 266 424
rect 206 368 266 390
rect 296 580 356 592
rect 296 546 309 580
rect 343 546 356 580
rect 296 508 356 546
rect 296 474 309 508
rect 343 474 356 508
rect 296 368 356 474
rect 386 531 448 592
rect 386 497 399 531
rect 433 497 448 531
rect 386 424 448 497
rect 386 390 399 424
rect 433 390 448 424
rect 386 368 448 390
rect 478 508 546 592
rect 478 474 499 508
rect 533 474 546 508
rect 478 368 546 474
rect 576 463 646 592
rect 576 429 599 463
rect 633 429 646 463
rect 576 368 646 429
rect 676 508 746 592
rect 676 474 699 508
rect 733 474 746 508
rect 676 368 746 474
rect 776 478 845 592
rect 776 444 799 478
rect 833 444 845 478
rect 776 410 845 444
rect 776 376 799 410
rect 833 376 845 410
rect 776 368 845 376
rect 899 418 1033 592
rect 899 384 911 418
rect 945 384 986 418
rect 1020 384 1033 418
rect 899 368 1033 384
rect 1063 580 1123 592
rect 1063 546 1076 580
rect 1110 546 1123 580
rect 1063 368 1123 546
rect 1153 423 1213 592
rect 1153 389 1166 423
rect 1200 389 1213 423
rect 1153 368 1213 389
rect 1243 580 1319 592
rect 1243 546 1259 580
rect 1293 546 1319 580
rect 1243 368 1319 546
rect 1349 580 1419 592
rect 1349 546 1362 580
rect 1396 546 1419 580
rect 1349 368 1419 546
rect 1449 580 1509 592
rect 1449 546 1462 580
rect 1496 546 1509 580
rect 1449 512 1509 546
rect 1449 478 1462 512
rect 1496 478 1509 512
rect 1449 368 1509 478
rect 1539 580 1619 592
rect 1539 546 1562 580
rect 1596 546 1619 580
rect 1539 368 1619 546
rect 1649 580 1709 592
rect 1649 546 1662 580
rect 1696 546 1709 580
rect 1649 512 1709 546
rect 1649 478 1662 512
rect 1696 478 1709 512
rect 1649 368 1709 478
rect 1739 536 1792 592
rect 1739 528 1810 536
rect 1739 494 1752 528
rect 1786 494 1810 528
rect 1739 444 1810 494
rect 1739 410 1752 444
rect 1786 410 1810 444
rect 1739 368 1810 410
rect 1840 524 1900 536
rect 1840 490 1853 524
rect 1887 490 1900 524
rect 1840 414 1900 490
rect 1840 380 1853 414
rect 1887 380 1900 414
rect 1840 368 1900 380
rect 1930 524 1989 536
rect 1930 490 1943 524
rect 1977 490 1989 524
rect 1930 456 1989 490
rect 1930 422 1943 456
rect 1977 422 1989 456
rect 1930 368 1989 422
<< ndiffc >>
rect 39 187 73 221
rect 39 97 73 131
rect 125 118 159 152
rect 211 147 245 181
rect 297 118 331 152
rect 400 191 434 225
rect 400 119 434 153
rect 500 119 534 153
rect 590 187 624 221
rect 681 119 715 153
rect 767 187 801 221
rect 1089 200 1123 234
rect 987 48 1021 82
rect 1293 184 1327 218
rect 1497 168 1531 202
rect 1497 94 1531 128
rect 1606 94 1640 128
rect 1715 168 1749 202
rect 1715 94 1749 128
rect 1815 168 1849 202
rect 1815 94 1849 128
rect 1915 168 1949 202
rect 1915 94 1949 128
rect 1191 48 1225 82
rect 1395 48 1429 82
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 129 546 163 580
rect 129 466 163 500
rect 219 497 253 531
rect 219 390 253 424
rect 309 546 343 580
rect 309 474 343 508
rect 399 497 433 531
rect 399 390 433 424
rect 499 474 533 508
rect 599 429 633 463
rect 699 474 733 508
rect 799 444 833 478
rect 799 376 833 410
rect 911 384 945 418
rect 986 384 1020 418
rect 1076 546 1110 580
rect 1166 389 1200 423
rect 1259 546 1293 580
rect 1362 546 1396 580
rect 1462 546 1496 580
rect 1462 478 1496 512
rect 1562 546 1596 580
rect 1662 546 1696 580
rect 1662 478 1696 512
rect 1752 494 1786 528
rect 1752 410 1786 444
rect 1853 490 1887 524
rect 1853 380 1887 414
rect 1943 490 1977 524
rect 1943 422 1977 456
<< poly >>
rect 86 592 116 618
rect 176 592 206 618
rect 266 592 296 618
rect 356 592 386 618
rect 448 592 478 618
rect 546 592 576 618
rect 646 592 676 618
rect 746 592 776 618
rect 1033 592 1063 618
rect 1123 592 1153 618
rect 1213 592 1243 618
rect 1319 592 1349 618
rect 1419 592 1449 618
rect 1509 592 1539 618
rect 1619 592 1649 618
rect 1709 592 1739 618
rect 1810 536 1840 562
rect 1900 536 1930 562
rect 86 353 116 368
rect 176 353 206 368
rect 266 353 296 368
rect 356 353 386 368
rect 448 353 478 368
rect 546 353 576 368
rect 646 353 676 368
rect 746 353 776 368
rect 1033 353 1063 368
rect 1123 353 1153 368
rect 1213 353 1243 368
rect 1319 353 1349 368
rect 1419 353 1449 368
rect 1509 353 1539 368
rect 1619 353 1649 368
rect 1709 353 1739 368
rect 1810 353 1840 368
rect 1900 353 1930 368
rect 83 336 119 353
rect 173 336 209 353
rect 263 336 299 353
rect 353 336 389 353
rect 83 320 389 336
rect 83 286 123 320
rect 157 286 191 320
rect 225 286 259 320
rect 293 286 327 320
rect 361 286 389 320
rect 83 270 389 286
rect 84 233 114 270
rect 170 233 200 270
rect 256 233 286 270
rect 359 233 389 270
rect 445 336 481 353
rect 543 336 579 353
rect 643 336 679 353
rect 445 320 679 336
rect 445 286 461 320
rect 495 286 529 320
rect 563 286 597 320
rect 631 300 679 320
rect 743 300 779 353
rect 631 286 779 300
rect 445 270 779 286
rect 1030 334 1066 353
rect 1120 334 1156 353
rect 1210 334 1246 353
rect 1316 334 1352 353
rect 1030 318 1368 334
rect 1030 284 1046 318
rect 1080 284 1114 318
rect 1148 284 1182 318
rect 1216 284 1250 318
rect 1284 284 1318 318
rect 1352 284 1368 318
rect 445 233 475 270
rect 545 233 575 270
rect 640 233 670 270
rect 726 233 756 270
rect 1030 268 1368 284
rect 1048 246 1078 268
rect 1134 246 1164 268
rect 1252 230 1282 268
rect 1338 230 1368 268
rect 1416 318 1452 353
rect 1506 318 1542 353
rect 1616 318 1652 353
rect 1706 318 1742 353
rect 1807 318 1843 353
rect 1897 318 1933 353
rect 1416 302 1933 318
rect 1416 268 1432 302
rect 1466 268 1500 302
rect 1534 268 1568 302
rect 1602 268 1636 302
rect 1670 268 1704 302
rect 1738 268 1772 302
rect 1806 268 1840 302
rect 1874 288 1933 302
rect 1874 268 1890 288
rect 1416 252 1890 268
rect 1456 230 1486 252
rect 1542 230 1572 252
rect 1674 230 1704 252
rect 1760 230 1790 252
rect 1860 230 1890 252
rect 84 59 114 85
rect 170 59 200 85
rect 256 59 286 85
rect 359 59 389 85
rect 445 59 475 85
rect 545 59 575 85
rect 640 59 670 85
rect 726 59 756 85
rect 1048 72 1078 98
rect 1134 72 1164 98
rect 1252 56 1282 82
rect 1338 56 1368 82
rect 1456 56 1486 82
rect 1542 56 1572 82
rect 1674 56 1704 82
rect 1760 56 1790 82
rect 1860 56 1890 82
<< polycont >>
rect 123 286 157 320
rect 191 286 225 320
rect 259 286 293 320
rect 327 286 361 320
rect 461 286 495 320
rect 529 286 563 320
rect 597 286 631 320
rect 1046 284 1080 318
rect 1114 284 1148 318
rect 1182 284 1216 318
rect 1250 284 1284 318
rect 1318 284 1352 318
rect 1432 268 1466 302
rect 1500 268 1534 302
rect 1568 268 1602 302
rect 1636 268 1670 302
rect 1704 268 1738 302
rect 1772 268 1806 302
rect 1840 268 1874 302
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 23 580 73 596
rect 23 546 39 580
rect 23 497 73 546
rect 23 463 39 497
rect 23 424 73 463
rect 113 581 1312 615
rect 113 580 179 581
rect 113 546 129 580
rect 163 546 179 580
rect 293 580 343 581
rect 113 500 179 546
rect 113 466 129 500
rect 163 466 179 500
rect 113 458 179 466
rect 219 531 253 547
rect 219 424 253 497
rect 293 546 309 580
rect 1060 580 1312 581
rect 293 508 343 546
rect 293 474 309 508
rect 293 458 343 474
rect 383 531 449 547
rect 383 497 399 531
rect 433 497 449 531
rect 383 424 449 497
rect 483 513 1026 547
rect 1060 546 1076 580
rect 1110 546 1259 580
rect 1293 546 1312 580
rect 1346 580 1412 649
rect 1346 546 1362 580
rect 1396 546 1412 580
rect 1446 580 1512 596
rect 1446 546 1462 580
rect 1496 546 1512 580
rect 1546 580 1612 649
rect 1546 546 1562 580
rect 1596 546 1612 580
rect 1646 580 1712 596
rect 1646 546 1662 580
rect 1696 546 1712 580
rect 483 508 549 513
rect 483 474 499 508
rect 533 474 549 508
rect 683 508 749 513
rect 483 458 549 474
rect 583 463 649 479
rect 583 429 599 463
rect 633 429 649 463
rect 683 474 699 508
rect 733 474 749 508
rect 992 512 1026 513
rect 1446 512 1512 546
rect 1646 512 1712 546
rect 683 458 749 474
rect 783 478 849 479
rect 992 478 1462 512
rect 1496 478 1662 512
rect 1696 478 1712 512
rect 1752 528 1802 649
rect 1786 494 1802 528
rect 583 424 649 429
rect 783 444 799 478
rect 833 444 849 478
rect 1752 444 1802 494
rect 783 424 849 444
rect 23 414 219 424
rect 23 380 39 414
rect 73 390 219 414
rect 253 390 399 424
rect 433 410 849 424
rect 433 390 799 410
rect 23 364 73 380
rect 697 376 799 390
rect 833 376 849 410
rect 107 320 377 356
rect 505 336 647 356
rect 107 286 123 320
rect 157 286 191 320
rect 225 286 259 320
rect 293 286 327 320
rect 361 286 377 320
rect 107 270 377 286
rect 445 320 647 336
rect 445 286 461 320
rect 495 286 529 320
rect 563 286 597 320
rect 631 286 647 320
rect 697 310 849 376
rect 895 423 1752 444
rect 895 418 1166 423
rect 895 384 911 418
rect 945 384 986 418
rect 1020 389 1166 418
rect 1200 410 1752 423
rect 1786 410 1802 444
rect 1837 524 1891 540
rect 1837 490 1853 524
rect 1887 490 1891 524
rect 1837 414 1891 490
rect 1200 389 1216 410
rect 1020 384 1216 389
rect 895 368 1216 384
rect 1837 380 1853 414
rect 1887 380 1891 414
rect 1927 524 1993 649
rect 1927 490 1943 524
rect 1977 490 1993 524
rect 1927 456 1993 490
rect 1927 422 1943 456
rect 1977 422 1993 456
rect 1927 410 1993 422
rect 1837 376 1891 380
rect 1334 342 1965 376
rect 1334 334 1368 342
rect 1030 318 1368 334
rect 445 270 647 286
rect 23 236 73 237
rect 783 236 817 310
rect 1030 284 1046 318
rect 1080 284 1114 318
rect 1148 284 1182 318
rect 1216 284 1250 318
rect 1284 284 1318 318
rect 1352 284 1368 318
rect 1030 268 1368 284
rect 1416 302 1895 308
rect 1416 268 1432 302
rect 1466 268 1500 302
rect 1534 268 1568 302
rect 1602 268 1636 302
rect 1670 268 1704 302
rect 1738 268 1772 302
rect 1806 268 1840 302
rect 1874 268 1895 302
rect 1416 236 1895 268
rect 23 225 817 236
rect 23 221 400 225
rect 23 187 39 221
rect 73 202 400 221
rect 23 131 73 187
rect 211 181 245 202
rect 23 97 39 131
rect 23 81 73 97
rect 109 152 175 168
rect 109 118 125 152
rect 159 118 175 152
rect 384 191 400 202
rect 434 221 817 225
rect 434 191 590 221
rect 384 187 590 191
rect 624 187 767 221
rect 801 187 817 221
rect 851 200 1089 234
rect 1123 218 1343 234
rect 1123 200 1293 218
rect 211 119 245 147
rect 281 152 347 168
rect 109 85 175 118
rect 281 118 297 152
rect 331 118 347 152
rect 384 153 450 187
rect 851 153 885 200
rect 1277 184 1293 200
rect 1327 184 1343 218
rect 1931 202 1965 342
rect 1481 168 1497 202
rect 1531 168 1715 202
rect 1749 168 1765 202
rect 384 119 400 153
rect 434 119 450 153
rect 484 119 500 153
rect 534 119 681 153
rect 715 119 885 153
rect 919 150 1105 166
rect 1481 150 1547 168
rect 919 132 1547 150
rect 281 85 347 118
rect 919 85 953 132
rect 1071 128 1547 132
rect 1699 128 1765 168
rect 1071 116 1497 128
rect 109 51 953 85
rect 987 82 1037 98
rect 1481 94 1497 116
rect 1531 94 1547 128
rect 1021 48 1037 82
rect 987 17 1037 48
rect 1175 48 1191 82
rect 1225 48 1241 82
rect 1175 17 1241 48
rect 1379 48 1395 82
rect 1429 48 1445 82
rect 1481 78 1547 94
rect 1581 94 1606 128
rect 1640 94 1665 128
rect 1379 17 1445 48
rect 1581 17 1665 94
rect 1699 94 1715 128
rect 1749 94 1765 128
rect 1699 78 1765 94
rect 1799 168 1815 202
rect 1849 168 1865 202
rect 1799 128 1865 168
rect 1799 94 1815 128
rect 1849 94 1865 128
rect 1799 17 1865 94
rect 1899 168 1915 202
rect 1949 168 1965 202
rect 1899 128 1965 168
rect 1899 94 1915 128
rect 1949 94 1965 128
rect 1899 78 1965 94
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
rlabel comment s 0 0 0 0 4 mux2i_4
flabel pwell s 0 0 2016 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 2016 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 2016 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 2016 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 1471 242 1505 276 0 FreeSans 340 0 0 0 S
port 3 nsew
flabel corelocali s 1567 242 1601 276 0 FreeSans 340 0 0 0 S
port 3 nsew
flabel corelocali s 1663 242 1697 276 0 FreeSans 340 0 0 0 S
port 3 nsew
flabel corelocali s 1759 242 1793 276 0 FreeSans 340 0 0 0 S
port 3 nsew
flabel corelocali s 1855 242 1889 276 0 FreeSans 340 0 0 0 S
port 3 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 A0
port 1 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 A0
port 1 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 A1
port 2 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A1
port 2 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A1
port 2 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 Y
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 2016 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 2005184
string GDS_START 1990824
<< end >>
