magic
tech sky130A
magscale 1 2
timestamp 1599588232
<< locali >>
rect 353 390 463 596
rect 217 352 263 356
rect 91 286 263 352
rect 313 270 395 356
rect 429 236 463 390
rect 354 96 463 236
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 78 420 144 516
rect 22 386 144 420
rect 185 390 251 649
rect 22 250 56 386
rect 22 112 154 250
rect 22 51 156 112
rect 190 17 256 252
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< metal1 >>
rect 0 683 480 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 0 617 480 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 480 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
rect 0 -49 480 -17
<< labels >>
rlabel locali s 313 270 395 356 6 A
port 1 nsew signal input
rlabel locali s 217 352 263 356 6 TE_B
port 2 nsew signal input
rlabel locali s 91 286 263 352 6 TE_B
port 2 nsew signal input
rlabel locali s 429 236 463 390 6 Z
port 3 nsew signal output
rlabel locali s 354 96 463 236 6 Z
port 3 nsew signal output
rlabel locali s 353 390 463 596 6 Z
port 3 nsew signal output
rlabel metal1 s 0 -49 480 49 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 5 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 617 480 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 480 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 2354780
string GDS_START 2349956
<< end >>
