magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1472 561
rect 103 435 169 527
rect 280 435 325 527
rect 439 435 505 527
rect 761 436 827 527
rect 1049 434 1117 527
rect 24 199 68 331
rect 230 298 532 332
rect 230 199 279 298
rect 489 264 532 298
rect 661 298 965 332
rect 661 264 720 298
rect 931 264 965 298
rect 1151 333 1185 493
rect 1219 367 1283 527
rect 1317 333 1355 493
rect 1389 367 1454 527
rect 1151 299 1455 333
rect 355 215 443 264
rect 489 216 564 264
rect 629 249 720 264
rect 826 249 897 264
rect 498 215 564 216
rect 627 215 720 249
rect 778 215 897 249
rect 931 215 997 264
rect 1401 173 1455 299
rect 622 17 688 97
rect 799 17 873 97
rect 1130 139 1455 173
rect 1007 17 1060 109
rect 1130 51 1175 139
rect 1215 17 1275 105
rect 1309 51 1349 139
rect 1383 17 1455 105
rect 0 -17 1472 17
<< obsli1 >>
rect 18 401 69 493
rect 203 401 246 493
rect 359 401 405 493
rect 539 401 657 493
rect 955 401 1013 493
rect 18 400 1013 401
rect 18 367 1110 400
rect 103 366 1110 367
rect 20 97 69 165
rect 103 131 172 366
rect 1076 264 1110 366
rect 1076 215 1352 264
rect 344 131 959 177
rect 20 51 588 97
rect 722 51 765 131
rect 907 51 959 131
<< metal1 >>
rect 0 496 1472 592
rect 0 -48 1472 48
<< labels >>
rlabel locali s 826 249 897 264 6 A1
port 1 nsew signal input
rlabel locali s 778 215 897 249 6 A1
port 1 nsew signal input
rlabel locali s 931 264 965 298 6 A2
port 2 nsew signal input
rlabel locali s 931 215 997 264 6 A2
port 2 nsew signal input
rlabel locali s 661 298 965 332 6 A2
port 2 nsew signal input
rlabel locali s 661 264 720 298 6 A2
port 2 nsew signal input
rlabel locali s 629 249 720 264 6 A2
port 2 nsew signal input
rlabel locali s 627 215 720 249 6 A2
port 2 nsew signal input
rlabel locali s 355 215 443 264 6 B1
port 3 nsew signal input
rlabel locali s 498 215 564 216 6 C1
port 4 nsew signal input
rlabel locali s 489 264 532 298 6 C1
port 4 nsew signal input
rlabel locali s 489 216 564 264 6 C1
port 4 nsew signal input
rlabel locali s 230 298 532 332 6 C1
port 4 nsew signal input
rlabel locali s 230 199 279 298 6 C1
port 4 nsew signal input
rlabel locali s 24 199 68 331 6 D1
port 5 nsew signal input
rlabel locali s 1401 173 1455 299 6 X
port 6 nsew signal output
rlabel locali s 1317 333 1355 493 6 X
port 6 nsew signal output
rlabel locali s 1309 51 1349 139 6 X
port 6 nsew signal output
rlabel locali s 1151 333 1185 493 6 X
port 6 nsew signal output
rlabel locali s 1151 299 1455 333 6 X
port 6 nsew signal output
rlabel locali s 1130 139 1455 173 6 X
port 6 nsew signal output
rlabel locali s 1130 51 1175 139 6 X
port 6 nsew signal output
rlabel locali s 1383 17 1455 105 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1215 17 1275 105 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1007 17 1060 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 799 17 873 97 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 622 17 688 97 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 1472 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1472 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1389 367 1454 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1219 367 1283 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1049 434 1117 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 761 436 827 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 439 435 505 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 280 435 325 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 103 435 169 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 1472 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 1472 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1472 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1248064
string GDS_START 1237138
<< end >>
