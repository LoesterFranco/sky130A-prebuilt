magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 1050 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 89 47 119 177
rect 183 47 213 177
rect 267 47 297 177
rect 371 47 401 177
rect 569 47 599 177
rect 663 47 693 177
rect 767 47 797 177
rect 871 47 901 177
<< pmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 561 297 597 497
rect 655 297 691 497
rect 769 297 805 497
rect 863 297 899 497
<< ndiff >>
rect 27 131 89 177
rect 27 97 35 131
rect 69 97 89 131
rect 27 47 89 97
rect 119 97 183 177
rect 119 63 129 97
rect 163 63 183 97
rect 119 47 183 63
rect 213 131 267 177
rect 213 97 223 131
rect 257 97 267 131
rect 213 47 267 97
rect 297 169 371 177
rect 297 135 317 169
rect 351 135 371 169
rect 297 47 371 135
rect 401 101 453 177
rect 401 67 411 101
rect 445 67 453 101
rect 401 47 453 67
rect 507 101 569 177
rect 507 67 515 101
rect 549 67 569 101
rect 507 47 569 67
rect 599 169 663 177
rect 599 135 609 169
rect 643 135 663 169
rect 599 47 663 135
rect 693 131 767 177
rect 693 97 723 131
rect 757 97 767 131
rect 693 47 767 97
rect 797 97 871 177
rect 797 63 817 97
rect 851 63 871 97
rect 797 47 871 63
rect 901 131 953 177
rect 901 97 911 131
rect 945 97 953 131
rect 901 47 953 97
<< pdiff >>
rect 27 445 81 497
rect 27 411 35 445
rect 69 411 81 445
rect 27 377 81 411
rect 27 343 35 377
rect 69 343 81 377
rect 27 297 81 343
rect 117 485 175 497
rect 117 451 129 485
rect 163 451 175 485
rect 117 417 175 451
rect 117 383 129 417
rect 163 383 175 417
rect 117 297 175 383
rect 211 417 269 497
rect 211 383 223 417
rect 257 383 269 417
rect 211 349 269 383
rect 211 315 223 349
rect 257 315 269 349
rect 211 297 269 315
rect 305 485 363 497
rect 305 451 317 485
rect 351 451 363 485
rect 305 417 363 451
rect 305 383 317 417
rect 351 383 363 417
rect 305 297 363 383
rect 399 417 453 497
rect 399 383 411 417
rect 445 383 453 417
rect 399 349 453 383
rect 399 315 411 349
rect 445 315 453 349
rect 399 297 453 315
rect 507 485 561 497
rect 507 451 515 485
rect 549 451 561 485
rect 507 417 561 451
rect 507 383 515 417
rect 549 383 561 417
rect 507 349 561 383
rect 507 315 515 349
rect 549 315 561 349
rect 507 297 561 315
rect 597 485 655 497
rect 597 451 609 485
rect 643 451 655 485
rect 597 417 655 451
rect 597 383 609 417
rect 643 383 655 417
rect 597 297 655 383
rect 691 485 769 497
rect 691 451 723 485
rect 757 451 769 485
rect 691 417 769 451
rect 691 383 723 417
rect 757 383 769 417
rect 691 349 769 383
rect 691 315 723 349
rect 757 315 769 349
rect 691 297 769 315
rect 805 485 863 497
rect 805 451 817 485
rect 851 451 863 485
rect 805 417 863 451
rect 805 383 817 417
rect 851 383 863 417
rect 805 297 863 383
rect 899 485 953 497
rect 899 451 911 485
rect 945 451 953 485
rect 899 417 953 451
rect 899 383 911 417
rect 945 383 953 417
rect 899 349 953 383
rect 899 315 911 349
rect 945 315 953 349
rect 899 297 953 315
<< ndiffc >>
rect 35 97 69 131
rect 129 63 163 97
rect 223 97 257 131
rect 317 135 351 169
rect 411 67 445 101
rect 515 67 549 101
rect 609 135 643 169
rect 723 97 757 131
rect 817 63 851 97
rect 911 97 945 131
<< pdiffc >>
rect 35 411 69 445
rect 35 343 69 377
rect 129 451 163 485
rect 129 383 163 417
rect 223 383 257 417
rect 223 315 257 349
rect 317 451 351 485
rect 317 383 351 417
rect 411 383 445 417
rect 411 315 445 349
rect 515 451 549 485
rect 515 383 549 417
rect 515 315 549 349
rect 609 451 643 485
rect 609 383 643 417
rect 723 451 757 485
rect 723 383 757 417
rect 723 315 757 349
rect 817 451 851 485
rect 817 383 851 417
rect 911 451 945 485
rect 911 383 945 417
rect 911 315 945 349
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 561 497 597 523
rect 655 497 691 523
rect 769 497 805 523
rect 863 497 899 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 561 282 597 297
rect 655 282 691 297
rect 769 282 805 297
rect 863 282 899 297
rect 79 265 119 282
rect 173 265 213 282
rect 55 249 213 265
rect 55 215 65 249
rect 99 215 213 249
rect 55 199 213 215
rect 89 177 119 199
rect 183 177 213 199
rect 267 265 307 282
rect 361 265 401 282
rect 559 265 599 282
rect 653 265 693 282
rect 267 249 401 265
rect 267 215 283 249
rect 317 215 401 249
rect 267 199 401 215
rect 535 249 693 265
rect 535 215 545 249
rect 579 215 693 249
rect 535 199 693 215
rect 267 177 297 199
rect 371 177 401 199
rect 569 177 599 199
rect 663 177 693 199
rect 767 265 807 282
rect 861 265 901 282
rect 767 249 901 265
rect 767 215 783 249
rect 817 215 901 249
rect 767 199 901 215
rect 767 177 797 199
rect 871 177 901 199
rect 89 21 119 47
rect 183 21 213 47
rect 267 21 297 47
rect 371 21 401 47
rect 569 21 599 47
rect 663 21 693 47
rect 767 21 797 47
rect 871 21 901 47
<< polycont >>
rect 65 215 99 249
rect 283 215 317 249
rect 545 215 579 249
rect 783 215 817 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 19 445 69 493
rect 19 411 35 445
rect 19 377 69 411
rect 19 343 35 377
rect 103 485 565 493
rect 103 451 129 485
rect 163 459 317 485
rect 103 417 163 451
rect 351 459 515 485
rect 103 383 129 417
rect 103 365 163 383
rect 197 417 273 425
rect 197 383 223 417
rect 257 383 273 417
rect 19 331 69 343
rect 197 349 273 383
rect 317 417 351 451
rect 549 451 565 485
rect 317 365 351 383
rect 385 417 472 425
rect 385 383 411 417
rect 445 383 472 417
rect 197 331 223 349
rect 19 315 223 331
rect 257 331 273 349
rect 385 349 472 383
rect 385 331 411 349
rect 257 315 411 331
rect 445 315 472 349
rect 19 297 472 315
rect 515 417 565 451
rect 549 383 565 417
rect 515 349 565 383
rect 609 485 643 527
rect 609 417 643 451
rect 609 365 643 383
rect 677 485 773 493
rect 677 451 723 485
rect 757 451 773 485
rect 677 417 773 451
rect 677 383 723 417
rect 757 383 773 417
rect 549 331 565 349
rect 677 349 773 383
rect 817 485 851 527
rect 817 417 851 451
rect 817 365 851 383
rect 885 485 961 493
rect 885 451 911 485
rect 945 451 961 485
rect 885 417 961 451
rect 885 383 911 417
rect 945 383 961 417
rect 677 331 723 349
rect 549 315 723 331
rect 757 331 773 349
rect 885 349 961 383
rect 885 331 911 349
rect 757 315 911 331
rect 945 315 961 349
rect 515 297 961 315
rect 30 249 166 255
rect 30 215 65 249
rect 99 215 166 249
rect 206 249 349 255
rect 206 215 283 249
rect 317 215 349 249
rect 19 136 257 170
rect 386 169 472 297
rect 529 249 707 255
rect 529 215 545 249
rect 579 215 707 249
rect 754 249 924 255
rect 754 215 783 249
rect 817 215 924 249
rect 19 131 69 136
rect 19 97 35 131
rect 223 131 257 136
rect 291 135 317 169
rect 351 135 609 169
rect 643 135 659 169
rect 723 136 975 170
rect 19 51 69 97
rect 103 97 179 102
rect 103 63 129 97
rect 163 63 179 97
rect 103 17 179 63
rect 723 131 757 136
rect 257 97 411 101
rect 223 67 411 97
rect 445 67 461 101
rect 223 51 461 67
rect 499 67 515 101
rect 549 97 723 101
rect 911 131 975 136
rect 549 67 757 97
rect 499 51 757 67
rect 796 97 872 102
rect 796 63 817 97
rect 851 63 872 97
rect 796 17 872 63
rect 945 97 975 131
rect 911 51 975 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
flabel corelocali s 664 221 698 255 0 FreeSans 200 0 0 0 A1
port 1 nsew
flabel corelocali s 585 221 619 255 0 FreeSans 200 0 0 0 A1
port 1 nsew
flabel corelocali s 758 221 792 255 0 FreeSans 200 0 0 0 A2
port 2 nsew
flabel corelocali s 860 221 894 255 0 FreeSans 200 0 0 0 A2
port 2 nsew
flabel corelocali s 304 221 338 255 0 FreeSans 200 0 0 0 B1
port 3 nsew
flabel corelocali s 121 221 155 255 0 FreeSans 200 0 0 0 B2
port 4 nsew
flabel corelocali s 397 153 431 187 0 FreeSans 200 0 0 0 Y
port 9 nsew
flabel corelocali s 397 221 431 255 0 FreeSans 200 0 0 0 Y
port 9 nsew
flabel corelocali s 397 357 431 391 0 FreeSans 200 0 0 0 Y
port 9 nsew
flabel corelocali s 397 289 431 323 0 FreeSans 200 0 0 0 Y
port 9 nsew
flabel corelocali s 132 527 166 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
flabel corelocali s 132 -17 166 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 200 0 0 0 B2
port 4 nsew
flabel corelocali s 217 221 251 255 0 FreeSans 200 0 0 0 B1
port 3 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
rlabel comment s 0 0 0 0 4 a22oi_2
<< properties >>
string FIXED_BBOX 0 0 1012 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1291754
string GDS_START 1282852
<< end >>
