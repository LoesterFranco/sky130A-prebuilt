magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 828 561
rect 120 427 186 527
rect 17 212 111 325
rect 510 427 576 527
rect 614 297 710 493
rect 744 297 811 527
rect 117 17 183 110
rect 671 128 710 297
rect 510 17 576 113
rect 610 51 710 128
rect 744 17 811 129
rect 0 -17 828 17
<< obsli1 >>
rect 17 393 86 493
rect 17 359 212 393
rect 178 249 212 359
rect 246 357 332 493
rect 366 393 420 493
rect 366 358 580 393
rect 298 297 332 357
rect 178 215 264 249
rect 298 215 483 297
rect 546 249 580 358
rect 546 215 637 249
rect 178 178 212 215
rect 298 181 332 215
rect 546 181 580 215
rect 17 144 212 178
rect 17 51 83 144
rect 256 51 332 181
rect 366 147 580 181
rect 366 51 420 147
<< metal1 >>
rect 0 496 828 592
rect 0 -48 828 48
<< labels >>
rlabel locali s 17 212 111 325 6 A
port 1 nsew signal input
rlabel locali s 671 128 710 297 6 X
port 2 nsew signal output
rlabel locali s 614 297 710 493 6 X
port 2 nsew signal output
rlabel locali s 610 51 710 128 6 X
port 2 nsew signal output
rlabel locali s 744 17 811 129 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 510 17 576 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 117 17 183 110 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 0 -17 828 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 828 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 744 297 811 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 510 427 576 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 120 427 186 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 0 527 828 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 496 828 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3148896
string GDS_START 3142330
<< end >>
