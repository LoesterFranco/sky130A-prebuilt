magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 1766 704
<< pwell >>
rect 0 0 1728 49
<< scnmos >>
rect 145 74 175 222
rect 231 74 261 222
rect 317 74 347 222
rect 403 74 433 222
rect 489 74 519 222
rect 575 74 605 222
rect 661 74 691 222
rect 747 74 777 222
rect 1137 74 1167 222
rect 1223 74 1253 222
rect 1309 74 1339 222
rect 1395 74 1425 222
<< pmoshvt >>
rect 132 368 162 592
rect 222 368 252 592
rect 312 368 342 592
rect 402 368 432 592
rect 492 368 522 592
rect 582 368 612 592
rect 672 368 702 592
rect 762 368 792 592
rect 956 368 986 592
rect 1046 368 1076 592
rect 1136 368 1166 592
rect 1226 368 1256 592
rect 1316 368 1346 592
rect 1406 368 1436 592
rect 1496 368 1526 592
rect 1586 368 1616 592
<< ndiff >>
rect 92 210 145 222
rect 92 176 100 210
rect 134 176 145 210
rect 92 120 145 176
rect 92 86 100 120
rect 134 86 145 120
rect 92 74 145 86
rect 175 152 231 222
rect 175 118 186 152
rect 220 118 231 152
rect 175 74 231 118
rect 261 210 317 222
rect 261 176 272 210
rect 306 176 317 210
rect 261 120 317 176
rect 261 86 272 120
rect 306 86 317 120
rect 261 74 317 86
rect 347 152 403 222
rect 347 118 358 152
rect 392 118 403 152
rect 347 74 403 118
rect 433 210 489 222
rect 433 176 444 210
rect 478 176 489 210
rect 433 120 489 176
rect 433 86 444 120
rect 478 86 489 120
rect 433 74 489 86
rect 519 207 575 222
rect 519 173 530 207
rect 564 173 575 207
rect 519 74 575 173
rect 605 120 661 222
rect 605 86 616 120
rect 650 86 661 120
rect 605 74 661 86
rect 691 207 747 222
rect 691 173 702 207
rect 736 173 747 207
rect 691 74 747 173
rect 777 120 834 222
rect 777 86 788 120
rect 822 86 834 120
rect 777 74 834 86
rect 1084 210 1137 222
rect 1084 176 1092 210
rect 1126 176 1137 210
rect 1084 120 1137 176
rect 1084 86 1092 120
rect 1126 86 1137 120
rect 1084 74 1137 86
rect 1167 142 1223 222
rect 1167 108 1178 142
rect 1212 108 1223 142
rect 1167 74 1223 108
rect 1253 210 1309 222
rect 1253 176 1264 210
rect 1298 176 1309 210
rect 1253 120 1309 176
rect 1253 86 1264 120
rect 1298 86 1309 120
rect 1253 74 1309 86
rect 1339 152 1395 222
rect 1339 118 1350 152
rect 1384 118 1395 152
rect 1339 74 1395 118
rect 1425 210 1478 222
rect 1425 176 1436 210
rect 1470 176 1478 210
rect 1425 120 1478 176
rect 1425 86 1436 120
rect 1470 86 1478 120
rect 1425 74 1478 86
<< pdiff >>
rect 77 580 132 592
rect 77 546 85 580
rect 119 546 132 580
rect 77 506 132 546
rect 77 472 85 506
rect 119 472 132 506
rect 77 424 132 472
rect 77 390 85 424
rect 119 390 132 424
rect 77 368 132 390
rect 162 580 222 592
rect 162 546 175 580
rect 209 546 222 580
rect 162 508 222 546
rect 162 474 175 508
rect 209 474 222 508
rect 162 368 222 474
rect 252 580 312 592
rect 252 546 265 580
rect 299 546 312 580
rect 252 506 312 546
rect 252 472 265 506
rect 299 472 312 506
rect 252 424 312 472
rect 252 390 265 424
rect 299 390 312 424
rect 252 368 312 390
rect 342 580 402 592
rect 342 546 355 580
rect 389 546 402 580
rect 342 499 402 546
rect 342 465 355 499
rect 389 465 402 499
rect 342 368 402 465
rect 432 580 492 592
rect 432 546 445 580
rect 479 546 492 580
rect 432 506 492 546
rect 432 472 445 506
rect 479 472 492 506
rect 432 424 492 472
rect 432 390 445 424
rect 479 390 492 424
rect 432 368 492 390
rect 522 580 582 592
rect 522 546 535 580
rect 569 546 582 580
rect 522 499 582 546
rect 522 465 535 499
rect 569 465 582 499
rect 522 368 582 465
rect 612 580 672 592
rect 612 546 625 580
rect 659 546 672 580
rect 612 506 672 546
rect 612 472 625 506
rect 659 472 672 506
rect 612 424 672 472
rect 612 390 625 424
rect 659 390 672 424
rect 612 368 672 390
rect 702 580 762 592
rect 702 546 715 580
rect 749 546 762 580
rect 702 499 762 546
rect 702 465 715 499
rect 749 465 762 499
rect 702 368 762 465
rect 792 580 847 592
rect 792 546 805 580
rect 839 546 847 580
rect 792 497 847 546
rect 792 463 805 497
rect 839 463 847 497
rect 792 414 847 463
rect 792 380 805 414
rect 839 380 847 414
rect 792 368 847 380
rect 901 580 956 592
rect 901 546 909 580
rect 943 546 956 580
rect 901 496 956 546
rect 901 462 909 496
rect 943 462 956 496
rect 901 368 956 462
rect 986 531 1046 592
rect 986 497 999 531
rect 1033 497 1046 531
rect 986 424 1046 497
rect 986 390 999 424
rect 1033 390 1046 424
rect 986 368 1046 390
rect 1076 584 1136 592
rect 1076 550 1089 584
rect 1123 550 1136 584
rect 1076 496 1136 550
rect 1076 462 1089 496
rect 1123 462 1136 496
rect 1076 368 1136 462
rect 1166 531 1226 592
rect 1166 497 1179 531
rect 1213 497 1226 531
rect 1166 424 1226 497
rect 1166 390 1179 424
rect 1213 390 1226 424
rect 1166 368 1226 390
rect 1256 580 1316 592
rect 1256 546 1269 580
rect 1303 546 1316 580
rect 1256 510 1316 546
rect 1256 476 1269 510
rect 1303 476 1316 510
rect 1256 440 1316 476
rect 1256 406 1269 440
rect 1303 406 1316 440
rect 1256 368 1316 406
rect 1346 531 1406 592
rect 1346 497 1359 531
rect 1393 497 1406 531
rect 1346 440 1406 497
rect 1346 406 1359 440
rect 1393 406 1406 440
rect 1346 368 1406 406
rect 1436 580 1496 592
rect 1436 546 1449 580
rect 1483 546 1496 580
rect 1436 508 1496 546
rect 1436 474 1449 508
rect 1483 474 1496 508
rect 1436 368 1496 474
rect 1526 531 1586 592
rect 1526 497 1539 531
rect 1573 497 1586 531
rect 1526 440 1586 497
rect 1526 406 1539 440
rect 1573 406 1586 440
rect 1526 368 1586 406
rect 1616 580 1671 592
rect 1616 546 1629 580
rect 1663 546 1671 580
rect 1616 474 1671 546
rect 1616 440 1629 474
rect 1663 440 1671 474
rect 1616 368 1671 440
<< ndiffc >>
rect 100 176 134 210
rect 100 86 134 120
rect 186 118 220 152
rect 272 176 306 210
rect 272 86 306 120
rect 358 118 392 152
rect 444 176 478 210
rect 444 86 478 120
rect 530 173 564 207
rect 616 86 650 120
rect 702 173 736 207
rect 788 86 822 120
rect 1092 176 1126 210
rect 1092 86 1126 120
rect 1178 108 1212 142
rect 1264 176 1298 210
rect 1264 86 1298 120
rect 1350 118 1384 152
rect 1436 176 1470 210
rect 1436 86 1470 120
<< pdiffc >>
rect 85 546 119 580
rect 85 472 119 506
rect 85 390 119 424
rect 175 546 209 580
rect 175 474 209 508
rect 265 546 299 580
rect 265 472 299 506
rect 265 390 299 424
rect 355 546 389 580
rect 355 465 389 499
rect 445 546 479 580
rect 445 472 479 506
rect 445 390 479 424
rect 535 546 569 580
rect 535 465 569 499
rect 625 546 659 580
rect 625 472 659 506
rect 625 390 659 424
rect 715 546 749 580
rect 715 465 749 499
rect 805 546 839 580
rect 805 463 839 497
rect 805 380 839 414
rect 909 546 943 580
rect 909 462 943 496
rect 999 497 1033 531
rect 999 390 1033 424
rect 1089 550 1123 584
rect 1089 462 1123 496
rect 1179 497 1213 531
rect 1179 390 1213 424
rect 1269 546 1303 580
rect 1269 476 1303 510
rect 1269 406 1303 440
rect 1359 497 1393 531
rect 1359 406 1393 440
rect 1449 546 1483 580
rect 1449 474 1483 508
rect 1539 497 1573 531
rect 1539 406 1573 440
rect 1629 546 1663 580
rect 1629 440 1663 474
<< poly >>
rect 132 592 162 618
rect 222 592 252 618
rect 312 592 342 618
rect 402 592 432 618
rect 492 592 522 618
rect 582 592 612 618
rect 672 592 702 618
rect 762 592 792 618
rect 956 592 986 618
rect 1046 592 1076 618
rect 1136 592 1166 618
rect 1226 592 1256 618
rect 1316 592 1346 618
rect 1406 592 1436 618
rect 1496 592 1526 618
rect 1586 592 1616 618
rect 132 353 162 368
rect 222 353 252 368
rect 312 353 342 368
rect 402 353 432 368
rect 492 353 522 368
rect 582 353 612 368
rect 672 353 702 368
rect 762 353 792 368
rect 956 353 986 368
rect 1046 353 1076 368
rect 1136 353 1166 368
rect 1226 353 1256 368
rect 1316 353 1346 368
rect 1406 353 1436 368
rect 1496 353 1526 368
rect 1586 353 1616 368
rect 129 336 165 353
rect 219 336 255 353
rect 309 336 345 353
rect 399 336 435 353
rect 129 320 435 336
rect 129 286 145 320
rect 179 286 213 320
rect 247 286 281 320
rect 315 286 349 320
rect 383 286 435 320
rect 129 270 435 286
rect 489 336 525 353
rect 579 336 615 353
rect 669 336 705 353
rect 759 336 795 353
rect 489 320 795 336
rect 489 286 517 320
rect 551 286 585 320
rect 619 286 653 320
rect 687 286 721 320
rect 755 286 795 320
rect 489 270 795 286
rect 953 326 989 353
rect 1043 326 1079 353
rect 1133 326 1169 353
rect 1223 326 1259 353
rect 1313 336 1349 353
rect 1403 336 1439 353
rect 1493 336 1529 353
rect 1583 336 1619 353
rect 953 310 1259 326
rect 953 276 969 310
rect 1003 276 1037 310
rect 1071 276 1105 310
rect 1139 276 1173 310
rect 1207 276 1259 310
rect 145 222 175 270
rect 231 222 261 270
rect 317 222 347 270
rect 403 222 433 270
rect 489 222 519 270
rect 575 222 605 270
rect 661 222 691 270
rect 747 222 777 270
rect 953 264 1259 276
rect 1309 320 1619 336
rect 1309 286 1325 320
rect 1359 286 1393 320
rect 1427 286 1461 320
rect 1495 286 1619 320
rect 1309 264 1619 286
rect 953 260 1253 264
rect 1137 222 1167 260
rect 1223 222 1253 260
rect 1309 222 1339 264
rect 1395 222 1425 264
rect 145 48 175 74
rect 231 48 261 74
rect 317 48 347 74
rect 403 48 433 74
rect 489 48 519 74
rect 575 48 605 74
rect 661 48 691 74
rect 747 48 777 74
rect 1137 48 1167 74
rect 1223 48 1253 74
rect 1309 48 1339 74
rect 1395 48 1425 74
<< polycont >>
rect 145 286 179 320
rect 213 286 247 320
rect 281 286 315 320
rect 349 286 383 320
rect 517 286 551 320
rect 585 286 619 320
rect 653 286 687 320
rect 721 286 755 320
rect 969 276 1003 310
rect 1037 276 1071 310
rect 1105 276 1139 310
rect 1173 276 1207 310
rect 1325 286 1359 320
rect 1393 286 1427 320
rect 1461 286 1495 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 69 580 135 596
rect 69 546 85 580
rect 119 546 135 580
rect 69 506 135 546
rect 69 472 85 506
rect 119 472 135 506
rect 69 424 135 472
rect 175 580 209 649
rect 175 508 209 546
rect 175 458 209 474
rect 249 580 299 596
rect 249 546 265 580
rect 249 506 299 546
rect 249 472 265 506
rect 249 424 299 472
rect 339 580 405 649
rect 339 546 355 580
rect 389 546 405 580
rect 339 499 405 546
rect 339 465 355 499
rect 389 465 405 499
rect 339 458 405 465
rect 445 580 479 596
rect 445 506 479 546
rect 445 424 479 472
rect 519 580 585 649
rect 519 546 535 580
rect 569 546 585 580
rect 519 499 585 546
rect 519 465 535 499
rect 569 465 585 499
rect 519 458 585 465
rect 625 580 659 596
rect 625 506 659 546
rect 625 424 659 472
rect 699 580 765 649
rect 699 546 715 580
rect 749 546 765 580
rect 699 499 765 546
rect 699 465 715 499
rect 749 465 765 499
rect 699 458 765 465
rect 805 580 855 596
rect 839 546 855 580
rect 805 497 855 546
rect 839 463 855 497
rect 805 424 855 463
rect 893 584 1679 615
rect 893 581 1089 584
rect 893 580 959 581
rect 893 546 909 580
rect 943 546 959 580
rect 1073 550 1089 581
rect 1123 581 1679 584
rect 1123 550 1139 581
rect 893 496 959 546
rect 893 462 909 496
rect 943 462 959 496
rect 893 458 959 462
rect 999 531 1033 547
rect 999 424 1033 497
rect 1073 496 1139 550
rect 1263 580 1319 581
rect 1073 462 1089 496
rect 1123 462 1139 496
rect 1073 458 1139 462
rect 1179 531 1229 547
rect 1213 497 1229 531
rect 1179 424 1229 497
rect 69 390 85 424
rect 119 390 265 424
rect 299 390 445 424
rect 479 390 625 424
rect 659 414 999 424
rect 659 390 805 414
rect 839 390 999 414
rect 1033 390 1179 424
rect 1213 390 1229 424
rect 1263 546 1269 580
rect 1303 546 1319 580
rect 1433 580 1499 581
rect 1263 510 1319 546
rect 1263 476 1269 510
rect 1303 476 1319 510
rect 1263 440 1319 476
rect 1263 406 1269 440
rect 1303 406 1319 440
rect 1263 390 1319 406
rect 1359 531 1393 547
rect 1359 440 1393 497
rect 1433 546 1449 580
rect 1483 546 1499 580
rect 1613 580 1679 581
rect 1433 508 1499 546
rect 1433 474 1449 508
rect 1483 474 1499 508
rect 1433 458 1499 474
rect 1539 531 1579 547
rect 1573 497 1579 531
rect 1539 440 1579 497
rect 1393 406 1539 424
rect 1573 406 1579 440
rect 1613 546 1629 580
rect 1663 546 1679 580
rect 1613 474 1679 546
rect 1613 440 1629 474
rect 1663 440 1679 474
rect 1613 424 1679 440
rect 1359 390 1579 406
rect 839 380 855 390
rect 805 364 855 380
rect 25 320 455 356
rect 25 286 145 320
rect 179 286 213 320
rect 247 286 281 320
rect 315 286 349 320
rect 383 286 455 320
rect 25 270 455 286
rect 501 320 771 356
rect 501 286 517 320
rect 551 286 585 320
rect 619 286 653 320
rect 687 286 721 320
rect 755 286 771 320
rect 501 270 771 286
rect 889 310 1223 356
rect 889 276 969 310
rect 1003 276 1037 310
rect 1071 276 1105 310
rect 1139 276 1173 310
rect 1207 276 1223 310
rect 889 260 1223 276
rect 1273 320 1511 356
rect 1273 286 1325 320
rect 1359 286 1393 320
rect 1427 286 1461 320
rect 1495 286 1511 320
rect 1273 270 1511 286
rect 1545 236 1703 390
rect 84 210 478 236
rect 1264 226 1703 236
rect 84 176 100 210
rect 134 202 272 210
rect 84 120 134 176
rect 306 202 444 210
rect 84 86 100 120
rect 84 70 134 86
rect 170 152 236 168
rect 170 118 186 152
rect 220 118 236 152
rect 170 17 236 118
rect 272 120 306 176
rect 272 70 306 86
rect 342 152 408 168
rect 342 118 358 152
rect 392 118 408 152
rect 342 17 408 118
rect 444 123 478 176
rect 514 210 1703 226
rect 514 207 1092 210
rect 514 173 530 207
rect 564 173 702 207
rect 736 192 1092 207
rect 736 173 752 192
rect 514 157 752 173
rect 1076 176 1092 192
rect 1126 192 1264 210
rect 444 120 838 123
rect 478 86 616 120
rect 650 86 788 120
rect 822 86 838 120
rect 444 70 838 86
rect 1076 120 1126 176
rect 1298 202 1436 210
rect 1076 86 1092 120
rect 1076 70 1126 86
rect 1162 142 1228 158
rect 1162 108 1178 142
rect 1212 108 1228 142
rect 1162 17 1228 108
rect 1264 120 1298 176
rect 1470 176 1703 210
rect 1264 70 1298 86
rect 1334 152 1400 168
rect 1334 118 1350 152
rect 1384 118 1400 152
rect 1334 17 1400 118
rect 1436 120 1703 176
rect 1470 86 1703 120
rect 1436 70 1703 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
<< metal1 >>
rect 0 683 1728 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 0 617 1728 649
rect 0 17 1728 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
rect 0 -49 1728 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a211oi_4
flabel pwell s 0 0 1728 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 1728 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 1728 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 1728 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 1567 94 1601 128 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 1567 168 1601 202 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 1567 242 1601 276 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 1567 316 1601 350 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 1663 94 1697 128 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 1663 168 1697 202 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 1663 242 1697 276 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 1663 316 1697 350 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 1279 316 1313 350 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 1375 316 1409 350 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 1471 316 1505 350 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 1087 316 1121 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 1183 316 1217 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 1728 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 4071700
string GDS_START 4057012
<< end >>
