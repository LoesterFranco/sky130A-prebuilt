magic
tech sky130A
magscale 1 2
timestamp 1599588244
<< locali >>
rect 25 364 180 596
rect 25 226 100 364
rect 275 270 359 356
rect 393 294 459 360
rect 505 291 597 356
rect 639 291 743 356
rect 25 70 173 226
rect 773 51 839 134
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 220 390 270 649
rect 307 428 357 596
rect 397 462 463 649
rect 501 581 737 615
rect 501 462 557 581
rect 591 428 657 547
rect 307 394 657 428
rect 307 390 357 394
rect 591 390 657 394
rect 697 390 737 581
rect 148 260 241 326
rect 207 236 241 260
rect 777 257 843 596
rect 493 236 843 257
rect 207 223 843 236
rect 207 202 572 223
rect 209 17 393 168
rect 484 75 572 202
rect 664 17 738 189
rect 772 168 843 223
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel locali s 393 294 459 360 6 A1
port 1 nsew signal input
rlabel locali s 275 270 359 356 6 A2
port 2 nsew signal input
rlabel locali s 505 291 597 356 6 B1
port 3 nsew signal input
rlabel locali s 639 291 743 356 6 B2
port 4 nsew signal input
rlabel locali s 773 51 839 134 6 C1
port 5 nsew signal input
rlabel locali s 25 364 180 596 6 X
port 6 nsew signal output
rlabel locali s 25 226 100 364 6 X
port 6 nsew signal output
rlabel locali s 25 70 173 226 6 X
port 6 nsew signal output
rlabel metal1 s 0 -49 864 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 8 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 9 nsew power bidirectional
rlabel metal1 s 0 617 864 715 6 VPWR
port 10 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 4026626
string GDS_START 4018346
<< end >>
