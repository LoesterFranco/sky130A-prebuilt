magic
tech sky130A
magscale 1 2
timestamp 1601050082
<< locali >>
rect 428 424 494 596
rect 876 424 942 596
rect 428 390 942 424
rect 409 270 839 356
rect 876 226 942 390
rect 1188 424 1254 596
rect 1464 424 1510 596
rect 1188 390 1579 424
rect 1193 310 1511 356
rect 1037 244 1511 310
rect 867 210 942 226
rect 1545 210 1579 390
rect 867 154 1579 210
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 132 390 394 649
rect 528 458 842 649
rect 21 236 372 271
rect 21 233 831 236
rect 21 70 71 233
rect 207 202 831 233
rect 976 364 1042 649
rect 1088 364 1154 649
rect 1288 458 1430 649
rect 1544 458 1610 649
rect 107 17 173 199
rect 207 70 245 202
rect 279 17 345 168
rect 379 70 431 202
rect 465 17 581 168
rect 615 70 661 202
rect 695 17 761 168
rect 797 120 831 202
rect 797 70 1609 120
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
rlabel locali s 1193 310 1511 356 6 A
port 1 nsew signal input
rlabel locali s 1037 244 1511 310 6 A
port 1 nsew signal input
rlabel locali s 409 270 839 356 6 B
port 2 nsew signal input
rlabel locali s 1545 210 1579 390 6 Y
port 3 nsew signal output
rlabel locali s 1464 424 1510 596 6 Y
port 3 nsew signal output
rlabel locali s 1188 424 1254 596 6 Y
port 3 nsew signal output
rlabel locali s 1188 390 1579 424 6 Y
port 3 nsew signal output
rlabel locali s 876 424 942 596 6 Y
port 3 nsew signal output
rlabel locali s 876 226 942 390 6 Y
port 3 nsew signal output
rlabel locali s 867 210 942 226 6 Y
port 3 nsew signal output
rlabel locali s 867 154 1579 210 6 Y
port 3 nsew signal output
rlabel locali s 428 424 494 596 6 Y
port 3 nsew signal output
rlabel locali s 428 390 942 424 6 Y
port 3 nsew signal output
rlabel metal1 s 0 -49 1632 49 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1632 715 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1645498
string GDS_START 1633406
<< end >>
