magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1196 561
rect 103 451 169 527
rect 282 451 348 527
rect 450 451 516 527
rect 666 451 732 527
rect 872 451 1074 527
rect 86 153 156 327
rect 192 309 432 343
rect 192 164 248 309
rect 192 130 416 164
rect 114 17 180 94
rect 214 51 248 130
rect 282 17 348 94
rect 382 51 416 130
rect 536 199 616 265
rect 650 151 709 265
rect 1097 199 1169 324
rect 454 17 520 89
rect 995 17 1061 93
rect 0 -17 1196 17
<< obsli1 >>
rect 17 417 69 493
rect 1127 417 1161 493
rect 17 383 898 417
rect 17 117 52 383
rect 466 309 830 343
rect 466 249 500 309
rect 864 265 898 383
rect 282 215 500 249
rect 17 51 69 117
rect 466 157 500 215
rect 466 123 588 157
rect 746 231 898 265
rect 990 383 1161 417
rect 746 199 780 231
rect 990 165 1024 383
rect 554 94 588 123
rect 851 94 922 162
rect 990 131 1161 165
rect 554 60 922 94
rect 1127 51 1161 131
<< metal1 >>
rect 0 496 1196 592
rect 0 -48 1196 48
<< labels >>
rlabel locali s 1097 199 1169 324 6 A_N
port 1 nsew signal input
rlabel locali s 86 153 156 327 6 B_N
port 2 nsew signal input
rlabel locali s 650 151 709 265 6 C
port 3 nsew signal input
rlabel locali s 536 199 616 265 6 D
port 4 nsew signal input
rlabel locali s 382 51 416 130 6 X
port 5 nsew signal output
rlabel locali s 214 51 248 130 6 X
port 5 nsew signal output
rlabel locali s 192 309 432 343 6 X
port 5 nsew signal output
rlabel locali s 192 164 248 309 6 X
port 5 nsew signal output
rlabel locali s 192 130 416 164 6 X
port 5 nsew signal output
rlabel locali s 995 17 1061 93 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 454 17 520 89 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 282 17 348 94 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 114 17 180 94 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 1196 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1196 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 872 451 1074 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 666 451 732 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 450 451 516 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 282 451 348 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 103 451 169 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 1196 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 1196 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3000766
string GDS_START 2992108
<< end >>
