magic
tech sky130A
magscale 1 2
timestamp 1604502705
<< nwell >>
rect -38 332 806 704
<< pwell >>
rect 0 0 768 49
<< scnmos >>
rect 84 100 114 248
rect 193 120 223 248
rect 271 120 301 248
rect 373 136 403 264
rect 451 136 481 264
rect 565 136 595 264
rect 649 136 679 264
<< pmoshvt >>
rect 95 368 125 592
rect 196 384 226 584
rect 280 384 310 584
rect 376 384 406 584
rect 460 384 490 584
rect 568 384 598 584
rect 652 384 682 584
<< ndiff >>
rect 323 248 373 264
rect 34 232 84 248
rect 27 220 84 232
rect 27 186 39 220
rect 73 186 84 220
rect 27 146 84 186
rect 27 112 39 146
rect 73 112 84 146
rect 27 100 84 112
rect 114 171 193 248
rect 114 137 143 171
rect 177 137 193 171
rect 114 120 193 137
rect 223 120 271 248
rect 301 236 373 248
rect 301 202 312 236
rect 346 202 373 236
rect 301 166 373 202
rect 301 132 312 166
rect 346 136 373 166
rect 403 136 451 264
rect 481 182 565 264
rect 481 148 506 182
rect 540 148 565 182
rect 481 136 565 148
rect 595 136 649 264
rect 679 248 729 264
rect 679 227 736 248
rect 679 193 690 227
rect 724 193 736 227
rect 679 172 736 193
rect 679 136 729 172
rect 346 132 358 136
rect 301 120 358 132
rect 114 100 164 120
<< pdiff >>
rect 36 580 95 592
rect 36 546 48 580
rect 82 546 95 580
rect 36 500 95 546
rect 36 466 48 500
rect 82 466 95 500
rect 36 420 95 466
rect 36 386 48 420
rect 82 386 95 420
rect 36 368 95 386
rect 125 584 178 592
rect 125 572 196 584
rect 125 538 148 572
rect 182 538 196 572
rect 125 504 196 538
rect 125 470 148 504
rect 182 470 196 504
rect 125 436 196 470
rect 125 402 148 436
rect 182 402 196 436
rect 125 384 196 402
rect 226 384 280 584
rect 310 572 376 584
rect 310 538 329 572
rect 363 538 376 572
rect 310 504 376 538
rect 310 470 329 504
rect 363 470 376 504
rect 310 436 376 470
rect 310 402 329 436
rect 363 402 376 436
rect 310 384 376 402
rect 406 384 460 584
rect 490 572 568 584
rect 490 538 511 572
rect 545 538 568 572
rect 490 492 568 538
rect 490 458 511 492
rect 545 458 568 492
rect 490 384 568 458
rect 598 384 652 584
rect 682 572 741 584
rect 682 538 695 572
rect 729 538 741 572
rect 682 504 741 538
rect 682 470 695 504
rect 729 470 741 504
rect 682 436 741 470
rect 682 402 695 436
rect 729 402 741 436
rect 682 384 741 402
rect 125 368 178 384
<< ndiffc >>
rect 39 186 73 220
rect 39 112 73 146
rect 143 137 177 171
rect 312 202 346 236
rect 312 132 346 166
rect 506 148 540 182
rect 690 193 724 227
<< pdiffc >>
rect 48 546 82 580
rect 48 466 82 500
rect 48 386 82 420
rect 148 538 182 572
rect 148 470 182 504
rect 148 402 182 436
rect 329 538 363 572
rect 329 470 363 504
rect 329 402 363 436
rect 511 538 545 572
rect 511 458 545 492
rect 695 538 729 572
rect 695 470 729 504
rect 695 402 729 436
<< poly >>
rect 95 592 125 618
rect 196 584 226 610
rect 280 584 310 610
rect 376 584 406 610
rect 460 584 490 610
rect 568 584 598 610
rect 652 584 682 610
rect 196 369 226 384
rect 280 369 310 384
rect 376 369 406 384
rect 460 369 490 384
rect 568 369 598 384
rect 652 369 682 384
rect 95 353 125 368
rect 92 336 128 353
rect 84 320 151 336
rect 84 286 101 320
rect 135 286 151 320
rect 84 270 151 286
rect 84 248 114 270
rect 193 263 229 369
rect 277 352 313 369
rect 373 352 409 369
rect 457 352 493 369
rect 271 336 409 352
rect 271 302 287 336
rect 321 302 409 336
rect 271 286 409 302
rect 451 336 523 352
rect 451 302 473 336
rect 507 302 523 336
rect 193 248 223 263
rect 271 248 301 286
rect 373 264 403 286
rect 451 280 523 302
rect 451 264 481 280
rect 565 279 601 369
rect 649 352 685 369
rect 649 336 715 352
rect 649 302 665 336
rect 699 302 715 336
rect 649 286 715 302
rect 565 264 595 279
rect 649 264 679 286
rect 84 74 114 100
rect 193 52 223 120
rect 271 94 301 120
rect 373 110 403 136
rect 451 110 481 136
rect 565 114 595 136
rect 529 98 595 114
rect 649 110 679 136
rect 529 64 545 98
rect 579 64 595 98
rect 529 52 595 64
rect 193 22 595 52
<< polycont >>
rect 101 286 135 320
rect 287 302 321 336
rect 473 302 507 336
rect 665 302 699 336
rect 545 64 579 98
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 17 580 98 596
rect 17 546 48 580
rect 82 546 98 580
rect 17 500 98 546
rect 17 466 48 500
rect 82 466 98 500
rect 17 420 98 466
rect 17 386 48 420
rect 82 386 98 420
rect 132 572 198 649
rect 132 538 148 572
rect 182 538 198 572
rect 132 504 198 538
rect 132 470 148 504
rect 182 470 198 504
rect 132 436 198 470
rect 132 402 148 436
rect 182 402 198 436
rect 132 390 198 402
rect 313 572 379 588
rect 313 538 329 572
rect 363 538 379 572
rect 313 504 379 538
rect 313 470 329 504
rect 363 470 379 504
rect 313 436 379 470
rect 487 572 568 649
rect 487 538 511 572
rect 545 538 568 572
rect 487 492 568 538
rect 487 458 511 492
rect 545 458 568 492
rect 679 572 745 588
rect 679 538 695 572
rect 729 538 745 572
rect 679 504 745 538
rect 679 470 695 504
rect 729 470 745 504
rect 313 402 329 436
rect 363 424 379 436
rect 679 436 745 470
rect 679 424 695 436
rect 363 402 695 424
rect 729 402 745 436
rect 313 390 745 402
rect 17 370 98 386
rect 17 236 51 370
rect 217 336 337 356
rect 85 320 157 336
rect 85 286 101 320
rect 135 286 157 320
rect 217 302 287 336
rect 321 302 337 336
rect 217 286 337 302
rect 85 270 157 286
rect 123 252 157 270
rect 379 252 413 390
rect 679 386 745 390
rect 457 352 551 356
rect 457 336 715 352
rect 457 302 473 336
rect 507 302 665 336
rect 699 302 715 336
rect 457 286 715 302
rect 123 236 740 252
rect 17 220 89 236
rect 17 186 39 220
rect 73 186 89 220
rect 123 218 312 236
rect 17 146 89 186
rect 296 202 312 218
rect 346 227 740 236
rect 346 218 690 227
rect 346 202 362 218
rect 17 112 39 146
rect 73 112 89 146
rect 17 96 89 112
rect 123 171 198 182
rect 123 137 143 171
rect 177 137 198 171
rect 123 17 198 137
rect 296 166 362 202
rect 674 193 690 218
rect 724 193 740 227
rect 296 132 312 166
rect 346 132 362 166
rect 296 116 362 132
rect 461 148 506 182
rect 540 148 570 182
rect 674 168 740 193
rect 461 17 495 148
rect 697 114 743 134
rect 529 98 743 114
rect 529 64 545 98
rect 579 64 743 98
rect 529 51 743 64
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel comment s 0 0 0 0 4 maj3_1
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 703 94 737 128 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 C
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 768 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2420170
string GDS_START 2413322
<< end >>
