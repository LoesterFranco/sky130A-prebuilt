magic
tech sky130A
magscale 1 2
timestamp 1604502705
<< nwell >>
rect -38 332 998 704
<< pwell >>
rect 0 0 960 49
<< scnmos >>
rect 118 74 148 222
rect 204 74 234 222
rect 304 74 334 222
rect 390 74 420 222
rect 528 74 558 222
rect 636 74 666 222
rect 722 74 752 222
rect 808 74 838 222
<< pmoshvt >>
rect 121 368 151 592
rect 211 368 241 592
rect 301 368 331 592
rect 453 368 483 592
rect 543 368 573 592
rect 639 368 669 592
rect 729 368 759 592
rect 819 368 849 592
<< ndiff >>
rect 65 210 118 222
rect 65 176 73 210
rect 107 176 118 210
rect 65 120 118 176
rect 65 86 73 120
rect 107 86 118 120
rect 65 74 118 86
rect 148 184 204 222
rect 148 150 159 184
rect 193 150 204 184
rect 148 116 204 150
rect 148 82 159 116
rect 193 82 204 116
rect 148 74 204 82
rect 234 116 304 222
rect 234 82 245 116
rect 279 82 304 116
rect 234 74 304 82
rect 334 124 390 222
rect 334 90 345 124
rect 379 90 390 124
rect 334 74 390 90
rect 420 210 528 222
rect 420 176 452 210
rect 486 176 528 210
rect 420 120 528 176
rect 420 86 452 120
rect 486 86 528 120
rect 420 74 528 86
rect 558 184 636 222
rect 558 150 583 184
rect 617 150 636 184
rect 558 116 636 150
rect 558 82 583 116
rect 617 82 636 116
rect 558 74 636 82
rect 666 116 722 222
rect 666 82 677 116
rect 711 82 722 116
rect 666 74 722 82
rect 752 184 808 222
rect 752 150 763 184
rect 797 150 808 184
rect 752 116 808 150
rect 752 82 763 116
rect 797 82 808 116
rect 752 74 808 82
rect 838 210 891 222
rect 838 176 849 210
rect 883 176 891 210
rect 838 120 891 176
rect 838 86 849 120
rect 883 86 891 120
rect 838 74 891 86
<< pdiff >>
rect 66 580 121 592
rect 66 546 74 580
rect 108 546 121 580
rect 66 510 121 546
rect 66 476 74 510
rect 108 476 121 510
rect 66 440 121 476
rect 66 406 74 440
rect 108 406 121 440
rect 66 368 121 406
rect 151 578 211 592
rect 151 544 164 578
rect 198 544 211 578
rect 151 368 211 544
rect 241 580 301 592
rect 241 546 254 580
rect 288 546 301 580
rect 241 492 301 546
rect 241 458 254 492
rect 288 458 301 492
rect 241 368 301 458
rect 331 578 453 592
rect 331 544 375 578
rect 409 544 453 578
rect 331 368 453 544
rect 483 583 543 592
rect 483 549 496 583
rect 530 549 543 583
rect 483 515 543 549
rect 483 481 496 515
rect 530 481 543 515
rect 483 447 543 481
rect 483 413 496 447
rect 530 413 543 447
rect 483 368 543 413
rect 573 531 639 592
rect 573 497 589 531
rect 623 497 639 531
rect 573 414 639 497
rect 573 380 589 414
rect 623 380 639 414
rect 573 368 639 380
rect 669 580 729 592
rect 669 546 682 580
rect 716 546 729 580
rect 669 494 729 546
rect 669 460 682 494
rect 716 460 729 494
rect 669 368 729 460
rect 759 531 819 592
rect 759 497 772 531
rect 806 497 819 531
rect 759 424 819 497
rect 759 390 772 424
rect 806 390 819 424
rect 759 368 819 390
rect 849 580 904 592
rect 849 546 862 580
rect 896 546 904 580
rect 849 494 904 546
rect 849 460 862 494
rect 896 460 904 494
rect 849 368 904 460
<< ndiffc >>
rect 73 176 107 210
rect 73 86 107 120
rect 159 150 193 184
rect 159 82 193 116
rect 245 82 279 116
rect 345 90 379 124
rect 452 176 486 210
rect 452 86 486 120
rect 583 150 617 184
rect 583 82 617 116
rect 677 82 711 116
rect 763 150 797 184
rect 763 82 797 116
rect 849 176 883 210
rect 849 86 883 120
<< pdiffc >>
rect 74 546 108 580
rect 74 476 108 510
rect 74 406 108 440
rect 164 544 198 578
rect 254 546 288 580
rect 254 458 288 492
rect 375 544 409 578
rect 496 549 530 583
rect 496 481 530 515
rect 496 413 530 447
rect 589 497 623 531
rect 589 380 623 414
rect 682 546 716 580
rect 682 460 716 494
rect 772 497 806 531
rect 772 390 806 424
rect 862 546 896 580
rect 862 460 896 494
<< poly >>
rect 121 592 151 618
rect 211 592 241 618
rect 301 592 331 618
rect 453 592 483 618
rect 543 592 573 618
rect 639 592 669 618
rect 729 592 759 618
rect 819 592 849 618
rect 121 353 151 368
rect 211 353 241 368
rect 301 353 331 368
rect 453 353 483 368
rect 543 353 573 368
rect 639 353 669 368
rect 729 353 759 368
rect 819 353 849 368
rect 118 336 154 353
rect 208 336 244 353
rect 298 336 334 353
rect 450 336 486 353
rect 88 320 154 336
rect 88 286 104 320
rect 138 286 154 320
rect 88 270 154 286
rect 204 320 334 336
rect 204 286 226 320
rect 260 286 334 320
rect 204 270 334 286
rect 376 320 486 336
rect 376 286 392 320
rect 426 286 486 320
rect 540 310 576 353
rect 636 336 672 353
rect 726 336 762 353
rect 636 320 762 336
rect 816 326 852 353
rect 376 270 486 286
rect 528 294 594 310
rect 118 222 148 270
rect 204 222 234 270
rect 304 222 334 270
rect 390 222 420 270
rect 528 260 544 294
rect 578 260 594 294
rect 528 244 594 260
rect 636 286 697 320
rect 731 286 762 320
rect 636 270 762 286
rect 808 310 874 326
rect 808 276 824 310
rect 858 276 874 310
rect 528 222 558 244
rect 636 222 666 270
rect 722 222 752 270
rect 808 260 874 276
rect 808 222 838 260
rect 118 48 148 74
rect 204 48 234 74
rect 304 48 334 74
rect 390 48 420 74
rect 528 48 558 74
rect 636 48 666 74
rect 722 48 752 74
rect 808 48 838 74
<< polycont >>
rect 104 286 138 320
rect 226 286 260 320
rect 392 286 426 320
rect 544 260 578 294
rect 697 286 731 320
rect 824 276 858 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 58 580 108 596
rect 58 546 74 580
rect 58 510 108 546
rect 148 578 198 649
rect 148 544 164 578
rect 148 526 198 544
rect 238 580 304 596
rect 238 546 254 580
rect 288 546 304 580
rect 58 476 74 510
rect 238 492 304 546
rect 338 578 446 649
rect 338 544 375 578
rect 409 544 446 578
rect 338 526 446 544
rect 480 583 912 615
rect 480 549 496 583
rect 530 581 912 583
rect 530 549 546 581
rect 480 515 546 549
rect 666 580 732 581
rect 480 492 496 515
rect 108 476 254 492
rect 58 458 254 476
rect 288 481 496 492
rect 530 481 546 515
rect 288 458 546 481
rect 58 440 108 458
rect 58 406 74 440
rect 480 447 546 458
rect 58 390 108 406
rect 142 390 442 424
rect 480 413 496 447
rect 530 413 546 447
rect 480 412 546 413
rect 586 531 626 547
rect 586 497 589 531
rect 623 497 626 531
rect 586 424 626 497
rect 666 546 682 580
rect 716 546 732 580
rect 846 580 912 581
rect 666 494 732 546
rect 666 460 682 494
rect 716 460 732 494
rect 666 458 732 460
rect 772 531 806 547
rect 772 424 806 497
rect 846 546 862 580
rect 896 546 912 580
rect 846 494 912 546
rect 846 460 862 494
rect 896 460 912 494
rect 846 458 912 460
rect 586 414 772 424
rect 142 356 176 390
rect 25 320 176 356
rect 25 286 104 320
rect 138 286 176 320
rect 210 320 284 356
rect 210 286 226 320
rect 260 286 284 320
rect 376 320 442 390
rect 586 380 589 414
rect 623 390 772 414
rect 806 390 942 424
rect 623 380 626 390
rect 586 378 626 380
rect 376 286 392 320
rect 426 286 442 320
rect 476 344 626 378
rect 476 252 510 344
rect 681 320 747 356
rect 57 218 510 252
rect 544 294 647 310
rect 578 260 647 294
rect 681 286 697 320
rect 731 286 747 320
rect 781 310 874 326
rect 544 252 647 260
rect 781 276 824 310
rect 858 276 874 310
rect 781 260 874 276
rect 781 252 815 260
rect 544 218 815 252
rect 908 226 942 390
rect 57 210 107 218
rect 57 176 73 210
rect 408 210 510 218
rect 57 120 107 176
rect 57 86 73 120
rect 57 70 107 86
rect 143 150 159 184
rect 193 150 363 184
rect 408 176 452 210
rect 486 176 510 210
rect 849 210 942 226
rect 408 162 510 176
rect 143 116 193 150
rect 329 128 363 150
rect 329 124 395 128
rect 143 82 159 116
rect 143 66 193 82
rect 229 82 245 116
rect 279 82 295 116
rect 229 17 295 82
rect 329 90 345 124
rect 379 90 395 124
rect 329 70 395 90
rect 429 120 510 162
rect 429 86 452 120
rect 486 86 510 120
rect 429 70 510 86
rect 567 150 583 184
rect 617 150 763 184
rect 797 150 813 184
rect 567 116 627 150
rect 763 116 813 150
rect 567 82 583 116
rect 617 82 627 116
rect 567 66 627 82
rect 661 82 677 116
rect 711 82 727 116
rect 661 17 727 82
rect 797 82 813 116
rect 763 66 813 82
rect 883 176 942 210
rect 849 120 942 176
rect 883 86 942 120
rect 849 70 942 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a22oi_2
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 415 168 449 202 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 607 242 641 276 0 FreeSans 340 0 0 0 B1
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 960 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3523080
string GDS_START 3514838
<< end >>
