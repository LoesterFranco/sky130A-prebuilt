magic
tech sky130A
magscale 1 2
timestamp 1599588218
<< nwell >>
rect -38 332 710 704
<< pwell >>
rect 0 0 672 49
<< scpmos >>
rect 99 392 135 592
rect 189 392 225 592
rect 285 392 321 592
rect 393 392 429 592
rect 539 368 575 592
<< nmoslvt >>
rect 105 123 135 251
rect 200 79 230 207
rect 272 79 302 207
rect 358 79 388 207
rect 560 74 590 222
<< ndiff >>
rect 52 228 105 251
rect 52 194 60 228
rect 94 194 105 228
rect 52 123 105 194
rect 135 207 185 251
rect 135 172 200 207
rect 135 138 150 172
rect 184 138 200 172
rect 135 123 200 138
rect 150 79 200 123
rect 230 79 272 207
rect 302 194 358 207
rect 302 160 313 194
rect 347 160 358 194
rect 302 79 358 160
rect 388 125 445 207
rect 388 91 399 125
rect 433 91 445 125
rect 388 79 445 91
rect 507 152 560 222
rect 507 118 515 152
rect 549 118 560 152
rect 507 74 560 118
rect 590 210 643 222
rect 590 176 601 210
rect 635 176 643 210
rect 590 120 643 176
rect 590 86 601 120
rect 635 86 643 120
rect 590 74 643 86
<< pdiff >>
rect 47 580 99 592
rect 47 546 55 580
rect 89 546 99 580
rect 47 512 99 546
rect 47 478 55 512
rect 89 478 99 512
rect 47 444 99 478
rect 47 410 55 444
rect 89 410 99 444
rect 47 392 99 410
rect 135 580 189 592
rect 135 546 145 580
rect 179 546 189 580
rect 135 512 189 546
rect 135 478 145 512
rect 179 478 189 512
rect 135 444 189 478
rect 135 410 145 444
rect 179 410 189 444
rect 135 392 189 410
rect 225 531 285 592
rect 225 497 235 531
rect 269 497 285 531
rect 225 444 285 497
rect 225 410 235 444
rect 269 410 285 444
rect 225 392 285 410
rect 321 580 393 592
rect 321 546 342 580
rect 376 546 393 580
rect 321 512 393 546
rect 321 478 342 512
rect 376 478 393 512
rect 321 392 393 478
rect 429 568 539 592
rect 429 534 440 568
rect 474 534 539 568
rect 429 503 539 534
rect 429 469 495 503
rect 529 469 539 503
rect 429 392 539 469
rect 487 368 539 392
rect 575 580 627 592
rect 575 546 585 580
rect 619 546 627 580
rect 575 497 627 546
rect 575 463 585 497
rect 619 463 627 497
rect 575 414 627 463
rect 575 380 585 414
rect 619 380 627 414
rect 575 368 627 380
<< ndiffc >>
rect 60 194 94 228
rect 150 138 184 172
rect 313 160 347 194
rect 399 91 433 125
rect 515 118 549 152
rect 601 176 635 210
rect 601 86 635 120
<< pdiffc >>
rect 55 546 89 580
rect 55 478 89 512
rect 55 410 89 444
rect 145 546 179 580
rect 145 478 179 512
rect 145 410 179 444
rect 235 497 269 531
rect 235 410 269 444
rect 342 546 376 580
rect 342 478 376 512
rect 440 534 474 568
rect 495 469 529 503
rect 585 546 619 580
rect 585 463 619 497
rect 585 380 619 414
<< poly >>
rect 99 592 135 618
rect 189 592 225 618
rect 285 592 321 618
rect 393 592 429 618
rect 539 592 575 618
rect 99 266 135 392
rect 189 360 225 392
rect 285 360 321 392
rect 177 344 243 360
rect 177 310 193 344
rect 227 310 243 344
rect 177 294 243 310
rect 285 344 351 360
rect 285 310 301 344
rect 335 310 351 344
rect 285 294 351 310
rect 393 336 429 392
rect 393 320 459 336
rect 539 326 575 368
rect 105 251 135 266
rect 200 207 230 294
rect 285 252 315 294
rect 393 286 409 320
rect 443 286 459 320
rect 393 270 459 286
rect 501 310 575 326
rect 501 276 517 310
rect 551 290 575 310
rect 551 276 590 290
rect 393 252 423 270
rect 501 260 590 276
rect 272 222 315 252
rect 358 222 423 252
rect 560 222 590 260
rect 272 207 302 222
rect 358 207 388 222
rect 105 101 135 123
rect 46 85 135 101
rect 46 51 62 85
rect 96 51 135 85
rect 200 53 230 79
rect 272 53 302 79
rect 358 53 388 79
rect 46 35 135 51
rect 560 48 590 74
<< polycont >>
rect 193 310 227 344
rect 301 310 335 344
rect 409 286 443 320
rect 517 276 551 310
rect 62 51 96 85
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 39 580 89 649
rect 39 546 55 580
rect 39 512 89 546
rect 39 478 55 512
rect 39 444 89 478
rect 39 410 55 444
rect 39 394 89 410
rect 129 581 399 615
rect 129 580 179 581
rect 129 546 145 580
rect 319 580 399 581
rect 129 512 179 546
rect 129 478 145 512
rect 129 444 179 478
rect 129 410 145 444
rect 129 394 179 410
rect 219 531 285 547
rect 219 497 235 531
rect 269 497 285 531
rect 219 444 285 497
rect 319 546 342 580
rect 376 546 399 580
rect 319 512 399 546
rect 319 478 342 512
rect 376 478 399 512
rect 319 462 399 478
rect 433 568 545 649
rect 433 534 440 568
rect 474 534 545 568
rect 433 503 545 534
rect 433 469 495 503
rect 529 469 545 503
rect 433 462 545 469
rect 585 580 651 596
rect 619 546 651 580
rect 585 497 651 546
rect 619 463 651 497
rect 219 410 235 444
rect 269 428 285 444
rect 269 410 551 428
rect 219 394 551 410
rect 25 344 243 360
rect 25 310 193 344
rect 227 310 243 344
rect 25 294 243 310
rect 285 344 359 360
rect 285 310 301 344
rect 335 310 359 344
rect 285 294 359 310
rect 393 320 459 356
rect 393 286 409 320
rect 443 286 459 320
rect 393 270 459 286
rect 501 310 551 394
rect 501 276 517 310
rect 44 228 257 260
rect 501 236 551 276
rect 44 194 60 228
rect 94 226 257 228
rect 94 194 110 226
rect 44 168 110 194
rect 146 172 189 192
rect 146 138 150 172
rect 184 138 189 172
rect 25 101 71 134
rect 25 85 112 101
rect 25 51 62 85
rect 96 51 112 85
rect 146 17 189 138
rect 223 125 257 226
rect 297 202 551 236
rect 585 414 651 463
rect 619 380 651 414
rect 585 210 651 380
rect 297 194 363 202
rect 297 160 313 194
rect 347 160 363 194
rect 585 176 601 210
rect 635 176 651 210
rect 297 159 363 160
rect 499 152 549 168
rect 223 91 399 125
rect 433 91 449 125
rect 223 75 449 91
rect 499 118 515 152
rect 499 17 549 118
rect 585 120 651 176
rect 585 86 601 120
rect 635 86 651 120
rect 585 70 651 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
rlabel comment s 0 0 0 0 4 a22o_1
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 607 94 641 128 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 607 168 641 202 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 607 242 641 276 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 607 390 641 424 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 607 464 641 498 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 607 538 641 572 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 31 94 65 128 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 672 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3547918
string GDS_START 3540618
<< end >>
