magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 118 424 184 596
rect 308 424 374 596
rect 498 424 564 596
rect 688 424 754 596
rect 878 424 944 596
rect 1068 424 1134 596
rect 57 390 1223 424
rect 57 236 91 390
rect 125 270 1143 356
rect 1177 236 1223 390
rect 57 202 1223 236
rect 123 92 525 202
rect 659 89 725 202
rect 859 89 925 202
rect 1059 89 1125 202
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 23 458 78 649
rect 224 458 274 649
rect 414 458 464 649
rect 604 458 654 649
rect 794 458 844 649
rect 984 458 1034 649
rect 1174 458 1224 649
rect 23 17 89 155
rect 559 17 625 155
rect 759 17 825 155
rect 959 17 1025 155
rect 1159 17 1225 155
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
<< metal1 >>
rect 0 683 1248 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 0 617 1248 649
rect 0 17 1248 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
rect 0 -49 1248 -17
<< labels >>
rlabel locali s 125 270 1143 356 6 A
port 1 nsew signal input
rlabel locali s 1177 236 1223 390 6 Y
port 2 nsew signal output
rlabel locali s 1068 424 1134 596 6 Y
port 2 nsew signal output
rlabel locali s 1059 89 1125 202 6 Y
port 2 nsew signal output
rlabel locali s 878 424 944 596 6 Y
port 2 nsew signal output
rlabel locali s 859 89 925 202 6 Y
port 2 nsew signal output
rlabel locali s 688 424 754 596 6 Y
port 2 nsew signal output
rlabel locali s 659 89 725 202 6 Y
port 2 nsew signal output
rlabel locali s 498 424 564 596 6 Y
port 2 nsew signal output
rlabel locali s 308 424 374 596 6 Y
port 2 nsew signal output
rlabel locali s 123 92 525 202 6 Y
port 2 nsew signal output
rlabel locali s 118 424 184 596 6 Y
port 2 nsew signal output
rlabel locali s 57 390 1223 424 6 Y
port 2 nsew signal output
rlabel locali s 57 236 91 390 6 Y
port 2 nsew signal output
rlabel locali s 57 202 1223 236 6 Y
port 2 nsew signal output
rlabel metal1 s 0 -49 1248 49 8 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 617 1248 715 6 VPWR
port 4 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1248 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 2795386
string GDS_START 2785516
<< end >>
