magic
tech sky130A
magscale 1 2
timestamp 1604502741
<< locali >>
rect 23 424 89 596
rect 23 390 167 424
rect 21 260 87 356
rect 121 226 167 390
rect 201 270 267 356
rect 313 270 391 356
rect 439 270 551 356
rect 585 260 651 356
rect 23 192 644 226
rect 23 70 89 192
rect 578 70 644 192
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 123 492 189 596
rect 223 526 357 649
rect 289 492 357 526
rect 481 492 549 649
rect 123 458 255 492
rect 583 458 649 596
rect 221 390 649 458
rect 123 17 252 136
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel locali s 585 260 651 356 6 A1
port 1 nsew signal input
rlabel locali s 439 270 551 356 6 A2
port 2 nsew signal input
rlabel locali s 313 270 391 356 6 A3
port 3 nsew signal input
rlabel locali s 201 270 267 356 6 A4
port 4 nsew signal input
rlabel locali s 21 260 87 356 6 B1
port 5 nsew signal input
rlabel locali s 578 70 644 192 6 Y
port 6 nsew signal output
rlabel locali s 121 226 167 390 6 Y
port 6 nsew signal output
rlabel locali s 23 424 89 596 6 Y
port 6 nsew signal output
rlabel locali s 23 390 167 424 6 Y
port 6 nsew signal output
rlabel locali s 23 192 644 226 6 Y
port 6 nsew signal output
rlabel locali s 23 70 89 192 6 Y
port 6 nsew signal output
rlabel metal1 s 0 -49 672 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 617 672 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3078518
string GDS_START 3072692
<< end >>
