magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 736 561
rect 103 467 169 527
rect 296 467 363 527
rect 397 425 534 483
rect 17 215 85 287
rect 187 299 250 365
rect 187 158 221 299
rect 351 215 464 255
rect 510 215 710 255
rect 187 136 249 158
rect 187 135 250 136
rect 126 17 160 113
rect 194 52 250 135
rect 287 17 363 97
rect 477 17 543 97
rect 645 17 711 117
rect 0 -17 736 17
<< obsli1 >>
rect 102 399 343 433
rect 572 443 669 477
rect 102 378 153 399
rect 17 321 153 378
rect 288 391 343 399
rect 572 391 606 443
rect 119 181 153 321
rect 17 147 153 181
rect 288 357 606 391
rect 645 323 712 363
rect 284 290 712 323
rect 283 289 712 290
rect 283 285 333 289
rect 283 284 331 285
rect 283 282 329 284
rect 283 280 326 282
rect 283 278 325 280
rect 283 276 324 278
rect 283 274 322 276
rect 283 271 320 274
rect 283 265 317 271
rect 258 199 317 265
rect 283 181 317 199
rect 17 65 70 147
rect 283 147 611 181
rect 397 61 431 147
rect 577 61 611 147
<< metal1 >>
rect 0 496 736 592
rect 0 -48 736 48
<< labels >>
rlabel locali s 351 215 464 255 6 A
port 1 nsew signal input
rlabel locali s 397 425 534 483 6 B
port 2 nsew signal input
rlabel locali s 510 215 710 255 6 C
port 3 nsew signal input
rlabel locali s 17 215 85 287 6 D_N
port 4 nsew signal input
rlabel locali s 194 52 250 135 6 X
port 5 nsew signal output
rlabel locali s 187 299 250 365 6 X
port 5 nsew signal output
rlabel locali s 187 158 221 299 6 X
port 5 nsew signal output
rlabel locali s 187 136 249 158 6 X
port 5 nsew signal output
rlabel locali s 187 135 250 136 6 X
port 5 nsew signal output
rlabel locali s 645 17 711 117 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 477 17 543 97 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 287 17 363 97 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 126 17 160 113 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 736 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 736 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 296 467 363 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 103 467 169 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 736 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 736 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1096794
string GDS_START 1090300
<< end >>
