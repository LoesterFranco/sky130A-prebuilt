magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1104 561
rect 119 359 161 527
rect 726 325 776 425
rect 998 427 1048 527
rect 726 291 807 325
rect 20 215 248 257
rect 284 215 527 257
rect 563 215 707 257
rect 743 215 807 291
rect 1037 257 1087 391
rect 961 215 1087 257
rect 743 181 784 215
rect 17 17 69 181
rect 103 145 784 181
rect 103 51 169 145
rect 203 17 237 111
rect 271 51 337 145
rect 371 17 516 111
rect 550 51 616 145
rect 650 17 684 111
rect 718 51 784 145
rect 818 17 859 179
rect 998 17 1048 165
rect 0 -17 1104 17
<< obsli1 >>
rect 17 325 85 493
rect 195 325 245 493
rect 279 459 608 493
rect 279 359 321 459
rect 355 325 421 425
rect 17 291 421 325
rect 455 325 532 425
rect 566 359 608 459
rect 642 459 859 493
rect 642 325 692 459
rect 455 291 692 325
rect 810 359 859 459
rect 893 407 964 490
rect 893 249 927 407
rect 864 215 927 249
rect 893 181 927 215
rect 893 76 964 181
<< metal1 >>
rect 0 496 1104 592
rect 0 -48 1104 48
<< labels >>
rlabel locali s 20 215 248 257 6 A
port 1 nsew signal input
rlabel locali s 284 215 527 257 6 B
port 2 nsew signal input
rlabel locali s 563 215 707 257 6 C
port 3 nsew signal input
rlabel locali s 1037 257 1087 391 6 D_N
port 4 nsew signal input
rlabel locali s 961 215 1087 257 6 D_N
port 4 nsew signal input
rlabel locali s 743 215 807 291 6 Y
port 5 nsew signal output
rlabel locali s 743 181 784 215 6 Y
port 5 nsew signal output
rlabel locali s 726 325 776 425 6 Y
port 5 nsew signal output
rlabel locali s 726 291 807 325 6 Y
port 5 nsew signal output
rlabel locali s 718 51 784 145 6 Y
port 5 nsew signal output
rlabel locali s 550 51 616 145 6 Y
port 5 nsew signal output
rlabel locali s 271 51 337 145 6 Y
port 5 nsew signal output
rlabel locali s 103 145 784 181 6 Y
port 5 nsew signal output
rlabel locali s 103 51 169 145 6 Y
port 5 nsew signal output
rlabel locali s 998 17 1048 165 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 818 17 859 179 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 650 17 684 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 371 17 516 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 203 17 237 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 17 17 69 181 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 1104 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1104 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 998 427 1048 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 119 359 161 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 1104 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 1104 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1104 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1177522
string GDS_START 1168252
<< end >>
