magic
tech sky130A
magscale 1 2
timestamp 1604502701
<< nwell >>
rect -38 332 1670 704
<< pwell >>
rect 0 0 1632 49
<< scpmos >>
rect 401 368 431 592
rect 501 368 531 592
rect 849 368 879 592
rect 939 368 969 592
rect 1161 368 1191 592
rect 1261 368 1291 592
rect 1427 368 1457 592
rect 1517 368 1547 592
<< nmoslvt >>
rect 82 74 112 222
rect 168 74 198 222
rect 254 74 284 222
rect 340 74 370 222
rect 426 74 456 222
rect 576 74 606 222
rect 670 74 700 222
rect 756 74 786 222
rect 842 74 872 222
rect 928 74 958 222
rect 1014 74 1044 222
rect 1100 74 1130 222
rect 1186 74 1216 222
rect 1272 74 1302 222
rect 1430 74 1460 222
rect 1516 74 1546 222
<< ndiff >>
rect 27 210 82 222
rect 27 176 37 210
rect 71 176 82 210
rect 27 120 82 176
rect 27 86 37 120
rect 71 86 82 120
rect 27 74 82 86
rect 112 199 168 222
rect 112 165 123 199
rect 157 165 168 199
rect 112 120 168 165
rect 112 86 123 120
rect 157 86 168 120
rect 112 74 168 86
rect 198 210 254 222
rect 198 176 209 210
rect 243 176 254 210
rect 198 120 254 176
rect 198 86 209 120
rect 243 86 254 120
rect 198 74 254 86
rect 284 152 340 222
rect 284 118 295 152
rect 329 118 340 152
rect 284 74 340 118
rect 370 210 426 222
rect 370 176 381 210
rect 415 176 426 210
rect 370 120 426 176
rect 370 86 381 120
rect 415 86 426 120
rect 370 74 426 86
rect 456 168 576 222
rect 456 134 531 168
rect 565 134 576 168
rect 456 116 576 134
rect 456 82 467 116
rect 501 82 576 116
rect 456 74 576 82
rect 606 210 670 222
rect 606 176 621 210
rect 655 176 670 210
rect 606 120 670 176
rect 606 86 621 120
rect 655 86 670 120
rect 606 74 670 86
rect 700 144 756 222
rect 700 110 711 144
rect 745 110 756 144
rect 700 74 756 110
rect 786 210 842 222
rect 786 176 797 210
rect 831 176 842 210
rect 786 120 842 176
rect 786 86 797 120
rect 831 86 842 120
rect 786 74 842 86
rect 872 207 928 222
rect 872 173 883 207
rect 917 173 928 207
rect 872 74 928 173
rect 958 120 1014 222
rect 958 86 969 120
rect 1003 86 1014 120
rect 958 74 1014 86
rect 1044 199 1100 222
rect 1044 165 1055 199
rect 1089 165 1100 199
rect 1044 74 1100 165
rect 1130 120 1186 222
rect 1130 86 1141 120
rect 1175 86 1186 120
rect 1130 74 1186 86
rect 1216 199 1272 222
rect 1216 165 1227 199
rect 1261 165 1272 199
rect 1216 74 1272 165
rect 1302 120 1430 222
rect 1302 86 1313 120
rect 1347 86 1385 120
rect 1419 86 1430 120
rect 1302 74 1430 86
rect 1460 199 1516 222
rect 1460 165 1471 199
rect 1505 165 1516 199
rect 1460 74 1516 165
rect 1546 132 1596 222
rect 1546 120 1605 132
rect 1546 86 1558 120
rect 1592 86 1605 120
rect 1546 74 1605 86
<< pdiff >>
rect 134 580 401 592
rect 134 546 148 580
rect 182 546 216 580
rect 250 546 285 580
rect 319 546 353 580
rect 387 546 401 580
rect 134 510 401 546
rect 134 476 148 510
rect 182 476 216 510
rect 250 476 285 510
rect 319 476 353 510
rect 387 476 401 510
rect 134 440 401 476
rect 134 406 148 440
rect 182 406 216 440
rect 250 406 285 440
rect 319 406 353 440
rect 387 406 401 440
rect 134 368 401 406
rect 431 580 501 592
rect 431 546 444 580
rect 478 546 501 580
rect 431 510 501 546
rect 431 476 444 510
rect 478 476 501 510
rect 431 440 501 476
rect 431 406 444 440
rect 478 406 501 440
rect 431 368 501 406
rect 531 580 849 592
rect 531 546 544 580
rect 578 546 629 580
rect 663 546 720 580
rect 754 546 801 580
rect 835 546 849 580
rect 531 508 849 546
rect 531 474 544 508
rect 578 474 629 508
rect 663 474 720 508
rect 754 474 801 508
rect 835 474 849 508
rect 531 368 849 474
rect 879 580 939 592
rect 879 546 892 580
rect 926 546 939 580
rect 879 497 939 546
rect 879 463 892 497
rect 926 463 939 497
rect 879 414 939 463
rect 879 380 892 414
rect 926 380 939 414
rect 879 368 939 380
rect 969 580 1038 592
rect 969 546 992 580
rect 1026 546 1038 580
rect 969 497 1038 546
rect 969 463 992 497
rect 1026 463 1038 497
rect 969 414 1038 463
rect 969 380 992 414
rect 1026 380 1038 414
rect 969 368 1038 380
rect 1092 580 1161 592
rect 1092 546 1104 580
rect 1138 546 1161 580
rect 1092 497 1161 546
rect 1092 463 1104 497
rect 1138 463 1161 497
rect 1092 414 1161 463
rect 1092 380 1104 414
rect 1138 380 1161 414
rect 1092 368 1161 380
rect 1191 580 1261 592
rect 1191 546 1204 580
rect 1238 546 1261 580
rect 1191 502 1261 546
rect 1191 468 1204 502
rect 1238 468 1261 502
rect 1191 424 1261 468
rect 1191 390 1204 424
rect 1238 390 1261 424
rect 1191 368 1261 390
rect 1291 580 1427 592
rect 1291 546 1304 580
rect 1338 546 1380 580
rect 1414 546 1427 580
rect 1291 492 1427 546
rect 1291 458 1304 492
rect 1338 458 1380 492
rect 1414 458 1427 492
rect 1291 368 1427 458
rect 1457 580 1517 592
rect 1457 546 1470 580
rect 1504 546 1517 580
rect 1457 502 1517 546
rect 1457 468 1470 502
rect 1504 468 1517 502
rect 1457 424 1517 468
rect 1457 390 1470 424
rect 1504 390 1517 424
rect 1457 368 1517 390
rect 1547 580 1605 592
rect 1547 546 1560 580
rect 1594 546 1605 580
rect 1547 492 1605 546
rect 1547 458 1560 492
rect 1594 458 1605 492
rect 1547 368 1605 458
<< ndiffc >>
rect 37 176 71 210
rect 37 86 71 120
rect 123 165 157 199
rect 123 86 157 120
rect 209 176 243 210
rect 209 86 243 120
rect 295 118 329 152
rect 381 176 415 210
rect 381 86 415 120
rect 531 134 565 168
rect 467 82 501 116
rect 621 176 655 210
rect 621 86 655 120
rect 711 110 745 144
rect 797 176 831 210
rect 797 86 831 120
rect 883 173 917 207
rect 969 86 1003 120
rect 1055 165 1089 199
rect 1141 86 1175 120
rect 1227 165 1261 199
rect 1313 86 1347 120
rect 1385 86 1419 120
rect 1471 165 1505 199
rect 1558 86 1592 120
<< pdiffc >>
rect 148 546 182 580
rect 216 546 250 580
rect 285 546 319 580
rect 353 546 387 580
rect 148 476 182 510
rect 216 476 250 510
rect 285 476 319 510
rect 353 476 387 510
rect 148 406 182 440
rect 216 406 250 440
rect 285 406 319 440
rect 353 406 387 440
rect 444 546 478 580
rect 444 476 478 510
rect 444 406 478 440
rect 544 546 578 580
rect 629 546 663 580
rect 720 546 754 580
rect 801 546 835 580
rect 544 474 578 508
rect 629 474 663 508
rect 720 474 754 508
rect 801 474 835 508
rect 892 546 926 580
rect 892 463 926 497
rect 892 380 926 414
rect 992 546 1026 580
rect 992 463 1026 497
rect 992 380 1026 414
rect 1104 546 1138 580
rect 1104 463 1138 497
rect 1104 380 1138 414
rect 1204 546 1238 580
rect 1204 468 1238 502
rect 1204 390 1238 424
rect 1304 546 1338 580
rect 1380 546 1414 580
rect 1304 458 1338 492
rect 1380 458 1414 492
rect 1470 546 1504 580
rect 1470 468 1504 502
rect 1470 390 1504 424
rect 1560 546 1594 580
rect 1560 458 1594 492
<< poly >>
rect 401 592 431 618
rect 501 592 531 618
rect 849 592 879 618
rect 939 592 969 618
rect 1161 592 1191 618
rect 1261 592 1291 618
rect 1427 592 1457 618
rect 1517 592 1547 618
rect 401 353 431 368
rect 501 353 531 368
rect 849 353 879 368
rect 939 353 969 368
rect 1161 353 1191 368
rect 1261 353 1291 368
rect 1427 353 1457 368
rect 1517 353 1547 368
rect 398 345 434 353
rect 498 345 534 353
rect 846 345 882 353
rect 936 345 972 353
rect 398 320 972 345
rect 398 286 425 320
rect 459 286 502 320
rect 536 286 580 320
rect 614 286 658 320
rect 692 286 736 320
rect 770 315 972 320
rect 770 286 786 315
rect 1158 310 1194 353
rect 1258 310 1294 353
rect 1424 310 1460 353
rect 1514 310 1550 353
rect 398 270 786 286
rect 398 267 456 270
rect 82 237 456 267
rect 82 222 112 237
rect 168 222 198 237
rect 254 222 284 237
rect 340 222 370 237
rect 426 222 456 237
rect 576 222 606 270
rect 670 222 700 270
rect 756 222 786 270
rect 1037 294 1550 310
rect 1037 267 1053 294
rect 842 260 1053 267
rect 1087 260 1121 294
rect 1155 260 1189 294
rect 1223 260 1257 294
rect 1291 260 1325 294
rect 1359 260 1393 294
rect 1427 260 1461 294
rect 1495 260 1550 294
rect 842 244 1550 260
rect 842 237 1216 244
rect 842 222 872 237
rect 928 222 958 237
rect 1014 222 1044 237
rect 1100 222 1130 237
rect 1186 222 1216 237
rect 1272 222 1302 244
rect 1430 222 1460 244
rect 1516 222 1546 244
rect 82 48 112 74
rect 168 48 198 74
rect 254 48 284 74
rect 340 48 370 74
rect 426 48 456 74
rect 576 48 606 74
rect 670 48 700 74
rect 756 48 786 74
rect 842 48 872 74
rect 928 48 958 74
rect 1014 48 1044 74
rect 1100 48 1130 74
rect 1186 48 1216 74
rect 1272 48 1302 74
rect 1430 48 1460 74
rect 1516 48 1546 74
<< polycont >>
rect 425 286 459 320
rect 502 286 536 320
rect 580 286 614 320
rect 658 286 692 320
rect 736 286 770 320
rect 1053 260 1087 294
rect 1121 260 1155 294
rect 1189 260 1223 294
rect 1257 260 1291 294
rect 1325 260 1359 294
rect 1393 260 1427 294
rect 1461 260 1495 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 132 580 394 649
rect 132 546 148 580
rect 182 546 216 580
rect 250 546 285 580
rect 319 546 353 580
rect 387 546 394 580
rect 132 510 394 546
rect 132 476 148 510
rect 182 476 216 510
rect 250 476 285 510
rect 319 476 353 510
rect 387 476 394 510
rect 132 440 394 476
rect 132 406 148 440
rect 182 406 216 440
rect 250 406 285 440
rect 319 406 353 440
rect 387 406 394 440
rect 132 390 394 406
rect 428 580 494 596
rect 428 546 444 580
rect 478 546 494 580
rect 428 510 494 546
rect 428 476 444 510
rect 478 476 494 510
rect 428 440 494 476
rect 528 580 842 649
rect 528 546 544 580
rect 578 546 629 580
rect 663 546 720 580
rect 754 546 801 580
rect 835 546 842 580
rect 528 508 842 546
rect 528 474 544 508
rect 578 474 629 508
rect 663 474 720 508
rect 754 474 801 508
rect 835 474 842 508
rect 528 458 842 474
rect 876 580 942 596
rect 876 546 892 580
rect 926 546 942 580
rect 876 497 942 546
rect 876 463 892 497
rect 926 463 942 497
rect 428 406 444 440
rect 478 424 494 440
rect 876 424 942 463
rect 478 414 942 424
rect 478 406 892 414
rect 428 390 892 406
rect 876 380 892 390
rect 926 380 942 414
rect 409 320 839 356
rect 409 286 425 320
rect 459 286 502 320
rect 536 286 580 320
rect 614 286 658 320
rect 692 286 736 320
rect 770 286 839 320
rect 21 236 372 271
rect 409 270 839 286
rect 21 233 831 236
rect 21 210 71 233
rect 21 176 37 210
rect 207 210 831 233
rect 876 226 942 380
rect 976 580 1042 649
rect 976 546 992 580
rect 1026 546 1042 580
rect 976 497 1042 546
rect 976 463 992 497
rect 1026 463 1042 497
rect 976 414 1042 463
rect 976 380 992 414
rect 1026 380 1042 414
rect 976 364 1042 380
rect 1088 580 1154 649
rect 1088 546 1104 580
rect 1138 546 1154 580
rect 1088 497 1154 546
rect 1088 463 1104 497
rect 1138 463 1154 497
rect 1088 414 1154 463
rect 1088 380 1104 414
rect 1138 380 1154 414
rect 1188 580 1254 596
rect 1188 546 1204 580
rect 1238 546 1254 580
rect 1188 502 1254 546
rect 1188 468 1204 502
rect 1238 468 1254 502
rect 1188 424 1254 468
rect 1288 580 1430 649
rect 1288 546 1304 580
rect 1338 546 1380 580
rect 1414 546 1430 580
rect 1288 492 1430 546
rect 1288 458 1304 492
rect 1338 458 1380 492
rect 1414 458 1430 492
rect 1464 580 1510 596
rect 1464 546 1470 580
rect 1504 546 1510 580
rect 1464 502 1510 546
rect 1464 468 1470 502
rect 1504 468 1510 502
rect 1464 424 1510 468
rect 1544 580 1610 649
rect 1544 546 1560 580
rect 1594 546 1610 580
rect 1544 492 1610 546
rect 1544 458 1560 492
rect 1594 458 1610 492
rect 1188 390 1204 424
rect 1238 390 1470 424
rect 1504 390 1579 424
rect 1088 364 1154 380
rect 1193 310 1511 356
rect 1037 294 1511 310
rect 1037 260 1053 294
rect 1087 260 1121 294
rect 1155 260 1189 294
rect 1223 260 1257 294
rect 1291 260 1325 294
rect 1359 260 1393 294
rect 1427 260 1461 294
rect 1495 260 1511 294
rect 1037 244 1511 260
rect 21 120 71 176
rect 21 86 37 120
rect 21 70 71 86
rect 107 165 123 199
rect 157 165 173 199
rect 107 120 173 165
rect 107 86 123 120
rect 157 86 173 120
rect 107 17 173 86
rect 207 176 209 210
rect 243 202 381 210
rect 243 176 245 202
rect 207 120 245 176
rect 379 176 381 202
rect 415 202 621 210
rect 415 176 431 202
rect 207 86 209 120
rect 243 86 245 120
rect 207 70 245 86
rect 279 152 345 168
rect 279 118 295 152
rect 329 118 345 152
rect 279 17 345 118
rect 379 120 431 176
rect 615 176 621 202
rect 655 202 797 210
rect 655 176 661 202
rect 379 86 381 120
rect 415 86 431 120
rect 379 70 431 86
rect 465 134 531 168
rect 565 134 581 168
rect 465 116 581 134
rect 465 82 467 116
rect 501 82 581 116
rect 465 17 581 82
rect 615 120 661 176
rect 615 86 621 120
rect 655 86 661 120
rect 615 70 661 86
rect 695 144 761 168
rect 695 110 711 144
rect 745 110 761 144
rect 695 17 761 110
rect 797 120 831 176
rect 867 210 942 226
rect 1545 210 1579 390
rect 867 207 1579 210
rect 867 173 883 207
rect 917 199 1579 207
rect 917 173 1055 199
rect 867 165 1055 173
rect 1089 165 1227 199
rect 1261 165 1471 199
rect 1505 165 1579 199
rect 867 154 1579 165
rect 831 86 969 120
rect 1003 86 1141 120
rect 1175 86 1313 120
rect 1347 86 1385 120
rect 1419 86 1558 120
rect 1592 86 1609 120
rect 797 70 1609 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
rlabel comment s 0 0 0 0 4 nand2_8
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 1279 316 1313 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 1375 316 1409 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 1471 316 1505 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 895 242 929 276 0 FreeSans 340 0 0 0 Y
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 1632 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 2074908
string GDS_START 2062816
<< end >>
