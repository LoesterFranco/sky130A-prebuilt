magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 2726 704
<< pwell >>
rect 0 0 2688 49
<< scnmos >>
rect 84 74 114 222
rect 170 74 200 222
rect 368 119 398 203
rect 493 119 523 203
rect 565 119 595 203
rect 651 119 681 203
rect 924 119 954 229
rect 1024 119 1054 229
rect 1124 119 1154 229
rect 1224 119 1254 229
rect 1319 114 1349 224
rect 1581 140 1611 224
rect 1659 140 1689 224
rect 1788 76 1818 224
rect 1874 76 1904 224
rect 1968 76 1998 224
rect 2173 149 2203 233
rect 2286 85 2316 233
rect 2478 74 2508 158
rect 2577 74 2607 222
<< pmoshvt >>
rect 84 368 114 592
rect 174 368 204 592
rect 387 503 417 587
rect 507 503 537 587
rect 591 503 621 587
rect 693 503 723 587
rect 903 424 933 592
rect 981 424 1011 592
rect 1071 424 1101 592
rect 1267 424 1297 592
rect 1345 424 1375 592
rect 1453 508 1483 592
rect 1537 508 1567 592
rect 1763 392 1793 592
rect 1887 392 1917 592
rect 1971 392 2001 592
rect 2167 368 2197 496
rect 2272 368 2302 592
rect 2469 410 2499 578
rect 2574 368 2604 592
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 142 170 222
rect 114 108 125 142
rect 159 108 170 142
rect 114 74 170 108
rect 200 210 257 222
rect 200 176 211 210
rect 245 176 257 210
rect 200 120 257 176
rect 200 86 211 120
rect 245 86 257 120
rect 311 175 368 203
rect 311 141 323 175
rect 357 141 368 175
rect 311 119 368 141
rect 398 119 493 203
rect 523 119 565 203
rect 595 172 651 203
rect 595 138 606 172
rect 640 138 651 172
rect 595 119 651 138
rect 681 123 813 203
rect 681 119 737 123
rect 413 118 478 119
rect 200 74 257 86
rect 413 84 428 118
rect 462 84 478 118
rect 413 72 478 84
rect 696 89 737 119
rect 771 89 813 123
rect 867 165 924 229
rect 867 131 879 165
rect 913 131 924 165
rect 867 119 924 131
rect 954 193 1024 229
rect 954 159 979 193
rect 1013 159 1024 193
rect 954 119 1024 159
rect 1054 191 1124 229
rect 1054 157 1079 191
rect 1113 157 1124 191
rect 1054 119 1124 157
rect 1154 191 1224 229
rect 1154 157 1179 191
rect 1213 157 1224 191
rect 1154 119 1224 157
rect 1254 224 1304 229
rect 1254 119 1319 224
rect 1269 114 1319 119
rect 1349 186 1581 224
rect 1349 152 1360 186
rect 1394 152 1440 186
rect 1474 152 1520 186
rect 1554 152 1581 186
rect 1349 140 1581 152
rect 1611 140 1659 224
rect 1689 140 1788 224
rect 1349 114 1566 140
rect 1731 129 1788 140
rect 696 77 813 89
rect 1731 95 1743 129
rect 1777 95 1788 129
rect 1731 76 1788 95
rect 1818 129 1874 224
rect 1818 95 1829 129
rect 1863 95 1874 129
rect 1818 76 1874 95
rect 1904 153 1968 224
rect 1904 119 1919 153
rect 1953 119 1968 153
rect 1904 76 1968 119
rect 1998 85 2065 224
rect 2119 221 2173 233
rect 2119 187 2128 221
rect 2162 187 2173 221
rect 2119 149 2173 187
rect 2203 149 2286 233
rect 1998 76 2022 85
rect 2013 51 2022 76
rect 2056 51 2065 85
rect 2013 39 2065 51
rect 2218 85 2286 149
rect 2316 214 2370 233
rect 2316 180 2327 214
rect 2361 180 2370 214
rect 2316 131 2370 180
rect 2523 158 2577 222
rect 2316 97 2327 131
rect 2361 97 2370 131
rect 2316 85 2370 97
rect 2424 133 2478 158
rect 2424 99 2433 133
rect 2467 99 2478 133
rect 2218 51 2227 85
rect 2261 51 2271 85
rect 2424 74 2478 99
rect 2508 133 2577 158
rect 2508 99 2532 133
rect 2566 99 2577 133
rect 2508 74 2577 99
rect 2607 210 2661 222
rect 2607 176 2618 210
rect 2652 176 2661 210
rect 2607 120 2661 176
rect 2607 86 2618 120
rect 2652 86 2661 120
rect 2607 74 2661 86
rect 2218 39 2271 51
<< pdiff >>
rect 1585 628 1650 639
rect 27 580 84 592
rect 27 546 37 580
rect 71 546 84 580
rect 27 510 84 546
rect 27 476 37 510
rect 71 476 84 510
rect 27 440 84 476
rect 27 406 37 440
rect 71 406 84 440
rect 27 368 84 406
rect 114 580 174 592
rect 114 546 127 580
rect 161 546 174 580
rect 114 508 174 546
rect 114 474 127 508
rect 161 474 174 508
rect 114 368 174 474
rect 204 580 260 592
rect 1585 594 1600 628
rect 1634 594 1650 628
rect 1811 628 1869 639
rect 1585 592 1650 594
rect 1811 594 1823 628
rect 1857 594 1869 628
rect 1811 592 1869 594
rect 204 546 217 580
rect 251 546 260 580
rect 204 497 260 546
rect 204 463 217 497
rect 251 463 260 497
rect 314 531 387 587
rect 314 497 323 531
rect 357 503 387 531
rect 417 565 507 587
rect 417 531 459 565
rect 493 531 507 565
rect 417 503 507 531
rect 537 503 591 587
rect 621 547 693 587
rect 621 513 640 547
rect 674 513 693 547
rect 621 503 693 513
rect 723 531 793 587
rect 723 503 750 531
rect 357 497 369 503
rect 314 485 369 497
rect 741 497 750 503
rect 784 497 793 531
rect 204 414 260 463
rect 204 380 217 414
rect 251 380 260 414
rect 204 368 260 380
rect 741 485 793 497
rect 847 580 903 592
rect 847 546 856 580
rect 890 546 903 580
rect 847 495 903 546
rect 847 461 856 495
rect 890 461 903 495
rect 847 424 903 461
rect 933 424 981 592
rect 1011 573 1071 592
rect 1011 539 1024 573
rect 1058 539 1071 573
rect 1011 424 1071 539
rect 1101 580 1157 592
rect 1101 546 1114 580
rect 1148 546 1157 580
rect 1101 498 1157 546
rect 1101 464 1114 498
rect 1148 464 1157 498
rect 1101 424 1157 464
rect 1211 573 1267 592
rect 1211 539 1220 573
rect 1254 539 1267 573
rect 1211 424 1267 539
rect 1297 424 1345 592
rect 1375 580 1453 592
rect 1375 546 1388 580
rect 1422 546 1453 580
rect 1375 508 1453 546
rect 1483 508 1537 592
rect 1567 508 1650 592
rect 1704 578 1763 592
rect 1704 544 1716 578
rect 1750 544 1763 578
rect 1375 470 1434 508
rect 1375 436 1388 470
rect 1422 436 1434 470
rect 1375 424 1434 436
rect 1704 392 1763 544
rect 1793 392 1887 592
rect 1917 392 1971 592
rect 2001 580 2057 592
rect 2001 546 2014 580
rect 2048 546 2057 580
rect 2001 508 2057 546
rect 2215 578 2272 592
rect 2215 544 2225 578
rect 2259 544 2272 578
rect 2001 474 2014 508
rect 2048 474 2057 508
rect 2215 496 2272 544
rect 2001 392 2057 474
rect 2111 424 2167 496
rect 2111 390 2120 424
rect 2154 390 2167 424
rect 2111 368 2167 390
rect 2197 368 2272 496
rect 2302 580 2358 592
rect 2302 546 2315 580
rect 2349 546 2358 580
rect 2517 580 2574 592
rect 2517 578 2527 580
rect 2302 497 2358 546
rect 2302 463 2315 497
rect 2349 463 2358 497
rect 2302 414 2358 463
rect 2302 380 2315 414
rect 2349 380 2358 414
rect 2412 566 2469 578
rect 2412 532 2422 566
rect 2456 532 2469 566
rect 2412 456 2469 532
rect 2412 422 2422 456
rect 2456 422 2469 456
rect 2412 410 2469 422
rect 2499 546 2527 578
rect 2561 546 2574 580
rect 2499 497 2574 546
rect 2499 463 2527 497
rect 2561 463 2574 497
rect 2499 414 2574 463
rect 2499 410 2527 414
rect 2302 368 2358 380
rect 2517 380 2527 410
rect 2561 380 2574 414
rect 2517 368 2574 380
rect 2604 580 2661 592
rect 2604 546 2617 580
rect 2651 546 2661 580
rect 2604 497 2661 546
rect 2604 463 2617 497
rect 2651 463 2661 497
rect 2604 414 2661 463
rect 2604 380 2617 414
rect 2651 380 2661 414
rect 2604 368 2661 380
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 125 108 159 142
rect 211 176 245 210
rect 211 86 245 120
rect 323 141 357 175
rect 606 138 640 172
rect 428 84 462 118
rect 737 89 771 123
rect 879 131 913 165
rect 979 159 1013 193
rect 1079 157 1113 191
rect 1179 157 1213 191
rect 1360 152 1394 186
rect 1440 152 1474 186
rect 1520 152 1554 186
rect 1743 95 1777 129
rect 1829 95 1863 129
rect 1919 119 1953 153
rect 2128 187 2162 221
rect 2022 51 2056 85
rect 2327 180 2361 214
rect 2327 97 2361 131
rect 2433 99 2467 133
rect 2227 51 2261 85
rect 2532 99 2566 133
rect 2618 176 2652 210
rect 2618 86 2652 120
<< pdiffc >>
rect 37 546 71 580
rect 37 476 71 510
rect 37 406 71 440
rect 127 546 161 580
rect 127 474 161 508
rect 1600 594 1634 628
rect 1823 594 1857 628
rect 217 546 251 580
rect 217 463 251 497
rect 323 497 357 531
rect 459 531 493 565
rect 640 513 674 547
rect 750 497 784 531
rect 217 380 251 414
rect 856 546 890 580
rect 856 461 890 495
rect 1024 539 1058 573
rect 1114 546 1148 580
rect 1114 464 1148 498
rect 1220 539 1254 573
rect 1388 546 1422 580
rect 1716 544 1750 578
rect 1388 436 1422 470
rect 2014 546 2048 580
rect 2225 544 2259 578
rect 2014 474 2048 508
rect 2120 390 2154 424
rect 2315 546 2349 580
rect 2315 463 2349 497
rect 2315 380 2349 414
rect 2422 532 2456 566
rect 2422 422 2456 456
rect 2527 546 2561 580
rect 2527 463 2561 497
rect 2527 380 2561 414
rect 2617 546 2651 580
rect 2617 463 2651 497
rect 2617 380 2651 414
<< poly >>
rect 84 592 114 618
rect 174 592 204 618
rect 387 587 417 613
rect 507 587 537 613
rect 591 587 621 613
rect 693 587 723 613
rect 903 592 933 618
rect 981 592 1011 618
rect 1071 592 1101 618
rect 1267 592 1297 618
rect 1345 592 1375 618
rect 1453 592 1483 618
rect 1537 592 1567 618
rect 1763 592 1793 618
rect 1887 592 1917 618
rect 1971 592 2001 618
rect 2272 592 2302 618
rect 387 488 417 503
rect 507 488 537 503
rect 591 488 621 503
rect 693 488 723 503
rect 84 353 114 368
rect 174 353 204 368
rect 81 326 117 353
rect 171 326 207 353
rect 33 310 117 326
rect 33 276 49 310
rect 83 276 117 310
rect 33 260 117 276
rect 159 310 225 326
rect 159 276 175 310
rect 209 276 225 310
rect 384 302 420 488
rect 504 471 540 488
rect 588 471 624 488
rect 474 455 540 471
rect 474 421 490 455
rect 524 421 540 455
rect 474 405 540 421
rect 582 455 648 471
rect 582 421 598 455
rect 632 421 648 455
rect 582 405 648 421
rect 159 260 225 276
rect 368 286 451 302
rect 84 222 114 260
rect 170 222 200 260
rect 368 252 401 286
rect 435 252 451 286
rect 368 236 451 252
rect 368 203 398 236
rect 493 203 523 405
rect 690 393 726 488
rect 1453 493 1483 508
rect 1537 493 1567 508
rect 903 409 933 424
rect 981 409 1011 424
rect 1071 409 1101 424
rect 1267 409 1297 424
rect 1345 409 1375 424
rect 690 363 720 393
rect 565 333 720 363
rect 565 203 595 333
rect 762 329 828 345
rect 762 295 778 329
rect 812 309 828 329
rect 900 309 936 409
rect 978 387 1014 409
rect 1068 405 1104 409
rect 978 357 1026 387
rect 1068 376 1170 405
rect 1264 392 1300 409
rect 1068 375 1120 376
rect 996 333 1026 357
rect 1104 342 1120 375
rect 1154 342 1170 376
rect 996 317 1062 333
rect 1104 326 1170 342
rect 1224 376 1300 392
rect 1224 342 1240 376
rect 1274 342 1300 376
rect 1224 326 1300 342
rect 1342 386 1378 409
rect 1342 370 1408 386
rect 1342 336 1358 370
rect 1392 336 1408 370
rect 812 295 954 309
rect 637 275 703 291
rect 762 279 954 295
rect 637 241 653 275
rect 687 241 703 275
rect 637 225 703 241
rect 924 229 954 279
rect 996 283 1012 317
rect 1046 283 1062 317
rect 996 267 1062 283
rect 1024 229 1054 267
rect 1124 229 1154 326
rect 1224 229 1254 326
rect 1342 320 1408 336
rect 1450 360 1486 493
rect 1534 476 1570 493
rect 1534 460 1689 476
rect 1534 446 1594 460
rect 1578 426 1594 446
rect 1628 426 1689 460
rect 1578 410 1689 426
rect 1450 269 1480 360
rect 1319 239 1480 269
rect 1522 296 1611 312
rect 1522 262 1538 296
rect 1572 262 1611 296
rect 1522 246 1611 262
rect 651 203 681 225
rect 368 93 398 119
rect 493 93 523 119
rect 84 48 114 74
rect 170 51 200 74
rect 565 51 595 119
rect 651 93 681 119
rect 1319 224 1349 239
rect 1581 224 1611 246
rect 1659 224 1689 410
rect 2167 496 2197 522
rect 1763 377 1793 392
rect 1887 377 1917 392
rect 1971 377 2001 392
rect 1760 316 1796 377
rect 1746 300 1812 316
rect 1884 312 1920 377
rect 1968 350 2004 377
rect 2469 578 2499 604
rect 2574 592 2604 618
rect 2469 395 2499 410
rect 2167 353 2197 368
rect 2272 353 2302 368
rect 2423 365 2502 395
rect 1968 334 2034 350
rect 2164 336 2200 353
rect 1746 266 1762 300
rect 1796 280 1812 300
rect 1860 296 1926 312
rect 1796 266 1818 280
rect 1746 250 1818 266
rect 1788 224 1818 250
rect 1860 262 1876 296
rect 1910 262 1926 296
rect 1860 246 1926 262
rect 1968 300 1984 334
rect 2018 300 2034 334
rect 1968 284 2034 300
rect 2137 320 2203 336
rect 2269 330 2305 353
rect 2137 286 2153 320
rect 2187 286 2203 320
rect 1874 224 1904 246
rect 1968 224 1998 284
rect 2137 270 2203 286
rect 2173 233 2203 270
rect 2251 327 2317 330
rect 2423 327 2453 365
rect 2574 353 2604 368
rect 2251 314 2453 327
rect 2571 317 2607 353
rect 2251 280 2267 314
rect 2301 280 2453 314
rect 2251 264 2453 280
rect 2286 233 2316 264
rect 924 93 954 119
rect 1024 93 1054 119
rect 1124 93 1154 119
rect 1224 93 1254 119
rect 1581 114 1611 140
rect 1659 114 1689 140
rect 1319 51 1349 114
rect 2173 123 2203 149
rect 170 21 1349 51
rect 1788 50 1818 76
rect 1874 50 1904 76
rect 1968 50 1998 76
rect 2423 203 2453 264
rect 2501 301 2607 317
rect 2501 267 2517 301
rect 2551 267 2607 301
rect 2501 251 2607 267
rect 2577 222 2607 251
rect 2423 173 2508 203
rect 2478 158 2508 173
rect 2286 59 2316 85
rect 2478 48 2508 74
rect 2577 48 2607 74
<< polycont >>
rect 49 276 83 310
rect 175 276 209 310
rect 490 421 524 455
rect 598 421 632 455
rect 401 252 435 286
rect 778 295 812 329
rect 1120 342 1154 376
rect 1240 342 1274 376
rect 1358 336 1392 370
rect 653 241 687 275
rect 1012 283 1046 317
rect 1594 426 1628 460
rect 1538 262 1572 296
rect 1762 266 1796 300
rect 1876 262 1910 296
rect 1984 300 2018 334
rect 2153 286 2187 320
rect 2267 280 2301 314
rect 2517 267 2551 301
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2688 683
rect 21 580 87 596
rect 21 546 37 580
rect 71 546 87 580
rect 21 510 87 546
rect 21 476 37 510
rect 71 476 87 510
rect 21 440 87 476
rect 127 580 161 649
rect 127 508 161 546
rect 127 458 161 474
rect 201 581 425 615
rect 201 580 283 581
rect 201 546 217 580
rect 251 546 283 580
rect 201 497 283 546
rect 201 463 217 497
rect 251 463 283 497
rect 21 406 37 440
rect 71 424 87 440
rect 71 406 167 424
rect 21 390 167 406
rect 25 310 99 356
rect 25 276 49 310
rect 83 276 99 310
rect 25 260 99 276
rect 133 326 167 390
rect 201 414 283 463
rect 201 380 217 414
rect 251 380 283 414
rect 201 364 283 380
rect 133 310 215 326
rect 133 276 175 310
rect 209 276 215 310
rect 133 260 215 276
rect 133 226 167 260
rect 249 226 283 364
rect 23 210 167 226
rect 23 176 39 210
rect 73 192 167 210
rect 211 210 283 226
rect 23 120 73 176
rect 245 176 283 210
rect 23 86 39 120
rect 23 70 73 86
rect 109 142 175 158
rect 109 108 125 142
rect 159 108 175 142
rect 109 17 175 108
rect 211 120 283 176
rect 245 86 283 120
rect 317 531 357 547
rect 317 497 323 531
rect 317 481 357 497
rect 317 202 351 481
rect 391 371 425 581
rect 459 565 493 649
rect 459 505 493 531
rect 527 581 906 615
rect 527 471 561 581
rect 840 580 906 581
rect 618 513 640 547
rect 674 513 716 547
rect 474 455 561 471
rect 474 421 490 455
rect 524 421 561 455
rect 474 405 561 421
rect 595 455 648 471
rect 595 421 598 455
rect 632 421 648 455
rect 595 371 648 421
rect 391 337 648 371
rect 385 286 551 302
rect 385 252 401 286
rect 435 252 551 286
rect 385 236 551 252
rect 595 291 648 337
rect 682 359 716 513
rect 750 531 800 547
rect 784 497 800 531
rect 750 427 800 497
rect 840 546 856 580
rect 890 546 906 580
rect 840 498 906 546
rect 1008 573 1074 649
rect 1008 539 1024 573
rect 1058 539 1074 573
rect 1008 532 1074 539
rect 1114 580 1164 596
rect 1148 546 1164 580
rect 1114 498 1164 546
rect 1204 573 1270 649
rect 1581 628 1654 649
rect 1204 539 1220 573
rect 1254 539 1270 573
rect 1204 532 1270 539
rect 1372 580 1483 596
rect 1581 594 1600 628
rect 1634 594 1654 628
rect 1807 628 1873 649
rect 1372 546 1388 580
rect 1422 546 1483 580
rect 1700 578 1766 596
rect 1807 594 1823 628
rect 1857 594 1873 628
rect 1700 560 1716 578
rect 840 495 1114 498
rect 840 461 856 495
rect 890 464 1114 495
rect 1148 464 1290 498
rect 890 461 963 464
rect 750 393 895 427
rect 682 329 827 359
rect 682 325 778 329
rect 727 295 778 325
rect 812 295 827 329
rect 595 276 693 291
rect 595 242 607 276
rect 641 275 693 276
rect 641 242 653 275
rect 595 241 653 242
rect 687 241 693 275
rect 595 225 693 241
rect 727 279 827 295
rect 317 175 550 202
rect 727 191 761 279
rect 861 233 895 393
rect 317 141 323 175
rect 357 168 550 175
rect 357 141 373 168
rect 317 115 373 141
rect 409 118 482 134
rect 211 70 283 86
rect 409 84 428 118
rect 462 84 482 118
rect 409 17 482 84
rect 516 85 550 168
rect 590 172 761 191
rect 590 138 606 172
rect 640 157 761 172
rect 795 199 895 233
rect 929 233 963 461
rect 1087 424 1127 430
rect 1121 392 1127 424
rect 1121 390 1170 392
rect 1087 376 1170 390
rect 1087 342 1120 376
rect 1154 342 1170 376
rect 1087 335 1170 342
rect 1224 376 1290 464
rect 1372 470 1483 546
rect 1372 436 1388 470
rect 1422 436 1483 470
rect 1372 420 1483 436
rect 1224 342 1240 376
rect 1274 342 1290 376
rect 1224 335 1290 342
rect 1342 370 1415 386
rect 1342 336 1358 370
rect 1392 336 1415 370
rect 1449 380 1483 420
rect 1578 544 1716 560
rect 1750 560 1766 578
rect 1998 580 2064 596
rect 1998 560 2014 580
rect 1750 546 2014 560
rect 2048 546 2064 580
rect 1750 544 2064 546
rect 1578 526 2064 544
rect 2209 578 2275 649
rect 2209 544 2225 578
rect 2259 544 2275 578
rect 2209 526 2275 544
rect 2315 580 2385 596
rect 2349 546 2385 580
rect 1578 460 1644 526
rect 1998 508 2064 526
rect 1578 426 1594 460
rect 1628 426 1644 460
rect 1578 414 1644 426
rect 1678 458 1880 492
rect 1998 474 2014 508
rect 2048 492 2064 508
rect 2315 497 2385 546
rect 2048 474 2277 492
rect 1998 458 2277 474
rect 1678 380 1712 458
rect 1846 424 1880 458
rect 1449 346 1712 380
rect 1746 390 1759 424
rect 1793 390 1812 424
rect 1846 390 2034 424
rect 997 317 1053 333
rect 997 283 1012 317
rect 1046 301 1053 317
rect 1342 312 1415 336
rect 1046 283 1297 301
rect 997 267 1297 283
rect 929 199 1029 233
rect 640 138 656 157
rect 590 119 656 138
rect 795 123 829 199
rect 963 193 1029 199
rect 692 89 737 123
rect 771 89 829 123
rect 692 85 829 89
rect 516 51 829 85
rect 863 131 879 165
rect 913 131 929 165
rect 963 159 979 193
rect 1013 159 1029 193
rect 963 143 1029 159
rect 1063 191 1129 207
rect 1063 157 1079 191
rect 1113 157 1129 191
rect 863 85 929 131
rect 1063 85 1129 157
rect 863 51 1129 85
rect 1163 191 1229 207
rect 1163 157 1179 191
rect 1213 157 1229 191
rect 1163 17 1229 157
rect 1263 102 1297 267
rect 1342 296 1573 312
rect 1342 276 1538 296
rect 1342 242 1375 276
rect 1409 262 1538 276
rect 1572 262 1573 296
rect 1409 242 1573 262
rect 1342 236 1573 242
rect 1607 202 1641 346
rect 1746 300 1812 390
rect 1968 334 2034 390
rect 1746 266 1762 300
rect 1796 266 1812 300
rect 1746 255 1812 266
rect 1860 296 1926 312
rect 1860 262 1876 296
rect 1910 262 1926 296
rect 1968 300 1984 334
rect 2018 300 2034 334
rect 1968 284 2034 300
rect 2069 390 2120 424
rect 2154 390 2170 424
rect 1860 221 1926 262
rect 2069 221 2103 390
rect 2137 320 2203 356
rect 2137 286 2153 320
rect 2187 286 2203 320
rect 2137 270 2203 286
rect 2243 330 2277 458
rect 2349 463 2385 497
rect 2315 414 2385 463
rect 2349 380 2385 414
rect 2315 364 2385 380
rect 2243 314 2317 330
rect 2243 280 2267 314
rect 2301 280 2317 314
rect 2243 264 2317 280
rect 1344 186 1641 202
rect 1344 152 1360 186
rect 1394 152 1440 186
rect 1474 152 1520 186
rect 1554 152 1641 186
rect 1344 136 1641 152
rect 1675 187 2128 221
rect 2162 187 2178 221
rect 1675 102 1709 187
rect 2243 153 2277 264
rect 2351 230 2385 364
rect 1263 68 1709 102
rect 1743 129 1777 153
rect 1743 17 1777 95
rect 1813 129 1863 153
rect 1813 95 1829 129
rect 1899 119 1919 153
rect 1953 119 2277 153
rect 2311 214 2385 230
rect 2311 180 2327 214
rect 2361 180 2385 214
rect 2311 131 2385 180
rect 1813 85 1863 95
rect 2311 97 2327 131
rect 2361 97 2385 131
rect 1813 51 2022 85
rect 2056 51 2072 85
rect 2211 51 2227 85
rect 2261 51 2277 85
rect 2311 81 2385 97
rect 2422 566 2472 582
rect 2456 532 2472 566
rect 2422 456 2472 532
rect 2456 422 2472 456
rect 2422 317 2472 422
rect 2511 580 2561 649
rect 2511 546 2527 580
rect 2511 497 2561 546
rect 2511 463 2527 497
rect 2511 414 2561 463
rect 2511 380 2527 414
rect 2511 364 2561 380
rect 2601 580 2668 596
rect 2601 546 2617 580
rect 2651 546 2668 580
rect 2601 497 2668 546
rect 2601 463 2617 497
rect 2651 463 2668 497
rect 2601 414 2668 463
rect 2601 380 2617 414
rect 2651 380 2668 414
rect 2422 301 2567 317
rect 2422 267 2517 301
rect 2551 267 2567 301
rect 2422 251 2567 267
rect 2422 133 2472 251
rect 2601 210 2668 380
rect 2601 176 2618 210
rect 2652 176 2668 210
rect 2422 99 2433 133
rect 2467 99 2472 133
rect 2422 70 2472 99
rect 2516 133 2566 162
rect 2516 99 2532 133
rect 2211 17 2277 51
rect 2516 17 2566 99
rect 2601 120 2668 176
rect 2601 86 2618 120
rect 2652 86 2668 120
rect 2601 70 2668 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2688 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 607 242 641 276
rect 1087 390 1121 424
rect 1759 390 1793 424
rect 1375 242 1409 276
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
<< metal1 >>
rect 0 683 2688 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2688 683
rect 0 617 2688 649
rect 1075 424 1133 430
rect 1075 390 1087 424
rect 1121 421 1133 424
rect 1747 424 1805 430
rect 1747 421 1759 424
rect 1121 393 1759 421
rect 1121 390 1133 393
rect 1075 384 1133 390
rect 1747 390 1759 393
rect 1793 390 1805 424
rect 1747 384 1805 390
rect 595 276 653 282
rect 595 242 607 276
rect 641 273 653 276
rect 1363 276 1421 282
rect 1363 273 1375 276
rect 641 245 1375 273
rect 641 242 653 245
rect 595 236 653 242
rect 1363 242 1375 245
rect 1409 242 1421 276
rect 1363 236 1421 242
rect 0 17 2688 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2688 17
rect 0 -49 2688 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dfbbn_1
flabel pwell s 0 0 2688 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nwell s 0 617 2688 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 1759 390 1793 424 0 FreeSans 340 0 0 0 SET_B
port 4 nsew
flabel metal1 s 0 617 2688 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 2688 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 2623 94 2657 128 0 FreeSans 340 0 0 0 Q
port 9 nsew
flabel corelocali s 2623 168 2657 202 0 FreeSans 340 0 0 0 Q
port 9 nsew
flabel corelocali s 2623 242 2657 276 0 FreeSans 340 0 0 0 Q
port 9 nsew
flabel corelocali s 2623 316 2657 350 0 FreeSans 340 0 0 0 Q
port 9 nsew
flabel corelocali s 2623 390 2657 424 0 FreeSans 340 0 0 0 Q
port 9 nsew
flabel corelocali s 2623 464 2657 498 0 FreeSans 340 0 0 0 Q
port 9 nsew
flabel corelocali s 2623 538 2657 572 0 FreeSans 340 0 0 0 Q
port 9 nsew
flabel corelocali s 415 242 449 276 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 511 242 545 276 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 2143 316 2177 350 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 CLK_N
port 1 nsew
flabel corelocali s 2335 390 2369 424 0 FreeSans 340 0 0 0 Q_N
port 10 nsew
flabel corelocali s 2335 464 2369 498 0 FreeSans 340 0 0 0 Q_N
port 10 nsew
flabel corelocali s 2335 538 2369 572 0 FreeSans 340 0 0 0 Q_N
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 2688 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2489012
string GDS_START 2468464
<< end >>
