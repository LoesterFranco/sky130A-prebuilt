magic
tech sky130A
magscale 1 2
timestamp 1601050039
<< nwell >>
rect -38 261 590 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 80 47 110 131
rect 177 47 207 131
rect 263 47 293 131
rect 349 47 379 131
rect 435 47 465 131
<< pmoshvt >>
rect 80 297 110 497
rect 176 297 206 497
rect 262 297 292 497
rect 348 297 378 497
rect 434 297 464 497
<< ndiff >>
rect 27 101 80 131
rect 27 67 35 101
rect 69 67 80 101
rect 27 47 80 67
rect 110 97 177 131
rect 110 63 121 97
rect 155 63 177 97
rect 110 47 177 63
rect 207 119 263 131
rect 207 85 218 119
rect 252 85 263 119
rect 207 47 263 85
rect 293 97 349 131
rect 293 63 304 97
rect 338 63 349 97
rect 293 47 349 63
rect 379 119 435 131
rect 379 85 390 119
rect 424 85 435 119
rect 379 47 435 85
rect 465 97 523 131
rect 465 63 476 97
rect 510 63 523 97
rect 465 47 523 63
<< pdiff >>
rect 27 477 80 497
rect 27 443 35 477
rect 69 443 80 477
rect 27 355 80 443
rect 27 321 35 355
rect 69 321 80 355
rect 27 297 80 321
rect 110 485 176 497
rect 110 451 121 485
rect 155 451 176 485
rect 110 417 176 451
rect 110 383 121 417
rect 155 383 176 417
rect 110 297 176 383
rect 206 450 262 497
rect 206 416 217 450
rect 251 416 262 450
rect 206 297 262 416
rect 292 485 348 497
rect 292 451 303 485
rect 337 451 348 485
rect 292 297 348 451
rect 378 477 434 497
rect 378 443 389 477
rect 423 443 434 477
rect 378 409 434 443
rect 378 375 389 409
rect 423 375 434 409
rect 378 341 434 375
rect 378 307 389 341
rect 423 307 434 341
rect 378 297 434 307
rect 464 471 524 497
rect 464 437 475 471
rect 509 437 524 471
rect 464 403 524 437
rect 464 369 475 403
rect 509 369 524 403
rect 464 297 524 369
<< ndiffc >>
rect 35 67 69 101
rect 121 63 155 97
rect 218 85 252 119
rect 304 63 338 97
rect 390 85 424 119
rect 476 63 510 97
<< pdiffc >>
rect 35 443 69 477
rect 35 321 69 355
rect 121 451 155 485
rect 121 383 155 417
rect 217 416 251 450
rect 303 451 337 485
rect 389 443 423 477
rect 389 375 423 409
rect 389 307 423 341
rect 475 437 509 471
rect 475 369 509 403
<< poly >>
rect 80 497 110 523
rect 176 497 206 523
rect 262 497 292 523
rect 348 497 378 523
rect 434 497 464 523
rect 80 265 110 297
rect 69 249 129 265
rect 69 215 85 249
rect 119 215 129 249
rect 69 199 129 215
rect 176 259 206 297
rect 262 259 292 297
rect 348 259 378 297
rect 434 259 464 297
rect 176 249 464 259
rect 176 215 231 249
rect 265 215 299 249
rect 333 215 367 249
rect 401 237 464 249
rect 401 215 465 237
rect 176 210 465 215
rect 177 204 465 210
rect 80 131 110 199
rect 177 131 207 204
rect 263 131 293 204
rect 349 131 379 204
rect 435 131 465 204
rect 80 21 110 47
rect 177 21 207 47
rect 263 21 293 47
rect 349 21 379 47
rect 435 21 465 47
<< polycont >>
rect 85 215 119 249
rect 231 215 265 249
rect 299 215 333 249
rect 367 215 401 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 17 477 79 493
rect 17 443 35 477
rect 69 443 79 477
rect 17 355 79 443
rect 113 485 175 527
rect 113 451 121 485
rect 155 451 175 485
rect 113 417 175 451
rect 113 383 121 417
rect 155 383 175 417
rect 113 367 175 383
rect 209 450 261 493
rect 209 416 217 450
rect 251 416 261 450
rect 295 485 346 527
rect 295 451 303 485
rect 337 451 346 485
rect 295 435 346 451
rect 381 477 433 493
rect 381 443 389 477
rect 423 443 433 477
rect 209 401 261 416
rect 381 409 433 443
rect 381 401 389 409
rect 209 375 389 401
rect 423 375 433 409
rect 209 367 433 375
rect 17 321 35 355
rect 69 333 79 355
rect 381 341 433 367
rect 467 471 524 527
rect 467 437 475 471
rect 509 437 524 471
rect 467 403 524 437
rect 467 369 475 403
rect 509 369 524 403
rect 467 353 524 369
rect 69 321 223 333
rect 17 299 223 321
rect 17 117 51 299
rect 85 249 155 265
rect 119 215 155 249
rect 189 249 223 299
rect 381 307 389 341
rect 423 317 433 341
rect 423 307 532 317
rect 381 283 532 307
rect 189 215 231 249
rect 265 215 299 249
rect 333 215 367 249
rect 401 215 417 249
rect 85 151 155 215
rect 451 181 532 283
rect 202 147 532 181
rect 202 119 261 147
rect 17 101 77 117
rect 17 67 35 101
rect 69 67 77 101
rect 17 51 77 67
rect 111 97 166 113
rect 111 63 121 97
rect 155 63 166 97
rect 202 85 218 119
rect 252 85 261 119
rect 381 119 433 147
rect 202 69 261 85
rect 295 97 346 113
rect 111 17 166 63
rect 295 63 304 97
rect 338 63 346 97
rect 381 85 390 119
rect 424 85 433 119
rect 381 69 433 85
rect 467 97 523 113
rect 295 17 346 63
rect 467 63 476 97
rect 510 63 523 97
rect 467 17 523 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
flabel corelocali s 397 289 431 323 0 FreeSans 200 0 0 0 X
port 6 nsew
flabel corelocali s 121 153 155 187 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 489 153 523 187 0 FreeSans 200 0 0 0 X
port 6 nsew
flabel corelocali s 121 221 155 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 489 221 523 255 0 FreeSans 200 0 0 0 X
port 6 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew
rlabel comment s 0 0 0 0 4 clkbuf_4
<< properties >>
string FIXED_BBOX 0 0 552 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3168094
string GDS_START 3162938
string path 0.000 13.600 13.800 13.600 
<< end >>
