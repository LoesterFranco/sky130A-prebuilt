magic
tech sky130A
magscale 1 2
timestamp 1601050082
<< locali >>
rect 474 424 524 547
rect 664 424 730 547
rect 876 424 942 596
rect 474 404 942 424
rect 1059 404 1125 596
rect 474 390 1125 404
rect 25 270 359 356
rect 505 270 743 356
rect 793 236 839 390
rect 876 370 1125 390
rect 1273 290 1415 356
rect 793 202 1119 236
rect 853 119 919 202
rect 1053 119 1119 202
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 24 424 74 596
rect 114 458 164 649
rect 204 424 254 596
rect 294 458 360 649
rect 400 581 830 615
rect 400 424 434 581
rect 24 390 434 424
rect 564 458 630 581
rect 764 458 830 581
rect 982 438 1016 649
rect 1171 458 1221 649
rect 1261 424 1311 596
rect 400 364 434 390
rect 1159 390 1311 424
rect 1351 420 1417 649
rect 1159 336 1193 390
rect 874 270 1193 336
rect 1159 256 1193 270
rect 23 202 615 236
rect 1159 222 1315 256
rect 23 70 73 202
rect 109 17 175 168
rect 221 70 255 202
rect 291 17 357 168
rect 393 70 427 202
rect 565 168 615 202
rect 463 17 529 168
rect 565 134 819 168
rect 565 70 615 134
rect 651 17 717 100
rect 753 85 819 134
rect 953 85 1019 168
rect 1153 85 1219 188
rect 1265 100 1315 222
rect 753 51 1219 85
rect 1351 17 1417 256
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 683 1440 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 0 617 1440 649
rect 0 17 1440 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -49 1440 -17
<< labels >>
rlabel locali s 25 270 359 356 6 A1
port 1 nsew signal input
rlabel locali s 505 270 743 356 6 A2
port 2 nsew signal input
rlabel locali s 1273 290 1415 356 6 B1_N
port 3 nsew signal input
rlabel locali s 1059 404 1125 596 6 Y
port 4 nsew signal output
rlabel locali s 1053 119 1119 202 6 Y
port 4 nsew signal output
rlabel locali s 876 424 942 596 6 Y
port 4 nsew signal output
rlabel locali s 876 370 1125 390 6 Y
port 4 nsew signal output
rlabel locali s 853 119 919 202 6 Y
port 4 nsew signal output
rlabel locali s 793 236 839 390 6 Y
port 4 nsew signal output
rlabel locali s 793 202 1119 236 6 Y
port 4 nsew signal output
rlabel locali s 664 424 730 547 6 Y
port 4 nsew signal output
rlabel locali s 474 424 524 547 6 Y
port 4 nsew signal output
rlabel locali s 474 404 942 424 6 Y
port 4 nsew signal output
rlabel locali s 474 390 1125 404 6 Y
port 4 nsew signal output
rlabel metal1 s 0 -49 1440 49 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1440 715 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1440 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1418522
string GDS_START 1406270
<< end >>
