magic
tech sky130A
magscale 1 2
timestamp 1604502741
<< locali >>
rect 310 424 365 596
rect 552 424 618 596
rect 752 424 818 596
rect 972 424 1038 596
rect 310 390 1038 424
rect 310 370 365 390
rect 552 364 647 390
rect 25 236 197 302
rect 409 270 518 356
rect 601 236 647 364
rect 697 270 839 356
rect 889 270 1127 356
rect 307 202 647 236
rect 307 160 379 202
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 101 370 167 572
rect 208 404 274 649
rect 399 458 518 649
rect 652 458 718 649
rect 864 458 930 649
rect 1072 390 1129 649
rect 101 336 265 370
rect 231 270 344 336
rect 231 202 265 270
rect 23 168 265 202
rect 23 70 73 168
rect 715 186 1129 236
rect 415 134 669 168
rect 109 17 175 134
rect 415 126 465 134
rect 221 70 465 126
rect 603 119 669 134
rect 715 119 765 186
rect 501 85 567 100
rect 801 85 867 152
rect 501 51 867 85
rect 901 80 939 186
rect 973 17 1039 152
rect 1079 80 1129 186
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
rlabel locali s 25 236 197 302 6 A_N
port 1 nsew signal input
rlabel locali s 409 270 518 356 6 B
port 2 nsew signal input
rlabel locali s 697 270 839 356 6 C
port 3 nsew signal input
rlabel locali s 889 270 1127 356 6 D
port 4 nsew signal input
rlabel locali s 972 424 1038 596 6 Y
port 5 nsew signal output
rlabel locali s 752 424 818 596 6 Y
port 5 nsew signal output
rlabel locali s 601 236 647 364 6 Y
port 5 nsew signal output
rlabel locali s 552 424 618 596 6 Y
port 5 nsew signal output
rlabel locali s 552 364 647 390 6 Y
port 5 nsew signal output
rlabel locali s 310 424 365 596 6 Y
port 5 nsew signal output
rlabel locali s 310 390 1038 424 6 Y
port 5 nsew signal output
rlabel locali s 310 370 365 390 6 Y
port 5 nsew signal output
rlabel locali s 307 202 647 236 6 Y
port 5 nsew signal output
rlabel locali s 307 160 379 202 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -49 1152 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 1152 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1425384
string GDS_START 1415482
<< end >>
