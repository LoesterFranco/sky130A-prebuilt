magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 216 340 252 493
rect 408 340 446 493
rect 17 287 446 340
rect 17 161 73 287
rect 558 289 920 337
rect 558 199 617 289
rect 651 207 818 255
rect 854 207 920 289
rect 965 299 1363 337
rect 965 207 1031 299
rect 1068 207 1223 265
rect 1260 207 1363 299
rect 17 127 351 161
rect 129 123 351 127
rect 129 51 163 123
rect 317 51 351 123
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 96 374 172 527
rect 288 374 364 527
rect 480 440 556 527
rect 600 405 672 493
rect 707 439 783 527
rect 817 405 883 493
rect 919 439 972 527
rect 1093 405 1169 493
rect 480 371 1169 405
rect 1285 383 1361 527
rect 480 253 524 371
rect 107 213 524 253
rect 480 163 524 213
rect 480 127 764 163
rect 895 139 1361 173
rect 19 17 85 93
rect 207 17 273 89
rect 895 93 961 139
rect 385 17 468 93
rect 516 51 961 93
rect 996 17 1059 105
rect 1093 51 1169 139
rect 1213 17 1251 105
rect 1285 51 1361 139
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
<< metal1 >>
rect 0 561 1380 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 0 496 1380 527
rect 0 17 1380 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
rect 0 -48 1380 -17
<< labels >>
rlabel locali s 1260 207 1363 299 6 A1
port 1 nsew signal input
rlabel locali s 965 299 1363 337 6 A1
port 1 nsew signal input
rlabel locali s 965 207 1031 299 6 A1
port 1 nsew signal input
rlabel locali s 1068 207 1223 265 6 A2
port 2 nsew signal input
rlabel locali s 854 207 920 289 6 B1
port 3 nsew signal input
rlabel locali s 558 289 920 337 6 B1
port 3 nsew signal input
rlabel locali s 558 199 617 289 6 B1
port 3 nsew signal input
rlabel locali s 651 207 818 255 6 C1
port 4 nsew signal input
rlabel locali s 408 340 446 493 6 X
port 5 nsew signal output
rlabel locali s 317 51 351 123 6 X
port 5 nsew signal output
rlabel locali s 216 340 252 493 6 X
port 5 nsew signal output
rlabel locali s 129 123 351 127 6 X
port 5 nsew signal output
rlabel locali s 129 51 163 123 6 X
port 5 nsew signal output
rlabel locali s 17 287 446 340 6 X
port 5 nsew signal output
rlabel locali s 17 161 73 287 6 X
port 5 nsew signal output
rlabel locali s 17 127 351 161 6 X
port 5 nsew signal output
rlabel metal1 s 0 -48 1380 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 1380 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1380 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2584542
string GDS_START 2575002
<< end >>
