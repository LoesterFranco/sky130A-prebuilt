magic
tech sky130A
magscale 1 2
timestamp 1604502705
<< nwell >>
rect -38 332 518 704
<< pwell >>
rect 0 0 480 49
<< scnmos >>
rect 83 94 113 222
rect 169 94 199 222
rect 270 74 300 222
rect 356 74 386 222
<< pmoshvt >>
rect 84 368 114 568
rect 162 368 192 568
rect 270 368 300 592
rect 364 368 394 592
<< ndiff >>
rect 27 184 83 222
rect 27 150 38 184
rect 72 150 83 184
rect 27 94 83 150
rect 113 210 169 222
rect 113 176 124 210
rect 158 176 169 210
rect 113 140 169 176
rect 113 106 124 140
rect 158 106 169 140
rect 113 94 169 106
rect 199 147 270 222
rect 199 113 225 147
rect 259 113 270 147
rect 199 94 270 113
rect 214 74 270 94
rect 300 210 356 222
rect 300 176 311 210
rect 345 176 356 210
rect 300 120 356 176
rect 300 86 311 120
rect 345 86 356 120
rect 300 74 356 86
rect 386 210 453 222
rect 386 176 410 210
rect 444 176 453 210
rect 386 120 453 176
rect 386 86 410 120
rect 444 86 453 120
rect 386 74 453 86
<< pdiff >>
rect 211 573 270 592
rect 211 568 223 573
rect 27 556 84 568
rect 27 522 37 556
rect 71 522 84 556
rect 27 485 84 522
rect 27 451 37 485
rect 71 451 84 485
rect 27 414 84 451
rect 27 380 37 414
rect 71 380 84 414
rect 27 368 84 380
rect 114 368 162 568
rect 192 539 223 568
rect 257 539 270 573
rect 192 368 270 539
rect 300 414 364 592
rect 300 380 315 414
rect 349 380 364 414
rect 300 368 364 380
rect 394 573 453 592
rect 394 539 407 573
rect 441 539 453 573
rect 394 368 453 539
<< ndiffc >>
rect 38 150 72 184
rect 124 176 158 210
rect 124 106 158 140
rect 225 113 259 147
rect 311 176 345 210
rect 311 86 345 120
rect 410 176 444 210
rect 410 86 444 120
<< pdiffc >>
rect 37 522 71 556
rect 37 451 71 485
rect 37 380 71 414
rect 223 539 257 573
rect 315 380 349 414
rect 407 539 441 573
<< poly >>
rect 84 568 114 594
rect 162 568 192 594
rect 270 592 300 618
rect 364 592 394 618
rect 84 353 114 368
rect 162 353 192 368
rect 270 353 300 368
rect 364 353 394 368
rect 81 310 117 353
rect 21 294 117 310
rect 21 260 37 294
rect 71 260 117 294
rect 159 336 195 353
rect 159 320 225 336
rect 159 286 175 320
rect 209 286 225 320
rect 159 270 225 286
rect 267 326 303 353
rect 361 326 397 353
rect 267 310 459 326
rect 267 276 409 310
rect 443 276 459 310
rect 21 244 117 260
rect 83 222 113 244
rect 169 222 199 270
rect 267 260 459 276
rect 270 222 300 260
rect 356 222 386 260
rect 83 68 113 94
rect 169 68 199 94
rect 270 48 300 74
rect 356 48 386 74
<< polycont >>
rect 37 260 71 294
rect 175 286 209 320
rect 409 276 443 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 207 573 273 649
rect 21 556 87 572
rect 21 522 37 556
rect 71 522 87 556
rect 207 539 223 573
rect 257 539 273 573
rect 207 532 273 539
rect 391 573 457 649
rect 391 539 407 573
rect 441 539 457 573
rect 391 532 457 539
rect 21 498 87 522
rect 21 485 459 498
rect 21 451 37 485
rect 71 464 459 485
rect 71 451 87 464
rect 21 414 87 451
rect 21 380 37 414
rect 71 380 87 414
rect 21 364 87 380
rect 121 320 209 430
rect 21 294 87 310
rect 21 260 37 294
rect 71 260 87 294
rect 121 286 175 320
rect 121 270 209 286
rect 21 236 87 260
rect 243 236 277 464
rect 124 210 277 236
rect 22 184 88 200
rect 22 150 38 184
rect 72 150 88 184
rect 22 17 88 150
rect 158 202 277 210
rect 311 414 367 430
rect 311 380 315 414
rect 349 380 367 414
rect 311 364 367 380
rect 311 210 359 364
rect 425 326 459 464
rect 393 310 459 326
rect 393 276 409 310
rect 443 276 459 310
rect 393 260 459 276
rect 158 176 174 202
rect 124 140 174 176
rect 345 176 359 210
rect 158 106 174 140
rect 124 90 174 106
rect 209 147 275 165
rect 209 113 225 147
rect 259 113 275 147
rect 209 17 275 113
rect 311 120 359 176
rect 345 86 359 120
rect 311 70 359 86
rect 394 210 460 226
rect 394 176 410 210
rect 444 176 460 210
rect 394 120 460 176
rect 394 86 410 120
rect 444 86 460 120
rect 394 17 460 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< metal1 >>
rect 0 683 480 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 0 617 480 649
rect 0 17 480 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
rect 0 -49 480 -17
<< labels >>
rlabel comment s 0 0 0 0 4 or2_2
flabel pwell s 0 0 480 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 0 617 480 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 0 617 480 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 480 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 319 94 353 128 0 FreeSans 340 0 0 0 X
port 7 nsew
flabel corelocali s 319 168 353 202 0 FreeSans 340 0 0 0 X
port 7 nsew
flabel corelocali s 319 242 353 276 0 FreeSans 340 0 0 0 X
port 7 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 X
port 7 nsew
flabel corelocali s 319 390 353 424 0 FreeSans 340 0 0 0 X
port 7 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 127 390 161 424 0 FreeSans 340 0 0 0 A
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 480 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1022090
string GDS_START 1016766
<< end >>
