magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 1694 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 89 47 119 177
rect 183 47 213 177
rect 277 47 307 177
rect 361 47 391 177
rect 455 47 485 177
rect 549 47 579 177
rect 653 47 683 177
rect 747 47 777 177
rect 831 47 861 177
rect 948 47 978 177
rect 1044 47 1074 177
rect 1139 47 1169 177
rect 1233 47 1263 177
rect 1327 47 1357 177
rect 1421 47 1451 177
rect 1517 47 1547 177
<< pmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 457 297 493 497
rect 551 297 587 497
rect 645 297 681 497
rect 739 297 775 497
rect 833 297 869 497
rect 927 297 963 497
rect 1021 297 1057 497
rect 1121 297 1157 497
rect 1217 297 1253 497
rect 1313 297 1349 497
rect 1413 297 1449 497
rect 1515 297 1551 497
<< ndiff >>
rect 27 93 89 177
rect 27 59 35 93
rect 69 59 89 93
rect 27 47 89 59
rect 119 157 183 177
rect 119 123 129 157
rect 163 123 183 157
rect 119 47 183 123
rect 213 89 277 177
rect 213 55 223 89
rect 257 55 277 89
rect 213 47 277 55
rect 307 89 361 177
rect 307 55 317 89
rect 351 55 361 89
rect 307 47 361 55
rect 391 169 455 177
rect 391 135 411 169
rect 445 135 455 169
rect 391 47 455 135
rect 485 89 549 177
rect 485 55 505 89
rect 539 55 549 89
rect 485 47 549 55
rect 579 169 653 177
rect 579 135 599 169
rect 633 135 653 169
rect 579 47 653 135
rect 683 89 747 177
rect 683 55 693 89
rect 727 55 747 89
rect 683 47 747 55
rect 777 89 831 177
rect 777 55 787 89
rect 821 55 831 89
rect 777 47 831 55
rect 861 169 948 177
rect 861 135 885 169
rect 919 135 948 169
rect 861 101 948 135
rect 861 67 885 101
rect 919 67 948 101
rect 861 47 948 67
rect 978 89 1044 177
rect 978 55 989 89
rect 1023 55 1044 89
rect 978 47 1044 55
rect 1074 169 1139 177
rect 1074 135 1085 169
rect 1119 135 1139 169
rect 1074 101 1139 135
rect 1074 67 1085 101
rect 1119 67 1139 101
rect 1074 47 1139 67
rect 1169 89 1233 177
rect 1169 55 1179 89
rect 1213 55 1233 89
rect 1169 47 1233 55
rect 1263 169 1327 177
rect 1263 135 1273 169
rect 1307 135 1327 169
rect 1263 101 1327 135
rect 1263 67 1273 101
rect 1307 67 1327 101
rect 1263 47 1327 67
rect 1357 89 1421 177
rect 1357 55 1367 89
rect 1401 55 1421 89
rect 1357 47 1421 55
rect 1451 165 1517 177
rect 1451 131 1463 165
rect 1497 131 1517 165
rect 1451 47 1517 131
rect 1547 89 1605 177
rect 1547 55 1559 89
rect 1593 55 1605 89
rect 1547 47 1605 55
<< pdiff >>
rect 27 477 81 497
rect 27 443 35 477
rect 69 443 81 477
rect 27 409 81 443
rect 27 375 35 409
rect 69 375 81 409
rect 27 297 81 375
rect 117 485 175 497
rect 117 451 129 485
rect 163 451 175 485
rect 117 297 175 451
rect 211 477 269 497
rect 211 443 223 477
rect 257 443 269 477
rect 211 409 269 443
rect 211 375 223 409
rect 257 375 269 409
rect 211 297 269 375
rect 305 489 363 497
rect 305 455 317 489
rect 351 455 363 489
rect 305 297 363 455
rect 399 477 457 497
rect 399 443 411 477
rect 445 443 457 477
rect 399 409 457 443
rect 399 375 411 409
rect 445 375 457 409
rect 399 297 457 375
rect 493 489 551 497
rect 493 455 505 489
rect 539 455 551 489
rect 493 297 551 455
rect 587 477 645 497
rect 587 443 599 477
rect 633 443 645 477
rect 587 409 645 443
rect 587 375 599 409
rect 633 375 645 409
rect 587 297 645 375
rect 681 489 739 497
rect 681 455 693 489
rect 727 455 739 489
rect 681 297 739 455
rect 775 477 833 497
rect 775 443 787 477
rect 821 443 833 477
rect 775 409 833 443
rect 775 375 787 409
rect 821 375 833 409
rect 775 297 833 375
rect 869 417 927 497
rect 869 383 881 417
rect 915 383 927 417
rect 869 297 927 383
rect 963 489 1021 497
rect 963 455 975 489
rect 1009 455 1021 489
rect 963 297 1021 455
rect 1057 297 1121 497
rect 1157 413 1217 497
rect 1157 379 1170 413
rect 1204 379 1217 413
rect 1157 297 1217 379
rect 1253 339 1313 497
rect 1253 305 1266 339
rect 1300 305 1313 339
rect 1253 297 1313 305
rect 1349 413 1413 497
rect 1349 379 1366 413
rect 1400 379 1413 413
rect 1349 297 1413 379
rect 1449 297 1515 497
rect 1551 485 1605 497
rect 1551 451 1563 485
rect 1597 451 1605 485
rect 1551 297 1605 451
<< ndiffc >>
rect 35 59 69 93
rect 129 123 163 157
rect 223 55 257 89
rect 317 55 351 89
rect 411 135 445 169
rect 505 55 539 89
rect 599 135 633 169
rect 693 55 727 89
rect 787 55 821 89
rect 885 135 919 169
rect 885 67 919 101
rect 989 55 1023 89
rect 1085 135 1119 169
rect 1085 67 1119 101
rect 1179 55 1213 89
rect 1273 135 1307 169
rect 1273 67 1307 101
rect 1367 55 1401 89
rect 1463 131 1497 165
rect 1559 55 1593 89
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 129 451 163 485
rect 223 443 257 477
rect 223 375 257 409
rect 317 455 351 489
rect 411 443 445 477
rect 411 375 445 409
rect 505 455 539 489
rect 599 443 633 477
rect 599 375 633 409
rect 693 455 727 489
rect 787 443 821 477
rect 787 375 821 409
rect 881 383 915 417
rect 975 455 1009 489
rect 1170 379 1204 413
rect 1266 305 1300 339
rect 1366 379 1400 413
rect 1563 451 1597 485
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 457 497 493 523
rect 551 497 587 523
rect 645 497 681 523
rect 739 497 775 523
rect 833 497 869 523
rect 927 497 963 523
rect 1021 497 1057 523
rect 1121 497 1157 523
rect 1217 497 1253 523
rect 1313 497 1349 523
rect 1413 497 1449 523
rect 1515 497 1551 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 457 282 493 297
rect 551 282 587 297
rect 645 282 681 297
rect 739 282 775 297
rect 833 282 869 297
rect 927 282 963 297
rect 1021 282 1057 297
rect 1121 282 1157 297
rect 1217 282 1253 297
rect 1313 282 1349 297
rect 1413 282 1449 297
rect 1515 282 1551 297
rect 79 259 119 282
rect 173 259 213 282
rect 267 259 307 282
rect 75 249 307 259
rect 75 215 91 249
rect 125 215 169 249
rect 203 215 247 249
rect 281 215 307 249
rect 75 205 307 215
rect 89 177 119 205
rect 183 177 213 205
rect 277 177 307 205
rect 361 259 401 282
rect 455 259 495 282
rect 549 259 589 282
rect 643 259 683 282
rect 737 265 777 282
rect 831 265 871 282
rect 925 265 965 282
rect 1019 265 1059 282
rect 1119 265 1159 282
rect 1215 265 1255 282
rect 1311 265 1351 282
rect 1411 265 1451 282
rect 1513 265 1553 282
rect 361 249 683 259
rect 361 215 377 249
rect 411 215 455 249
rect 489 215 533 249
rect 567 215 611 249
rect 645 215 683 249
rect 361 205 683 215
rect 361 177 391 205
rect 455 177 485 205
rect 549 177 579 205
rect 653 177 683 205
rect 725 249 789 265
rect 725 215 735 249
rect 769 215 789 249
rect 725 199 789 215
rect 831 249 1074 265
rect 831 215 845 249
rect 879 215 923 249
rect 957 215 1001 249
rect 1035 215 1074 249
rect 831 199 1074 215
rect 1116 249 1451 265
rect 1116 215 1126 249
rect 1160 215 1204 249
rect 1238 215 1282 249
rect 1316 215 1360 249
rect 1394 215 1451 249
rect 1116 199 1451 215
rect 1493 249 1558 265
rect 1493 215 1503 249
rect 1537 215 1558 249
rect 1493 199 1558 215
rect 747 177 777 199
rect 831 177 861 199
rect 948 177 978 199
rect 1044 177 1074 199
rect 1139 177 1169 199
rect 1233 177 1263 199
rect 1327 177 1357 199
rect 1421 177 1451 199
rect 1517 177 1547 199
rect 89 21 119 47
rect 183 21 213 47
rect 277 21 307 47
rect 361 21 391 47
rect 455 21 485 47
rect 549 21 579 47
rect 653 21 683 47
rect 747 21 777 47
rect 831 21 861 47
rect 948 21 978 47
rect 1044 21 1074 47
rect 1139 21 1169 47
rect 1233 21 1263 47
rect 1327 21 1357 47
rect 1421 21 1451 47
rect 1517 21 1547 47
<< polycont >>
rect 91 215 125 249
rect 169 215 203 249
rect 247 215 281 249
rect 377 215 411 249
rect 455 215 489 249
rect 533 215 567 249
rect 611 215 645 249
rect 735 215 769 249
rect 845 215 879 249
rect 923 215 957 249
rect 1001 215 1035 249
rect 1126 215 1160 249
rect 1204 215 1238 249
rect 1282 215 1316 249
rect 1360 215 1394 249
rect 1503 215 1537 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 19 477 69 493
rect 19 443 35 477
rect 103 485 179 527
rect 103 451 129 485
rect 163 451 179 485
rect 223 477 257 493
rect 19 417 69 443
rect 291 489 367 527
rect 291 455 317 489
rect 351 455 367 489
rect 411 477 445 493
rect 223 421 257 443
rect 479 489 555 527
rect 479 455 505 489
rect 539 455 555 489
rect 599 477 633 493
rect 411 421 445 443
rect 667 489 743 527
rect 667 455 693 489
rect 727 455 743 489
rect 787 489 1614 493
rect 787 477 975 489
rect 599 421 633 443
rect 821 455 975 477
rect 1009 485 1614 489
rect 1009 455 1563 485
rect 821 451 1563 455
rect 1597 451 1614 485
rect 787 421 821 443
rect 223 417 821 421
rect 19 409 821 417
rect 19 375 35 409
rect 69 375 223 409
rect 257 375 411 409
rect 445 375 599 409
rect 633 375 787 409
rect 19 359 821 375
rect 855 383 881 417
rect 915 383 1092 417
rect 855 357 1092 383
rect 1144 413 1632 417
rect 1144 379 1170 413
rect 1204 379 1366 413
rect 1400 379 1632 413
rect 1144 373 1632 379
rect 1026 339 1092 357
rect 20 289 795 325
rect 20 249 307 289
rect 20 215 91 249
rect 125 215 169 249
rect 203 215 247 249
rect 281 215 307 249
rect 20 207 307 215
rect 361 249 661 255
rect 361 215 377 249
rect 411 215 455 249
rect 489 215 533 249
rect 567 215 611 249
rect 645 215 661 249
rect 361 207 661 215
rect 719 249 795 289
rect 719 215 735 249
rect 769 215 795 249
rect 719 207 795 215
rect 829 289 857 323
rect 891 289 992 323
rect 1026 305 1266 339
rect 1300 305 1322 339
rect 1026 289 1322 305
rect 829 255 992 289
rect 1366 255 1410 339
rect 829 249 1061 255
rect 829 215 845 249
rect 879 215 923 249
rect 957 215 1001 249
rect 1035 215 1061 249
rect 829 207 1061 215
rect 1110 249 1410 255
rect 1110 215 1126 249
rect 1160 215 1204 249
rect 1238 215 1282 249
rect 1316 215 1360 249
rect 1394 215 1410 249
rect 1110 207 1410 215
rect 1460 323 1502 331
rect 1460 289 1468 323
rect 1536 299 1632 373
rect 1460 265 1502 289
rect 1460 249 1547 265
rect 1460 215 1503 249
rect 1537 215 1547 249
rect 1460 199 1547 215
rect 123 157 351 173
rect 123 123 129 157
rect 163 139 351 157
rect 163 123 165 139
rect 19 93 79 117
rect 123 106 165 123
rect 19 59 35 93
rect 69 59 79 93
rect 19 17 79 59
rect 200 89 257 105
rect 200 55 223 89
rect 200 17 257 55
rect 291 101 351 139
rect 385 169 1411 173
rect 385 135 411 169
rect 445 135 599 169
rect 633 139 885 169
rect 633 135 736 139
rect 855 135 885 139
rect 919 135 1085 169
rect 1119 135 1273 169
rect 1307 165 1411 169
rect 1581 165 1632 299
rect 1307 135 1463 165
rect 855 131 1463 135
rect 1497 131 1632 165
rect 855 125 1632 131
rect 855 123 1119 125
rect 291 89 743 101
rect 291 55 317 89
rect 351 55 505 89
rect 539 55 693 89
rect 727 55 743 89
rect 291 51 743 55
rect 787 89 821 105
rect 787 17 821 55
rect 855 101 929 123
rect 855 67 885 101
rect 919 67 929 101
rect 1085 101 1119 123
rect 855 51 929 67
rect 973 55 989 89
rect 1023 55 1039 89
rect 973 17 1039 55
rect 1273 123 1632 125
rect 1273 101 1307 123
rect 1085 51 1119 67
rect 1163 55 1179 89
rect 1213 55 1229 89
rect 1163 17 1229 55
rect 1273 51 1307 67
rect 1351 55 1367 89
rect 1401 55 1417 89
rect 1351 17 1417 55
rect 1533 55 1559 89
rect 1593 55 1614 89
rect 1533 17 1614 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 857 289 891 323
rect 1468 289 1502 323
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
<< metal1 >>
rect 0 561 1656 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 0 496 1656 527
rect 845 323 903 329
rect 845 289 857 323
rect 891 320 903 323
rect 1456 323 1514 329
rect 1456 320 1468 323
rect 891 292 1468 320
rect 891 289 903 292
rect 845 283 903 289
rect 1456 289 1468 292
rect 1502 289 1514 323
rect 1456 283 1514 289
rect 0 17 1656 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
rect 0 -48 1656 -17
<< labels >>
flabel corelocali s 214 289 248 323 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 397 221 431 255 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 1133 221 1167 255 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 1570 374 1570 374 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel metal1 s 857 289 891 323 0 FreeSans 400 0 0 0 B1
port 3 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 1656 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1127076
string GDS_START 1115802
<< end >>
