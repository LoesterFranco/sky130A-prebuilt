magic
tech sky130A
magscale 1 2
timestamp 1601050056
<< nwell >>
rect -38 332 1958 704
<< pwell >>
rect 0 0 1920 49
<< scpmos >>
rect 84 368 120 592
rect 174 368 210 592
rect 264 368 300 592
rect 354 368 390 592
rect 446 368 482 592
rect 536 368 572 592
rect 626 368 662 592
rect 716 368 752 592
rect 806 368 842 592
rect 896 368 932 592
rect 986 368 1022 592
rect 1076 368 1112 592
rect 1166 368 1202 592
rect 1256 368 1292 592
rect 1346 368 1382 592
rect 1436 368 1472 592
rect 1526 368 1562 592
rect 1616 368 1652 592
rect 1710 368 1746 592
rect 1800 368 1836 592
<< nmoslvt >>
rect 84 74 114 158
rect 170 74 200 158
rect 260 74 290 158
rect 346 74 376 158
rect 446 74 476 158
rect 532 74 562 158
rect 618 74 648 158
rect 704 74 734 158
rect 790 74 820 158
rect 876 74 906 158
rect 976 74 1006 158
rect 1062 74 1092 158
rect 1162 74 1192 158
rect 1248 74 1278 158
rect 1348 74 1378 158
rect 1434 74 1464 158
rect 1534 74 1564 158
rect 1620 74 1650 158
rect 1720 74 1750 158
rect 1806 74 1836 158
<< ndiff >>
rect 27 133 84 158
rect 27 99 39 133
rect 73 99 84 133
rect 27 74 84 99
rect 114 133 170 158
rect 114 99 125 133
rect 159 99 170 133
rect 114 74 170 99
rect 200 133 260 158
rect 200 99 211 133
rect 245 99 260 133
rect 200 74 260 99
rect 290 133 346 158
rect 290 99 301 133
rect 335 99 346 133
rect 290 74 346 99
rect 376 133 446 158
rect 376 99 387 133
rect 421 99 446 133
rect 376 74 446 99
rect 476 133 532 158
rect 476 99 487 133
rect 521 99 532 133
rect 476 74 532 99
rect 562 120 618 158
rect 562 86 573 120
rect 607 86 618 120
rect 562 74 618 86
rect 648 133 704 158
rect 648 99 659 133
rect 693 99 704 133
rect 648 74 704 99
rect 734 129 790 158
rect 734 95 745 129
rect 779 95 790 129
rect 734 74 790 95
rect 820 133 876 158
rect 820 99 831 133
rect 865 99 876 133
rect 820 74 876 99
rect 906 132 976 158
rect 906 98 917 132
rect 951 98 976 132
rect 906 74 976 98
rect 1006 133 1062 158
rect 1006 99 1017 133
rect 1051 99 1062 133
rect 1006 74 1062 99
rect 1092 120 1162 158
rect 1092 86 1103 120
rect 1137 86 1162 120
rect 1092 74 1162 86
rect 1192 133 1248 158
rect 1192 99 1203 133
rect 1237 99 1248 133
rect 1192 74 1248 99
rect 1278 120 1348 158
rect 1278 86 1289 120
rect 1323 86 1348 120
rect 1278 74 1348 86
rect 1378 133 1434 158
rect 1378 99 1389 133
rect 1423 99 1434 133
rect 1378 74 1434 99
rect 1464 120 1534 158
rect 1464 86 1475 120
rect 1509 86 1534 120
rect 1464 74 1534 86
rect 1564 133 1620 158
rect 1564 99 1575 133
rect 1609 99 1620 133
rect 1564 74 1620 99
rect 1650 120 1720 158
rect 1650 86 1661 120
rect 1695 86 1720 120
rect 1650 74 1720 86
rect 1750 133 1806 158
rect 1750 99 1761 133
rect 1795 99 1806 133
rect 1750 74 1806 99
rect 1836 133 1893 158
rect 1836 99 1847 133
rect 1881 99 1893 133
rect 1836 74 1893 99
<< pdiff >>
rect 28 580 84 592
rect 28 546 40 580
rect 74 546 84 580
rect 28 510 84 546
rect 28 476 40 510
rect 74 476 84 510
rect 28 440 84 476
rect 28 406 40 440
rect 74 406 84 440
rect 28 368 84 406
rect 120 580 174 592
rect 120 546 130 580
rect 164 546 174 580
rect 120 510 174 546
rect 120 476 130 510
rect 164 476 174 510
rect 120 440 174 476
rect 120 406 130 440
rect 164 406 174 440
rect 120 368 174 406
rect 210 580 264 592
rect 210 546 220 580
rect 254 546 264 580
rect 210 508 264 546
rect 210 474 220 508
rect 254 474 264 508
rect 210 368 264 474
rect 300 580 354 592
rect 300 546 310 580
rect 344 546 354 580
rect 300 510 354 546
rect 300 476 310 510
rect 344 476 354 510
rect 300 440 354 476
rect 300 406 310 440
rect 344 406 354 440
rect 300 368 354 406
rect 390 580 446 592
rect 390 546 400 580
rect 434 546 446 580
rect 390 508 446 546
rect 390 474 400 508
rect 434 474 446 508
rect 390 368 446 474
rect 482 580 536 592
rect 482 546 492 580
rect 526 546 536 580
rect 482 497 536 546
rect 482 463 492 497
rect 526 463 536 497
rect 482 414 536 463
rect 482 380 492 414
rect 526 380 536 414
rect 482 368 536 380
rect 572 580 626 592
rect 572 546 582 580
rect 616 546 626 580
rect 572 508 626 546
rect 572 474 582 508
rect 616 474 626 508
rect 572 440 626 474
rect 572 406 582 440
rect 616 406 626 440
rect 572 368 626 406
rect 662 580 716 592
rect 662 546 672 580
rect 706 546 716 580
rect 662 497 716 546
rect 662 463 672 497
rect 706 463 716 497
rect 662 414 716 463
rect 662 380 672 414
rect 706 380 716 414
rect 662 368 716 380
rect 752 580 806 592
rect 752 546 762 580
rect 796 546 806 580
rect 752 510 806 546
rect 752 476 762 510
rect 796 476 806 510
rect 752 440 806 476
rect 752 406 762 440
rect 796 406 806 440
rect 752 368 806 406
rect 842 580 896 592
rect 842 546 852 580
rect 886 546 896 580
rect 842 497 896 546
rect 842 463 852 497
rect 886 463 896 497
rect 842 414 896 463
rect 842 380 852 414
rect 886 380 896 414
rect 842 368 896 380
rect 932 580 986 592
rect 932 546 942 580
rect 976 546 986 580
rect 932 510 986 546
rect 932 476 942 510
rect 976 476 986 510
rect 932 440 986 476
rect 932 406 942 440
rect 976 406 986 440
rect 932 368 986 406
rect 1022 580 1076 592
rect 1022 546 1032 580
rect 1066 546 1076 580
rect 1022 497 1076 546
rect 1022 463 1032 497
rect 1066 463 1076 497
rect 1022 414 1076 463
rect 1022 380 1032 414
rect 1066 380 1076 414
rect 1022 368 1076 380
rect 1112 580 1166 592
rect 1112 546 1122 580
rect 1156 546 1166 580
rect 1112 510 1166 546
rect 1112 476 1122 510
rect 1156 476 1166 510
rect 1112 440 1166 476
rect 1112 406 1122 440
rect 1156 406 1166 440
rect 1112 368 1166 406
rect 1202 580 1256 592
rect 1202 546 1212 580
rect 1246 546 1256 580
rect 1202 497 1256 546
rect 1202 463 1212 497
rect 1246 463 1256 497
rect 1202 414 1256 463
rect 1202 380 1212 414
rect 1246 380 1256 414
rect 1202 368 1256 380
rect 1292 580 1346 592
rect 1292 546 1302 580
rect 1336 546 1346 580
rect 1292 510 1346 546
rect 1292 476 1302 510
rect 1336 476 1346 510
rect 1292 440 1346 476
rect 1292 406 1302 440
rect 1336 406 1346 440
rect 1292 368 1346 406
rect 1382 580 1436 592
rect 1382 546 1392 580
rect 1426 546 1436 580
rect 1382 497 1436 546
rect 1382 463 1392 497
rect 1426 463 1436 497
rect 1382 414 1436 463
rect 1382 380 1392 414
rect 1426 380 1436 414
rect 1382 368 1436 380
rect 1472 580 1526 592
rect 1472 546 1482 580
rect 1516 546 1526 580
rect 1472 510 1526 546
rect 1472 476 1482 510
rect 1516 476 1526 510
rect 1472 440 1526 476
rect 1472 406 1482 440
rect 1516 406 1526 440
rect 1472 368 1526 406
rect 1562 580 1616 592
rect 1562 546 1572 580
rect 1606 546 1616 580
rect 1562 497 1616 546
rect 1562 463 1572 497
rect 1606 463 1616 497
rect 1562 414 1616 463
rect 1562 380 1572 414
rect 1606 380 1616 414
rect 1562 368 1616 380
rect 1652 580 1710 592
rect 1652 546 1662 580
rect 1696 546 1710 580
rect 1652 510 1710 546
rect 1652 476 1662 510
rect 1696 476 1710 510
rect 1652 440 1710 476
rect 1652 406 1662 440
rect 1696 406 1710 440
rect 1652 368 1710 406
rect 1746 580 1800 592
rect 1746 546 1756 580
rect 1790 546 1800 580
rect 1746 497 1800 546
rect 1746 463 1756 497
rect 1790 463 1800 497
rect 1746 414 1800 463
rect 1746 380 1756 414
rect 1790 380 1800 414
rect 1746 368 1800 380
rect 1836 580 1892 592
rect 1836 546 1846 580
rect 1880 546 1892 580
rect 1836 510 1892 546
rect 1836 476 1846 510
rect 1880 476 1892 510
rect 1836 440 1892 476
rect 1836 406 1846 440
rect 1880 406 1892 440
rect 1836 368 1892 406
<< ndiffc >>
rect 39 99 73 133
rect 125 99 159 133
rect 211 99 245 133
rect 301 99 335 133
rect 387 99 421 133
rect 487 99 521 133
rect 573 86 607 120
rect 659 99 693 133
rect 745 95 779 129
rect 831 99 865 133
rect 917 98 951 132
rect 1017 99 1051 133
rect 1103 86 1137 120
rect 1203 99 1237 133
rect 1289 86 1323 120
rect 1389 99 1423 133
rect 1475 86 1509 120
rect 1575 99 1609 133
rect 1661 86 1695 120
rect 1761 99 1795 133
rect 1847 99 1881 133
<< pdiffc >>
rect 40 546 74 580
rect 40 476 74 510
rect 40 406 74 440
rect 130 546 164 580
rect 130 476 164 510
rect 130 406 164 440
rect 220 546 254 580
rect 220 474 254 508
rect 310 546 344 580
rect 310 476 344 510
rect 310 406 344 440
rect 400 546 434 580
rect 400 474 434 508
rect 492 546 526 580
rect 492 463 526 497
rect 492 380 526 414
rect 582 546 616 580
rect 582 474 616 508
rect 582 406 616 440
rect 672 546 706 580
rect 672 463 706 497
rect 672 380 706 414
rect 762 546 796 580
rect 762 476 796 510
rect 762 406 796 440
rect 852 546 886 580
rect 852 463 886 497
rect 852 380 886 414
rect 942 546 976 580
rect 942 476 976 510
rect 942 406 976 440
rect 1032 546 1066 580
rect 1032 463 1066 497
rect 1032 380 1066 414
rect 1122 546 1156 580
rect 1122 476 1156 510
rect 1122 406 1156 440
rect 1212 546 1246 580
rect 1212 463 1246 497
rect 1212 380 1246 414
rect 1302 546 1336 580
rect 1302 476 1336 510
rect 1302 406 1336 440
rect 1392 546 1426 580
rect 1392 463 1426 497
rect 1392 380 1426 414
rect 1482 546 1516 580
rect 1482 476 1516 510
rect 1482 406 1516 440
rect 1572 546 1606 580
rect 1572 463 1606 497
rect 1572 380 1606 414
rect 1662 546 1696 580
rect 1662 476 1696 510
rect 1662 406 1696 440
rect 1756 546 1790 580
rect 1756 463 1790 497
rect 1756 380 1790 414
rect 1846 546 1880 580
rect 1846 476 1880 510
rect 1846 406 1880 440
<< poly >>
rect 84 592 120 618
rect 174 592 210 618
rect 264 592 300 618
rect 354 592 390 618
rect 446 592 482 618
rect 536 592 572 618
rect 626 592 662 618
rect 716 592 752 618
rect 806 592 842 618
rect 896 592 932 618
rect 986 592 1022 618
rect 1076 592 1112 618
rect 1166 592 1202 618
rect 1256 592 1292 618
rect 1346 592 1382 618
rect 1436 592 1472 618
rect 1526 592 1562 618
rect 1616 592 1652 618
rect 1710 592 1746 618
rect 1800 592 1836 618
rect 84 336 120 368
rect 174 336 210 368
rect 264 336 300 368
rect 354 336 390 368
rect 84 320 390 336
rect 84 286 100 320
rect 134 286 168 320
rect 202 286 236 320
rect 270 286 304 320
rect 338 286 390 320
rect 84 270 390 286
rect 446 304 482 368
rect 536 304 572 368
rect 626 304 662 368
rect 716 304 752 368
rect 806 304 842 368
rect 896 304 932 368
rect 986 304 1022 368
rect 1076 304 1112 368
rect 1166 304 1202 368
rect 1256 304 1292 368
rect 1346 304 1382 368
rect 1436 304 1472 368
rect 1526 304 1562 368
rect 1616 304 1652 368
rect 1710 304 1746 368
rect 1800 304 1836 368
rect 446 288 1836 304
rect 84 158 114 270
rect 170 158 200 270
rect 260 158 290 270
rect 346 158 376 270
rect 446 254 578 288
rect 612 254 750 288
rect 784 254 918 288
rect 952 254 1101 288
rect 1135 254 1289 288
rect 1323 254 1475 288
rect 1509 254 1661 288
rect 1695 254 1836 288
rect 446 238 1836 254
rect 446 158 476 238
rect 532 158 562 238
rect 618 158 648 238
rect 704 158 734 238
rect 790 158 820 238
rect 876 158 906 238
rect 976 158 1006 238
rect 1062 158 1092 238
rect 1162 158 1192 238
rect 1248 158 1278 238
rect 1348 158 1378 238
rect 1434 158 1464 238
rect 1534 158 1564 238
rect 1620 158 1650 238
rect 1720 158 1750 238
rect 1806 158 1836 238
rect 84 48 114 74
rect 170 48 200 74
rect 260 48 290 74
rect 346 48 376 74
rect 446 48 476 74
rect 532 48 562 74
rect 618 48 648 74
rect 704 48 734 74
rect 790 48 820 74
rect 876 48 906 74
rect 976 48 1006 74
rect 1062 48 1092 74
rect 1162 48 1192 74
rect 1248 48 1278 74
rect 1348 48 1378 74
rect 1434 48 1464 74
rect 1534 48 1564 74
rect 1620 48 1650 74
rect 1720 48 1750 74
rect 1806 48 1836 74
<< polycont >>
rect 100 286 134 320
rect 168 286 202 320
rect 236 286 270 320
rect 304 286 338 320
rect 578 254 612 288
rect 750 254 784 288
rect 918 254 952 288
rect 1101 254 1135 288
rect 1289 254 1323 288
rect 1475 254 1509 288
rect 1661 254 1695 288
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 24 580 74 649
rect 24 546 40 580
rect 24 510 74 546
rect 24 476 40 510
rect 24 440 74 476
rect 24 406 40 440
rect 24 390 74 406
rect 114 580 180 596
rect 114 546 130 580
rect 164 546 180 580
rect 114 510 180 546
rect 114 476 130 510
rect 164 476 180 510
rect 114 440 180 476
rect 220 580 254 649
rect 220 508 254 546
rect 220 458 254 474
rect 294 580 360 596
rect 294 546 310 580
rect 344 546 360 580
rect 294 510 360 546
rect 294 476 310 510
rect 344 476 360 510
rect 114 406 130 440
rect 164 424 180 440
rect 294 440 360 476
rect 400 580 450 649
rect 434 546 450 580
rect 400 508 450 546
rect 434 474 450 508
rect 400 458 450 474
rect 486 580 532 596
rect 486 546 492 580
rect 526 546 532 580
rect 486 497 532 546
rect 486 463 492 497
rect 526 463 532 497
rect 294 424 310 440
rect 164 406 310 424
rect 344 424 360 440
rect 486 424 532 463
rect 344 406 427 424
rect 114 390 427 406
rect 25 320 359 356
rect 25 286 100 320
rect 134 286 168 320
rect 202 286 236 320
rect 270 286 304 320
rect 338 286 359 320
rect 25 270 359 286
rect 393 282 427 390
rect 478 380 492 424
rect 526 380 532 424
rect 566 580 632 649
rect 566 546 582 580
rect 616 546 632 580
rect 566 508 632 546
rect 566 474 582 508
rect 616 474 632 508
rect 566 440 632 474
rect 566 406 582 440
rect 616 406 632 440
rect 668 580 709 596
rect 668 546 672 580
rect 706 546 709 580
rect 668 497 709 546
rect 668 463 672 497
rect 706 463 709 497
rect 668 424 709 463
rect 393 276 442 282
rect 393 242 402 276
rect 436 242 442 276
rect 393 236 442 242
rect 393 230 427 236
rect 109 196 427 230
rect 23 133 73 162
rect 23 99 39 133
rect 23 17 73 99
rect 109 133 159 196
rect 109 99 125 133
rect 109 70 159 99
rect 195 133 245 162
rect 195 99 211 133
rect 195 17 245 99
rect 285 133 335 196
rect 285 99 301 133
rect 285 70 335 99
rect 371 133 437 162
rect 371 99 387 133
rect 421 99 437 133
rect 371 17 437 99
rect 478 133 532 380
rect 668 380 672 424
rect 706 380 709 424
rect 746 580 812 649
rect 746 546 762 580
rect 796 546 812 580
rect 746 510 812 546
rect 746 476 762 510
rect 796 476 812 510
rect 746 440 812 476
rect 746 406 762 440
rect 796 406 812 440
rect 846 580 886 596
rect 846 546 852 580
rect 846 497 886 546
rect 846 463 852 497
rect 846 424 886 463
rect 668 372 709 380
rect 846 390 849 424
rect 883 414 886 424
rect 926 580 992 649
rect 926 546 942 580
rect 976 546 992 580
rect 926 510 992 546
rect 926 476 942 510
rect 976 476 992 510
rect 926 440 992 476
rect 926 406 942 440
rect 976 406 992 440
rect 1028 580 1070 596
rect 1028 546 1032 580
rect 1066 546 1070 580
rect 1028 497 1070 546
rect 1028 463 1032 497
rect 1066 463 1070 497
rect 1028 424 1070 463
rect 846 380 852 390
rect 846 372 886 380
rect 1028 380 1032 424
rect 1066 380 1070 424
rect 1106 580 1172 649
rect 1106 546 1122 580
rect 1156 546 1172 580
rect 1106 510 1172 546
rect 1106 476 1122 510
rect 1156 476 1172 510
rect 1106 440 1172 476
rect 1106 406 1122 440
rect 1156 406 1172 440
rect 1208 580 1249 596
rect 1208 546 1212 580
rect 1246 546 1249 580
rect 1208 497 1249 546
rect 1208 463 1212 497
rect 1246 463 1249 497
rect 1208 424 1249 463
rect 1028 372 1070 380
rect 1208 380 1212 424
rect 1246 380 1249 424
rect 1286 580 1352 649
rect 1286 546 1302 580
rect 1336 546 1352 580
rect 1286 510 1352 546
rect 1286 476 1302 510
rect 1336 476 1352 510
rect 1286 440 1352 476
rect 1286 406 1302 440
rect 1336 406 1352 440
rect 1389 580 1430 596
rect 1389 546 1392 580
rect 1426 546 1430 580
rect 1389 497 1430 546
rect 1389 463 1392 497
rect 1426 463 1430 497
rect 1389 424 1430 463
rect 1208 372 1249 380
rect 1389 380 1392 424
rect 1426 380 1430 424
rect 1466 580 1532 649
rect 1466 546 1482 580
rect 1516 546 1532 580
rect 1466 510 1532 546
rect 1466 476 1482 510
rect 1516 476 1532 510
rect 1466 440 1532 476
rect 1466 406 1482 440
rect 1516 406 1532 440
rect 1568 580 1610 596
rect 1568 546 1572 580
rect 1606 546 1610 580
rect 1568 497 1610 546
rect 1568 463 1572 497
rect 1606 463 1610 497
rect 1568 424 1610 463
rect 1389 372 1430 380
rect 1568 380 1572 424
rect 1606 380 1610 424
rect 1646 580 1712 649
rect 1646 546 1662 580
rect 1696 546 1712 580
rect 1646 510 1712 546
rect 1646 476 1662 510
rect 1696 476 1712 510
rect 1646 440 1712 476
rect 1646 406 1662 440
rect 1696 406 1712 440
rect 1750 580 1794 596
rect 1750 546 1756 580
rect 1790 546 1794 580
rect 1750 497 1794 546
rect 1750 463 1756 497
rect 1790 463 1794 497
rect 1750 424 1794 463
rect 1568 372 1610 380
rect 1750 380 1756 424
rect 1790 380 1794 424
rect 1830 580 1896 649
rect 1830 546 1846 580
rect 1880 546 1896 580
rect 1830 510 1896 546
rect 1830 476 1846 510
rect 1880 476 1896 510
rect 1830 440 1896 476
rect 1830 406 1846 440
rect 1880 406 1896 440
rect 1750 372 1794 380
rect 655 338 709 372
rect 834 338 886 372
rect 1005 338 1070 372
rect 1187 338 1249 372
rect 1373 338 1430 372
rect 1559 338 1610 372
rect 1745 366 1794 372
rect 567 288 621 304
rect 567 242 578 288
rect 612 242 621 288
rect 567 238 621 242
rect 478 99 487 133
rect 521 99 532 133
rect 478 70 532 99
rect 573 120 607 136
rect 573 17 607 86
rect 655 133 700 338
rect 734 288 800 304
rect 734 242 750 288
rect 784 242 800 288
rect 734 238 800 242
rect 834 149 868 338
rect 902 288 968 304
rect 902 242 918 288
rect 952 242 968 288
rect 902 238 968 242
rect 655 99 659 133
rect 693 99 700 133
rect 655 70 700 99
rect 734 129 779 145
rect 734 95 745 129
rect 734 17 779 95
rect 815 133 868 149
rect 815 99 831 133
rect 865 99 868 133
rect 815 70 868 99
rect 902 132 967 148
rect 902 98 917 132
rect 951 98 967 132
rect 902 17 967 98
rect 1005 133 1051 338
rect 1085 288 1151 304
rect 1085 242 1101 288
rect 1135 242 1151 288
rect 1085 238 1151 242
rect 1005 99 1017 133
rect 1005 70 1051 99
rect 1087 120 1153 136
rect 1087 86 1103 120
rect 1137 86 1153 120
rect 1087 17 1153 86
rect 1187 133 1237 338
rect 1273 288 1339 304
rect 1273 242 1289 288
rect 1323 242 1339 288
rect 1273 238 1339 242
rect 1187 99 1203 133
rect 1187 70 1237 99
rect 1273 120 1339 136
rect 1273 86 1289 120
rect 1323 86 1339 120
rect 1273 17 1339 86
rect 1373 133 1423 338
rect 1459 288 1525 304
rect 1459 242 1475 288
rect 1509 242 1525 288
rect 1459 238 1525 242
rect 1373 99 1389 133
rect 1373 70 1423 99
rect 1459 120 1525 136
rect 1459 86 1475 120
rect 1509 86 1525 120
rect 1459 17 1525 86
rect 1559 133 1609 338
rect 1645 288 1711 304
rect 1645 242 1661 288
rect 1695 242 1711 288
rect 1645 238 1711 242
rect 1559 99 1575 133
rect 1559 70 1609 99
rect 1645 120 1711 136
rect 1645 86 1661 120
rect 1695 86 1711 120
rect 1645 17 1711 86
rect 1745 133 1795 366
rect 1745 99 1761 133
rect 1745 70 1795 99
rect 1831 133 1897 149
rect 1831 99 1847 133
rect 1881 99 1897 133
rect 1831 17 1897 99
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 492 414 526 424
rect 492 390 526 414
rect 402 242 436 276
rect 672 414 706 424
rect 672 390 706 414
rect 849 414 883 424
rect 849 390 852 414
rect 852 390 883 414
rect 1032 414 1066 424
rect 1032 390 1066 414
rect 1212 414 1246 424
rect 1212 390 1246 414
rect 1392 414 1426 424
rect 1392 390 1426 414
rect 1572 414 1606 424
rect 1572 390 1606 414
rect 1756 414 1790 424
rect 1756 390 1790 414
rect 578 254 612 276
rect 578 242 612 254
rect 750 254 784 276
rect 750 242 784 254
rect 918 254 952 276
rect 918 242 952 254
rect 1101 254 1135 276
rect 1101 242 1135 254
rect 1289 254 1323 276
rect 1289 242 1323 254
rect 1475 254 1509 276
rect 1475 242 1509 254
rect 1661 254 1695 276
rect 1661 242 1695 254
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
<< metal1 >>
rect 0 683 1920 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 0 617 1920 649
rect 478 424 1818 430
rect 478 390 492 424
rect 526 390 672 424
rect 706 390 849 424
rect 883 390 1032 424
rect 1066 390 1212 424
rect 1246 390 1392 424
rect 1426 390 1572 424
rect 1606 390 1756 424
rect 1790 390 1818 424
rect 478 384 1818 390
rect 388 276 1728 282
rect 388 242 402 276
rect 436 242 578 276
rect 612 242 750 276
rect 784 242 918 276
rect 952 242 1101 276
rect 1135 242 1289 276
rect 1323 242 1475 276
rect 1509 242 1661 276
rect 1695 242 1728 276
rect 388 236 1728 242
rect 0 17 1920 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
rect 0 -49 1920 -17
<< labels >>
flabel pwell s 0 0 1920 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew
flabel nbase s 0 617 1920 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew
rlabel comment s 0 0 0 0 4 clkbuf_16
flabel metal1 s 0 617 1920 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew
flabel metal1 s 0 0 1920 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew
flabel metal1 s 478 384 1818 430 0 FreeSans 400 0 0 0 X
port 6 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 1920 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3394684
string GDS_START 3379398
<< end >>
