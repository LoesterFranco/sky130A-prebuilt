magic
tech sky130A
magscale 1 2
timestamp 1601050058
<< locali >>
rect 112 391 162 493
rect 468 391 518 425
rect 820 391 870 425
rect 112 357 870 391
rect 112 289 170 357
rect 17 215 87 255
rect 121 173 170 289
rect 204 289 652 323
rect 204 215 407 289
rect 441 215 552 255
rect 586 215 652 289
rect 686 289 963 323
rect 686 215 752 289
rect 929 255 963 289
rect 796 215 895 255
rect 929 215 1087 255
rect 104 129 170 173
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 28 291 78 527
rect 196 425 350 527
rect 384 459 602 493
rect 384 425 434 459
rect 552 425 602 459
rect 636 425 702 527
rect 736 459 954 493
rect 736 425 786 459
rect 904 357 954 459
rect 20 95 70 179
rect 997 291 1038 527
rect 204 129 610 181
rect 644 147 1046 181
rect 204 95 254 129
rect 644 95 710 147
rect 812 145 1046 147
rect 20 51 254 95
rect 292 51 710 95
rect 744 17 778 111
rect 812 51 878 145
rect 912 17 946 111
rect 980 51 1046 145
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
rlabel locali s 929 255 963 289 6 A1
port 1 nsew signal input
rlabel locali s 929 215 1087 255 6 A1
port 1 nsew signal input
rlabel locali s 686 289 963 323 6 A1
port 1 nsew signal input
rlabel locali s 686 215 752 289 6 A1
port 1 nsew signal input
rlabel locali s 796 215 895 255 6 A2
port 2 nsew signal input
rlabel locali s 586 215 652 289 6 B1
port 3 nsew signal input
rlabel locali s 204 289 652 323 6 B1
port 3 nsew signal input
rlabel locali s 204 215 407 289 6 B1
port 3 nsew signal input
rlabel locali s 441 215 552 255 6 B2
port 4 nsew signal input
rlabel locali s 17 215 87 255 6 C1
port 5 nsew signal input
rlabel locali s 820 391 870 425 6 Y
port 6 nsew signal output
rlabel locali s 468 391 518 425 6 Y
port 6 nsew signal output
rlabel locali s 121 173 170 289 6 Y
port 6 nsew signal output
rlabel locali s 112 391 162 493 6 Y
port 6 nsew signal output
rlabel locali s 112 357 870 391 6 Y
port 6 nsew signal output
rlabel locali s 112 289 170 357 6 Y
port 6 nsew signal output
rlabel locali s 104 129 170 173 6 Y
port 6 nsew signal output
rlabel metal1 s 0 -48 1104 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1104 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1104 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1453250
string GDS_START 1444584
<< end >>
