magic
tech sky130A
magscale 1 2
timestamp 1599588244
<< locali >>
rect 23 364 89 596
rect 23 70 73 364
rect 217 289 287 356
rect 343 289 455 356
rect 489 260 555 356
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 123 458 236 649
rect 272 424 338 559
rect 139 390 338 424
rect 487 390 553 649
rect 139 310 173 390
rect 107 255 173 310
rect 107 221 279 255
rect 109 17 175 187
rect 229 70 279 221
rect 315 192 553 226
rect 315 70 365 192
rect 401 17 467 158
rect 503 70 553 192
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
rlabel locali s 489 260 555 356 6 A1
port 1 nsew signal input
rlabel locali s 343 289 455 356 6 A2
port 2 nsew signal input
rlabel locali s 217 289 287 356 6 B1
port 3 nsew signal input
rlabel locali s 23 364 89 596 6 X
port 4 nsew signal output
rlabel locali s 23 70 73 364 6 X
port 4 nsew signal output
rlabel metal1 s 0 -49 576 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 6 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 617 576 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 576 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1040682
string GDS_START 1034210
<< end >>
