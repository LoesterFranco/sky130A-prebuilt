magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 17 191 66 333
rect 178 191 259 391
rect 1394 331 1444 493
rect 1394 297 1535 331
rect 1498 177 1535 297
rect 1394 143 1535 177
rect 1394 89 1434 143
rect 1368 51 1434 89
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 17 367 69 527
rect 103 425 256 493
rect 322 425 460 493
rect 103 157 144 425
rect 293 241 392 391
rect 426 275 460 425
rect 504 415 621 527
rect 665 417 709 493
rect 777 451 1151 527
rect 1195 417 1229 493
rect 1279 451 1345 527
rect 665 383 1151 417
rect 665 381 709 383
rect 494 327 709 381
rect 494 315 533 327
rect 426 241 641 275
rect 17 123 259 157
rect 293 141 360 241
rect 394 141 461 207
rect 495 199 641 241
rect 17 51 69 123
rect 103 17 179 89
rect 223 51 259 123
rect 495 107 529 199
rect 293 51 529 107
rect 582 17 616 165
rect 675 51 709 327
rect 747 315 829 349
rect 747 187 781 315
rect 873 299 1043 349
rect 873 255 934 299
rect 815 221 934 255
rect 747 153 832 187
rect 876 157 934 221
rect 993 255 1037 265
rect 993 221 1002 255
rect 1036 221 1037 255
rect 993 199 1037 221
rect 1081 199 1151 383
rect 1195 299 1350 417
rect 1195 255 1281 265
rect 1195 221 1200 255
rect 1234 221 1281 255
rect 1195 199 1281 221
rect 1316 263 1350 299
rect 1488 365 1538 527
rect 1316 211 1454 263
rect 1316 157 1350 211
rect 747 51 813 153
rect 876 123 1017 157
rect 857 17 923 89
rect 967 51 1017 123
rect 1101 123 1350 157
rect 1101 51 1135 123
rect 1267 17 1334 89
rect 1478 17 1512 109
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1002 221 1036 255
rect 1200 221 1234 255
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
<< metal1 >>
rect 0 561 1564 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 0 496 1564 527
rect 990 255 1048 261
rect 990 221 1002 255
rect 1036 252 1048 255
rect 1188 255 1246 261
rect 1188 252 1200 255
rect 1036 224 1200 252
rect 1036 221 1048 224
rect 990 215 1048 221
rect 1188 221 1200 224
rect 1234 221 1246 255
rect 1188 215 1246 221
rect 0 17 1564 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
rect 0 -48 1564 -17
<< obsm1 >>
rect 313 320 371 329
rect 888 320 946 329
rect 313 292 946 320
rect 313 283 371 292
rect 888 283 946 292
rect 415 184 473 193
rect 786 184 844 193
rect 415 156 844 184
rect 415 147 473 156
rect 786 147 844 156
<< labels >>
rlabel metal1 s 1188 252 1246 261 6 CLK
port 1 nsew signal input
rlabel metal1 s 1188 215 1246 224 6 CLK
port 1 nsew signal input
rlabel metal1 s 990 252 1048 261 6 CLK
port 1 nsew signal input
rlabel metal1 s 990 224 1246 252 6 CLK
port 1 nsew signal input
rlabel metal1 s 990 215 1048 224 6 CLK
port 1 nsew signal input
rlabel locali s 178 191 259 391 6 GATE
port 2 nsew signal input
rlabel locali s 1498 177 1535 297 6 GCLK
port 3 nsew signal output
rlabel locali s 1394 331 1444 493 6 GCLK
port 3 nsew signal output
rlabel locali s 1394 297 1535 331 6 GCLK
port 3 nsew signal output
rlabel locali s 1394 143 1535 177 6 GCLK
port 3 nsew signal output
rlabel locali s 1394 89 1434 143 6 GCLK
port 3 nsew signal output
rlabel locali s 1368 51 1434 89 6 GCLK
port 3 nsew signal output
rlabel locali s 17 191 66 333 6 SCE
port 4 nsew signal input
rlabel metal1 s 0 -48 1564 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 1564 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1564 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 393366
string GDS_START 381334
<< end >>
