magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 1190 704
<< pwell >>
rect 0 0 1152 49
<< scnmos >>
rect 88 136 118 264
rect 477 74 507 222
rect 577 74 607 222
rect 663 74 693 222
rect 765 74 795 222
rect 856 74 886 222
rect 952 74 982 222
rect 1038 74 1068 222
<< pmoshvt >>
rect 85 392 115 592
rect 187 392 217 592
rect 277 392 307 592
rect 379 392 409 592
rect 474 392 504 592
rect 564 392 594 592
rect 666 392 696 592
rect 768 368 798 592
rect 858 368 888 592
rect 948 368 978 592
rect 1038 368 1068 592
<< ndiff >>
rect 31 232 88 264
rect 31 198 43 232
rect 77 198 88 232
rect 31 136 88 198
rect 118 136 278 264
rect 193 112 278 136
rect 193 78 218 112
rect 252 78 278 112
rect 193 66 278 78
rect 421 196 477 222
rect 421 162 432 196
rect 466 162 477 196
rect 421 120 477 162
rect 421 86 432 120
rect 466 86 477 120
rect 421 74 477 86
rect 507 124 577 222
rect 507 90 532 124
rect 566 90 577 124
rect 507 74 577 90
rect 607 196 663 222
rect 607 162 618 196
rect 652 162 663 196
rect 607 120 663 162
rect 607 86 618 120
rect 652 86 663 120
rect 607 74 663 86
rect 693 120 765 222
rect 693 86 719 120
rect 753 86 765 120
rect 693 74 765 86
rect 795 210 856 222
rect 795 176 811 210
rect 845 176 856 210
rect 795 120 856 176
rect 795 86 811 120
rect 845 86 856 120
rect 795 74 856 86
rect 886 136 952 222
rect 886 102 897 136
rect 931 102 952 136
rect 886 74 952 102
rect 982 210 1038 222
rect 982 176 993 210
rect 1027 176 1038 210
rect 982 120 1038 176
rect 982 86 993 120
rect 1027 86 1038 120
rect 982 74 1038 86
rect 1068 142 1125 222
rect 1068 108 1079 142
rect 1113 108 1125 142
rect 1068 74 1125 108
<< pdiff >>
rect 27 580 85 592
rect 27 546 38 580
rect 72 546 85 580
rect 27 509 85 546
rect 27 475 38 509
rect 72 475 85 509
rect 27 438 85 475
rect 27 404 38 438
rect 72 404 85 438
rect 27 392 85 404
rect 115 580 187 592
rect 115 546 128 580
rect 162 546 187 580
rect 115 509 187 546
rect 115 475 128 509
rect 162 475 187 509
rect 115 438 187 475
rect 115 404 128 438
rect 162 404 187 438
rect 115 392 187 404
rect 217 580 277 592
rect 217 546 230 580
rect 264 546 277 580
rect 217 512 277 546
rect 217 478 230 512
rect 264 478 277 512
rect 217 444 277 478
rect 217 410 230 444
rect 264 410 277 444
rect 217 392 277 410
rect 307 577 379 592
rect 307 543 332 577
rect 366 543 379 577
rect 307 392 379 543
rect 409 438 474 592
rect 409 404 424 438
rect 458 404 474 438
rect 409 392 474 404
rect 504 577 564 592
rect 504 543 517 577
rect 551 543 564 577
rect 504 392 564 543
rect 594 580 666 592
rect 594 546 617 580
rect 651 546 666 580
rect 594 512 666 546
rect 594 478 617 512
rect 651 478 666 512
rect 594 392 666 478
rect 696 580 768 592
rect 696 546 717 580
rect 751 546 768 580
rect 696 512 768 546
rect 696 478 717 512
rect 751 478 768 512
rect 696 392 768 478
rect 715 368 768 392
rect 798 580 858 592
rect 798 546 811 580
rect 845 546 858 580
rect 798 497 858 546
rect 798 463 811 497
rect 845 463 858 497
rect 798 414 858 463
rect 798 380 811 414
rect 845 380 858 414
rect 798 368 858 380
rect 888 580 948 592
rect 888 546 901 580
rect 935 546 948 580
rect 888 478 948 546
rect 888 444 901 478
rect 935 444 948 478
rect 888 368 948 444
rect 978 580 1038 592
rect 978 546 991 580
rect 1025 546 1038 580
rect 978 497 1038 546
rect 978 463 991 497
rect 1025 463 1038 497
rect 978 414 1038 463
rect 978 380 991 414
rect 1025 380 1038 414
rect 978 368 1038 380
rect 1068 580 1125 592
rect 1068 546 1081 580
rect 1115 546 1125 580
rect 1068 478 1125 546
rect 1068 444 1081 478
rect 1115 444 1125 478
rect 1068 368 1125 444
<< ndiffc >>
rect 43 198 77 232
rect 218 78 252 112
rect 432 162 466 196
rect 432 86 466 120
rect 532 90 566 124
rect 618 162 652 196
rect 618 86 652 120
rect 719 86 753 120
rect 811 176 845 210
rect 811 86 845 120
rect 897 102 931 136
rect 993 176 1027 210
rect 993 86 1027 120
rect 1079 108 1113 142
<< pdiffc >>
rect 38 546 72 580
rect 38 475 72 509
rect 38 404 72 438
rect 128 546 162 580
rect 128 475 162 509
rect 128 404 162 438
rect 230 546 264 580
rect 230 478 264 512
rect 230 410 264 444
rect 332 543 366 577
rect 424 404 458 438
rect 517 543 551 577
rect 617 546 651 580
rect 617 478 651 512
rect 717 546 751 580
rect 717 478 751 512
rect 811 546 845 580
rect 811 463 845 497
rect 811 380 845 414
rect 901 546 935 580
rect 901 444 935 478
rect 991 546 1025 580
rect 991 463 1025 497
rect 991 380 1025 414
rect 1081 546 1115 580
rect 1081 444 1115 478
<< poly >>
rect 85 592 115 618
rect 187 592 217 618
rect 277 592 307 618
rect 379 592 409 618
rect 474 592 504 618
rect 564 592 594 618
rect 666 592 696 618
rect 768 592 798 618
rect 858 592 888 618
rect 948 592 978 618
rect 1038 592 1068 618
rect 85 377 115 392
rect 187 377 217 392
rect 277 377 307 392
rect 379 377 409 392
rect 474 377 504 392
rect 564 377 594 392
rect 666 377 696 392
rect 82 279 118 377
rect 184 352 220 377
rect 274 360 310 377
rect 160 336 226 352
rect 160 302 176 336
rect 210 302 226 336
rect 160 286 226 302
rect 268 344 334 360
rect 268 310 284 344
rect 318 310 334 344
rect 268 294 334 310
rect 88 264 118 279
rect 376 267 412 377
rect 471 267 507 377
rect 561 360 597 377
rect 549 344 615 360
rect 549 310 565 344
rect 599 310 615 344
rect 663 310 699 377
rect 768 353 798 368
rect 858 353 888 368
rect 948 353 978 368
rect 1038 353 1068 368
rect 765 326 801 353
rect 855 326 891 353
rect 945 326 981 353
rect 1035 326 1071 353
rect 765 310 1071 326
rect 549 294 615 310
rect 657 294 723 310
rect 376 237 507 267
rect 376 196 406 237
rect 477 222 507 237
rect 577 222 607 294
rect 657 260 673 294
rect 707 260 723 294
rect 657 244 723 260
rect 765 276 781 310
rect 815 276 849 310
rect 883 276 917 310
rect 951 276 985 310
rect 1019 276 1071 310
rect 765 260 1071 276
rect 663 222 693 244
rect 765 222 795 260
rect 856 222 886 260
rect 952 222 982 260
rect 1038 222 1068 260
rect 88 114 118 136
rect 21 98 155 114
rect 21 64 37 98
rect 71 64 105 98
rect 139 64 155 98
rect 316 180 406 196
rect 316 146 332 180
rect 366 146 406 180
rect 316 112 406 146
rect 316 78 332 112
rect 366 78 406 112
rect 21 48 155 64
rect 316 62 406 78
rect 477 48 507 74
rect 577 48 607 74
rect 663 48 693 74
rect 765 48 795 74
rect 856 48 886 74
rect 952 48 982 74
rect 1038 48 1068 74
<< polycont >>
rect 176 302 210 336
rect 284 310 318 344
rect 565 310 599 344
rect 673 260 707 294
rect 781 276 815 310
rect 849 276 883 310
rect 917 276 951 310
rect 985 276 1019 310
rect 37 64 71 98
rect 105 64 139 98
rect 332 146 366 180
rect 332 78 366 112
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 22 580 72 596
rect 22 546 38 580
rect 22 509 72 546
rect 22 475 38 509
rect 22 438 72 475
rect 22 404 38 438
rect 22 268 72 404
rect 112 580 178 649
rect 112 546 128 580
rect 162 546 178 580
rect 112 509 178 546
rect 112 475 128 509
rect 162 475 178 509
rect 112 438 178 475
rect 112 404 128 438
rect 162 404 178 438
rect 112 388 178 404
rect 214 580 280 596
rect 214 546 230 580
rect 264 546 280 580
rect 214 512 280 546
rect 316 577 567 596
rect 316 543 332 577
rect 366 543 517 577
rect 551 543 567 577
rect 316 540 567 543
rect 601 580 667 596
rect 601 546 617 580
rect 651 546 667 580
rect 214 478 230 512
rect 264 506 280 512
rect 601 512 667 546
rect 601 506 617 512
rect 264 478 617 506
rect 651 478 667 512
rect 214 472 667 478
rect 214 444 280 472
rect 601 462 667 472
rect 701 580 767 649
rect 701 546 717 580
rect 751 546 767 580
rect 701 512 767 546
rect 701 478 717 512
rect 751 478 767 512
rect 701 462 767 478
rect 811 580 845 596
rect 811 497 845 546
rect 214 410 230 444
rect 264 410 280 444
rect 214 394 280 410
rect 406 404 424 438
rect 458 428 477 438
rect 458 404 777 428
rect 406 394 777 404
rect 160 336 226 352
rect 160 302 176 336
rect 210 302 226 336
rect 22 232 93 268
rect 22 198 43 232
rect 77 198 93 232
rect 160 264 226 302
rect 268 344 615 360
rect 268 310 284 344
rect 318 310 565 344
rect 599 310 615 344
rect 743 326 777 394
rect 811 414 845 463
rect 885 580 935 649
rect 885 546 901 580
rect 885 478 935 546
rect 885 444 901 478
rect 885 428 935 444
rect 975 580 1041 596
rect 975 546 991 580
rect 1025 546 1041 580
rect 975 497 1041 546
rect 975 463 991 497
rect 1025 463 1041 497
rect 975 414 1041 463
rect 1081 580 1131 649
rect 1115 546 1131 580
rect 1081 478 1131 546
rect 1115 444 1131 478
rect 1081 428 1131 444
rect 975 394 991 414
rect 845 380 991 394
rect 1025 394 1041 414
rect 1025 380 1127 394
rect 811 360 1127 380
rect 743 310 1035 326
rect 268 298 334 310
rect 657 294 709 310
rect 657 276 673 294
rect 601 264 673 276
rect 160 260 673 264
rect 707 260 709 294
rect 160 230 709 260
rect 743 276 781 310
rect 815 276 849 310
rect 883 276 917 310
rect 951 276 985 310
rect 1019 276 1035 310
rect 743 260 1035 276
rect 22 196 93 198
rect 743 196 777 260
rect 1081 226 1127 360
rect 22 180 382 196
rect 22 162 332 180
rect 316 146 332 162
rect 366 146 382 180
rect 21 98 155 128
rect 21 64 37 98
rect 71 64 105 98
rect 139 64 155 98
rect 21 51 155 64
rect 189 112 282 128
rect 189 78 218 112
rect 252 78 282 112
rect 189 17 282 78
rect 316 112 382 146
rect 316 78 332 112
rect 366 78 382 112
rect 316 62 382 78
rect 416 162 432 196
rect 466 162 618 196
rect 652 162 777 196
rect 811 210 1127 226
rect 845 192 993 210
rect 416 120 482 162
rect 416 86 432 120
rect 466 86 482 120
rect 416 70 482 86
rect 516 124 582 128
rect 516 90 532 124
rect 566 90 582 124
rect 516 17 582 90
rect 618 120 668 162
rect 811 120 845 176
rect 977 176 993 192
rect 1027 192 1127 210
rect 652 86 668 120
rect 618 70 668 86
rect 702 86 719 120
rect 753 86 770 120
rect 702 17 770 86
rect 811 70 845 86
rect 881 136 931 158
rect 881 102 897 136
rect 881 17 931 102
rect 977 120 1027 176
rect 977 86 993 120
rect 977 70 1027 86
rect 1063 142 1129 158
rect 1063 108 1079 142
rect 1113 108 1129 142
rect 1063 17 1129 108
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
rlabel comment s 0 0 0 0 4 or3b_4
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 607 242 641 276 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 31 94 65 128 0 FreeSans 340 0 0 0 C_N
port 3 nsew
flabel corelocali s 1087 242 1121 276 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 1087 316 1121 350 0 FreeSans 340 0 0 0 X
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 1152 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1060000
string GDS_START 1049840
<< end >>
