magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 1878 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 89 47 119 131
rect 183 47 213 131
rect 280 47 310 119
rect 395 47 425 119
rect 537 47 567 131
rect 667 47 697 177
rect 865 47 895 131
rect 959 47 989 131
rect 1187 47 1217 177
rect 1259 47 1289 177
rect 1376 47 1406 177
rect 1470 47 1500 177
rect 1564 47 1594 177
rect 1695 47 1725 177
<< pmoshvt >>
rect 81 369 117 497
rect 163 369 199 497
rect 279 413 315 497
rect 385 413 421 497
rect 507 413 543 497
rect 659 297 695 497
rect 857 303 893 431
rect 977 303 1013 431
rect 1179 297 1215 497
rect 1273 297 1309 497
rect 1378 297 1414 497
rect 1472 297 1508 497
rect 1566 297 1602 497
rect 1687 297 1723 497
<< ndiff >>
rect 27 103 89 131
rect 27 69 35 103
rect 69 69 89 103
rect 27 47 89 69
rect 119 89 183 131
rect 119 55 129 89
rect 163 55 183 89
rect 119 47 183 55
rect 213 119 265 131
rect 582 131 667 177
rect 477 119 537 131
rect 213 101 280 119
rect 213 67 223 101
rect 257 67 280 101
rect 213 47 280 67
rect 310 89 395 119
rect 310 55 340 89
rect 374 55 395 89
rect 310 47 395 55
rect 425 47 537 119
rect 567 119 667 131
rect 567 85 596 119
rect 630 85 667 119
rect 567 47 667 85
rect 697 101 749 177
rect 697 67 707 101
rect 741 67 749 101
rect 697 47 749 67
rect 803 110 865 131
rect 803 76 811 110
rect 845 76 865 110
rect 803 47 865 76
rect 895 89 959 131
rect 895 55 905 89
rect 939 55 959 89
rect 895 47 959 55
rect 989 110 1041 131
rect 989 76 999 110
rect 1033 76 1041 110
rect 989 47 1041 76
rect 1125 109 1187 177
rect 1125 75 1133 109
rect 1167 75 1187 109
rect 1125 47 1187 75
rect 1217 47 1259 177
rect 1289 89 1376 177
rect 1289 55 1316 89
rect 1350 55 1376 89
rect 1289 47 1376 55
rect 1406 89 1470 177
rect 1406 55 1426 89
rect 1460 55 1470 89
rect 1406 47 1470 55
rect 1500 93 1564 177
rect 1500 59 1520 93
rect 1554 59 1564 93
rect 1500 47 1564 59
rect 1594 101 1695 177
rect 1594 67 1641 101
rect 1675 67 1695 101
rect 1594 47 1695 67
rect 1725 161 1799 177
rect 1725 127 1753 161
rect 1787 127 1799 161
rect 1725 93 1799 127
rect 1725 59 1753 93
rect 1787 59 1799 93
rect 1725 47 1799 59
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 369 81 383
rect 117 369 163 497
rect 199 475 279 497
rect 199 441 222 475
rect 256 441 279 475
rect 199 413 279 441
rect 315 480 385 497
rect 315 446 333 480
rect 367 446 385 480
rect 315 413 385 446
rect 421 413 507 497
rect 543 489 659 497
rect 543 455 592 489
rect 626 455 659 489
rect 543 413 659 455
rect 199 369 262 413
rect 607 297 659 413
rect 695 458 749 497
rect 695 424 707 458
rect 741 424 749 458
rect 910 485 960 497
rect 910 451 918 485
rect 952 451 960 485
rect 1121 489 1179 497
rect 910 431 960 451
rect 1121 455 1133 489
rect 1167 455 1179 489
rect 695 297 749 424
rect 803 349 857 431
rect 803 315 811 349
rect 845 315 857 349
rect 803 303 857 315
rect 893 303 977 431
rect 1013 349 1067 431
rect 1013 315 1025 349
rect 1059 315 1067 349
rect 1013 303 1067 315
rect 1121 297 1179 455
rect 1215 442 1273 497
rect 1215 408 1227 442
rect 1261 408 1273 442
rect 1215 297 1273 408
rect 1309 489 1378 497
rect 1309 455 1327 489
rect 1361 455 1378 489
rect 1309 297 1378 455
rect 1414 448 1472 497
rect 1414 414 1426 448
rect 1460 414 1472 448
rect 1414 380 1472 414
rect 1414 346 1426 380
rect 1460 346 1472 380
rect 1414 297 1472 346
rect 1508 485 1566 497
rect 1508 451 1520 485
rect 1554 451 1566 485
rect 1508 417 1566 451
rect 1508 383 1520 417
rect 1554 383 1566 417
rect 1508 297 1566 383
rect 1602 448 1687 497
rect 1602 414 1641 448
rect 1675 414 1687 448
rect 1602 380 1687 414
rect 1602 346 1641 380
rect 1675 346 1687 380
rect 1602 297 1687 346
rect 1723 485 1799 497
rect 1723 451 1753 485
rect 1787 451 1799 485
rect 1723 417 1799 451
rect 1723 383 1753 417
rect 1787 383 1799 417
rect 1723 349 1799 383
rect 1723 315 1753 349
rect 1787 315 1799 349
rect 1723 297 1799 315
<< ndiffc >>
rect 35 69 69 103
rect 129 55 163 89
rect 223 67 257 101
rect 340 55 374 89
rect 596 85 630 119
rect 707 67 741 101
rect 811 76 845 110
rect 905 55 939 89
rect 999 76 1033 110
rect 1133 75 1167 109
rect 1316 55 1350 89
rect 1426 55 1460 89
rect 1520 59 1554 93
rect 1641 67 1675 101
rect 1753 127 1787 161
rect 1753 59 1787 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 222 441 256 475
rect 333 446 367 480
rect 592 455 626 489
rect 707 424 741 458
rect 918 451 952 485
rect 1133 455 1167 489
rect 811 315 845 349
rect 1025 315 1059 349
rect 1227 408 1261 442
rect 1327 455 1361 489
rect 1426 414 1460 448
rect 1426 346 1460 380
rect 1520 451 1554 485
rect 1520 383 1554 417
rect 1641 414 1675 448
rect 1641 346 1675 380
rect 1753 451 1787 485
rect 1753 383 1787 417
rect 1753 315 1787 349
<< poly >>
rect 81 497 117 523
rect 163 497 199 523
rect 279 497 315 523
rect 385 497 421 523
rect 507 497 543 523
rect 659 497 695 523
rect 279 398 315 413
rect 385 398 421 413
rect 507 398 543 413
rect 81 354 117 369
rect 163 354 199 369
rect 79 265 119 354
rect 22 249 119 265
rect 22 215 32 249
rect 66 215 119 249
rect 22 199 119 215
rect 161 265 201 354
rect 277 273 317 398
rect 383 381 423 398
rect 359 365 423 381
rect 359 331 369 365
rect 403 331 423 365
rect 359 315 423 331
rect 505 381 545 398
rect 505 365 567 381
rect 505 331 515 365
rect 549 331 567 365
rect 505 315 567 331
rect 161 249 235 265
rect 161 215 181 249
rect 215 215 235 249
rect 277 243 435 273
rect 161 199 235 215
rect 395 207 435 243
rect 89 131 119 199
rect 183 131 213 199
rect 280 191 353 201
rect 280 157 296 191
rect 330 157 353 191
rect 280 147 353 157
rect 395 191 459 207
rect 395 157 405 191
rect 439 157 459 191
rect 280 119 310 147
rect 395 141 459 157
rect 395 119 425 141
rect 537 131 567 315
rect 855 457 895 523
rect 857 431 893 457
rect 975 457 1015 523
rect 1179 497 1215 523
rect 1273 497 1309 523
rect 1378 497 1414 523
rect 1472 497 1508 523
rect 1566 497 1602 523
rect 1687 497 1723 523
rect 977 431 1013 457
rect 659 282 695 297
rect 857 288 893 303
rect 977 288 1013 303
rect 657 265 697 282
rect 855 265 895 288
rect 975 265 1015 288
rect 1179 282 1215 297
rect 1273 282 1309 297
rect 1378 282 1414 297
rect 1472 282 1508 297
rect 1566 282 1602 297
rect 1687 282 1723 297
rect 1177 265 1217 282
rect 1271 265 1311 282
rect 609 249 697 265
rect 609 215 619 249
rect 653 215 697 249
rect 609 199 697 215
rect 847 255 923 265
rect 847 221 863 255
rect 897 221 923 255
rect 847 211 923 221
rect 975 249 1069 265
rect 975 215 1025 249
rect 1059 215 1069 249
rect 667 177 697 199
rect 865 131 895 211
rect 975 176 1069 215
rect 1131 249 1217 265
rect 1131 215 1141 249
rect 1175 215 1217 249
rect 1131 199 1217 215
rect 1187 177 1217 199
rect 1259 249 1323 265
rect 1259 215 1269 249
rect 1303 215 1323 249
rect 1259 199 1323 215
rect 1376 259 1416 282
rect 1470 259 1510 282
rect 1564 259 1604 282
rect 1685 259 1725 282
rect 1376 249 1725 259
rect 1376 215 1392 249
rect 1426 215 1725 249
rect 1376 205 1725 215
rect 1259 177 1289 199
rect 1376 177 1406 205
rect 1470 177 1500 205
rect 1564 177 1594 205
rect 1695 177 1725 205
rect 959 146 1069 176
rect 959 131 989 146
rect 89 21 119 47
rect 183 21 213 47
rect 280 21 310 47
rect 395 21 425 47
rect 537 21 567 47
rect 667 21 697 47
rect 865 21 895 47
rect 959 21 989 47
rect 1187 21 1217 47
rect 1259 21 1289 47
rect 1376 21 1406 47
rect 1470 21 1500 47
rect 1564 21 1594 47
rect 1695 21 1725 47
<< polycont >>
rect 32 215 66 249
rect 369 331 403 365
rect 515 331 549 365
rect 181 215 215 249
rect 296 157 330 191
rect 405 157 439 191
rect 619 215 653 249
rect 863 221 897 255
rect 1025 215 1059 249
rect 1141 215 1175 249
rect 1269 215 1303 249
rect 1392 215 1426 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 17 485 69 527
rect 17 451 35 485
rect 17 417 69 451
rect 17 383 35 417
rect 17 367 69 383
rect 103 475 272 493
rect 103 441 222 475
rect 256 441 272 475
rect 103 425 272 441
rect 306 480 481 493
rect 306 446 333 480
rect 367 446 481 480
rect 306 425 481 446
rect 17 249 69 333
rect 17 215 32 249
rect 66 215 69 249
rect 17 191 69 215
rect 103 157 147 425
rect 181 289 268 391
rect 302 365 403 391
rect 302 331 369 365
rect 302 323 403 331
rect 302 289 336 323
rect 370 289 403 323
rect 181 249 259 289
rect 302 265 403 289
rect 215 215 259 249
rect 181 191 259 215
rect 293 241 403 265
rect 447 275 481 425
rect 515 489 653 527
rect 515 455 592 489
rect 626 455 653 489
rect 515 415 653 455
rect 697 458 741 493
rect 697 424 707 458
rect 779 489 1183 527
rect 779 485 1133 489
rect 779 451 918 485
rect 952 455 1133 485
rect 1167 455 1183 489
rect 952 451 1183 455
rect 697 417 741 424
rect 1227 442 1261 493
rect 1311 489 1377 527
rect 1311 455 1327 489
rect 1361 455 1377 489
rect 1311 451 1377 455
rect 697 383 1183 417
rect 697 381 741 383
rect 515 365 741 381
rect 549 331 741 365
rect 515 327 741 331
rect 515 315 559 327
rect 447 249 653 275
rect 447 241 619 249
rect 293 191 371 241
rect 506 215 619 241
rect 293 157 296 191
rect 330 157 371 191
rect 17 123 259 157
rect 293 141 371 157
rect 405 191 472 207
rect 439 187 472 191
rect 405 153 438 157
rect 405 141 472 153
rect 506 199 653 215
rect 17 103 69 123
rect 17 69 35 103
rect 223 101 259 123
rect 506 107 540 199
rect 17 51 69 69
rect 103 55 129 89
rect 163 55 179 89
rect 103 17 179 55
rect 257 67 259 101
rect 223 51 259 67
rect 293 89 540 107
rect 293 55 340 89
rect 374 55 540 89
rect 293 51 540 55
rect 584 119 653 165
rect 584 85 596 119
rect 630 85 653 119
rect 584 17 653 85
rect 697 101 741 327
rect 697 67 707 101
rect 697 51 741 67
rect 779 315 811 349
rect 845 315 861 349
rect 905 323 1025 349
rect 779 187 813 315
rect 905 289 932 323
rect 966 315 1025 323
rect 1059 315 1075 349
rect 966 299 1075 315
rect 905 255 966 289
rect 847 221 863 255
rect 897 221 966 255
rect 779 153 830 187
rect 908 157 966 221
rect 1011 255 1069 265
rect 1011 221 1023 255
rect 1057 249 1069 255
rect 1011 215 1025 221
rect 1059 215 1069 249
rect 1011 199 1069 215
rect 1113 249 1183 383
rect 1426 448 1476 493
rect 1261 408 1382 417
rect 1227 299 1382 408
rect 1113 215 1141 249
rect 1175 215 1183 249
rect 1113 199 1183 215
rect 1227 255 1313 265
rect 1227 221 1232 255
rect 1266 249 1313 255
rect 1266 221 1269 249
rect 1227 215 1269 221
rect 1303 215 1313 249
rect 1227 199 1313 215
rect 1348 263 1382 299
rect 1460 414 1476 448
rect 1426 380 1476 414
rect 1460 346 1476 380
rect 1520 485 1570 527
rect 1554 451 1570 485
rect 1520 417 1570 451
rect 1554 383 1570 417
rect 1520 365 1570 383
rect 1641 448 1719 493
rect 1675 414 1719 448
rect 1641 380 1719 414
rect 1426 331 1476 346
rect 1675 346 1719 380
rect 1426 297 1564 331
rect 1530 263 1564 297
rect 1641 263 1719 346
rect 1753 485 1807 527
rect 1787 451 1807 485
rect 1753 417 1807 451
rect 1787 383 1807 417
rect 1753 349 1807 383
rect 1787 315 1807 349
rect 1753 297 1807 315
rect 1348 249 1486 263
rect 1348 215 1392 249
rect 1426 215 1486 249
rect 1348 211 1486 215
rect 1530 211 1811 263
rect 1348 157 1382 211
rect 1530 177 1564 211
rect 779 110 845 153
rect 908 123 1049 157
rect 779 76 811 110
rect 999 110 1049 123
rect 779 51 845 76
rect 879 55 905 89
rect 939 55 955 89
rect 879 17 955 55
rect 1033 76 1049 110
rect 999 51 1049 76
rect 1083 123 1382 157
rect 1426 143 1564 177
rect 1083 109 1167 123
rect 1083 75 1133 109
rect 1426 89 1476 143
rect 1083 51 1167 75
rect 1201 55 1316 89
rect 1350 55 1366 89
rect 1201 17 1366 55
rect 1400 55 1426 89
rect 1460 55 1476 89
rect 1400 51 1476 55
rect 1520 93 1570 109
rect 1554 59 1570 93
rect 1520 17 1570 59
rect 1641 101 1719 211
rect 1675 67 1719 101
rect 1641 51 1719 67
rect 1753 161 1807 177
rect 1787 127 1807 161
rect 1753 93 1807 127
rect 1787 59 1807 93
rect 1753 17 1807 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 336 289 370 323
rect 438 157 439 187
rect 439 157 472 187
rect 438 153 472 157
rect 932 289 966 323
rect 830 153 864 187
rect 1023 249 1057 255
rect 1023 221 1025 249
rect 1025 221 1057 249
rect 1232 221 1266 255
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
<< metal1 >>
rect 0 561 1840 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 0 496 1840 527
rect 324 323 382 329
rect 324 289 336 323
rect 370 320 382 323
rect 920 323 978 329
rect 920 320 932 323
rect 370 292 932 320
rect 370 289 382 292
rect 324 283 382 289
rect 920 289 932 292
rect 966 289 978 323
rect 920 283 978 289
rect 1011 255 1069 261
rect 1011 221 1023 255
rect 1057 252 1069 255
rect 1220 255 1278 261
rect 1220 252 1232 255
rect 1057 224 1232 252
rect 1057 221 1069 224
rect 1011 215 1069 221
rect 1220 221 1232 224
rect 1266 221 1278 255
rect 1220 215 1278 221
rect 426 187 484 193
rect 426 153 438 187
rect 472 184 484 187
rect 818 187 876 193
rect 818 184 830 187
rect 472 156 830 184
rect 472 153 484 156
rect 426 147 484 153
rect 818 153 830 156
rect 864 153 876 187
rect 818 147 876 153
rect 0 17 1840 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
rect 0 -48 1840 -17
<< labels >>
flabel corelocali s 30 289 64 323 0 FreeSans 200 0 0 0 SCE
port 3 nsew
flabel corelocali s 214 357 248 391 0 FreeSans 200 0 0 0 GATE
port 2 nsew
flabel corelocali s 214 289 248 323 0 FreeSans 200 0 0 0 GATE
port 2 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 200 0 0 0 SCE
port 3 nsew
flabel corelocali s 1685 221 1719 255 0 FreeSans 200 0 0 0 GCLK
port 8 nsew
flabel corelocali s 1685 425 1719 459 0 FreeSans 200 0 0 0 GCLK
port 8 nsew
flabel corelocali s 1685 357 1719 391 0 FreeSans 200 0 0 0 GCLK
port 8 nsew
flabel corelocali s 1685 289 1719 323 0 FreeSans 200 0 0 0 GCLK
port 8 nsew
flabel corelocali s 1593 221 1627 255 0 FreeSans 200 0 0 0 GCLK
port 8 nsew
flabel corelocali s 1777 221 1811 255 0 FreeSans 200 0 0 0 GCLK
port 8 nsew
flabel corelocali s 1685 153 1719 187 0 FreeSans 200 0 0 0 GCLK
port 8 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
flabel metal1 s 1015 221 1049 255 0 FreeSans 200 0 0 0 CLK
port 1 nsew
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
rlabel comment s 0 0 0 0 4 sdlclkp_4
<< properties >>
string FIXED_BBOX 0 0 1840 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 407202
string GDS_START 393426
<< end >>
