magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 18 199 66 323
rect 301 333 377 493
rect 489 333 565 493
rect 771 333 847 493
rect 977 333 1053 493
rect 301 289 1053 333
rect 301 127 377 289
rect 432 215 670 255
rect 722 215 937 255
rect 1004 215 1177 255
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 18 417 69 493
rect 103 451 267 527
rect 18 383 144 417
rect 100 249 144 383
rect 217 289 267 451
rect 421 367 455 527
rect 609 367 737 527
rect 891 367 943 527
rect 1097 299 1176 527
rect 100 215 267 249
rect 100 161 144 215
rect 18 127 144 161
rect 18 51 69 127
rect 217 93 267 181
rect 421 127 659 181
rect 697 143 1158 181
rect 697 127 961 143
rect 421 93 455 127
rect 901 123 961 127
rect 103 17 179 93
rect 217 51 455 93
rect 489 51 857 93
rect 901 51 953 123
rect 1013 17 1047 109
rect 1091 51 1158 143
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
rlabel locali s 18 199 66 323 6 A_N
port 1 nsew signal input
rlabel locali s 432 215 670 255 6 B
port 2 nsew signal input
rlabel locali s 722 215 937 255 6 C
port 3 nsew signal input
rlabel locali s 1004 215 1177 255 6 D
port 4 nsew signal input
rlabel locali s 977 333 1053 493 6 Y
port 5 nsew signal output
rlabel locali s 771 333 847 493 6 Y
port 5 nsew signal output
rlabel locali s 489 333 565 493 6 Y
port 5 nsew signal output
rlabel locali s 301 333 377 493 6 Y
port 5 nsew signal output
rlabel locali s 301 289 1053 333 6 Y
port 5 nsew signal output
rlabel locali s 301 127 377 289 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -48 1196 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 1196 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2331924
string GDS_START 2321864
<< end >>
