magic
tech sky130A
magscale 1 2
timestamp 1604502741
<< locali >>
rect 65 424 115 596
rect 405 424 471 596
rect 65 390 471 424
rect 21 260 87 356
rect 121 226 155 390
rect 193 270 327 356
rect 375 270 455 356
rect 505 336 555 578
rect 489 270 555 336
rect 601 260 743 356
rect 23 192 155 226
rect 23 70 89 192
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 149 458 312 649
rect 633 390 699 649
rect 235 226 501 236
rect 235 202 745 226
rect 235 160 301 202
rect 435 192 745 202
rect 123 104 189 154
rect 335 104 401 159
rect 123 70 401 104
rect 435 70 501 192
rect 535 17 645 158
rect 679 70 745 192
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel locali s 601 260 743 356 6 A1
port 1 nsew signal input
rlabel locali s 505 336 555 578 6 A2
port 2 nsew signal input
rlabel locali s 489 270 555 336 6 A2
port 2 nsew signal input
rlabel locali s 193 270 327 356 6 B1
port 3 nsew signal input
rlabel locali s 375 270 455 356 6 B2
port 4 nsew signal input
rlabel locali s 21 260 87 356 6 C1
port 5 nsew signal input
rlabel locali s 405 424 471 596 6 Y
port 6 nsew signal output
rlabel locali s 121 226 155 390 6 Y
port 6 nsew signal output
rlabel locali s 65 424 115 596 6 Y
port 6 nsew signal output
rlabel locali s 65 390 471 424 6 Y
port 6 nsew signal output
rlabel locali s 23 192 155 226 6 Y
port 6 nsew signal output
rlabel locali s 23 70 89 192 6 Y
port 6 nsew signal output
rlabel metal1 s 0 -49 768 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 617 768 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1163018
string GDS_START 1155714
<< end >>
