magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 87 199 165 339
rect 199 199 267 265
rect 569 199 629 475
rect 837 325 887 493
rect 1025 325 1075 493
rect 663 280 735 323
rect 837 291 1171 325
rect 691 199 735 280
rect 1125 181 1171 291
rect 845 145 1171 181
rect 845 51 895 145
rect 1007 51 1083 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 19 414 69 491
rect 103 448 179 527
rect 245 459 513 493
rect 245 414 279 459
rect 19 380 279 414
rect 322 391 445 425
rect 19 165 53 380
rect 208 312 339 346
rect 301 265 339 312
rect 301 199 359 265
rect 301 165 339 199
rect 19 90 80 165
rect 141 17 175 165
rect 235 131 339 165
rect 407 165 445 391
rect 479 199 513 459
rect 732 359 782 527
rect 931 359 981 527
rect 1119 359 1169 527
rect 769 215 1089 249
rect 769 165 803 215
rect 407 131 803 165
rect 235 90 269 131
rect 323 17 389 96
rect 449 61 483 131
rect 517 17 593 97
rect 637 61 671 131
rect 723 17 799 97
rect 939 17 973 111
rect 1127 17 1161 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
rlabel locali s 691 199 735 280 6 A
port 1 nsew signal input
rlabel locali s 663 280 735 323 6 A
port 1 nsew signal input
rlabel locali s 569 199 629 475 6 B
port 2 nsew signal input
rlabel locali s 87 199 165 339 6 C_N
port 3 nsew signal input
rlabel locali s 199 199 267 265 6 D_N
port 4 nsew signal input
rlabel locali s 1125 181 1171 291 6 X
port 5 nsew signal output
rlabel locali s 1025 325 1075 493 6 X
port 5 nsew signal output
rlabel locali s 1007 51 1083 145 6 X
port 5 nsew signal output
rlabel locali s 845 145 1171 181 6 X
port 5 nsew signal output
rlabel locali s 845 51 895 145 6 X
port 5 nsew signal output
rlabel locali s 837 325 887 493 6 X
port 5 nsew signal output
rlabel locali s 837 291 1171 325 6 X
port 5 nsew signal output
rlabel metal1 s 0 -48 1196 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 1196 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 165908
string GDS_START 156888
<< end >>
