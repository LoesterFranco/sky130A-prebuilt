magic
tech sky130A
magscale 1 2
timestamp 1599588209
<< nwell >>
rect -38 332 1670 704
<< pwell >>
rect 0 0 1632 49
<< scpmos >>
rect 87 368 117 592
rect 177 368 207 592
rect 277 368 307 592
rect 367 368 397 592
rect 467 368 497 592
rect 557 368 587 592
rect 647 368 677 592
rect 737 368 767 592
rect 847 368 877 592
rect 937 368 967 592
rect 1027 368 1057 592
rect 1127 368 1157 592
rect 1217 368 1247 592
rect 1307 368 1337 592
rect 1399 368 1429 592
rect 1497 368 1527 592
<< nmoslvt >>
rect 84 74 114 222
rect 184 74 214 222
rect 270 74 300 222
rect 370 74 400 222
rect 456 74 486 222
rect 556 74 586 222
rect 650 74 680 222
rect 756 74 786 222
rect 844 74 874 222
rect 942 74 972 222
rect 1030 74 1060 222
rect 1116 74 1146 222
rect 1202 74 1232 222
rect 1302 74 1332 222
rect 1402 74 1432 222
rect 1502 74 1532 222
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 141 184 222
rect 114 107 139 141
rect 173 107 184 141
rect 114 74 184 107
rect 214 210 270 222
rect 214 176 225 210
rect 259 176 270 210
rect 214 120 270 176
rect 214 86 225 120
rect 259 86 270 120
rect 214 74 270 86
rect 300 127 370 222
rect 300 93 325 127
rect 359 93 370 127
rect 300 74 370 93
rect 400 202 456 222
rect 400 168 411 202
rect 445 168 456 202
rect 400 120 456 168
rect 400 86 411 120
rect 445 86 456 120
rect 400 74 456 86
rect 486 127 556 222
rect 486 93 511 127
rect 545 93 556 127
rect 486 74 556 93
rect 586 202 650 222
rect 586 168 597 202
rect 631 168 650 202
rect 586 120 650 168
rect 586 86 597 120
rect 631 86 650 120
rect 586 74 650 86
rect 680 127 756 222
rect 680 93 697 127
rect 731 93 756 127
rect 680 74 756 93
rect 786 210 844 222
rect 786 176 797 210
rect 831 176 844 210
rect 786 120 844 176
rect 786 86 797 120
rect 831 86 844 120
rect 786 74 844 86
rect 874 205 942 222
rect 874 171 897 205
rect 931 171 942 205
rect 874 74 942 171
rect 972 116 1030 222
rect 972 82 984 116
rect 1018 82 1030 116
rect 972 74 1030 82
rect 1060 184 1116 222
rect 1060 150 1071 184
rect 1105 150 1116 184
rect 1060 74 1116 150
rect 1146 116 1202 222
rect 1146 82 1157 116
rect 1191 82 1202 116
rect 1146 74 1202 82
rect 1232 160 1302 222
rect 1232 126 1257 160
rect 1291 126 1302 160
rect 1232 74 1302 126
rect 1332 116 1402 222
rect 1332 82 1357 116
rect 1391 82 1402 116
rect 1332 74 1402 82
rect 1432 160 1502 222
rect 1432 126 1457 160
rect 1491 126 1502 160
rect 1432 74 1502 126
rect 1532 100 1605 222
rect 1532 74 1559 100
rect 1547 66 1559 74
rect 1593 66 1605 100
rect 1547 54 1605 66
<< pdiff >>
rect 28 580 87 592
rect 28 546 40 580
rect 74 546 87 580
rect 28 497 87 546
rect 28 463 40 497
rect 74 463 87 497
rect 28 414 87 463
rect 28 380 40 414
rect 74 380 87 414
rect 28 368 87 380
rect 117 580 177 592
rect 117 546 130 580
rect 164 546 177 580
rect 117 497 177 546
rect 117 463 130 497
rect 164 463 177 497
rect 117 414 177 463
rect 117 380 130 414
rect 164 380 177 414
rect 117 368 177 380
rect 207 582 277 592
rect 207 548 220 582
rect 254 548 277 582
rect 207 514 277 548
rect 207 480 220 514
rect 254 480 277 514
rect 207 368 277 480
rect 307 580 367 592
rect 307 546 320 580
rect 354 546 367 580
rect 307 462 367 546
rect 307 428 320 462
rect 354 428 367 462
rect 307 368 367 428
rect 397 472 467 592
rect 397 438 420 472
rect 454 438 467 472
rect 397 368 467 438
rect 497 573 557 592
rect 497 539 510 573
rect 544 539 557 573
rect 497 368 557 539
rect 587 498 647 592
rect 587 464 600 498
rect 634 464 647 498
rect 587 368 647 464
rect 677 573 737 592
rect 677 539 690 573
rect 724 539 737 573
rect 677 368 737 539
rect 767 573 847 592
rect 767 539 790 573
rect 824 539 847 573
rect 767 368 847 539
rect 877 580 937 592
rect 877 546 890 580
rect 924 546 937 580
rect 877 488 937 546
rect 877 454 890 488
rect 924 454 937 488
rect 877 368 937 454
rect 967 568 1027 592
rect 967 534 980 568
rect 1014 534 1027 568
rect 967 368 1027 534
rect 1057 580 1127 592
rect 1057 546 1080 580
rect 1114 546 1127 580
rect 1057 488 1127 546
rect 1057 454 1080 488
rect 1114 454 1127 488
rect 1057 368 1127 454
rect 1157 531 1217 592
rect 1157 497 1170 531
rect 1204 497 1217 531
rect 1157 420 1217 497
rect 1157 386 1170 420
rect 1204 386 1217 420
rect 1157 368 1217 386
rect 1247 580 1307 592
rect 1247 546 1260 580
rect 1294 546 1307 580
rect 1247 508 1307 546
rect 1247 474 1260 508
rect 1294 474 1307 508
rect 1247 368 1307 474
rect 1337 531 1399 592
rect 1337 497 1350 531
rect 1384 497 1399 531
rect 1337 440 1399 497
rect 1337 406 1350 440
rect 1384 406 1399 440
rect 1337 368 1399 406
rect 1429 580 1497 592
rect 1429 546 1450 580
rect 1484 546 1497 580
rect 1429 508 1497 546
rect 1429 474 1450 508
rect 1484 474 1497 508
rect 1429 368 1497 474
rect 1527 580 1596 592
rect 1527 546 1550 580
rect 1584 546 1596 580
rect 1527 508 1596 546
rect 1527 474 1550 508
rect 1584 474 1596 508
rect 1527 368 1596 474
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 139 107 173 141
rect 225 176 259 210
rect 225 86 259 120
rect 325 93 359 127
rect 411 168 445 202
rect 411 86 445 120
rect 511 93 545 127
rect 597 168 631 202
rect 597 86 631 120
rect 697 93 731 127
rect 797 176 831 210
rect 797 86 831 120
rect 897 171 931 205
rect 984 82 1018 116
rect 1071 150 1105 184
rect 1157 82 1191 116
rect 1257 126 1291 160
rect 1357 82 1391 116
rect 1457 126 1491 160
rect 1559 66 1593 100
<< pdiffc >>
rect 40 546 74 580
rect 40 463 74 497
rect 40 380 74 414
rect 130 546 164 580
rect 130 463 164 497
rect 130 380 164 414
rect 220 548 254 582
rect 220 480 254 514
rect 320 546 354 580
rect 320 428 354 462
rect 420 438 454 472
rect 510 539 544 573
rect 600 464 634 498
rect 690 539 724 573
rect 790 539 824 573
rect 890 546 924 580
rect 890 454 924 488
rect 980 534 1014 568
rect 1080 546 1114 580
rect 1080 454 1114 488
rect 1170 497 1204 531
rect 1170 386 1204 420
rect 1260 546 1294 580
rect 1260 474 1294 508
rect 1350 497 1384 531
rect 1350 406 1384 440
rect 1450 546 1484 580
rect 1450 474 1484 508
rect 1550 546 1584 580
rect 1550 474 1584 508
<< poly >>
rect 87 592 117 618
rect 177 592 207 618
rect 277 592 307 618
rect 367 592 397 618
rect 467 592 497 618
rect 557 592 587 618
rect 647 592 677 618
rect 737 592 767 618
rect 847 592 877 618
rect 937 592 967 618
rect 1027 592 1057 618
rect 1127 592 1157 618
rect 1217 592 1247 618
rect 1307 592 1337 618
rect 1399 592 1429 618
rect 1497 592 1527 618
rect 87 353 117 368
rect 177 353 207 368
rect 277 353 307 368
rect 367 353 397 368
rect 467 353 497 368
rect 557 353 587 368
rect 647 353 677 368
rect 737 353 767 368
rect 847 353 877 368
rect 937 353 967 368
rect 1027 353 1057 368
rect 1127 353 1157 368
rect 1217 353 1247 368
rect 1307 353 1337 368
rect 1399 353 1429 368
rect 1497 353 1527 368
rect 84 330 120 353
rect 174 330 210 353
rect 274 330 310 353
rect 84 314 310 330
rect 84 280 124 314
rect 158 280 192 314
rect 226 280 260 314
rect 294 280 310 314
rect 364 310 400 353
rect 464 310 500 353
rect 554 310 590 353
rect 644 310 680 353
rect 734 336 770 353
rect 84 264 310 280
rect 370 294 680 310
rect 84 222 114 264
rect 184 222 214 264
rect 270 222 300 264
rect 370 260 393 294
rect 427 260 461 294
rect 495 260 529 294
rect 563 260 597 294
rect 631 260 680 294
rect 728 320 794 336
rect 728 286 744 320
rect 778 286 794 320
rect 728 270 794 286
rect 844 326 880 353
rect 934 326 970 353
rect 1024 326 1060 353
rect 1124 336 1160 353
rect 1214 336 1250 353
rect 1304 336 1340 353
rect 1396 336 1432 353
rect 844 310 1060 326
rect 844 276 874 310
rect 908 276 942 310
rect 976 276 1010 310
rect 1044 276 1060 310
rect 370 244 680 260
rect 370 222 400 244
rect 456 222 486 244
rect 556 222 586 244
rect 650 222 680 244
rect 756 222 786 270
rect 844 260 1060 276
rect 844 222 874 260
rect 942 222 972 260
rect 1030 222 1060 260
rect 1116 320 1432 336
rect 1116 286 1177 320
rect 1211 286 1245 320
rect 1279 286 1313 320
rect 1347 286 1381 320
rect 1415 286 1432 320
rect 1494 310 1530 353
rect 1116 270 1432 286
rect 1116 222 1146 270
rect 1202 222 1232 270
rect 1302 222 1332 270
rect 1402 222 1432 270
rect 1480 294 1546 310
rect 1480 260 1496 294
rect 1530 260 1546 294
rect 1480 244 1546 260
rect 1502 222 1532 244
rect 84 48 114 74
rect 184 48 214 74
rect 270 48 300 74
rect 370 48 400 74
rect 456 48 486 74
rect 556 48 586 74
rect 650 48 680 74
rect 756 48 786 74
rect 844 48 874 74
rect 942 48 972 74
rect 1030 48 1060 74
rect 1116 48 1146 74
rect 1202 48 1232 74
rect 1302 48 1332 74
rect 1402 48 1432 74
rect 1502 48 1532 74
<< polycont >>
rect 124 280 158 314
rect 192 280 226 314
rect 260 280 294 314
rect 393 260 427 294
rect 461 260 495 294
rect 529 260 563 294
rect 597 260 631 294
rect 744 286 778 320
rect 874 276 908 310
rect 942 276 976 310
rect 1010 276 1044 310
rect 1177 286 1211 320
rect 1245 286 1279 320
rect 1313 286 1347 320
rect 1381 286 1415 320
rect 1496 260 1530 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 24 580 74 649
rect 24 546 40 580
rect 24 497 74 546
rect 24 463 40 497
rect 24 414 74 463
rect 24 380 40 414
rect 24 364 74 380
rect 114 580 170 596
rect 114 546 130 580
rect 164 546 170 580
rect 114 497 170 546
rect 114 463 130 497
rect 164 463 170 497
rect 204 582 270 649
rect 204 548 220 582
rect 254 548 270 582
rect 204 514 270 548
rect 204 480 220 514
rect 254 480 270 514
rect 304 580 740 596
rect 304 546 320 580
rect 354 573 740 580
rect 354 546 510 573
rect 304 539 510 546
rect 544 539 690 573
rect 724 539 740 573
rect 304 532 740 539
rect 774 573 840 649
rect 774 539 790 573
rect 824 539 840 573
rect 774 532 840 539
rect 874 580 940 596
rect 874 546 890 580
rect 924 546 940 580
rect 114 446 170 463
rect 304 462 370 532
rect 304 446 320 462
rect 114 428 320 446
rect 354 428 370 462
rect 114 414 370 428
rect 114 380 130 414
rect 164 412 370 414
rect 404 472 600 498
rect 404 438 420 472
rect 454 464 600 472
rect 634 464 830 498
rect 454 438 470 464
rect 404 412 470 438
rect 164 380 180 412
rect 114 364 180 380
rect 505 378 647 430
rect 796 404 830 464
rect 874 488 940 546
rect 980 568 1030 649
rect 1014 534 1030 568
rect 980 506 1030 534
rect 1064 581 1500 615
rect 1064 580 1114 581
rect 1064 546 1080 580
rect 1260 580 1294 581
rect 874 454 890 488
rect 924 472 940 488
rect 1064 488 1114 546
rect 1064 472 1080 488
rect 924 454 1080 472
rect 874 438 1114 454
rect 1154 531 1220 547
rect 1154 497 1170 531
rect 1204 497 1220 531
rect 1154 424 1220 497
rect 1434 580 1500 581
rect 1260 508 1294 546
rect 1260 458 1294 474
rect 1334 531 1400 547
rect 1334 497 1350 531
rect 1384 497 1400 531
rect 1334 440 1400 497
rect 1434 546 1450 580
rect 1484 546 1500 580
rect 1434 508 1500 546
rect 1434 474 1450 508
rect 1484 474 1500 508
rect 1434 458 1500 474
rect 1534 580 1600 649
rect 1534 546 1550 580
rect 1584 546 1600 580
rect 1534 508 1600 546
rect 1534 474 1550 508
rect 1584 474 1600 508
rect 1534 458 1600 474
rect 1334 424 1350 440
rect 1154 420 1350 424
rect 1154 404 1170 420
rect 796 386 1170 404
rect 1204 406 1350 420
rect 1384 424 1400 440
rect 1384 406 1614 424
rect 1204 390 1614 406
rect 1204 386 1220 390
rect 276 344 762 378
rect 796 370 1220 386
rect 276 330 310 344
rect 108 314 310 330
rect 108 280 124 314
rect 158 280 192 314
rect 226 280 260 314
rect 294 280 310 314
rect 728 336 762 344
rect 1273 336 1431 356
rect 728 320 794 336
rect 108 264 310 280
rect 377 294 647 310
rect 377 260 393 294
rect 427 260 461 294
rect 495 260 529 294
rect 563 260 597 294
rect 631 260 647 294
rect 728 286 744 320
rect 778 286 794 320
rect 728 270 794 286
rect 858 310 1127 326
rect 858 276 874 310
rect 908 276 942 310
rect 976 276 1010 310
rect 1044 276 1127 310
rect 1161 320 1431 336
rect 1161 286 1177 320
rect 1211 286 1245 320
rect 1279 286 1313 320
rect 1347 286 1381 320
rect 1415 286 1431 320
rect 1480 294 1546 310
rect 858 260 1127 276
rect 377 236 647 260
rect 1081 252 1127 260
rect 1480 260 1496 294
rect 1530 260 1546 294
rect 1480 252 1546 260
rect 23 210 275 230
rect 23 176 39 210
rect 73 196 225 210
rect 73 176 89 196
rect 23 120 89 176
rect 259 202 275 210
rect 781 210 847 226
rect 781 202 797 210
rect 259 176 411 202
rect 225 168 411 176
rect 445 168 597 202
rect 631 176 797 202
rect 831 176 847 210
rect 631 168 847 176
rect 23 86 39 120
rect 73 86 89 120
rect 23 70 89 86
rect 123 141 189 162
rect 123 107 139 141
rect 173 107 189 141
rect 123 17 189 107
rect 225 120 275 168
rect 259 86 275 120
rect 225 70 275 86
rect 309 127 375 134
rect 309 93 325 127
rect 359 93 375 127
rect 309 17 375 93
rect 411 120 461 168
rect 445 86 461 120
rect 411 70 461 86
rect 495 127 561 134
rect 495 93 511 127
rect 545 93 561 127
rect 495 17 561 93
rect 597 120 647 168
rect 631 86 647 120
rect 597 70 647 86
rect 681 127 747 134
rect 681 93 697 127
rect 731 93 747 127
rect 681 17 747 93
rect 781 120 847 168
rect 881 205 1031 226
rect 1081 218 1546 252
rect 881 171 897 205
rect 931 184 1031 205
rect 1580 184 1614 390
rect 931 171 1071 184
rect 881 150 1071 171
rect 1105 160 1614 184
rect 1105 150 1257 160
rect 781 86 797 120
rect 831 116 847 120
rect 1241 126 1257 150
rect 1291 150 1457 160
rect 1291 126 1307 150
rect 1241 119 1307 126
rect 1441 126 1457 150
rect 1491 150 1614 160
rect 1491 126 1507 150
rect 1441 119 1507 126
rect 831 86 984 116
rect 781 82 984 86
rect 1018 82 1157 116
rect 1191 85 1207 116
rect 1341 85 1357 116
rect 1191 82 1357 85
rect 1391 85 1407 116
rect 1543 100 1609 116
rect 1543 85 1559 100
rect 1391 82 1559 85
rect 781 66 1559 82
rect 1593 66 1609 100
rect 781 51 1609 66
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o22ai_4
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nwell s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 1087 242 1121 276 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 1279 316 1313 350 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 1375 316 1409 350 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 895 168 929 202 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 991 168 1025 202 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 415 242 449 276 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 511 242 545 276 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 607 242 641 276 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 511 390 545 424 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 607 390 641 424 0 FreeSans 340 0 0 0 A1
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 1632 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1273554
string GDS_START 1260856
<< end >>
