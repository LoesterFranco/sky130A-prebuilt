magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 0 1071 29 1105
rect 63 1071 121 1105
rect 155 1071 213 1105
rect 247 1071 305 1105
rect 339 1071 397 1105
rect 431 1071 489 1105
rect 523 1071 581 1105
rect 615 1071 673 1105
rect 707 1071 765 1105
rect 799 1071 857 1105
rect 891 1071 949 1105
rect 983 1071 1041 1105
rect 1075 1071 1133 1105
rect 1167 1071 1225 1105
rect 1259 1071 1317 1105
rect 1351 1071 1409 1105
rect 1443 1071 1501 1105
rect 1535 1071 1593 1105
rect 1627 1071 1685 1105
rect 1719 1071 1777 1105
rect 1811 1071 1869 1105
rect 1903 1071 1961 1105
rect 1995 1071 2053 1105
rect 2087 1071 2145 1105
rect 2179 1071 2237 1105
rect 2271 1071 2329 1105
rect 2363 1071 2421 1105
rect 2455 1071 2513 1105
rect 2547 1071 2605 1105
rect 2639 1071 2697 1105
rect 2731 1071 2789 1105
rect 2823 1071 2881 1105
rect 2915 1071 2973 1105
rect 3007 1071 3065 1105
rect 3099 1071 3157 1105
rect 3191 1071 3249 1105
rect 3283 1071 3341 1105
rect 3375 1071 3433 1105
rect 3467 1071 3525 1105
rect 3559 1071 3617 1105
rect 3651 1071 3709 1105
rect 3743 1071 3801 1105
rect 3835 1071 3893 1105
rect 3927 1071 3985 1105
rect 4019 1071 4077 1105
rect 4111 1071 4169 1105
rect 4203 1071 4261 1105
rect 4295 1071 4353 1105
rect 4387 1071 4445 1105
rect 4479 1071 4537 1105
rect 4571 1071 4629 1105
rect 4663 1071 4721 1105
rect 4755 1071 4813 1105
rect 4847 1071 4905 1105
rect 4939 1071 4997 1105
rect 5031 1071 5089 1105
rect 5123 1071 5152 1105
rect 129 979 172 1071
rect 301 911 367 969
rect 619 956 669 1071
rect 19 823 183 877
rect 113 667 179 721
rect 119 561 179 667
rect 317 737 351 911
rect 558 829 625 883
rect 663 829 730 883
rect 1116 979 1159 1071
rect 1417 979 1460 1071
rect 1907 956 1957 1071
rect 293 731 379 737
rect 293 697 305 731
rect 339 697 379 731
rect 293 663 379 697
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 283 561
rect 119 421 179 527
rect 113 367 179 421
rect 317 425 351 663
rect 1105 823 1269 877
rect 1307 823 1471 877
rect 293 391 379 425
rect 293 357 305 391
rect 339 357 379 391
rect 293 351 379 357
rect 19 211 183 265
rect 317 177 351 351
rect 1109 667 1175 721
rect 1109 561 1169 667
rect 1401 667 1467 721
rect 1407 561 1467 667
rect 1846 829 1913 883
rect 1951 829 2018 883
rect 2404 979 2447 1071
rect 2705 979 2748 1071
rect 3195 956 3245 1071
rect 1005 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1571 561
rect 129 17 172 109
rect 301 119 367 177
rect 558 205 625 259
rect 663 205 730 259
rect 1109 421 1169 527
rect 1109 367 1175 421
rect 1407 421 1467 527
rect 1401 367 1467 421
rect 2393 823 2557 877
rect 2595 823 2759 877
rect 1105 211 1269 265
rect 1307 211 1471 265
rect 2397 667 2463 721
rect 2397 561 2457 667
rect 2689 667 2755 721
rect 2695 561 2755 667
rect 3134 829 3201 883
rect 3239 829 3306 883
rect 3692 979 3735 1071
rect 3993 979 4036 1071
rect 4483 956 4533 1071
rect 2293 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2859 561
rect 619 17 669 132
rect 1116 17 1159 109
rect 1417 17 1460 109
rect 1846 205 1913 259
rect 1951 205 2018 259
rect 2397 421 2457 527
rect 2397 367 2463 421
rect 2695 421 2755 527
rect 2689 367 2755 421
rect 3681 823 3845 877
rect 3883 823 4047 877
rect 2393 211 2557 265
rect 2595 211 2759 265
rect 3685 667 3751 721
rect 3685 561 3745 667
rect 3977 667 4043 721
rect 3983 561 4043 667
rect 4422 829 4489 883
rect 4527 829 4594 883
rect 4980 979 5023 1071
rect 3581 527 3617 561
rect 3651 527 3709 561
rect 3743 527 3801 561
rect 3835 527 3893 561
rect 3927 527 3985 561
rect 4019 527 4077 561
rect 4111 527 4147 561
rect 1907 17 1957 132
rect 2404 17 2447 109
rect 2705 17 2748 109
rect 3134 205 3201 259
rect 3239 205 3306 259
rect 3685 421 3745 527
rect 3685 367 3751 421
rect 3983 421 4043 527
rect 3977 367 4043 421
rect 4969 823 5133 877
rect 3681 211 3845 265
rect 3883 211 4047 265
rect 4973 667 5039 721
rect 4973 561 5033 667
rect 4869 527 4905 561
rect 4939 527 4997 561
rect 5031 527 5089 561
rect 5123 527 5152 561
rect 3195 17 3245 132
rect 3692 17 3735 109
rect 3993 17 4036 109
rect 4422 205 4489 259
rect 4527 205 4594 259
rect 4973 421 5033 527
rect 4973 367 5039 421
rect 4969 211 5133 265
rect 4483 17 4533 132
rect 4980 17 5023 109
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3341 17
rect 3375 -17 3433 17
rect 3467 -17 3525 17
rect 3559 -17 3617 17
rect 3651 -17 3709 17
rect 3743 -17 3801 17
rect 3835 -17 3893 17
rect 3927 -17 3985 17
rect 4019 -17 4077 17
rect 4111 -17 4169 17
rect 4203 -17 4261 17
rect 4295 -17 4353 17
rect 4387 -17 4445 17
rect 4479 -17 4537 17
rect 4571 -17 4629 17
rect 4663 -17 4721 17
rect 4755 -17 4813 17
rect 4847 -17 4905 17
rect 4939 -17 4997 17
rect 5031 -17 5089 17
rect 5123 -17 5152 17
<< viali >>
rect 29 1071 63 1105
rect 121 1071 155 1105
rect 213 1071 247 1105
rect 305 1071 339 1105
rect 397 1071 431 1105
rect 489 1071 523 1105
rect 581 1071 615 1105
rect 673 1071 707 1105
rect 765 1071 799 1105
rect 857 1071 891 1105
rect 949 1071 983 1105
rect 1041 1071 1075 1105
rect 1133 1071 1167 1105
rect 1225 1071 1259 1105
rect 1317 1071 1351 1105
rect 1409 1071 1443 1105
rect 1501 1071 1535 1105
rect 1593 1071 1627 1105
rect 1685 1071 1719 1105
rect 1777 1071 1811 1105
rect 1869 1071 1903 1105
rect 1961 1071 1995 1105
rect 2053 1071 2087 1105
rect 2145 1071 2179 1105
rect 2237 1071 2271 1105
rect 2329 1071 2363 1105
rect 2421 1071 2455 1105
rect 2513 1071 2547 1105
rect 2605 1071 2639 1105
rect 2697 1071 2731 1105
rect 2789 1071 2823 1105
rect 2881 1071 2915 1105
rect 2973 1071 3007 1105
rect 3065 1071 3099 1105
rect 3157 1071 3191 1105
rect 3249 1071 3283 1105
rect 3341 1071 3375 1105
rect 3433 1071 3467 1105
rect 3525 1071 3559 1105
rect 3617 1071 3651 1105
rect 3709 1071 3743 1105
rect 3801 1071 3835 1105
rect 3893 1071 3927 1105
rect 3985 1071 4019 1105
rect 4077 1071 4111 1105
rect 4169 1071 4203 1105
rect 4261 1071 4295 1105
rect 4353 1071 4387 1105
rect 4445 1071 4479 1105
rect 4537 1071 4571 1105
rect 4629 1071 4663 1105
rect 4721 1071 4755 1105
rect 4813 1071 4847 1105
rect 4905 1071 4939 1105
rect 4997 1071 5031 1105
rect 5089 1071 5123 1105
rect 305 697 339 731
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 357 339 391
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 3617 527 3651 561
rect 3709 527 3743 561
rect 3801 527 3835 561
rect 3893 527 3927 561
rect 3985 527 4019 561
rect 4077 527 4111 561
rect 4905 527 4939 561
rect 4997 527 5031 561
rect 5089 527 5123 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
rect 2881 -17 2915 17
rect 2973 -17 3007 17
rect 3065 -17 3099 17
rect 3157 -17 3191 17
rect 3249 -17 3283 17
rect 3341 -17 3375 17
rect 3433 -17 3467 17
rect 3525 -17 3559 17
rect 3617 -17 3651 17
rect 3709 -17 3743 17
rect 3801 -17 3835 17
rect 3893 -17 3927 17
rect 3985 -17 4019 17
rect 4077 -17 4111 17
rect 4169 -17 4203 17
rect 4261 -17 4295 17
rect 4353 -17 4387 17
rect 4445 -17 4479 17
rect 4537 -17 4571 17
rect 4629 -17 4663 17
rect 4721 -17 4755 17
rect 4813 -17 4847 17
rect 4905 -17 4939 17
rect 4997 -17 5031 17
rect 5089 -17 5123 17
<< obsli1 >>
rect 29 945 95 1037
rect 206 1003 435 1037
rect 206 945 267 1003
rect 29 911 267 945
rect 401 934 435 1003
rect 535 971 585 1022
rect 469 937 585 971
rect 703 971 753 1022
rect 853 1003 1082 1037
rect 703 937 819 971
rect 206 903 267 911
rect 19 755 257 789
rect 19 646 79 755
rect 19 595 85 646
rect 223 629 257 755
rect 469 847 503 937
rect 420 827 503 847
rect 785 847 819 937
rect 853 934 887 1003
rect 921 911 987 969
rect 1021 945 1082 1003
rect 1193 945 1259 1037
rect 1021 911 1259 945
rect 1317 945 1383 1037
rect 1494 1003 1723 1037
rect 1494 945 1555 1003
rect 1317 911 1555 945
rect 1589 911 1655 969
rect 1689 934 1723 1003
rect 1823 971 1873 1022
rect 1757 937 1873 971
rect 1991 971 2041 1022
rect 2141 1003 2370 1037
rect 1991 937 2107 971
rect 785 827 868 847
rect 420 795 524 827
rect 764 795 868 827
rect 420 793 576 795
rect 490 761 576 793
rect 223 595 283 629
rect 19 442 85 493
rect 19 333 79 442
rect 223 459 283 493
rect 223 333 257 459
rect 422 629 456 759
rect 385 595 456 629
rect 510 595 576 761
rect 611 561 677 795
rect 712 793 868 795
rect 712 761 798 793
rect 712 595 778 761
rect 832 629 866 759
rect 937 737 971 911
rect 1021 903 1082 911
rect 1494 903 1555 911
rect 1031 755 1269 789
rect 909 731 995 737
rect 909 697 949 731
rect 983 697 995 731
rect 909 663 995 697
rect 832 595 903 629
rect 385 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 903 561
rect 385 459 456 493
rect 19 299 257 333
rect 206 177 267 185
rect 422 329 456 459
rect 510 327 576 493
rect 490 295 576 327
rect 420 293 576 295
rect 611 293 677 527
rect 712 327 778 493
rect 832 459 903 493
rect 832 329 866 459
rect 937 425 971 663
rect 1031 629 1065 755
rect 1005 595 1065 629
rect 1209 646 1269 755
rect 1203 595 1269 646
rect 1307 755 1545 789
rect 1307 646 1367 755
rect 1307 595 1373 646
rect 1511 629 1545 755
rect 1605 737 1639 911
rect 1757 847 1791 937
rect 1708 827 1791 847
rect 2073 847 2107 937
rect 2141 934 2175 1003
rect 2209 911 2275 969
rect 2309 945 2370 1003
rect 2481 945 2547 1037
rect 2309 911 2547 945
rect 2605 945 2671 1037
rect 2782 1003 3011 1037
rect 2782 945 2843 1003
rect 2605 911 2843 945
rect 2877 911 2943 969
rect 2977 934 3011 1003
rect 3111 971 3161 1022
rect 3045 937 3161 971
rect 3279 971 3329 1022
rect 3429 1003 3658 1037
rect 3279 937 3395 971
rect 2073 827 2156 847
rect 1708 795 1812 827
rect 2052 795 2156 827
rect 1708 793 1864 795
rect 1778 761 1864 793
rect 1581 731 1667 737
rect 1581 697 1593 731
rect 1627 697 1667 731
rect 1581 663 1667 697
rect 1511 595 1571 629
rect 1005 459 1065 493
rect 909 391 995 425
rect 909 357 949 391
rect 983 357 995 391
rect 909 351 995 357
rect 712 295 798 327
rect 712 293 868 295
rect 420 261 524 293
rect 764 261 868 293
rect 420 241 503 261
rect 29 143 267 177
rect 29 51 95 143
rect 206 85 267 143
rect 401 85 435 154
rect 469 151 503 241
rect 785 241 868 261
rect 785 151 819 241
rect 937 177 971 351
rect 1031 333 1065 459
rect 1203 442 1269 493
rect 1209 333 1269 442
rect 1031 299 1269 333
rect 1307 442 1373 493
rect 1307 333 1367 442
rect 1511 459 1571 493
rect 1511 333 1545 459
rect 1605 425 1639 663
rect 1710 629 1744 759
rect 1673 595 1744 629
rect 1798 595 1864 761
rect 1899 561 1965 795
rect 2000 793 2156 795
rect 2000 761 2086 793
rect 2000 595 2066 761
rect 2120 629 2154 759
rect 2225 737 2259 911
rect 2309 903 2370 911
rect 2782 903 2843 911
rect 2319 755 2557 789
rect 2197 731 2283 737
rect 2197 697 2237 731
rect 2271 697 2283 731
rect 2197 663 2283 697
rect 2120 595 2191 629
rect 1673 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2191 561
rect 1673 459 1744 493
rect 1581 391 1667 425
rect 1581 357 1593 391
rect 1627 357 1667 391
rect 1581 351 1667 357
rect 1307 299 1545 333
rect 1021 177 1082 185
rect 1494 177 1555 185
rect 1605 177 1639 351
rect 1710 329 1744 459
rect 1798 327 1864 493
rect 1778 295 1864 327
rect 1708 293 1864 295
rect 1899 293 1965 527
rect 2000 327 2066 493
rect 2120 459 2191 493
rect 2120 329 2154 459
rect 2225 425 2259 663
rect 2319 629 2353 755
rect 2293 595 2353 629
rect 2497 646 2557 755
rect 2491 595 2557 646
rect 2595 755 2833 789
rect 2595 646 2655 755
rect 2595 595 2661 646
rect 2799 629 2833 755
rect 2893 737 2927 911
rect 3045 847 3079 937
rect 2996 827 3079 847
rect 3361 847 3395 937
rect 3429 934 3463 1003
rect 3497 911 3563 969
rect 3597 945 3658 1003
rect 3769 945 3835 1037
rect 3597 911 3835 945
rect 3893 945 3959 1037
rect 4070 1003 4299 1037
rect 4070 945 4131 1003
rect 3893 911 4131 945
rect 4165 911 4231 969
rect 4265 934 4299 1003
rect 4399 971 4449 1022
rect 4333 937 4449 971
rect 4567 971 4617 1022
rect 4717 1003 4946 1037
rect 4567 937 4683 971
rect 3361 827 3444 847
rect 2996 795 3100 827
rect 3340 795 3444 827
rect 2996 793 3152 795
rect 3066 761 3152 793
rect 2869 731 2955 737
rect 2869 697 2881 731
rect 2915 697 2955 731
rect 2869 663 2955 697
rect 2799 595 2859 629
rect 2293 459 2353 493
rect 2197 391 2283 425
rect 2197 357 2237 391
rect 2271 357 2283 391
rect 2197 351 2283 357
rect 2000 295 2086 327
rect 2000 293 2156 295
rect 1708 261 1812 293
rect 2052 261 2156 293
rect 1708 241 1791 261
rect 469 117 585 151
rect 206 51 435 85
rect 535 66 585 117
rect 703 117 819 151
rect 703 66 753 117
rect 853 85 887 154
rect 921 119 987 177
rect 1021 143 1259 177
rect 1021 85 1082 143
rect 853 51 1082 85
rect 1193 51 1259 143
rect 1317 143 1555 177
rect 1317 51 1383 143
rect 1494 85 1555 143
rect 1589 119 1655 177
rect 1689 85 1723 154
rect 1757 151 1791 241
rect 2073 241 2156 261
rect 2073 151 2107 241
rect 2225 177 2259 351
rect 2319 333 2353 459
rect 2491 442 2557 493
rect 2497 333 2557 442
rect 2319 299 2557 333
rect 2595 442 2661 493
rect 2595 333 2655 442
rect 2799 459 2859 493
rect 2799 333 2833 459
rect 2893 425 2927 663
rect 2998 629 3032 759
rect 2961 595 3032 629
rect 3086 595 3152 761
rect 3187 561 3253 795
rect 3288 793 3444 795
rect 3288 761 3374 793
rect 3288 595 3354 761
rect 3408 629 3442 759
rect 3513 737 3547 911
rect 3597 903 3658 911
rect 4070 903 4131 911
rect 3607 755 3845 789
rect 3485 731 3571 737
rect 3485 697 3525 731
rect 3559 697 3571 731
rect 3485 663 3571 697
rect 3408 595 3479 629
rect 2961 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3157 561
rect 3191 527 3249 561
rect 3283 527 3341 561
rect 3375 527 3433 561
rect 3467 527 3479 561
rect 2961 459 3032 493
rect 2869 391 2955 425
rect 2869 357 2881 391
rect 2915 357 2955 391
rect 2869 351 2955 357
rect 2595 299 2833 333
rect 2309 177 2370 185
rect 2782 177 2843 185
rect 2893 177 2927 351
rect 2998 329 3032 459
rect 3086 327 3152 493
rect 3066 295 3152 327
rect 2996 293 3152 295
rect 3187 293 3253 527
rect 3288 327 3354 493
rect 3408 459 3479 493
rect 3408 329 3442 459
rect 3513 425 3547 663
rect 3607 629 3641 755
rect 3581 595 3641 629
rect 3785 646 3845 755
rect 3779 595 3845 646
rect 3883 755 4121 789
rect 3883 646 3943 755
rect 3883 595 3949 646
rect 4087 629 4121 755
rect 4181 737 4215 911
rect 4333 847 4367 937
rect 4284 827 4367 847
rect 4649 847 4683 937
rect 4717 934 4751 1003
rect 4785 911 4851 969
rect 4885 945 4946 1003
rect 5057 945 5123 1037
rect 4885 911 5123 945
rect 4649 827 4732 847
rect 4284 795 4388 827
rect 4628 795 4732 827
rect 4284 793 4440 795
rect 4354 761 4440 793
rect 4157 731 4243 737
rect 4157 697 4169 731
rect 4203 697 4243 731
rect 4157 663 4243 697
rect 4087 595 4147 629
rect 3581 459 3641 493
rect 3485 391 3571 425
rect 3485 357 3525 391
rect 3559 357 3571 391
rect 3485 351 3571 357
rect 3288 295 3374 327
rect 3288 293 3444 295
rect 2996 261 3100 293
rect 3340 261 3444 293
rect 2996 241 3079 261
rect 1757 117 1873 151
rect 1494 51 1723 85
rect 1823 66 1873 117
rect 1991 117 2107 151
rect 1991 66 2041 117
rect 2141 85 2175 154
rect 2209 119 2275 177
rect 2309 143 2547 177
rect 2309 85 2370 143
rect 2141 51 2370 85
rect 2481 51 2547 143
rect 2605 143 2843 177
rect 2605 51 2671 143
rect 2782 85 2843 143
rect 2877 119 2943 177
rect 2977 85 3011 154
rect 3045 151 3079 241
rect 3361 241 3444 261
rect 3361 151 3395 241
rect 3513 177 3547 351
rect 3607 333 3641 459
rect 3779 442 3845 493
rect 3785 333 3845 442
rect 3607 299 3845 333
rect 3883 442 3949 493
rect 3883 333 3943 442
rect 4087 459 4147 493
rect 4087 333 4121 459
rect 4181 425 4215 663
rect 4286 629 4320 759
rect 4249 595 4320 629
rect 4374 595 4440 761
rect 4475 561 4541 795
rect 4576 793 4732 795
rect 4576 761 4662 793
rect 4576 595 4642 761
rect 4696 629 4730 759
rect 4801 737 4835 911
rect 4885 903 4946 911
rect 4895 755 5133 789
rect 4773 731 4859 737
rect 4773 697 4813 731
rect 4847 697 4859 731
rect 4773 663 4859 697
rect 4696 595 4767 629
rect 4249 527 4261 561
rect 4295 527 4353 561
rect 4387 527 4445 561
rect 4479 527 4537 561
rect 4571 527 4629 561
rect 4663 527 4721 561
rect 4755 527 4767 561
rect 4249 459 4320 493
rect 4157 391 4243 425
rect 4157 357 4169 391
rect 4203 357 4243 391
rect 4157 351 4243 357
rect 3883 299 4121 333
rect 3597 177 3658 185
rect 4070 177 4131 185
rect 4181 177 4215 351
rect 4286 329 4320 459
rect 4374 327 4440 493
rect 4354 295 4440 327
rect 4284 293 4440 295
rect 4475 293 4541 527
rect 4576 327 4642 493
rect 4696 459 4767 493
rect 4696 329 4730 459
rect 4801 425 4835 663
rect 4895 629 4929 755
rect 4869 595 4929 629
rect 5073 646 5133 755
rect 5067 595 5133 646
rect 4869 459 4929 493
rect 4773 391 4859 425
rect 4773 357 4813 391
rect 4847 357 4859 391
rect 4773 351 4859 357
rect 4576 295 4662 327
rect 4576 293 4732 295
rect 4284 261 4388 293
rect 4628 261 4732 293
rect 4284 241 4367 261
rect 3045 117 3161 151
rect 2782 51 3011 85
rect 3111 66 3161 117
rect 3279 117 3395 151
rect 3279 66 3329 117
rect 3429 85 3463 154
rect 3497 119 3563 177
rect 3597 143 3835 177
rect 3597 85 3658 143
rect 3429 51 3658 85
rect 3769 51 3835 143
rect 3893 143 4131 177
rect 3893 51 3959 143
rect 4070 85 4131 143
rect 4165 119 4231 177
rect 4265 85 4299 154
rect 4333 151 4367 241
rect 4649 241 4732 261
rect 4649 151 4683 241
rect 4801 177 4835 351
rect 4895 333 4929 459
rect 5067 442 5133 493
rect 5073 333 5133 442
rect 4895 299 5133 333
rect 4885 177 4946 185
rect 4333 117 4449 151
rect 4070 51 4299 85
rect 4399 66 4449 117
rect 4567 117 4683 151
rect 4567 66 4617 117
rect 4717 85 4751 154
rect 4785 119 4851 177
rect 4885 143 5123 177
rect 4885 85 4946 143
rect 4717 51 4946 85
rect 5057 51 5123 143
<< obsli1c >>
rect 949 697 983 731
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 1593 697 1627 731
rect 949 357 983 391
rect 2237 697 2271 731
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 1593 357 1627 391
rect 2881 697 2915 731
rect 2237 357 2271 391
rect 3525 697 3559 731
rect 2973 527 3007 561
rect 3065 527 3099 561
rect 3157 527 3191 561
rect 3249 527 3283 561
rect 3341 527 3375 561
rect 3433 527 3467 561
rect 2881 357 2915 391
rect 4169 697 4203 731
rect 3525 357 3559 391
rect 4813 697 4847 731
rect 4261 527 4295 561
rect 4353 527 4387 561
rect 4445 527 4479 561
rect 4537 527 4571 561
rect 4629 527 4663 561
rect 4721 527 4755 561
rect 4169 357 4203 391
rect 4813 357 4847 391
<< metal1 >>
rect 0 1105 5152 1136
rect 0 1071 29 1105
rect 63 1071 121 1105
rect 155 1071 213 1105
rect 247 1071 305 1105
rect 339 1071 397 1105
rect 431 1071 489 1105
rect 523 1071 581 1105
rect 615 1071 673 1105
rect 707 1071 765 1105
rect 799 1071 857 1105
rect 891 1071 949 1105
rect 983 1071 1041 1105
rect 1075 1071 1133 1105
rect 1167 1071 1225 1105
rect 1259 1071 1317 1105
rect 1351 1071 1409 1105
rect 1443 1071 1501 1105
rect 1535 1071 1593 1105
rect 1627 1071 1685 1105
rect 1719 1071 1777 1105
rect 1811 1071 1869 1105
rect 1903 1071 1961 1105
rect 1995 1071 2053 1105
rect 2087 1071 2145 1105
rect 2179 1071 2237 1105
rect 2271 1071 2329 1105
rect 2363 1071 2421 1105
rect 2455 1071 2513 1105
rect 2547 1071 2605 1105
rect 2639 1071 2697 1105
rect 2731 1071 2789 1105
rect 2823 1071 2881 1105
rect 2915 1071 2973 1105
rect 3007 1071 3065 1105
rect 3099 1071 3157 1105
rect 3191 1071 3249 1105
rect 3283 1071 3341 1105
rect 3375 1071 3433 1105
rect 3467 1071 3525 1105
rect 3559 1071 3617 1105
rect 3651 1071 3709 1105
rect 3743 1071 3801 1105
rect 3835 1071 3893 1105
rect 3927 1071 3985 1105
rect 4019 1071 4077 1105
rect 4111 1071 4169 1105
rect 4203 1071 4261 1105
rect 4295 1071 4353 1105
rect 4387 1071 4445 1105
rect 4479 1071 4537 1105
rect 4571 1071 4629 1105
rect 4663 1071 4721 1105
rect 4755 1071 4813 1105
rect 4847 1071 4905 1105
rect 4939 1071 4997 1105
rect 5031 1071 5089 1105
rect 5123 1071 5152 1105
rect 0 1040 5152 1071
rect 293 731 351 737
rect 293 697 305 731
rect 339 728 351 731
rect 937 731 995 737
rect 937 728 949 731
rect 339 700 949 728
rect 339 697 351 700
rect 293 691 351 697
rect 937 697 949 700
rect 983 728 995 731
rect 1581 731 1639 737
rect 1581 728 1593 731
rect 983 700 1593 728
rect 983 697 995 700
rect 937 691 995 697
rect 1581 697 1593 700
rect 1627 728 1639 731
rect 2225 731 2283 737
rect 2225 728 2237 731
rect 1627 700 2237 728
rect 1627 697 1639 700
rect 1581 691 1639 697
rect 2225 697 2237 700
rect 2271 728 2283 731
rect 2869 731 2927 737
rect 2869 728 2881 731
rect 2271 700 2881 728
rect 2271 697 2283 700
rect 2225 691 2283 697
rect 2869 697 2881 700
rect 2915 728 2927 731
rect 3513 731 3571 737
rect 3513 728 3525 731
rect 2915 700 3525 728
rect 2915 697 2927 700
rect 2869 691 2927 697
rect 3513 697 3525 700
rect 3559 728 3571 731
rect 4157 731 4215 737
rect 4157 728 4169 731
rect 3559 700 4169 728
rect 3559 697 3571 700
rect 3513 691 3571 697
rect 4157 697 4169 700
rect 4203 728 4215 731
rect 4801 731 4859 737
rect 4801 728 4813 731
rect 4203 700 4813 728
rect 4203 697 4215 700
rect 4157 691 4215 697
rect 4801 697 4813 700
rect 4847 697 4859 731
rect 4801 691 4859 697
rect 0 561 5152 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3157 561
rect 3191 527 3249 561
rect 3283 527 3341 561
rect 3375 527 3433 561
rect 3467 527 3617 561
rect 3651 527 3709 561
rect 3743 527 3801 561
rect 3835 527 3893 561
rect 3927 527 3985 561
rect 4019 527 4077 561
rect 4111 527 4261 561
rect 4295 527 4353 561
rect 4387 527 4445 561
rect 4479 527 4537 561
rect 4571 527 4629 561
rect 4663 527 4721 561
rect 4755 527 4905 561
rect 4939 527 4997 561
rect 5031 527 5089 561
rect 5123 527 5152 561
rect 0 496 5152 527
rect 293 391 351 397
rect 293 357 305 391
rect 339 388 351 391
rect 937 391 995 397
rect 937 388 949 391
rect 339 360 949 388
rect 339 357 351 360
rect 293 351 351 357
rect 937 357 949 360
rect 983 388 995 391
rect 1581 391 1639 397
rect 1581 388 1593 391
rect 983 360 1593 388
rect 983 357 995 360
rect 937 351 995 357
rect 1581 357 1593 360
rect 1627 388 1639 391
rect 2225 391 2283 397
rect 2225 388 2237 391
rect 1627 360 2237 388
rect 1627 357 1639 360
rect 1581 351 1639 357
rect 2225 357 2237 360
rect 2271 388 2283 391
rect 2869 391 2927 397
rect 2869 388 2881 391
rect 2271 360 2881 388
rect 2271 357 2283 360
rect 2225 351 2283 357
rect 2869 357 2881 360
rect 2915 388 2927 391
rect 3513 391 3571 397
rect 3513 388 3525 391
rect 2915 360 3525 388
rect 2915 357 2927 360
rect 2869 351 2927 357
rect 3513 357 3525 360
rect 3559 388 3571 391
rect 4157 391 4215 397
rect 4157 388 4169 391
rect 3559 360 4169 388
rect 3559 357 3571 360
rect 3513 351 3571 357
rect 4157 357 4169 360
rect 4203 388 4215 391
rect 4801 391 4859 397
rect 4801 388 4813 391
rect 4203 360 4813 388
rect 4203 357 4215 360
rect 4157 351 4215 357
rect 4801 357 4813 360
rect 4847 357 4859 391
rect 4801 351 4859 357
rect 0 17 5152 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3341 17
rect 3375 -17 3433 17
rect 3467 -17 3525 17
rect 3559 -17 3617 17
rect 3651 -17 3709 17
rect 3743 -17 3801 17
rect 3835 -17 3893 17
rect 3927 -17 3985 17
rect 4019 -17 4077 17
rect 4111 -17 4169 17
rect 4203 -17 4261 17
rect 4295 -17 4353 17
rect 4387 -17 4445 17
rect 4479 -17 4537 17
rect 4571 -17 4629 17
rect 4663 -17 4721 17
rect 4755 -17 4813 17
rect 4847 -17 4905 17
rect 4939 -17 4997 17
rect 5031 -17 5089 17
rect 5123 -17 5152 17
rect 0 -48 5152 -17
<< obsm1 >>
rect 23 657 81 666
rect 211 657 269 666
rect 410 657 468 666
rect 23 629 468 657
rect 23 620 81 629
rect 211 620 269 629
rect 410 620 468 629
rect 820 657 878 666
rect 1019 657 1077 666
rect 1207 657 1265 666
rect 820 629 1265 657
rect 820 620 878 629
rect 1019 620 1077 629
rect 1207 620 1265 629
rect 1311 657 1369 666
rect 1499 657 1557 666
rect 1698 657 1756 666
rect 1311 629 1756 657
rect 1311 620 1369 629
rect 1499 620 1557 629
rect 1698 620 1756 629
rect 2108 657 2166 666
rect 2307 657 2365 666
rect 2495 657 2553 666
rect 2108 629 2553 657
rect 2108 620 2166 629
rect 2307 620 2365 629
rect 2495 620 2553 629
rect 2599 657 2657 666
rect 2787 657 2845 666
rect 2986 657 3044 666
rect 2599 629 3044 657
rect 2599 620 2657 629
rect 2787 620 2845 629
rect 2986 620 3044 629
rect 3396 657 3454 666
rect 3595 657 3653 666
rect 3783 657 3841 666
rect 3396 629 3841 657
rect 3396 620 3454 629
rect 3595 620 3653 629
rect 3783 620 3841 629
rect 3887 657 3945 666
rect 4075 657 4133 666
rect 4274 657 4332 666
rect 3887 629 4332 657
rect 3887 620 3945 629
rect 4075 620 4133 629
rect 4274 620 4332 629
rect 4684 657 4742 666
rect 4883 657 4941 666
rect 5071 657 5129 666
rect 4684 629 5129 657
rect 4684 620 4742 629
rect 4883 620 4941 629
rect 5071 620 5129 629
rect 23 459 81 468
rect 211 459 269 468
rect 410 459 468 468
rect 23 431 468 459
rect 23 422 81 431
rect 211 422 269 431
rect 410 422 468 431
rect 820 459 878 468
rect 1019 459 1077 468
rect 1207 459 1265 468
rect 820 431 1265 459
rect 820 422 878 431
rect 1019 422 1077 431
rect 1207 422 1265 431
rect 1311 459 1369 468
rect 1499 459 1557 468
rect 1698 459 1756 468
rect 1311 431 1756 459
rect 1311 422 1369 431
rect 1499 422 1557 431
rect 1698 422 1756 431
rect 2108 459 2166 468
rect 2307 459 2365 468
rect 2495 459 2553 468
rect 2108 431 2553 459
rect 2108 422 2166 431
rect 2307 422 2365 431
rect 2495 422 2553 431
rect 2599 459 2657 468
rect 2787 459 2845 468
rect 2986 459 3044 468
rect 2599 431 3044 459
rect 2599 422 2657 431
rect 2787 422 2845 431
rect 2986 422 3044 431
rect 3396 459 3454 468
rect 3595 459 3653 468
rect 3783 459 3841 468
rect 3396 431 3841 459
rect 3396 422 3454 431
rect 3595 422 3653 431
rect 3783 422 3841 431
rect 3887 459 3945 468
rect 4075 459 4133 468
rect 4274 459 4332 468
rect 3887 431 4332 459
rect 3887 422 3945 431
rect 4075 422 4133 431
rect 4274 422 4332 431
rect 4684 459 4742 468
rect 4883 459 4941 468
rect 5071 459 5129 468
rect 4684 431 5129 459
rect 4684 422 4742 431
rect 4883 422 4941 431
rect 5071 422 5129 431
<< labels >>
rlabel locali s 19 211 183 265 6 D[0]
port 1 nsew signal input
rlabel locali s 1105 211 1269 265 6 D[1]
port 2 nsew signal input
rlabel locali s 1307 211 1471 265 6 D[2]
port 3 nsew signal input
rlabel locali s 2393 211 2557 265 6 D[3]
port 4 nsew signal input
rlabel locali s 2595 211 2759 265 6 D[4]
port 5 nsew signal input
rlabel locali s 3681 211 3845 265 6 D[5]
port 6 nsew signal input
rlabel locali s 3883 211 4047 265 6 D[6]
port 7 nsew signal input
rlabel locali s 4969 211 5133 265 6 D[7]
port 8 nsew signal input
rlabel locali s 19 823 183 877 6 D[8]
port 9 nsew signal input
rlabel locali s 1105 823 1269 877 6 D[9]
port 10 nsew signal input
rlabel locali s 1307 823 1471 877 6 D[10]
port 11 nsew signal input
rlabel locali s 2393 823 2557 877 6 D[11]
port 12 nsew signal input
rlabel locali s 2595 823 2759 877 6 D[12]
port 13 nsew signal input
rlabel locali s 3681 823 3845 877 6 D[13]
port 14 nsew signal input
rlabel locali s 3883 823 4047 877 6 D[14]
port 15 nsew signal input
rlabel locali s 4969 823 5133 877 6 D[15]
port 16 nsew signal input
rlabel locali s 558 205 625 259 6 S[0]
port 17 nsew signal input
rlabel locali s 663 205 730 259 6 S[1]
port 18 nsew signal input
rlabel locali s 1846 205 1913 259 6 S[2]
port 19 nsew signal input
rlabel locali s 1951 205 2018 259 6 S[3]
port 20 nsew signal input
rlabel locali s 3134 205 3201 259 6 S[4]
port 21 nsew signal input
rlabel locali s 3239 205 3306 259 6 S[5]
port 22 nsew signal input
rlabel locali s 4422 205 4489 259 6 S[6]
port 23 nsew signal input
rlabel locali s 4527 205 4594 259 6 S[7]
port 24 nsew signal input
rlabel locali s 558 829 625 883 6 S[8]
port 25 nsew signal input
rlabel locali s 663 829 730 883 6 S[9]
port 26 nsew signal input
rlabel locali s 1846 829 1913 883 6 S[10]
port 27 nsew signal input
rlabel locali s 1951 829 2018 883 6 S[11]
port 28 nsew signal input
rlabel locali s 3134 829 3201 883 6 S[12]
port 29 nsew signal input
rlabel locali s 3239 829 3306 883 6 S[13]
port 30 nsew signal input
rlabel locali s 4422 829 4489 883 6 S[14]
port 31 nsew signal input
rlabel locali s 4527 829 4594 883 6 S[15]
port 32 nsew signal input
rlabel viali s 305 697 339 731 6 Z
port 33 nsew signal output
rlabel viali s 305 357 339 391 6 Z
port 33 nsew signal output
rlabel locali s 317 737 351 911 6 Z
port 33 nsew signal output
rlabel locali s 317 425 351 663 6 Z
port 33 nsew signal output
rlabel locali s 317 177 351 351 6 Z
port 33 nsew signal output
rlabel locali s 301 911 367 969 6 Z
port 33 nsew signal output
rlabel locali s 301 119 367 177 6 Z
port 33 nsew signal output
rlabel locali s 293 663 379 737 6 Z
port 33 nsew signal output
rlabel locali s 293 351 379 425 6 Z
port 33 nsew signal output
rlabel metal1 s 4801 728 4859 737 6 Z
port 33 nsew signal output
rlabel metal1 s 4801 691 4859 700 6 Z
port 33 nsew signal output
rlabel metal1 s 4801 388 4859 397 6 Z
port 33 nsew signal output
rlabel metal1 s 4801 351 4859 360 6 Z
port 33 nsew signal output
rlabel metal1 s 4157 728 4215 737 6 Z
port 33 nsew signal output
rlabel metal1 s 4157 691 4215 700 6 Z
port 33 nsew signal output
rlabel metal1 s 4157 388 4215 397 6 Z
port 33 nsew signal output
rlabel metal1 s 4157 351 4215 360 6 Z
port 33 nsew signal output
rlabel metal1 s 3513 728 3571 737 6 Z
port 33 nsew signal output
rlabel metal1 s 3513 691 3571 700 6 Z
port 33 nsew signal output
rlabel metal1 s 3513 388 3571 397 6 Z
port 33 nsew signal output
rlabel metal1 s 3513 351 3571 360 6 Z
port 33 nsew signal output
rlabel metal1 s 2869 728 2927 737 6 Z
port 33 nsew signal output
rlabel metal1 s 2869 691 2927 700 6 Z
port 33 nsew signal output
rlabel metal1 s 2869 388 2927 397 6 Z
port 33 nsew signal output
rlabel metal1 s 2869 351 2927 360 6 Z
port 33 nsew signal output
rlabel metal1 s 2225 728 2283 737 6 Z
port 33 nsew signal output
rlabel metal1 s 2225 691 2283 700 6 Z
port 33 nsew signal output
rlabel metal1 s 2225 388 2283 397 6 Z
port 33 nsew signal output
rlabel metal1 s 2225 351 2283 360 6 Z
port 33 nsew signal output
rlabel metal1 s 1581 728 1639 737 6 Z
port 33 nsew signal output
rlabel metal1 s 1581 691 1639 700 6 Z
port 33 nsew signal output
rlabel metal1 s 1581 388 1639 397 6 Z
port 33 nsew signal output
rlabel metal1 s 1581 351 1639 360 6 Z
port 33 nsew signal output
rlabel metal1 s 937 728 995 737 6 Z
port 33 nsew signal output
rlabel metal1 s 937 691 995 700 6 Z
port 33 nsew signal output
rlabel metal1 s 937 388 995 397 6 Z
port 33 nsew signal output
rlabel metal1 s 937 351 995 360 6 Z
port 33 nsew signal output
rlabel metal1 s 293 728 351 737 6 Z
port 33 nsew signal output
rlabel metal1 s 293 700 4859 728 6 Z
port 33 nsew signal output
rlabel metal1 s 293 691 351 700 6 Z
port 33 nsew signal output
rlabel metal1 s 293 388 351 397 6 Z
port 33 nsew signal output
rlabel metal1 s 293 360 4859 388 6 Z
port 33 nsew signal output
rlabel metal1 s 293 351 351 360 6 Z
port 33 nsew signal output
rlabel viali s 5089 -17 5123 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 4997 -17 5031 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 4905 -17 4939 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 4813 -17 4847 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 4721 -17 4755 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 4629 -17 4663 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 4537 -17 4571 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 4445 -17 4479 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 4353 -17 4387 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 4261 -17 4295 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 4169 -17 4203 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 4077 -17 4111 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 3985 -17 4019 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 3893 -17 3927 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 3801 -17 3835 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 3709 -17 3743 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 3617 -17 3651 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 3525 -17 3559 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 3433 -17 3467 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 3341 -17 3375 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 3249 -17 3283 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 3157 -17 3191 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 3065 -17 3099 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 2973 -17 3007 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 2881 -17 2915 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 2789 -17 2823 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 2697 -17 2731 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 2605 -17 2639 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 2513 -17 2547 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 2421 -17 2455 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 2329 -17 2363 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 2237 -17 2271 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 2145 -17 2179 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 2053 -17 2087 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 1961 -17 1995 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 1869 -17 1903 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 1777 -17 1811 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 1685 -17 1719 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 1593 -17 1627 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 1501 -17 1535 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 1409 -17 1443 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 1317 -17 1351 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 1225 -17 1259 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 1133 -17 1167 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 1041 -17 1075 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 949 -17 983 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 857 -17 891 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 765 -17 799 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 673 -17 707 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 581 -17 615 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 489 -17 523 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 397 -17 431 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 305 -17 339 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 213 -17 247 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 121 -17 155 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 29 -17 63 17 8 VGND
port 34 nsew ground bidirectional
rlabel locali s 4980 17 5023 109 6 VGND
port 34 nsew ground bidirectional
rlabel locali s 4483 17 4533 132 6 VGND
port 34 nsew ground bidirectional
rlabel locali s 3993 17 4036 109 6 VGND
port 34 nsew ground bidirectional
rlabel locali s 3692 17 3735 109 6 VGND
port 34 nsew ground bidirectional
rlabel locali s 3195 17 3245 132 6 VGND
port 34 nsew ground bidirectional
rlabel locali s 2705 17 2748 109 6 VGND
port 34 nsew ground bidirectional
rlabel locali s 2404 17 2447 109 6 VGND
port 34 nsew ground bidirectional
rlabel locali s 1907 17 1957 132 6 VGND
port 34 nsew ground bidirectional
rlabel locali s 1417 17 1460 109 6 VGND
port 34 nsew ground bidirectional
rlabel locali s 1116 17 1159 109 6 VGND
port 34 nsew ground bidirectional
rlabel locali s 619 17 669 132 6 VGND
port 34 nsew ground bidirectional
rlabel locali s 129 17 172 109 6 VGND
port 34 nsew ground bidirectional
rlabel locali s 0 -17 5152 17 8 VGND
port 34 nsew ground bidirectional
rlabel viali s 5089 1071 5123 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 4997 1071 5031 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 4905 1071 4939 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 4813 1071 4847 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 4721 1071 4755 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 4629 1071 4663 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 4537 1071 4571 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 4445 1071 4479 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 4353 1071 4387 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 4261 1071 4295 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 4169 1071 4203 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 4077 1071 4111 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 3985 1071 4019 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 3893 1071 3927 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 3801 1071 3835 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 3709 1071 3743 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 3617 1071 3651 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 3525 1071 3559 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 3433 1071 3467 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 3341 1071 3375 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 3249 1071 3283 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 3157 1071 3191 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 3065 1071 3099 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 2973 1071 3007 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 2881 1071 2915 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 2789 1071 2823 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 2697 1071 2731 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 2605 1071 2639 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 2513 1071 2547 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 2421 1071 2455 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 2329 1071 2363 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 2237 1071 2271 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 2145 1071 2179 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 2053 1071 2087 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 1961 1071 1995 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 1869 1071 1903 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 1777 1071 1811 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 1685 1071 1719 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 1593 1071 1627 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 1501 1071 1535 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 1409 1071 1443 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 1317 1071 1351 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 1225 1071 1259 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 1133 1071 1167 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 1041 1071 1075 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 949 1071 983 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 857 1071 891 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 765 1071 799 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 673 1071 707 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 581 1071 615 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 489 1071 523 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 397 1071 431 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 305 1071 339 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 213 1071 247 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 121 1071 155 1105 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 29 1071 63 1105 6 VGND
port 34 nsew ground bidirectional
rlabel locali s 4980 979 5023 1071 6 VGND
port 34 nsew ground bidirectional
rlabel locali s 4483 956 4533 1071 6 VGND
port 34 nsew ground bidirectional
rlabel locali s 3993 979 4036 1071 6 VGND
port 34 nsew ground bidirectional
rlabel locali s 3692 979 3735 1071 6 VGND
port 34 nsew ground bidirectional
rlabel locali s 3195 956 3245 1071 6 VGND
port 34 nsew ground bidirectional
rlabel locali s 2705 979 2748 1071 6 VGND
port 34 nsew ground bidirectional
rlabel locali s 2404 979 2447 1071 6 VGND
port 34 nsew ground bidirectional
rlabel locali s 1907 956 1957 1071 6 VGND
port 34 nsew ground bidirectional
rlabel locali s 1417 979 1460 1071 6 VGND
port 34 nsew ground bidirectional
rlabel locali s 1116 979 1159 1071 6 VGND
port 34 nsew ground bidirectional
rlabel locali s 619 956 669 1071 6 VGND
port 34 nsew ground bidirectional
rlabel locali s 129 979 172 1071 6 VGND
port 34 nsew ground bidirectional
rlabel locali s 0 1071 5152 1105 6 VGND
port 34 nsew ground bidirectional
rlabel metal1 s 0 -48 5152 48 8 VGND
port 34 nsew ground bidirectional
rlabel metal1 s 0 1040 5152 1136 6 VGND
port 34 nsew ground bidirectional
rlabel viali s 213 527 247 561 6 VPWR
port 35 nsew power bidirectional
rlabel viali s 121 527 155 561 6 VPWR
port 35 nsew power bidirectional
rlabel viali s 29 527 63 561 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 119 561 179 667 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 119 421 179 527 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 113 667 179 721 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 113 367 179 421 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 0 527 283 561 6 VPWR
port 35 nsew power bidirectional
rlabel viali s 2789 527 2823 561 6 VPWR
port 35 nsew power bidirectional
rlabel viali s 2697 527 2731 561 6 VPWR
port 35 nsew power bidirectional
rlabel viali s 2605 527 2639 561 6 VPWR
port 35 nsew power bidirectional
rlabel viali s 2513 527 2547 561 6 VPWR
port 35 nsew power bidirectional
rlabel viali s 2421 527 2455 561 6 VPWR
port 35 nsew power bidirectional
rlabel viali s 2329 527 2363 561 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 2695 561 2755 667 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 2695 421 2755 527 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 2689 667 2755 721 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 2689 367 2755 421 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 2397 667 2463 721 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 2397 561 2457 667 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 2397 421 2457 527 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 2397 367 2463 421 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 2293 527 2859 561 6 VPWR
port 35 nsew power bidirectional
rlabel viali s 4077 527 4111 561 6 VPWR
port 35 nsew power bidirectional
rlabel viali s 3985 527 4019 561 6 VPWR
port 35 nsew power bidirectional
rlabel viali s 3893 527 3927 561 6 VPWR
port 35 nsew power bidirectional
rlabel viali s 3801 527 3835 561 6 VPWR
port 35 nsew power bidirectional
rlabel viali s 3709 527 3743 561 6 VPWR
port 35 nsew power bidirectional
rlabel viali s 3617 527 3651 561 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 3983 561 4043 667 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 3983 421 4043 527 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 3977 667 4043 721 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 3977 367 4043 421 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 3685 667 3751 721 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 3685 561 3745 667 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 3685 421 3745 527 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 3685 367 3751 421 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 3581 527 4147 561 6 VPWR
port 35 nsew power bidirectional
rlabel viali s 5089 527 5123 561 6 VPWR
port 35 nsew power bidirectional
rlabel viali s 4997 527 5031 561 6 VPWR
port 35 nsew power bidirectional
rlabel viali s 4905 527 4939 561 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 4973 667 5039 721 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 4973 561 5033 667 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 4973 421 5033 527 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 4973 367 5039 421 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 4869 527 5152 561 6 VPWR
port 35 nsew power bidirectional
rlabel viali s 1501 527 1535 561 6 VPWR
port 35 nsew power bidirectional
rlabel viali s 1409 527 1443 561 6 VPWR
port 35 nsew power bidirectional
rlabel viali s 1317 527 1351 561 6 VPWR
port 35 nsew power bidirectional
rlabel viali s 1225 527 1259 561 6 VPWR
port 35 nsew power bidirectional
rlabel viali s 1133 527 1167 561 6 VPWR
port 35 nsew power bidirectional
rlabel viali s 1041 527 1075 561 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 1407 561 1467 667 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 1407 421 1467 527 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 1401 667 1467 721 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 1401 367 1467 421 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 1109 667 1175 721 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 1109 561 1169 667 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 1109 421 1169 527 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 1109 367 1175 421 6 VPWR
port 35 nsew power bidirectional
rlabel locali s 1005 527 1571 561 6 VPWR
port 35 nsew power bidirectional
rlabel metal1 s 0 496 5152 592 6 VPWR
port 35 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 5152 1088
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3118222
string GDS_START 3026152
<< end >>
