magic
tech sky130A
magscale 1 2
timestamp 1601050058
<< locali >>
rect 1483 343 1547 395
rect 1595 343 1661 417
rect 1763 343 1829 417
rect 24 199 347 265
rect 387 199 710 265
rect 761 199 1084 265
rect 1134 199 1371 326
rect 1483 309 1829 343
rect 1483 161 1547 309
rect 1595 306 1661 309
rect 1587 199 1906 265
rect 795 127 1897 161
rect 1315 51 1349 127
rect 1483 51 1517 127
rect 1695 51 1729 127
rect 1863 51 1897 127
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 19 315 85 527
rect 119 333 153 493
rect 187 383 253 527
rect 287 333 321 493
rect 355 383 421 527
rect 455 333 489 493
rect 523 383 589 527
rect 623 333 657 493
rect 691 383 757 527
rect 791 333 825 493
rect 859 383 925 527
rect 959 417 993 493
rect 1027 451 1093 527
rect 1131 451 1913 485
rect 959 383 1449 417
rect 959 333 993 383
rect 119 299 993 333
rect 1863 367 1913 451
rect 35 127 757 161
rect 35 51 69 127
rect 103 17 169 93
rect 203 51 237 127
rect 271 17 337 93
rect 371 51 405 127
rect 439 59 1113 93
rect 1215 17 1281 93
rect 1383 17 1449 93
rect 1595 17 1661 93
rect 1763 17 1829 93
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< labels >>
rlabel locali s 761 199 1084 265 6 A1
port 1 nsew signal input
rlabel locali s 387 199 710 265 6 A2
port 2 nsew signal input
rlabel locali s 24 199 347 265 6 A3
port 3 nsew signal input
rlabel locali s 1134 199 1371 326 6 B1
port 4 nsew signal input
rlabel locali s 1587 199 1906 265 6 C1
port 5 nsew signal input
rlabel locali s 1863 51 1897 127 6 Y
port 6 nsew signal output
rlabel locali s 1763 343 1829 417 6 Y
port 6 nsew signal output
rlabel locali s 1695 51 1729 127 6 Y
port 6 nsew signal output
rlabel locali s 1595 343 1661 417 6 Y
port 6 nsew signal output
rlabel locali s 1595 306 1661 309 6 Y
port 6 nsew signal output
rlabel locali s 1483 343 1547 395 6 Y
port 6 nsew signal output
rlabel locali s 1483 309 1829 343 6 Y
port 6 nsew signal output
rlabel locali s 1483 161 1547 309 6 Y
port 6 nsew signal output
rlabel locali s 1483 51 1517 127 6 Y
port 6 nsew signal output
rlabel locali s 1315 51 1349 127 6 Y
port 6 nsew signal output
rlabel locali s 795 127 1897 161 6 Y
port 6 nsew signal output
rlabel metal1 s 0 -48 1932 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1932 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1932 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3584904
string GDS_START 3569358
<< end >>
