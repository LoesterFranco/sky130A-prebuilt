magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 2706 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 89 47 119 131
rect 171 47 201 131
rect 265 47 295 131
rect 349 47 379 131
rect 563 47 593 131
rect 761 47 791 131
rect 855 47 885 131
rect 1053 47 1083 131
rect 1147 47 1177 131
rect 1229 47 1259 131
rect 1437 47 1467 131
rect 1509 47 1539 131
rect 1615 47 1645 175
rect 1803 47 1833 175
rect 1925 47 1955 131
rect 1997 47 2027 131
rect 2103 47 2133 131
rect 2221 47 2251 131
rect 2433 47 2463 131
rect 2548 47 2578 177
<< pmoshvt >>
rect 81 369 117 497
rect 175 369 211 497
rect 257 369 293 497
rect 351 369 387 497
rect 549 369 585 497
rect 747 369 783 497
rect 841 369 877 497
rect 1039 413 1075 497
rect 1133 413 1169 497
rect 1245 413 1281 497
rect 1383 413 1419 497
rect 1501 413 1537 497
rect 1607 329 1643 497
rect 1689 329 1725 497
rect 1805 413 1841 497
rect 1923 413 1959 497
rect 2034 413 2070 497
rect 2237 413 2273 497
rect 2435 369 2471 497
rect 2540 297 2576 497
<< ndiff >>
rect 1554 131 1615 175
rect 27 103 89 131
rect 27 69 35 103
rect 69 69 89 103
rect 27 47 89 69
rect 119 47 171 131
rect 201 93 265 131
rect 201 59 211 93
rect 245 59 265 93
rect 201 47 265 59
rect 295 47 349 131
rect 379 93 447 131
rect 379 59 405 93
rect 439 59 447 93
rect 379 47 447 59
rect 501 105 563 131
rect 501 71 509 105
rect 543 71 563 105
rect 501 47 563 71
rect 593 93 645 131
rect 593 59 603 93
rect 637 59 645 93
rect 593 47 645 59
rect 699 105 761 131
rect 699 71 707 105
rect 741 71 761 105
rect 699 47 761 71
rect 791 89 855 131
rect 791 55 801 89
rect 835 55 855 89
rect 791 47 855 55
rect 885 101 937 131
rect 885 67 895 101
rect 929 67 937 101
rect 885 47 937 67
rect 991 101 1053 131
rect 991 67 999 101
rect 1033 67 1053 101
rect 991 47 1053 67
rect 1083 101 1147 131
rect 1083 67 1093 101
rect 1127 67 1147 101
rect 1083 47 1147 67
rect 1177 47 1229 131
rect 1259 93 1311 131
rect 1259 59 1269 93
rect 1303 59 1311 93
rect 1259 47 1311 59
rect 1365 119 1437 131
rect 1365 85 1373 119
rect 1407 85 1437 119
rect 1365 47 1437 85
rect 1467 47 1509 131
rect 1539 89 1615 131
rect 1539 55 1561 89
rect 1595 55 1615 89
rect 1539 47 1615 55
rect 1645 47 1803 175
rect 1833 131 1883 175
rect 2488 131 2548 177
rect 1833 89 1925 131
rect 1833 55 1843 89
rect 1877 55 1925 89
rect 1833 47 1925 55
rect 1955 47 1997 131
rect 2027 47 2103 131
rect 2133 89 2221 131
rect 2133 55 2167 89
rect 2201 55 2221 89
rect 2133 47 2221 55
rect 2251 101 2327 131
rect 2251 67 2285 101
rect 2319 67 2327 101
rect 2251 47 2327 67
rect 2381 102 2433 131
rect 2381 68 2389 102
rect 2423 68 2433 102
rect 2381 47 2433 68
rect 2463 89 2548 131
rect 2463 55 2488 89
rect 2522 55 2548 89
rect 2463 47 2548 55
rect 2578 105 2630 177
rect 2578 71 2588 105
rect 2622 71 2630 105
rect 2578 47 2630 71
<< pdiff >>
rect 27 431 81 497
rect 27 397 35 431
rect 69 397 81 431
rect 27 369 81 397
rect 117 489 175 497
rect 117 455 129 489
rect 163 455 175 489
rect 117 369 175 455
rect 211 369 257 497
rect 293 411 351 497
rect 293 377 305 411
rect 339 377 351 411
rect 293 369 351 377
rect 387 485 441 497
rect 387 451 399 485
rect 433 451 441 485
rect 387 369 441 451
rect 495 415 549 497
rect 495 381 503 415
rect 537 381 549 415
rect 495 369 549 381
rect 585 485 639 497
rect 585 451 597 485
rect 631 451 639 485
rect 585 369 639 451
rect 693 449 747 497
rect 693 415 701 449
rect 735 415 747 449
rect 693 369 747 415
rect 783 489 841 497
rect 783 455 795 489
rect 829 455 841 489
rect 783 369 841 455
rect 877 477 931 497
rect 877 443 889 477
rect 923 443 931 477
rect 877 369 931 443
rect 985 477 1039 497
rect 985 443 993 477
rect 1027 443 1039 477
rect 985 413 1039 443
rect 1075 477 1133 497
rect 1075 443 1087 477
rect 1121 443 1133 477
rect 1075 413 1133 443
rect 1169 413 1245 497
rect 1281 489 1383 497
rect 1281 455 1305 489
rect 1339 455 1383 489
rect 1281 413 1383 455
rect 1419 474 1501 497
rect 1419 440 1436 474
rect 1470 440 1501 474
rect 1419 413 1501 440
rect 1537 489 1607 497
rect 1537 455 1558 489
rect 1592 455 1607 489
rect 1537 413 1607 455
rect 1555 329 1607 413
rect 1643 329 1689 497
rect 1725 475 1805 497
rect 1725 441 1759 475
rect 1793 441 1805 475
rect 1725 413 1805 441
rect 1841 413 1923 497
rect 1959 489 2034 497
rect 1959 455 1988 489
rect 2022 455 2034 489
rect 1959 413 2034 455
rect 2070 474 2124 497
rect 2070 440 2082 474
rect 2116 440 2124 474
rect 2070 413 2124 440
rect 2183 485 2237 497
rect 2183 451 2191 485
rect 2225 451 2237 485
rect 2183 413 2237 451
rect 2273 474 2327 497
rect 2273 440 2285 474
rect 2319 440 2327 474
rect 2273 413 2327 440
rect 2381 483 2435 497
rect 2381 449 2389 483
rect 2423 449 2435 483
rect 2381 415 2435 449
rect 1725 329 1777 413
rect 2381 381 2389 415
rect 2423 381 2435 415
rect 2381 369 2435 381
rect 2471 489 2540 497
rect 2471 455 2488 489
rect 2522 455 2540 489
rect 2471 421 2540 455
rect 2471 387 2488 421
rect 2522 387 2540 421
rect 2471 369 2540 387
rect 2488 297 2540 369
rect 2576 474 2630 497
rect 2576 440 2588 474
rect 2622 440 2630 474
rect 2576 297 2630 440
<< ndiffc >>
rect 35 69 69 103
rect 211 59 245 93
rect 405 59 439 93
rect 509 71 543 105
rect 603 59 637 93
rect 707 71 741 105
rect 801 55 835 89
rect 895 67 929 101
rect 999 67 1033 101
rect 1093 67 1127 101
rect 1269 59 1303 93
rect 1373 85 1407 119
rect 1561 55 1595 89
rect 1843 55 1877 89
rect 2167 55 2201 89
rect 2285 67 2319 101
rect 2389 68 2423 102
rect 2488 55 2522 89
rect 2588 71 2622 105
<< pdiffc >>
rect 35 397 69 431
rect 129 455 163 489
rect 305 377 339 411
rect 399 451 433 485
rect 503 381 537 415
rect 597 451 631 485
rect 701 415 735 449
rect 795 455 829 489
rect 889 443 923 477
rect 993 443 1027 477
rect 1087 443 1121 477
rect 1305 455 1339 489
rect 1436 440 1470 474
rect 1558 455 1592 489
rect 1759 441 1793 475
rect 1988 455 2022 489
rect 2082 440 2116 474
rect 2191 451 2225 485
rect 2285 440 2319 474
rect 2389 449 2423 483
rect 2389 381 2423 415
rect 2488 455 2522 489
rect 2488 387 2522 421
rect 2588 440 2622 474
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 257 497 293 523
rect 351 497 387 523
rect 549 497 585 523
rect 747 497 783 523
rect 841 497 877 523
rect 1039 497 1075 523
rect 1133 497 1169 523
rect 1245 497 1281 523
rect 1383 497 1419 523
rect 1501 497 1537 523
rect 1607 497 1643 523
rect 1689 497 1725 523
rect 1805 497 1841 523
rect 1923 497 1959 523
rect 2034 497 2070 523
rect 2237 497 2273 523
rect 2435 497 2471 523
rect 2540 497 2576 523
rect 1039 398 1075 413
rect 1133 398 1169 413
rect 1245 398 1281 413
rect 1383 398 1419 413
rect 1501 398 1537 413
rect 81 354 117 369
rect 175 354 211 369
rect 257 354 293 369
rect 351 354 387 369
rect 549 354 585 369
rect 747 354 783 369
rect 841 354 877 369
rect 978 368 1077 398
rect 1131 381 1171 398
rect 1243 381 1283 398
rect 48 324 119 354
rect 48 265 78 324
rect 173 283 213 354
rect 21 249 78 265
rect 21 215 34 249
rect 68 215 78 249
rect 130 267 213 283
rect 130 233 140 267
rect 174 253 213 267
rect 174 233 201 253
rect 130 217 201 233
rect 255 219 295 354
rect 349 265 389 354
rect 547 265 587 354
rect 733 324 785 354
rect 733 284 763 324
rect 839 284 879 354
rect 978 284 1008 368
rect 1119 365 1183 381
rect 1119 331 1129 365
rect 1163 331 1183 365
rect 1119 315 1183 331
rect 1243 365 1329 381
rect 1243 331 1285 365
rect 1319 331 1329 365
rect 1243 315 1329 331
rect 709 268 763 284
rect 349 249 478 265
rect 21 199 78 215
rect 48 176 78 199
rect 48 146 119 176
rect 89 131 119 146
rect 171 131 201 217
rect 243 203 307 219
rect 243 169 253 203
rect 287 169 307 203
rect 243 153 307 169
rect 349 215 413 249
rect 447 215 478 249
rect 349 199 478 215
rect 520 249 593 265
rect 520 215 530 249
rect 564 215 593 249
rect 709 234 719 268
rect 753 234 763 268
rect 709 218 763 234
rect 815 268 879 284
rect 815 234 825 268
rect 859 234 879 268
rect 815 218 879 234
rect 924 268 1008 284
rect 924 234 934 268
rect 968 248 1008 268
rect 968 234 1177 248
rect 924 218 1177 234
rect 520 199 593 215
rect 265 131 295 153
rect 349 131 379 199
rect 563 131 593 199
rect 733 176 763 218
rect 842 176 879 218
rect 733 146 791 176
rect 842 146 1083 176
rect 761 131 791 146
rect 855 131 885 146
rect 1053 131 1083 146
rect 1147 131 1177 218
rect 1243 213 1283 315
rect 1381 273 1421 398
rect 1499 369 1539 398
rect 1463 353 1539 369
rect 1463 319 1473 353
rect 1507 319 1539 353
rect 1805 398 1841 413
rect 1923 398 1959 413
rect 2034 398 2070 413
rect 2237 398 2273 413
rect 1803 381 1843 398
rect 1803 365 1868 381
rect 1803 331 1824 365
rect 1858 331 1868 365
rect 1463 303 1539 319
rect 1607 314 1643 329
rect 1689 314 1725 329
rect 1803 315 1868 331
rect 1921 325 1961 398
rect 2032 397 2072 398
rect 2032 367 2133 397
rect 2079 343 2133 367
rect 2235 365 2275 398
rect 1345 263 1421 273
rect 1345 229 1361 263
rect 1395 229 1421 263
rect 1345 219 1421 229
rect 1229 203 1295 213
rect 1229 169 1245 203
rect 1279 169 1295 203
rect 1229 159 1295 169
rect 1381 176 1421 219
rect 1229 131 1259 159
rect 1381 146 1467 176
rect 1437 131 1467 146
rect 1509 131 1539 303
rect 1605 265 1645 314
rect 1591 249 1645 265
rect 1591 215 1601 249
rect 1635 215 1645 249
rect 1591 199 1645 215
rect 1687 265 1727 314
rect 1687 249 1741 265
rect 1687 215 1697 249
rect 1731 215 1741 249
rect 1687 199 1741 215
rect 1615 175 1645 199
rect 1803 175 1833 315
rect 1921 295 2037 325
rect 1901 235 1955 251
rect 1901 201 1911 235
rect 1945 201 1955 235
rect 1901 185 1955 201
rect 1925 131 1955 185
rect 1997 237 2037 295
rect 2079 309 2089 343
rect 2123 309 2133 343
rect 2175 355 2275 365
rect 2175 321 2191 355
rect 2225 321 2275 355
rect 2435 354 2471 369
rect 2175 311 2275 321
rect 2079 293 2133 309
rect 1997 221 2061 237
rect 1997 187 2007 221
rect 2041 187 2061 221
rect 1997 171 2061 187
rect 1997 131 2027 171
rect 2103 131 2133 293
rect 2187 271 2275 311
rect 2433 307 2473 354
rect 2433 271 2463 307
rect 2540 282 2576 297
rect 2187 241 2463 271
rect 2538 265 2578 282
rect 2187 203 2251 241
rect 2187 169 2197 203
rect 2231 169 2251 203
rect 2187 153 2251 169
rect 2221 131 2251 153
rect 2433 131 2463 241
rect 2505 249 2578 265
rect 2505 215 2515 249
rect 2549 215 2578 249
rect 2505 199 2578 215
rect 2548 177 2578 199
rect 89 21 119 47
rect 171 21 201 47
rect 265 21 295 47
rect 349 21 379 47
rect 563 21 593 47
rect 761 21 791 47
rect 855 21 885 47
rect 1053 21 1083 47
rect 1147 21 1177 47
rect 1229 21 1259 47
rect 1437 21 1467 47
rect 1509 21 1539 47
rect 1615 21 1645 47
rect 1803 21 1833 47
rect 1925 21 1955 47
rect 1997 21 2027 47
rect 2103 21 2133 47
rect 2221 21 2251 47
rect 2433 21 2463 47
rect 2548 21 2578 47
<< polycont >>
rect 34 215 68 249
rect 140 233 174 267
rect 1129 331 1163 365
rect 1285 331 1319 365
rect 253 169 287 203
rect 413 215 447 249
rect 530 215 564 249
rect 719 234 753 268
rect 825 234 859 268
rect 934 234 968 268
rect 1473 319 1507 353
rect 1824 331 1858 365
rect 1361 229 1395 263
rect 1245 169 1279 203
rect 1601 215 1635 249
rect 1697 215 1731 249
rect 1911 201 1945 235
rect 2089 309 2123 343
rect 2191 321 2225 355
rect 2007 187 2041 221
rect 2197 169 2231 203
rect 2515 215 2549 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2668 561
rect 17 431 69 493
rect 103 489 167 527
rect 103 455 129 489
rect 163 455 167 489
rect 103 439 167 455
rect 211 485 449 493
rect 211 451 399 485
rect 433 451 449 485
rect 17 397 35 431
rect 211 405 245 451
rect 494 417 544 493
rect 588 485 647 527
rect 588 451 597 485
rect 631 451 647 485
rect 769 489 845 527
rect 588 428 647 451
rect 701 449 735 465
rect 769 455 795 489
rect 829 455 845 489
rect 889 477 958 493
rect 69 397 245 405
rect 17 369 245 397
rect 279 411 369 417
rect 279 377 305 411
rect 339 377 369 411
rect 279 369 369 377
rect 17 249 68 335
rect 17 215 34 249
rect 17 153 68 215
rect 108 267 174 335
rect 108 255 140 267
rect 108 221 128 255
rect 162 221 174 233
rect 108 153 174 221
rect 208 203 297 335
rect 208 169 253 203
rect 287 169 297 203
rect 208 153 297 169
rect 331 323 369 369
rect 331 289 335 323
rect 331 119 369 289
rect 413 415 544 417
rect 413 381 503 415
rect 537 381 544 415
rect 413 354 544 381
rect 923 443 958 477
rect 889 427 958 443
rect 701 400 735 415
rect 701 391 859 400
rect 701 366 825 391
rect 807 357 825 366
rect 413 249 480 354
rect 447 215 480 249
rect 514 255 590 320
rect 514 221 529 255
rect 563 249 590 255
rect 514 215 530 221
rect 564 215 590 249
rect 631 268 763 330
rect 631 234 719 268
rect 753 234 763 268
rect 413 181 480 215
rect 631 211 763 234
rect 807 268 859 357
rect 807 234 825 268
rect 413 143 544 181
rect 807 177 859 234
rect 17 103 150 119
rect 17 69 35 103
rect 69 69 150 103
rect 17 17 150 69
rect 184 93 369 119
rect 184 59 211 93
rect 245 59 369 93
rect 184 51 369 59
rect 405 93 458 109
rect 439 59 458 93
rect 405 17 458 59
rect 492 105 544 143
rect 704 143 859 177
rect 895 284 958 427
rect 993 477 1036 493
rect 1027 443 1036 477
rect 993 323 1036 443
rect 1087 477 1241 493
rect 1121 443 1241 477
rect 1289 489 1366 527
rect 1289 455 1305 489
rect 1339 455 1366 489
rect 1431 474 1484 490
rect 1087 427 1241 443
rect 993 318 1002 323
rect 1155 365 1173 391
rect 1121 331 1129 357
rect 1163 331 1173 365
rect 1121 315 1173 331
rect 895 268 968 284
rect 895 254 934 268
rect 895 220 927 254
rect 961 220 968 234
rect 895 217 968 220
rect 492 71 509 105
rect 543 71 544 105
rect 492 51 544 71
rect 588 93 670 111
rect 588 59 603 93
rect 637 59 670 93
rect 588 17 670 59
rect 704 105 741 143
rect 704 71 707 105
rect 704 51 741 71
rect 785 89 851 109
rect 785 55 801 89
rect 835 55 851 89
rect 785 17 851 55
rect 895 101 937 217
rect 1002 156 1036 289
rect 1207 279 1241 427
rect 1431 440 1436 474
rect 1470 440 1484 474
rect 1431 421 1484 440
rect 1542 489 1725 527
rect 1542 455 1558 489
rect 1592 455 1725 489
rect 1542 425 1725 455
rect 1759 475 1938 492
rect 1793 441 1938 475
rect 1972 489 2038 527
rect 1972 455 1988 489
rect 2022 455 2038 489
rect 1972 447 2038 455
rect 2079 474 2119 490
rect 1759 425 1938 441
rect 1285 387 1484 421
rect 1904 413 1938 425
rect 2079 440 2082 474
rect 2116 440 2119 474
rect 2175 485 2251 527
rect 2175 451 2191 485
rect 2225 451 2251 485
rect 2175 447 2251 451
rect 2285 474 2337 493
rect 2079 413 2119 440
rect 2319 440 2337 474
rect 1285 365 1319 387
rect 1577 357 1642 391
rect 1676 357 1757 391
rect 1285 315 1319 331
rect 1438 319 1473 353
rect 1507 323 1543 353
rect 1577 334 1757 357
rect 1438 289 1487 319
rect 1521 289 1543 323
rect 929 67 937 101
rect 895 51 937 67
rect 971 101 1036 156
rect 971 67 999 101
rect 1033 67 1036 101
rect 971 51 1036 67
rect 1093 263 1395 279
rect 1093 245 1361 263
rect 1093 101 1178 245
rect 1581 255 1663 265
rect 1395 249 1663 255
rect 1395 229 1601 249
rect 1361 215 1601 229
rect 1635 215 1663 249
rect 1219 169 1245 203
rect 1279 169 1295 203
rect 1361 195 1663 215
rect 1697 249 1757 334
rect 1731 215 1757 249
rect 1791 365 1858 381
rect 1904 379 2251 413
rect 1791 331 1824 365
rect 2175 355 2251 379
rect 1791 255 1858 331
rect 1916 343 2139 345
rect 1916 323 2089 343
rect 1916 289 1925 323
rect 1959 309 2089 323
rect 2123 309 2139 343
rect 2175 321 2191 355
rect 2225 321 2251 355
rect 1959 289 1972 309
rect 1916 285 1972 289
rect 2285 273 2337 440
rect 1791 221 1810 255
rect 1844 221 1858 255
rect 1791 215 1858 221
rect 1904 235 1970 251
rect 1219 161 1295 169
rect 1697 181 1757 215
rect 1904 201 1911 235
rect 1945 201 1970 235
rect 1904 181 1970 201
rect 1219 127 1407 161
rect 1127 67 1178 101
rect 1357 119 1407 127
rect 1093 51 1178 67
rect 1212 59 1269 93
rect 1303 59 1319 93
rect 1212 17 1319 59
rect 1357 85 1373 119
rect 1357 51 1407 85
rect 1451 89 1663 161
rect 1697 144 1970 181
rect 2007 239 2337 273
rect 2007 221 2056 239
rect 2041 187 2056 221
rect 2007 171 2056 187
rect 2090 169 2197 203
rect 2231 169 2257 203
rect 2090 157 2257 169
rect 2090 109 2130 157
rect 2291 117 2337 239
rect 1451 55 1561 89
rect 1595 55 1663 89
rect 1805 89 2130 109
rect 1805 55 1843 89
rect 1877 55 2130 89
rect 2167 89 2217 109
rect 2201 55 2217 89
rect 1451 17 1663 55
rect 2167 17 2217 55
rect 2269 101 2337 117
rect 2269 67 2285 101
rect 2319 67 2337 101
rect 2269 51 2337 67
rect 2371 483 2439 493
rect 2371 449 2389 483
rect 2423 449 2439 483
rect 2371 415 2439 449
rect 2371 381 2389 415
rect 2423 381 2439 415
rect 2371 265 2439 381
rect 2487 489 2538 527
rect 2487 455 2488 489
rect 2522 455 2538 489
rect 2487 421 2538 455
rect 2487 387 2488 421
rect 2522 387 2538 421
rect 2487 369 2538 387
rect 2583 474 2648 490
rect 2583 440 2588 474
rect 2622 440 2648 474
rect 2371 249 2549 265
rect 2371 215 2515 249
rect 2371 199 2549 215
rect 2371 102 2423 199
rect 2371 68 2389 102
rect 2371 51 2423 68
rect 2457 89 2538 110
rect 2457 55 2488 89
rect 2522 55 2538 89
rect 2583 105 2648 440
rect 2583 71 2588 105
rect 2622 71 2648 105
rect 2583 55 2648 71
rect 2457 17 2538 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2668 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 128 233 140 255
rect 140 233 162 255
rect 128 221 162 233
rect 335 289 369 323
rect 825 357 859 391
rect 529 249 563 255
rect 529 221 530 249
rect 530 221 563 249
rect 1002 289 1036 323
rect 1121 365 1155 391
rect 1121 357 1129 365
rect 1129 357 1155 365
rect 927 234 934 254
rect 934 234 961 254
rect 927 220 961 234
rect 1642 357 1676 391
rect 1487 319 1507 323
rect 1507 319 1521 323
rect 1487 289 1521 319
rect 1925 289 1959 323
rect 1810 221 1844 255
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
<< metal1 >>
rect 0 561 2668 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2668 561
rect 0 496 2668 527
rect 813 391 881 397
rect 813 357 825 391
rect 859 388 881 391
rect 1109 391 1177 397
rect 1109 388 1121 391
rect 859 360 1121 388
rect 859 357 881 360
rect 813 351 881 357
rect 1109 357 1121 360
rect 1155 388 1177 391
rect 1630 391 1698 397
rect 1630 388 1642 391
rect 1155 360 1642 388
rect 1155 357 1177 360
rect 1109 351 1177 357
rect 1630 357 1642 360
rect 1676 357 1698 391
rect 1630 351 1698 357
rect 323 323 391 329
rect 323 289 335 323
rect 369 320 391 323
rect 990 323 1048 329
rect 990 320 1002 323
rect 369 292 1002 320
rect 369 289 391 292
rect 323 283 391 289
rect 990 289 1002 292
rect 1036 289 1048 323
rect 990 283 1048 289
rect 1475 323 1543 329
rect 1475 289 1487 323
rect 1521 320 1543 323
rect 1913 323 1981 329
rect 1913 320 1925 323
rect 1521 292 1925 320
rect 1521 289 1543 292
rect 1475 283 1543 289
rect 1913 289 1925 292
rect 1959 289 1981 323
rect 1913 283 1981 289
rect 116 255 174 261
rect 116 221 128 255
rect 162 252 174 255
rect 517 255 575 261
rect 517 252 529 255
rect 162 224 529 252
rect 162 221 174 224
rect 116 215 174 221
rect 517 221 529 224
rect 563 221 575 255
rect 517 215 575 221
rect 915 254 973 260
rect 915 220 927 254
rect 961 252 973 254
rect 1788 255 1866 261
rect 1788 252 1810 255
rect 961 224 1810 252
rect 961 220 973 224
rect 915 214 973 220
rect 1788 221 1810 224
rect 1844 221 1866 255
rect 1788 215 1866 221
rect 0 17 2668 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2668 17
rect 0 -48 2668 -17
<< labels >>
flabel comment s 1263 286 1263 286 0 FreeSans 200 0 0 0 no_jumper_check
rlabel comment s 0 0 0 0 4 sdfstp_4
flabel comment s 2233 287 2233 287 0 FreeSans 200 0 0 0 no_jumper_check
flabel metal1 s 121 221 155 255 0 FreeSans 200 0 0 0 SCE
port 4 nsew
flabel metal1 s 1501 289 1535 323 0 FreeSans 200 0 0 0 SET_B
port 5 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew
flabel corelocali s 673 221 707 255 0 FreeSans 200 0 0 0 CLK
port 1 nsew
flabel corelocali s 213 153 247 187 0 FreeSans 200 0 0 0 D
port 2 nsew
flabel corelocali s 29 289 63 323 0 FreeSans 200 0 0 0 SCD
port 3 nsew
flabel corelocali s 213 289 247 323 0 FreeSans 200 0 0 0 D
port 2 nsew
flabel corelocali s 29 153 63 187 0 FreeSans 200 0 0 0 SCD
port 3 nsew
flabel corelocali s 2607 357 2641 391 0 FreeSans 200 0 0 0 Q
port 10 nsew
flabel corelocali s 2607 425 2641 459 0 FreeSans 200 0 0 0 Q
port 10 nsew
flabel corelocali s 2607 221 2641 255 0 FreeSans 200 0 0 0 Q
port 10 nsew
flabel corelocali s 2607 153 2641 187 0 FreeSans 200 0 0 0 Q
port 10 nsew
flabel corelocali s 2607 85 2641 119 0 FreeSans 200 0 0 0 Q
port 10 nsew
flabel corelocali s 2607 289 2641 323 0 FreeSans 200 0 0 0 Q
port 10 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 2668 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 243194
string GDS_START 223698
<< end >>
