magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 920 561
rect 123 367 157 527
rect 467 333 533 425
rect 635 333 701 493
rect 735 367 801 527
rect 835 333 903 493
rect 467 299 903 333
rect 18 211 248 265
rect 282 211 444 265
rect 478 211 641 265
rect 123 17 157 109
rect 291 17 393 109
rect 535 17 601 109
rect 735 119 801 299
rect 835 151 903 265
rect 0 -17 920 17
<< obsli1 >>
rect 18 333 89 493
rect 191 333 257 493
rect 291 459 601 493
rect 291 367 325 459
rect 359 333 425 425
rect 18 299 425 333
rect 567 367 601 459
rect 18 143 701 177
rect 18 51 89 143
rect 191 51 257 143
rect 435 51 501 143
rect 635 85 701 143
rect 835 85 903 117
rect 635 51 903 85
<< metal1 >>
rect 0 496 920 592
rect 0 -48 920 48
<< labels >>
rlabel locali s 18 211 248 265 6 A1
port 1 nsew signal input
rlabel locali s 282 211 444 265 6 A2
port 2 nsew signal input
rlabel locali s 478 211 641 265 6 A3
port 3 nsew signal input
rlabel locali s 835 151 903 265 6 B1
port 4 nsew signal input
rlabel locali s 835 333 903 493 6 Y
port 5 nsew signal output
rlabel locali s 735 119 801 299 6 Y
port 5 nsew signal output
rlabel locali s 635 333 701 493 6 Y
port 5 nsew signal output
rlabel locali s 467 333 533 425 6 Y
port 5 nsew signal output
rlabel locali s 467 299 903 333 6 Y
port 5 nsew signal output
rlabel locali s 535 17 601 109 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 291 17 393 109 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 123 17 157 109 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 920 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 920 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 735 367 801 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 123 367 157 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 920 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 920 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 920 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 849346
string GDS_START 840418
<< end >>
