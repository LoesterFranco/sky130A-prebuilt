magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 129 325 171 425
rect 309 325 359 425
rect 497 325 547 425
rect 685 325 735 425
rect 129 289 735 325
rect 18 215 419 255
rect 479 177 539 289
rect 573 215 888 255
rect 935 215 1257 257
rect 1302 215 1707 257
rect 479 129 1223 177
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 18 459 933 493
rect 18 291 85 459
rect 215 359 265 459
rect 403 359 453 459
rect 591 359 641 459
rect 779 325 933 459
rect 977 359 1027 527
rect 1071 325 1121 493
rect 1165 359 1215 527
rect 1259 325 1309 493
rect 1353 359 1403 527
rect 1447 325 1497 493
rect 1541 359 1591 527
rect 1635 325 1685 493
rect 779 291 1685 325
rect 19 145 445 181
rect 19 51 85 145
rect 129 17 163 111
rect 197 51 273 145
rect 317 17 351 111
rect 385 95 445 145
rect 1267 145 1693 181
rect 1267 95 1317 145
rect 385 51 837 95
rect 875 51 1317 95
rect 1361 17 1395 111
rect 1429 51 1505 145
rect 1549 17 1583 111
rect 1617 51 1693 145
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
<< metal1 >>
rect 0 561 1748 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 0 496 1748 527
rect 0 17 1748 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
rect 0 -48 1748 -17
<< labels >>
rlabel locali s 935 215 1257 257 6 A1
port 1 nsew signal input
rlabel locali s 1302 215 1707 257 6 A2
port 2 nsew signal input
rlabel locali s 573 215 888 255 6 B1
port 3 nsew signal input
rlabel locali s 18 215 419 255 6 B2
port 4 nsew signal input
rlabel locali s 685 325 735 425 6 Y
port 5 nsew signal output
rlabel locali s 497 325 547 425 6 Y
port 5 nsew signal output
rlabel locali s 479 177 539 289 6 Y
port 5 nsew signal output
rlabel locali s 479 129 1223 177 6 Y
port 5 nsew signal output
rlabel locali s 309 325 359 425 6 Y
port 5 nsew signal output
rlabel locali s 129 325 171 425 6 Y
port 5 nsew signal output
rlabel locali s 129 289 735 325 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -48 1748 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 1748 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1748 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1304530
string GDS_START 1291812
<< end >>
