magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 736 561
rect 19 451 85 527
rect 25 151 66 415
rect 214 383 280 527
rect 447 367 513 527
rect 547 299 614 493
rect 649 367 715 527
rect 178 84 249 265
rect 284 261 318 265
rect 284 83 344 261
rect 380 83 432 265
rect 466 17 513 178
rect 579 161 614 299
rect 547 68 614 161
rect 547 59 613 68
rect 651 17 717 162
rect 0 -17 736 17
<< obsli1 >>
rect 120 333 170 493
rect 317 333 367 493
rect 100 299 511 333
rect 100 117 134 299
rect 35 51 134 117
rect 466 263 511 299
rect 466 215 545 263
<< metal1 >>
rect 0 496 736 592
rect 0 -48 736 48
<< labels >>
rlabel locali s 25 151 66 415 6 A
port 1 nsew signal input
rlabel locali s 178 84 249 265 6 B
port 2 nsew signal input
rlabel locali s 284 261 318 265 6 C
port 3 nsew signal input
rlabel locali s 284 83 344 261 6 C
port 3 nsew signal input
rlabel locali s 380 83 432 265 6 D
port 4 nsew signal input
rlabel locali s 579 161 614 299 6 X
port 5 nsew signal output
rlabel locali s 547 299 614 493 6 X
port 5 nsew signal output
rlabel locali s 547 68 614 161 6 X
port 5 nsew signal output
rlabel locali s 547 59 613 68 6 X
port 5 nsew signal output
rlabel locali s 651 17 717 162 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 466 17 513 178 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 736 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 736 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 649 367 715 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 447 367 513 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 214 383 280 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 19 451 85 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 736 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 736 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3814836
string GDS_START 3807618
<< end >>
