magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 920 561
rect 115 357 181 421
rect 20 199 81 323
rect 115 171 171 357
rect 487 367 533 527
rect 659 367 705 527
rect 831 367 877 527
rect 207 257 251 323
rect 835 257 900 331
rect 207 207 357 257
rect 474 207 616 257
rect 748 207 900 257
rect 29 17 79 163
rect 115 131 629 171
rect 115 51 167 131
rect 201 17 267 95
rect 301 57 339 131
rect 373 17 439 95
rect 735 17 801 91
rect 0 -17 920 17
<< obsli1 >>
rect 29 457 443 491
rect 29 357 81 457
rect 215 451 443 457
rect 215 357 253 451
rect 287 331 353 415
rect 387 367 443 451
rect 569 331 623 493
rect 741 331 795 493
rect 287 291 795 331
rect 665 127 887 171
rect 665 95 699 127
rect 477 53 699 95
rect 837 53 887 127
<< metal1 >>
rect 0 496 920 592
rect 0 -48 920 48
<< labels >>
rlabel locali s 474 207 616 257 6 A1
port 1 nsew signal input
rlabel locali s 835 257 900 331 6 A2
port 2 nsew signal input
rlabel locali s 748 207 900 257 6 A2
port 2 nsew signal input
rlabel locali s 207 257 251 323 6 B1
port 3 nsew signal input
rlabel locali s 207 207 357 257 6 B1
port 3 nsew signal input
rlabel locali s 20 199 81 323 6 C1
port 4 nsew signal input
rlabel locali s 301 57 339 131 6 Y
port 5 nsew signal output
rlabel locali s 115 357 181 421 6 Y
port 5 nsew signal output
rlabel locali s 115 171 171 357 6 Y
port 5 nsew signal output
rlabel locali s 115 131 629 171 6 Y
port 5 nsew signal output
rlabel locali s 115 51 167 131 6 Y
port 5 nsew signal output
rlabel locali s 735 17 801 91 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 373 17 439 95 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 201 17 267 95 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 29 17 79 163 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 920 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 920 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 831 367 877 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 659 367 705 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 487 367 533 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 920 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 920 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 920 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3964922
string GDS_START 3955980
<< end >>
