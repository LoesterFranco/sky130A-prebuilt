magic
tech sky130A
timestamp 1601049429
<< properties >>
string gencell sky130_fd_pr__cap_vpp_08p6x07p8_m1m2_lishield
string parameter m=1
string library sky130
<< end >>
