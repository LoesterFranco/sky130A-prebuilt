magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 87 252 167 380
rect 201 252 267 380
rect 1338 344 1423 570
rect 1175 236 1236 310
rect 1389 210 1423 344
rect 1313 70 1423 210
rect 1639 364 1706 596
rect 1672 226 1706 364
rect 1649 70 1706 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 19 448 73 596
rect 113 482 179 649
rect 501 580 567 649
rect 624 581 858 615
rect 213 546 403 580
rect 213 448 247 546
rect 369 512 582 546
rect 19 414 247 448
rect 281 478 335 512
rect 281 444 511 478
rect 281 420 335 444
rect 19 218 53 414
rect 301 218 335 420
rect 19 108 90 218
rect 126 17 192 218
rect 226 70 335 218
rect 369 344 443 410
rect 369 192 403 344
rect 477 310 511 444
rect 437 260 511 310
rect 548 360 582 512
rect 624 428 658 581
rect 692 481 758 547
rect 624 394 690 428
rect 548 294 614 360
rect 656 290 690 394
rect 724 358 758 481
rect 792 410 858 581
rect 936 504 1089 649
rect 1123 458 1189 570
rect 906 392 1189 458
rect 1223 412 1289 649
rect 1058 378 1189 392
rect 724 324 945 358
rect 875 310 945 324
rect 1058 344 1304 378
rect 656 260 722 290
rect 437 226 722 260
rect 656 224 722 226
rect 369 190 435 192
rect 775 190 841 290
rect 369 156 841 190
rect 875 244 1024 310
rect 369 70 435 156
rect 875 122 909 244
rect 1058 210 1092 344
rect 1270 310 1304 344
rect 1270 244 1355 310
rect 469 17 583 120
rect 681 72 909 122
rect 946 17 996 206
rect 1042 70 1092 210
rect 1206 17 1272 202
rect 1457 326 1507 556
rect 1549 364 1602 649
rect 1457 260 1638 326
rect 1457 108 1512 260
rect 1549 17 1615 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
<< metal1 >>
rect 0 683 1728 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 0 617 1728 649
rect 0 17 1728 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
rect 0 -49 1728 -17
<< labels >>
rlabel locali s 87 252 167 380 6 D
port 1 nsew signal input
rlabel locali s 1389 210 1423 344 6 Q
port 2 nsew signal output
rlabel locali s 1338 344 1423 570 6 Q
port 2 nsew signal output
rlabel locali s 1313 70 1423 210 6 Q
port 2 nsew signal output
rlabel locali s 1672 226 1706 364 6 Q_N
port 3 nsew signal output
rlabel locali s 1649 70 1706 226 6 Q_N
port 3 nsew signal output
rlabel locali s 1639 364 1706 596 6 Q_N
port 3 nsew signal output
rlabel locali s 1175 236 1236 310 6 RESET_B
port 4 nsew signal input
rlabel locali s 201 252 267 380 6 GATE_N
port 5 nsew clock input
rlabel metal1 s 0 -49 1728 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 1728 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1728 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3057024
string GDS_START 3043414
<< end >>
