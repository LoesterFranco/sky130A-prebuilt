magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 5190 582
<< pwell >>
rect 29 -17 63 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 3801 -17 3835 17
rect 3893 -17 3927 17
rect 5089 -17 5123 17
<< scnmos >>
rect 89 47 119 177
rect 173 47 203 177
rect 277 69 307 173
rect 361 69 391 173
rect 587 47 617 151
rect 671 47 701 151
rect 897 69 927 173
rect 981 69 1011 173
rect 1085 47 1115 177
rect 1169 47 1199 177
rect 1377 47 1407 177
rect 1461 47 1491 177
rect 1565 69 1595 173
rect 1649 69 1679 173
rect 1875 47 1905 151
rect 1959 47 1989 151
rect 2185 69 2215 173
rect 2269 69 2299 173
rect 2373 47 2403 177
rect 2457 47 2487 177
rect 2665 47 2695 177
rect 2749 47 2779 177
rect 2853 69 2883 173
rect 2937 69 2967 173
rect 3163 47 3193 151
rect 3247 47 3277 151
rect 3473 69 3503 173
rect 3557 69 3587 173
rect 3661 47 3691 177
rect 3745 47 3775 177
rect 3953 47 3983 177
rect 4037 47 4067 177
rect 4141 69 4171 173
rect 4225 69 4255 173
rect 4451 47 4481 151
rect 4535 47 4565 151
rect 4761 69 4791 173
rect 4845 69 4875 173
rect 4949 47 4979 177
rect 5033 47 5063 177
<< pmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 280 333 316 497
rect 374 333 410 497
rect 572 297 608 497
rect 680 297 716 497
rect 878 333 914 497
rect 972 333 1008 497
rect 1077 297 1113 497
rect 1171 297 1207 497
rect 1369 297 1405 497
rect 1463 297 1499 497
rect 1568 333 1604 497
rect 1662 333 1698 497
rect 1860 297 1896 497
rect 1968 297 2004 497
rect 2166 333 2202 497
rect 2260 333 2296 497
rect 2365 297 2401 497
rect 2459 297 2495 497
rect 2657 297 2693 497
rect 2751 297 2787 497
rect 2856 333 2892 497
rect 2950 333 2986 497
rect 3148 297 3184 497
rect 3256 297 3292 497
rect 3454 333 3490 497
rect 3548 333 3584 497
rect 3653 297 3689 497
rect 3747 297 3783 497
rect 3945 297 3981 497
rect 4039 297 4075 497
rect 4144 333 4180 497
rect 4238 333 4274 497
rect 4436 297 4472 497
rect 4544 297 4580 497
rect 4742 333 4778 497
rect 4836 333 4872 497
rect 4941 297 4977 497
rect 5035 297 5071 497
<< ndiff >>
rect 27 161 89 177
rect 27 127 45 161
rect 79 127 89 161
rect 27 93 89 127
rect 27 59 45 93
rect 79 59 89 93
rect 27 47 89 59
rect 119 93 173 177
rect 119 59 129 93
rect 163 59 173 93
rect 119 47 173 59
rect 203 173 262 177
rect 203 169 277 173
rect 203 135 218 169
rect 252 135 277 169
rect 203 101 277 135
rect 203 67 218 101
rect 252 69 277 101
rect 307 153 361 173
rect 307 119 317 153
rect 351 119 361 153
rect 307 69 361 119
rect 391 138 443 173
rect 391 104 401 138
rect 435 104 443 138
rect 391 69 443 104
rect 252 67 262 69
rect 203 47 262 67
rect 1026 173 1085 177
rect 535 116 587 151
rect 535 82 543 116
rect 577 82 587 116
rect 535 47 587 82
rect 617 116 671 151
rect 617 82 627 116
rect 661 82 671 116
rect 617 47 671 82
rect 701 116 753 151
rect 701 82 711 116
rect 745 82 753 116
rect 701 47 753 82
rect 845 138 897 173
rect 845 104 853 138
rect 887 104 897 138
rect 845 69 897 104
rect 927 153 981 173
rect 927 119 937 153
rect 971 119 981 153
rect 927 69 981 119
rect 1011 169 1085 173
rect 1011 135 1036 169
rect 1070 135 1085 169
rect 1011 101 1085 135
rect 1011 69 1036 101
rect 1026 67 1036 69
rect 1070 67 1085 101
rect 1026 47 1085 67
rect 1115 93 1169 177
rect 1115 59 1125 93
rect 1159 59 1169 93
rect 1115 47 1169 59
rect 1199 161 1261 177
rect 1199 127 1209 161
rect 1243 127 1261 161
rect 1199 93 1261 127
rect 1199 59 1209 93
rect 1243 59 1261 93
rect 1199 47 1261 59
rect 1315 161 1377 177
rect 1315 127 1333 161
rect 1367 127 1377 161
rect 1315 93 1377 127
rect 1315 59 1333 93
rect 1367 59 1377 93
rect 1315 47 1377 59
rect 1407 93 1461 177
rect 1407 59 1417 93
rect 1451 59 1461 93
rect 1407 47 1461 59
rect 1491 173 1550 177
rect 1491 169 1565 173
rect 1491 135 1506 169
rect 1540 135 1565 169
rect 1491 101 1565 135
rect 1491 67 1506 101
rect 1540 69 1565 101
rect 1595 153 1649 173
rect 1595 119 1605 153
rect 1639 119 1649 153
rect 1595 69 1649 119
rect 1679 138 1731 173
rect 1679 104 1689 138
rect 1723 104 1731 138
rect 1679 69 1731 104
rect 1540 67 1550 69
rect 1491 47 1550 67
rect 2314 173 2373 177
rect 1823 116 1875 151
rect 1823 82 1831 116
rect 1865 82 1875 116
rect 1823 47 1875 82
rect 1905 116 1959 151
rect 1905 82 1915 116
rect 1949 82 1959 116
rect 1905 47 1959 82
rect 1989 116 2041 151
rect 1989 82 1999 116
rect 2033 82 2041 116
rect 1989 47 2041 82
rect 2133 138 2185 173
rect 2133 104 2141 138
rect 2175 104 2185 138
rect 2133 69 2185 104
rect 2215 153 2269 173
rect 2215 119 2225 153
rect 2259 119 2269 153
rect 2215 69 2269 119
rect 2299 169 2373 173
rect 2299 135 2324 169
rect 2358 135 2373 169
rect 2299 101 2373 135
rect 2299 69 2324 101
rect 2314 67 2324 69
rect 2358 67 2373 101
rect 2314 47 2373 67
rect 2403 93 2457 177
rect 2403 59 2413 93
rect 2447 59 2457 93
rect 2403 47 2457 59
rect 2487 161 2549 177
rect 2487 127 2497 161
rect 2531 127 2549 161
rect 2487 93 2549 127
rect 2487 59 2497 93
rect 2531 59 2549 93
rect 2487 47 2549 59
rect 2603 161 2665 177
rect 2603 127 2621 161
rect 2655 127 2665 161
rect 2603 93 2665 127
rect 2603 59 2621 93
rect 2655 59 2665 93
rect 2603 47 2665 59
rect 2695 93 2749 177
rect 2695 59 2705 93
rect 2739 59 2749 93
rect 2695 47 2749 59
rect 2779 173 2838 177
rect 2779 169 2853 173
rect 2779 135 2794 169
rect 2828 135 2853 169
rect 2779 101 2853 135
rect 2779 67 2794 101
rect 2828 69 2853 101
rect 2883 153 2937 173
rect 2883 119 2893 153
rect 2927 119 2937 153
rect 2883 69 2937 119
rect 2967 138 3019 173
rect 2967 104 2977 138
rect 3011 104 3019 138
rect 2967 69 3019 104
rect 2828 67 2838 69
rect 2779 47 2838 67
rect 3602 173 3661 177
rect 3111 116 3163 151
rect 3111 82 3119 116
rect 3153 82 3163 116
rect 3111 47 3163 82
rect 3193 116 3247 151
rect 3193 82 3203 116
rect 3237 82 3247 116
rect 3193 47 3247 82
rect 3277 116 3329 151
rect 3277 82 3287 116
rect 3321 82 3329 116
rect 3277 47 3329 82
rect 3421 138 3473 173
rect 3421 104 3429 138
rect 3463 104 3473 138
rect 3421 69 3473 104
rect 3503 153 3557 173
rect 3503 119 3513 153
rect 3547 119 3557 153
rect 3503 69 3557 119
rect 3587 169 3661 173
rect 3587 135 3612 169
rect 3646 135 3661 169
rect 3587 101 3661 135
rect 3587 69 3612 101
rect 3602 67 3612 69
rect 3646 67 3661 101
rect 3602 47 3661 67
rect 3691 93 3745 177
rect 3691 59 3701 93
rect 3735 59 3745 93
rect 3691 47 3745 59
rect 3775 161 3837 177
rect 3775 127 3785 161
rect 3819 127 3837 161
rect 3775 93 3837 127
rect 3775 59 3785 93
rect 3819 59 3837 93
rect 3775 47 3837 59
rect 3891 161 3953 177
rect 3891 127 3909 161
rect 3943 127 3953 161
rect 3891 93 3953 127
rect 3891 59 3909 93
rect 3943 59 3953 93
rect 3891 47 3953 59
rect 3983 93 4037 177
rect 3983 59 3993 93
rect 4027 59 4037 93
rect 3983 47 4037 59
rect 4067 173 4126 177
rect 4067 169 4141 173
rect 4067 135 4082 169
rect 4116 135 4141 169
rect 4067 101 4141 135
rect 4067 67 4082 101
rect 4116 69 4141 101
rect 4171 153 4225 173
rect 4171 119 4181 153
rect 4215 119 4225 153
rect 4171 69 4225 119
rect 4255 138 4307 173
rect 4255 104 4265 138
rect 4299 104 4307 138
rect 4255 69 4307 104
rect 4116 67 4126 69
rect 4067 47 4126 67
rect 4890 173 4949 177
rect 4399 116 4451 151
rect 4399 82 4407 116
rect 4441 82 4451 116
rect 4399 47 4451 82
rect 4481 116 4535 151
rect 4481 82 4491 116
rect 4525 82 4535 116
rect 4481 47 4535 82
rect 4565 116 4617 151
rect 4565 82 4575 116
rect 4609 82 4617 116
rect 4565 47 4617 82
rect 4709 138 4761 173
rect 4709 104 4717 138
rect 4751 104 4761 138
rect 4709 69 4761 104
rect 4791 153 4845 173
rect 4791 119 4801 153
rect 4835 119 4845 153
rect 4791 69 4845 119
rect 4875 169 4949 173
rect 4875 135 4900 169
rect 4934 135 4949 169
rect 4875 101 4949 135
rect 4875 69 4900 101
rect 4890 67 4900 69
rect 4934 67 4949 101
rect 4890 47 4949 67
rect 4979 93 5033 177
rect 4979 59 4989 93
rect 5023 59 5033 93
rect 4979 47 5033 59
rect 5063 161 5125 177
rect 5063 127 5073 161
rect 5107 127 5125 161
rect 5063 93 5125 127
rect 5063 59 5073 93
rect 5107 59 5125 93
rect 5063 47 5125 59
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 485 175 497
rect 117 451 129 485
rect 163 451 175 485
rect 117 405 175 451
rect 117 371 129 405
rect 163 371 175 405
rect 117 297 175 371
rect 211 477 280 497
rect 211 443 223 477
rect 257 443 280 477
rect 211 373 280 443
rect 211 339 223 373
rect 257 339 280 373
rect 211 333 280 339
rect 316 421 374 497
rect 316 387 328 421
rect 362 387 374 421
rect 316 333 374 387
rect 410 477 464 497
rect 410 443 422 477
rect 456 443 464 477
rect 410 379 464 443
rect 410 345 422 379
rect 456 345 464 379
rect 410 333 464 345
rect 518 479 572 497
rect 518 445 526 479
rect 560 445 572 479
rect 518 411 572 445
rect 518 377 526 411
rect 560 377 572 411
rect 518 343 572 377
rect 211 297 263 333
rect 518 309 526 343
rect 560 309 572 343
rect 518 297 572 309
rect 608 479 680 497
rect 608 445 627 479
rect 661 445 680 479
rect 608 411 680 445
rect 608 377 627 411
rect 661 377 680 411
rect 608 343 680 377
rect 608 309 627 343
rect 661 309 680 343
rect 608 297 680 309
rect 716 479 770 497
rect 716 445 728 479
rect 762 445 770 479
rect 716 411 770 445
rect 716 377 728 411
rect 762 377 770 411
rect 716 343 770 377
rect 716 309 728 343
rect 762 309 770 343
rect 824 477 878 497
rect 824 443 832 477
rect 866 443 878 477
rect 824 379 878 443
rect 824 345 832 379
rect 866 345 878 379
rect 824 333 878 345
rect 914 421 972 497
rect 914 387 926 421
rect 960 387 972 421
rect 914 333 972 387
rect 1008 477 1077 497
rect 1008 443 1031 477
rect 1065 443 1077 477
rect 1008 373 1077 443
rect 1008 339 1031 373
rect 1065 339 1077 373
rect 1008 333 1077 339
rect 716 297 770 309
rect 1025 297 1077 333
rect 1113 485 1171 497
rect 1113 451 1125 485
rect 1159 451 1171 485
rect 1113 405 1171 451
rect 1113 371 1125 405
rect 1159 371 1171 405
rect 1113 297 1171 371
rect 1207 485 1261 497
rect 1207 451 1219 485
rect 1253 451 1261 485
rect 1207 417 1261 451
rect 1207 383 1219 417
rect 1253 383 1261 417
rect 1207 349 1261 383
rect 1207 315 1219 349
rect 1253 315 1261 349
rect 1207 297 1261 315
rect 1315 485 1369 497
rect 1315 451 1323 485
rect 1357 451 1369 485
rect 1315 417 1369 451
rect 1315 383 1323 417
rect 1357 383 1369 417
rect 1315 349 1369 383
rect 1315 315 1323 349
rect 1357 315 1369 349
rect 1315 297 1369 315
rect 1405 485 1463 497
rect 1405 451 1417 485
rect 1451 451 1463 485
rect 1405 405 1463 451
rect 1405 371 1417 405
rect 1451 371 1463 405
rect 1405 297 1463 371
rect 1499 477 1568 497
rect 1499 443 1511 477
rect 1545 443 1568 477
rect 1499 373 1568 443
rect 1499 339 1511 373
rect 1545 339 1568 373
rect 1499 333 1568 339
rect 1604 421 1662 497
rect 1604 387 1616 421
rect 1650 387 1662 421
rect 1604 333 1662 387
rect 1698 477 1752 497
rect 1698 443 1710 477
rect 1744 443 1752 477
rect 1698 379 1752 443
rect 1698 345 1710 379
rect 1744 345 1752 379
rect 1698 333 1752 345
rect 1806 479 1860 497
rect 1806 445 1814 479
rect 1848 445 1860 479
rect 1806 411 1860 445
rect 1806 377 1814 411
rect 1848 377 1860 411
rect 1806 343 1860 377
rect 1499 297 1551 333
rect 1806 309 1814 343
rect 1848 309 1860 343
rect 1806 297 1860 309
rect 1896 479 1968 497
rect 1896 445 1915 479
rect 1949 445 1968 479
rect 1896 411 1968 445
rect 1896 377 1915 411
rect 1949 377 1968 411
rect 1896 343 1968 377
rect 1896 309 1915 343
rect 1949 309 1968 343
rect 1896 297 1968 309
rect 2004 479 2058 497
rect 2004 445 2016 479
rect 2050 445 2058 479
rect 2004 411 2058 445
rect 2004 377 2016 411
rect 2050 377 2058 411
rect 2004 343 2058 377
rect 2004 309 2016 343
rect 2050 309 2058 343
rect 2112 477 2166 497
rect 2112 443 2120 477
rect 2154 443 2166 477
rect 2112 379 2166 443
rect 2112 345 2120 379
rect 2154 345 2166 379
rect 2112 333 2166 345
rect 2202 421 2260 497
rect 2202 387 2214 421
rect 2248 387 2260 421
rect 2202 333 2260 387
rect 2296 477 2365 497
rect 2296 443 2319 477
rect 2353 443 2365 477
rect 2296 373 2365 443
rect 2296 339 2319 373
rect 2353 339 2365 373
rect 2296 333 2365 339
rect 2004 297 2058 309
rect 2313 297 2365 333
rect 2401 485 2459 497
rect 2401 451 2413 485
rect 2447 451 2459 485
rect 2401 405 2459 451
rect 2401 371 2413 405
rect 2447 371 2459 405
rect 2401 297 2459 371
rect 2495 485 2549 497
rect 2495 451 2507 485
rect 2541 451 2549 485
rect 2495 417 2549 451
rect 2495 383 2507 417
rect 2541 383 2549 417
rect 2495 349 2549 383
rect 2495 315 2507 349
rect 2541 315 2549 349
rect 2495 297 2549 315
rect 2603 485 2657 497
rect 2603 451 2611 485
rect 2645 451 2657 485
rect 2603 417 2657 451
rect 2603 383 2611 417
rect 2645 383 2657 417
rect 2603 349 2657 383
rect 2603 315 2611 349
rect 2645 315 2657 349
rect 2603 297 2657 315
rect 2693 485 2751 497
rect 2693 451 2705 485
rect 2739 451 2751 485
rect 2693 405 2751 451
rect 2693 371 2705 405
rect 2739 371 2751 405
rect 2693 297 2751 371
rect 2787 477 2856 497
rect 2787 443 2799 477
rect 2833 443 2856 477
rect 2787 373 2856 443
rect 2787 339 2799 373
rect 2833 339 2856 373
rect 2787 333 2856 339
rect 2892 421 2950 497
rect 2892 387 2904 421
rect 2938 387 2950 421
rect 2892 333 2950 387
rect 2986 477 3040 497
rect 2986 443 2998 477
rect 3032 443 3040 477
rect 2986 379 3040 443
rect 2986 345 2998 379
rect 3032 345 3040 379
rect 2986 333 3040 345
rect 3094 479 3148 497
rect 3094 445 3102 479
rect 3136 445 3148 479
rect 3094 411 3148 445
rect 3094 377 3102 411
rect 3136 377 3148 411
rect 3094 343 3148 377
rect 2787 297 2839 333
rect 3094 309 3102 343
rect 3136 309 3148 343
rect 3094 297 3148 309
rect 3184 479 3256 497
rect 3184 445 3203 479
rect 3237 445 3256 479
rect 3184 411 3256 445
rect 3184 377 3203 411
rect 3237 377 3256 411
rect 3184 343 3256 377
rect 3184 309 3203 343
rect 3237 309 3256 343
rect 3184 297 3256 309
rect 3292 479 3346 497
rect 3292 445 3304 479
rect 3338 445 3346 479
rect 3292 411 3346 445
rect 3292 377 3304 411
rect 3338 377 3346 411
rect 3292 343 3346 377
rect 3292 309 3304 343
rect 3338 309 3346 343
rect 3400 477 3454 497
rect 3400 443 3408 477
rect 3442 443 3454 477
rect 3400 379 3454 443
rect 3400 345 3408 379
rect 3442 345 3454 379
rect 3400 333 3454 345
rect 3490 421 3548 497
rect 3490 387 3502 421
rect 3536 387 3548 421
rect 3490 333 3548 387
rect 3584 477 3653 497
rect 3584 443 3607 477
rect 3641 443 3653 477
rect 3584 373 3653 443
rect 3584 339 3607 373
rect 3641 339 3653 373
rect 3584 333 3653 339
rect 3292 297 3346 309
rect 3601 297 3653 333
rect 3689 485 3747 497
rect 3689 451 3701 485
rect 3735 451 3747 485
rect 3689 405 3747 451
rect 3689 371 3701 405
rect 3735 371 3747 405
rect 3689 297 3747 371
rect 3783 485 3837 497
rect 3783 451 3795 485
rect 3829 451 3837 485
rect 3783 417 3837 451
rect 3783 383 3795 417
rect 3829 383 3837 417
rect 3783 349 3837 383
rect 3783 315 3795 349
rect 3829 315 3837 349
rect 3783 297 3837 315
rect 3891 485 3945 497
rect 3891 451 3899 485
rect 3933 451 3945 485
rect 3891 417 3945 451
rect 3891 383 3899 417
rect 3933 383 3945 417
rect 3891 349 3945 383
rect 3891 315 3899 349
rect 3933 315 3945 349
rect 3891 297 3945 315
rect 3981 485 4039 497
rect 3981 451 3993 485
rect 4027 451 4039 485
rect 3981 405 4039 451
rect 3981 371 3993 405
rect 4027 371 4039 405
rect 3981 297 4039 371
rect 4075 477 4144 497
rect 4075 443 4087 477
rect 4121 443 4144 477
rect 4075 373 4144 443
rect 4075 339 4087 373
rect 4121 339 4144 373
rect 4075 333 4144 339
rect 4180 421 4238 497
rect 4180 387 4192 421
rect 4226 387 4238 421
rect 4180 333 4238 387
rect 4274 477 4328 497
rect 4274 443 4286 477
rect 4320 443 4328 477
rect 4274 379 4328 443
rect 4274 345 4286 379
rect 4320 345 4328 379
rect 4274 333 4328 345
rect 4382 479 4436 497
rect 4382 445 4390 479
rect 4424 445 4436 479
rect 4382 411 4436 445
rect 4382 377 4390 411
rect 4424 377 4436 411
rect 4382 343 4436 377
rect 4075 297 4127 333
rect 4382 309 4390 343
rect 4424 309 4436 343
rect 4382 297 4436 309
rect 4472 479 4544 497
rect 4472 445 4491 479
rect 4525 445 4544 479
rect 4472 411 4544 445
rect 4472 377 4491 411
rect 4525 377 4544 411
rect 4472 343 4544 377
rect 4472 309 4491 343
rect 4525 309 4544 343
rect 4472 297 4544 309
rect 4580 479 4634 497
rect 4580 445 4592 479
rect 4626 445 4634 479
rect 4580 411 4634 445
rect 4580 377 4592 411
rect 4626 377 4634 411
rect 4580 343 4634 377
rect 4580 309 4592 343
rect 4626 309 4634 343
rect 4688 477 4742 497
rect 4688 443 4696 477
rect 4730 443 4742 477
rect 4688 379 4742 443
rect 4688 345 4696 379
rect 4730 345 4742 379
rect 4688 333 4742 345
rect 4778 421 4836 497
rect 4778 387 4790 421
rect 4824 387 4836 421
rect 4778 333 4836 387
rect 4872 477 4941 497
rect 4872 443 4895 477
rect 4929 443 4941 477
rect 4872 373 4941 443
rect 4872 339 4895 373
rect 4929 339 4941 373
rect 4872 333 4941 339
rect 4580 297 4634 309
rect 4889 297 4941 333
rect 4977 485 5035 497
rect 4977 451 4989 485
rect 5023 451 5035 485
rect 4977 405 5035 451
rect 4977 371 4989 405
rect 5023 371 5035 405
rect 4977 297 5035 371
rect 5071 485 5125 497
rect 5071 451 5083 485
rect 5117 451 5125 485
rect 5071 417 5125 451
rect 5071 383 5083 417
rect 5117 383 5125 417
rect 5071 349 5125 383
rect 5071 315 5083 349
rect 5117 315 5125 349
rect 5071 297 5125 315
<< ndiffc >>
rect 45 127 79 161
rect 45 59 79 93
rect 129 59 163 93
rect 218 135 252 169
rect 218 67 252 101
rect 317 119 351 153
rect 401 104 435 138
rect 543 82 577 116
rect 627 82 661 116
rect 711 82 745 116
rect 853 104 887 138
rect 937 119 971 153
rect 1036 135 1070 169
rect 1036 67 1070 101
rect 1125 59 1159 93
rect 1209 127 1243 161
rect 1209 59 1243 93
rect 1333 127 1367 161
rect 1333 59 1367 93
rect 1417 59 1451 93
rect 1506 135 1540 169
rect 1506 67 1540 101
rect 1605 119 1639 153
rect 1689 104 1723 138
rect 1831 82 1865 116
rect 1915 82 1949 116
rect 1999 82 2033 116
rect 2141 104 2175 138
rect 2225 119 2259 153
rect 2324 135 2358 169
rect 2324 67 2358 101
rect 2413 59 2447 93
rect 2497 127 2531 161
rect 2497 59 2531 93
rect 2621 127 2655 161
rect 2621 59 2655 93
rect 2705 59 2739 93
rect 2794 135 2828 169
rect 2794 67 2828 101
rect 2893 119 2927 153
rect 2977 104 3011 138
rect 3119 82 3153 116
rect 3203 82 3237 116
rect 3287 82 3321 116
rect 3429 104 3463 138
rect 3513 119 3547 153
rect 3612 135 3646 169
rect 3612 67 3646 101
rect 3701 59 3735 93
rect 3785 127 3819 161
rect 3785 59 3819 93
rect 3909 127 3943 161
rect 3909 59 3943 93
rect 3993 59 4027 93
rect 4082 135 4116 169
rect 4082 67 4116 101
rect 4181 119 4215 153
rect 4265 104 4299 138
rect 4407 82 4441 116
rect 4491 82 4525 116
rect 4575 82 4609 116
rect 4717 104 4751 138
rect 4801 119 4835 153
rect 4900 135 4934 169
rect 4900 67 4934 101
rect 4989 59 5023 93
rect 5073 127 5107 161
rect 5073 59 5107 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 451 163 485
rect 129 371 163 405
rect 223 443 257 477
rect 223 339 257 373
rect 328 387 362 421
rect 422 443 456 477
rect 422 345 456 379
rect 526 445 560 479
rect 526 377 560 411
rect 526 309 560 343
rect 627 445 661 479
rect 627 377 661 411
rect 627 309 661 343
rect 728 445 762 479
rect 728 377 762 411
rect 728 309 762 343
rect 832 443 866 477
rect 832 345 866 379
rect 926 387 960 421
rect 1031 443 1065 477
rect 1031 339 1065 373
rect 1125 451 1159 485
rect 1125 371 1159 405
rect 1219 451 1253 485
rect 1219 383 1253 417
rect 1219 315 1253 349
rect 1323 451 1357 485
rect 1323 383 1357 417
rect 1323 315 1357 349
rect 1417 451 1451 485
rect 1417 371 1451 405
rect 1511 443 1545 477
rect 1511 339 1545 373
rect 1616 387 1650 421
rect 1710 443 1744 477
rect 1710 345 1744 379
rect 1814 445 1848 479
rect 1814 377 1848 411
rect 1814 309 1848 343
rect 1915 445 1949 479
rect 1915 377 1949 411
rect 1915 309 1949 343
rect 2016 445 2050 479
rect 2016 377 2050 411
rect 2016 309 2050 343
rect 2120 443 2154 477
rect 2120 345 2154 379
rect 2214 387 2248 421
rect 2319 443 2353 477
rect 2319 339 2353 373
rect 2413 451 2447 485
rect 2413 371 2447 405
rect 2507 451 2541 485
rect 2507 383 2541 417
rect 2507 315 2541 349
rect 2611 451 2645 485
rect 2611 383 2645 417
rect 2611 315 2645 349
rect 2705 451 2739 485
rect 2705 371 2739 405
rect 2799 443 2833 477
rect 2799 339 2833 373
rect 2904 387 2938 421
rect 2998 443 3032 477
rect 2998 345 3032 379
rect 3102 445 3136 479
rect 3102 377 3136 411
rect 3102 309 3136 343
rect 3203 445 3237 479
rect 3203 377 3237 411
rect 3203 309 3237 343
rect 3304 445 3338 479
rect 3304 377 3338 411
rect 3304 309 3338 343
rect 3408 443 3442 477
rect 3408 345 3442 379
rect 3502 387 3536 421
rect 3607 443 3641 477
rect 3607 339 3641 373
rect 3701 451 3735 485
rect 3701 371 3735 405
rect 3795 451 3829 485
rect 3795 383 3829 417
rect 3795 315 3829 349
rect 3899 451 3933 485
rect 3899 383 3933 417
rect 3899 315 3933 349
rect 3993 451 4027 485
rect 3993 371 4027 405
rect 4087 443 4121 477
rect 4087 339 4121 373
rect 4192 387 4226 421
rect 4286 443 4320 477
rect 4286 345 4320 379
rect 4390 445 4424 479
rect 4390 377 4424 411
rect 4390 309 4424 343
rect 4491 445 4525 479
rect 4491 377 4525 411
rect 4491 309 4525 343
rect 4592 445 4626 479
rect 4592 377 4626 411
rect 4592 309 4626 343
rect 4696 443 4730 477
rect 4696 345 4730 379
rect 4790 387 4824 421
rect 4895 443 4929 477
rect 4895 339 4929 373
rect 4989 451 5023 485
rect 4989 371 5023 405
rect 5083 451 5117 485
rect 5083 383 5117 417
rect 5083 315 5117 349
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 280 497 316 523
rect 374 497 410 523
rect 572 497 608 523
rect 680 497 716 523
rect 878 497 914 523
rect 972 497 1008 523
rect 1077 497 1113 523
rect 1171 497 1207 523
rect 1369 497 1405 523
rect 1463 497 1499 523
rect 1568 497 1604 523
rect 1662 497 1698 523
rect 1860 497 1896 523
rect 1968 497 2004 523
rect 2166 497 2202 523
rect 2260 497 2296 523
rect 2365 497 2401 523
rect 2459 497 2495 523
rect 2657 497 2693 523
rect 2751 497 2787 523
rect 2856 497 2892 523
rect 2950 497 2986 523
rect 3148 497 3184 523
rect 3256 497 3292 523
rect 3454 497 3490 523
rect 3548 497 3584 523
rect 3653 497 3689 523
rect 3747 497 3783 523
rect 3945 497 3981 523
rect 4039 497 4075 523
rect 4144 497 4180 523
rect 4238 497 4274 523
rect 4436 497 4472 523
rect 4544 497 4580 523
rect 4742 497 4778 523
rect 4836 497 4872 523
rect 4941 497 4977 523
rect 5035 497 5071 523
rect 81 259 117 297
rect 175 259 211 297
rect 280 295 316 333
rect 374 295 410 333
rect 278 285 486 295
rect 278 265 436 285
rect 49 249 213 259
rect 49 215 65 249
rect 99 215 133 249
rect 167 215 213 249
rect 420 251 436 265
rect 470 251 486 285
rect 572 282 608 297
rect 680 282 716 297
rect 878 295 914 333
rect 972 295 1008 333
rect 802 285 1010 295
rect 570 265 610 282
rect 678 265 718 282
rect 420 241 486 251
rect 564 249 618 265
rect 49 205 213 215
rect 564 215 574 249
rect 608 215 618 249
rect 89 177 119 205
rect 173 177 203 205
rect 564 199 618 215
rect 670 249 724 265
rect 670 215 680 249
rect 714 215 724 249
rect 802 251 818 285
rect 852 265 1010 285
rect 852 251 868 265
rect 1077 259 1113 297
rect 1171 259 1207 297
rect 1369 259 1405 297
rect 1463 259 1499 297
rect 1568 295 1604 333
rect 1662 295 1698 333
rect 1566 285 1774 295
rect 1566 265 1724 285
rect 802 241 868 251
rect 1075 249 1239 259
rect 670 199 724 215
rect 1075 215 1121 249
rect 1155 215 1189 249
rect 1223 215 1239 249
rect 1075 205 1239 215
rect 1337 249 1501 259
rect 1337 215 1353 249
rect 1387 215 1421 249
rect 1455 215 1501 249
rect 1708 251 1724 265
rect 1758 251 1774 285
rect 1860 282 1896 297
rect 1968 282 2004 297
rect 2166 295 2202 333
rect 2260 295 2296 333
rect 2090 285 2298 295
rect 1858 265 1898 282
rect 1966 265 2006 282
rect 1708 241 1774 251
rect 1852 249 1906 265
rect 1337 205 1501 215
rect 1852 215 1862 249
rect 1896 215 1906 249
rect 277 173 307 199
rect 361 173 391 199
rect 458 169 617 199
rect 277 51 307 69
rect 361 51 391 69
rect 458 51 488 169
rect 587 151 617 169
rect 671 169 830 199
rect 897 173 927 199
rect 981 173 1011 199
rect 1085 177 1115 205
rect 1169 177 1199 205
rect 1377 177 1407 205
rect 1461 177 1491 205
rect 1852 199 1906 215
rect 1958 249 2012 265
rect 1958 215 1968 249
rect 2002 215 2012 249
rect 2090 251 2106 285
rect 2140 265 2298 285
rect 2140 251 2156 265
rect 2365 259 2401 297
rect 2459 259 2495 297
rect 2657 259 2693 297
rect 2751 259 2787 297
rect 2856 295 2892 333
rect 2950 295 2986 333
rect 2854 285 3062 295
rect 2854 265 3012 285
rect 2090 241 2156 251
rect 2363 249 2527 259
rect 1958 199 2012 215
rect 2363 215 2409 249
rect 2443 215 2477 249
rect 2511 215 2527 249
rect 2363 205 2527 215
rect 2625 249 2789 259
rect 2625 215 2641 249
rect 2675 215 2709 249
rect 2743 215 2789 249
rect 2996 251 3012 265
rect 3046 251 3062 285
rect 3148 282 3184 297
rect 3256 282 3292 297
rect 3454 295 3490 333
rect 3548 295 3584 333
rect 3378 285 3586 295
rect 3146 265 3186 282
rect 3254 265 3294 282
rect 2996 241 3062 251
rect 3140 249 3194 265
rect 2625 205 2789 215
rect 3140 215 3150 249
rect 3184 215 3194 249
rect 671 151 701 169
rect 89 19 119 47
rect 173 21 203 47
rect 277 21 488 51
rect 800 51 830 169
rect 897 51 927 69
rect 981 51 1011 69
rect 587 21 617 47
rect 671 21 701 47
rect 800 21 1011 51
rect 1565 173 1595 199
rect 1649 173 1679 199
rect 1746 169 1905 199
rect 1565 51 1595 69
rect 1649 51 1679 69
rect 1746 51 1776 169
rect 1875 151 1905 169
rect 1959 169 2118 199
rect 2185 173 2215 199
rect 2269 173 2299 199
rect 2373 177 2403 205
rect 2457 177 2487 205
rect 2665 177 2695 205
rect 2749 177 2779 205
rect 3140 199 3194 215
rect 3246 249 3300 265
rect 3246 215 3256 249
rect 3290 215 3300 249
rect 3378 251 3394 285
rect 3428 265 3586 285
rect 3428 251 3444 265
rect 3653 259 3689 297
rect 3747 259 3783 297
rect 3945 259 3981 297
rect 4039 259 4075 297
rect 4144 295 4180 333
rect 4238 295 4274 333
rect 4142 285 4350 295
rect 4142 265 4300 285
rect 3378 241 3444 251
rect 3651 249 3815 259
rect 3246 199 3300 215
rect 3651 215 3697 249
rect 3731 215 3765 249
rect 3799 215 3815 249
rect 3651 205 3815 215
rect 3913 249 4077 259
rect 3913 215 3929 249
rect 3963 215 3997 249
rect 4031 215 4077 249
rect 4284 251 4300 265
rect 4334 251 4350 285
rect 4436 282 4472 297
rect 4544 282 4580 297
rect 4742 295 4778 333
rect 4836 295 4872 333
rect 4666 285 4874 295
rect 4434 265 4474 282
rect 4542 265 4582 282
rect 4284 241 4350 251
rect 4428 249 4482 265
rect 3913 205 4077 215
rect 4428 215 4438 249
rect 4472 215 4482 249
rect 1959 151 1989 169
rect 1085 21 1115 47
rect 1169 19 1199 47
rect 1377 19 1407 47
rect 1461 21 1491 47
rect 1565 21 1776 51
rect 2088 51 2118 169
rect 2185 51 2215 69
rect 2269 51 2299 69
rect 1875 21 1905 47
rect 1959 21 1989 47
rect 2088 21 2299 51
rect 2853 173 2883 199
rect 2937 173 2967 199
rect 3034 169 3193 199
rect 2853 51 2883 69
rect 2937 51 2967 69
rect 3034 51 3064 169
rect 3163 151 3193 169
rect 3247 169 3406 199
rect 3473 173 3503 199
rect 3557 173 3587 199
rect 3661 177 3691 205
rect 3745 177 3775 205
rect 3953 177 3983 205
rect 4037 177 4067 205
rect 4428 199 4482 215
rect 4534 249 4588 265
rect 4534 215 4544 249
rect 4578 215 4588 249
rect 4666 251 4682 285
rect 4716 265 4874 285
rect 4716 251 4732 265
rect 4941 259 4977 297
rect 5035 259 5071 297
rect 4666 241 4732 251
rect 4939 249 5103 259
rect 4534 199 4588 215
rect 4939 215 4985 249
rect 5019 215 5053 249
rect 5087 215 5103 249
rect 4939 205 5103 215
rect 3247 151 3277 169
rect 2373 21 2403 47
rect 2457 19 2487 47
rect 2665 19 2695 47
rect 2749 21 2779 47
rect 2853 21 3064 51
rect 3376 51 3406 169
rect 3473 51 3503 69
rect 3557 51 3587 69
rect 3163 21 3193 47
rect 3247 21 3277 47
rect 3376 21 3587 51
rect 4141 173 4171 199
rect 4225 173 4255 199
rect 4322 169 4481 199
rect 4141 51 4171 69
rect 4225 51 4255 69
rect 4322 51 4352 169
rect 4451 151 4481 169
rect 4535 169 4694 199
rect 4761 173 4791 199
rect 4845 173 4875 199
rect 4949 177 4979 205
rect 5033 177 5063 205
rect 4535 151 4565 169
rect 3661 21 3691 47
rect 3745 19 3775 47
rect 3953 19 3983 47
rect 4037 21 4067 47
rect 4141 21 4352 51
rect 4664 51 4694 169
rect 4761 51 4791 69
rect 4845 51 4875 69
rect 4451 21 4481 47
rect 4535 21 4565 47
rect 4664 21 4875 51
rect 4949 21 4979 47
rect 5033 19 5063 47
<< polycont >>
rect 65 215 99 249
rect 133 215 167 249
rect 436 251 470 285
rect 574 215 608 249
rect 680 215 714 249
rect 818 251 852 285
rect 1121 215 1155 249
rect 1189 215 1223 249
rect 1353 215 1387 249
rect 1421 215 1455 249
rect 1724 251 1758 285
rect 1862 215 1896 249
rect 1968 215 2002 249
rect 2106 251 2140 285
rect 2409 215 2443 249
rect 2477 215 2511 249
rect 2641 215 2675 249
rect 2709 215 2743 249
rect 3012 251 3046 285
rect 3150 215 3184 249
rect 3256 215 3290 249
rect 3394 251 3428 285
rect 3697 215 3731 249
rect 3765 215 3799 249
rect 3929 215 3963 249
rect 3997 215 4031 249
rect 4300 251 4334 285
rect 4438 215 4472 249
rect 4544 215 4578 249
rect 4682 251 4716 285
rect 4985 215 5019 249
rect 5053 215 5087 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3157 561
rect 3191 527 3249 561
rect 3283 527 3341 561
rect 3375 527 3433 561
rect 3467 527 3525 561
rect 3559 527 3617 561
rect 3651 527 3709 561
rect 3743 527 3801 561
rect 3835 527 3893 561
rect 3927 527 3985 561
rect 4019 527 4077 561
rect 4111 527 4169 561
rect 4203 527 4261 561
rect 4295 527 4353 561
rect 4387 527 4445 561
rect 4479 527 4537 561
rect 4571 527 4629 561
rect 4663 527 4721 561
rect 4755 527 4813 561
rect 4847 527 4905 561
rect 4939 527 4997 561
rect 5031 527 5089 561
rect 5123 527 5152 561
rect 19 485 85 493
rect 19 451 35 485
rect 69 451 85 485
rect 19 442 85 451
rect 119 485 179 527
rect 119 451 129 485
rect 163 451 179 485
rect 19 417 79 442
rect 119 421 179 451
rect 19 383 35 417
rect 69 383 79 417
rect 19 349 79 383
rect 113 405 179 421
rect 113 371 129 405
rect 163 371 179 405
rect 113 367 179 371
rect 223 477 456 493
rect 257 459 422 477
rect 223 373 257 443
rect 19 315 35 349
rect 69 333 79 349
rect 293 421 379 425
rect 293 391 328 421
rect 293 357 305 391
rect 362 387 379 421
rect 339 357 379 387
rect 293 351 379 357
rect 422 379 456 443
rect 223 333 257 339
rect 69 315 257 333
rect 19 299 257 315
rect 19 249 183 265
rect 19 215 65 249
rect 99 215 133 249
rect 167 215 183 249
rect 19 211 183 215
rect 206 177 267 185
rect 317 177 351 351
rect 422 329 456 345
rect 510 479 576 493
rect 510 445 526 479
rect 560 445 576 479
rect 510 411 576 445
rect 510 377 526 411
rect 560 377 576 411
rect 510 343 576 377
rect 510 327 526 343
rect 490 309 526 327
rect 560 309 576 343
rect 490 295 576 309
rect 420 293 576 295
rect 611 479 677 527
rect 611 445 627 479
rect 661 445 677 479
rect 611 411 677 445
rect 611 377 627 411
rect 661 377 677 411
rect 611 343 677 377
rect 611 309 627 343
rect 661 309 677 343
rect 611 293 677 309
rect 712 479 778 493
rect 712 445 728 479
rect 762 445 778 479
rect 712 411 778 445
rect 712 377 728 411
rect 762 377 778 411
rect 712 343 778 377
rect 712 309 728 343
rect 762 327 778 343
rect 832 477 1065 493
rect 866 459 1031 477
rect 832 379 866 443
rect 909 421 995 425
rect 909 387 926 421
rect 960 391 995 421
rect 909 357 949 387
rect 983 357 995 391
rect 909 351 995 357
rect 1031 373 1065 443
rect 832 329 866 345
rect 762 309 798 327
rect 712 295 798 309
rect 712 293 868 295
rect 420 285 524 293
rect 420 251 436 285
rect 470 261 524 285
rect 764 285 868 293
rect 764 261 818 285
rect 470 251 503 261
rect 420 241 503 251
rect 29 169 267 177
rect 29 161 218 169
rect 29 127 45 161
rect 79 143 218 161
rect 79 127 95 143
rect 29 93 95 127
rect 206 135 218 143
rect 252 135 267 169
rect 29 59 45 93
rect 79 59 95 93
rect 29 51 95 59
rect 129 93 172 109
rect 163 59 172 93
rect 129 17 172 59
rect 206 101 267 135
rect 301 153 367 177
rect 301 119 317 153
rect 351 119 367 153
rect 401 138 435 154
rect 206 67 218 101
rect 252 85 267 101
rect 469 151 503 241
rect 558 249 625 259
rect 558 215 574 249
rect 608 215 625 249
rect 558 205 625 215
rect 663 249 730 259
rect 663 215 680 249
rect 714 215 730 249
rect 663 205 730 215
rect 785 251 818 261
rect 852 251 868 285
rect 785 241 868 251
rect 785 151 819 241
rect 937 177 971 351
rect 1109 485 1169 527
rect 1109 451 1125 485
rect 1159 451 1169 485
rect 1109 421 1169 451
rect 1203 485 1269 493
rect 1203 451 1219 485
rect 1253 451 1269 485
rect 1203 442 1269 451
rect 1109 405 1175 421
rect 1109 371 1125 405
rect 1159 371 1175 405
rect 1109 367 1175 371
rect 1209 417 1269 442
rect 1209 383 1219 417
rect 1253 383 1269 417
rect 1031 333 1065 339
rect 1209 349 1269 383
rect 1209 333 1219 349
rect 1031 315 1219 333
rect 1253 315 1269 349
rect 1031 299 1269 315
rect 1307 485 1373 493
rect 1307 451 1323 485
rect 1357 451 1373 485
rect 1307 442 1373 451
rect 1407 485 1467 527
rect 1407 451 1417 485
rect 1451 451 1467 485
rect 1307 417 1367 442
rect 1407 421 1467 451
rect 1307 383 1323 417
rect 1357 383 1367 417
rect 1307 349 1367 383
rect 1401 405 1467 421
rect 1401 371 1417 405
rect 1451 371 1467 405
rect 1401 367 1467 371
rect 1511 477 1744 493
rect 1545 459 1710 477
rect 1511 373 1545 443
rect 1307 315 1323 349
rect 1357 333 1367 349
rect 1581 421 1667 425
rect 1581 391 1616 421
rect 1581 357 1593 391
rect 1650 387 1667 421
rect 1627 357 1667 387
rect 1581 351 1667 357
rect 1710 379 1744 443
rect 1511 333 1545 339
rect 1357 315 1545 333
rect 1307 299 1545 315
rect 1105 249 1269 265
rect 1105 215 1121 249
rect 1155 215 1189 249
rect 1223 215 1269 249
rect 1105 211 1269 215
rect 1307 249 1471 265
rect 1307 215 1353 249
rect 1387 215 1421 249
rect 1455 215 1471 249
rect 1307 211 1471 215
rect 1021 177 1082 185
rect 1494 177 1555 185
rect 1605 177 1639 351
rect 1710 329 1744 345
rect 1798 479 1864 493
rect 1798 445 1814 479
rect 1848 445 1864 479
rect 1798 411 1864 445
rect 1798 377 1814 411
rect 1848 377 1864 411
rect 1798 343 1864 377
rect 1798 327 1814 343
rect 1778 309 1814 327
rect 1848 309 1864 343
rect 1778 295 1864 309
rect 1708 293 1864 295
rect 1899 479 1965 527
rect 1899 445 1915 479
rect 1949 445 1965 479
rect 1899 411 1965 445
rect 1899 377 1915 411
rect 1949 377 1965 411
rect 1899 343 1965 377
rect 1899 309 1915 343
rect 1949 309 1965 343
rect 1899 293 1965 309
rect 2000 479 2066 493
rect 2000 445 2016 479
rect 2050 445 2066 479
rect 2000 411 2066 445
rect 2000 377 2016 411
rect 2050 377 2066 411
rect 2000 343 2066 377
rect 2000 309 2016 343
rect 2050 327 2066 343
rect 2120 477 2353 493
rect 2154 459 2319 477
rect 2120 379 2154 443
rect 2197 421 2283 425
rect 2197 387 2214 421
rect 2248 391 2283 421
rect 2197 357 2237 387
rect 2271 357 2283 391
rect 2197 351 2283 357
rect 2319 373 2353 443
rect 2120 329 2154 345
rect 2050 309 2086 327
rect 2000 295 2086 309
rect 2000 293 2156 295
rect 1708 285 1812 293
rect 1708 251 1724 285
rect 1758 261 1812 285
rect 2052 285 2156 293
rect 2052 261 2106 285
rect 1758 251 1791 261
rect 1708 241 1791 251
rect 469 117 585 151
rect 401 85 435 104
rect 252 67 435 85
rect 206 51 435 67
rect 535 116 585 117
rect 535 82 543 116
rect 577 82 585 116
rect 535 66 585 82
rect 619 116 669 132
rect 619 82 627 116
rect 661 82 669 116
rect 619 17 669 82
rect 703 117 819 151
rect 853 138 887 154
rect 703 116 753 117
rect 703 82 711 116
rect 745 82 753 116
rect 703 66 753 82
rect 921 153 987 177
rect 921 119 937 153
rect 971 119 987 153
rect 1021 169 1259 177
rect 1021 135 1036 169
rect 1070 161 1259 169
rect 1070 143 1209 161
rect 1070 135 1082 143
rect 853 85 887 104
rect 1021 101 1082 135
rect 1193 127 1209 143
rect 1243 127 1259 161
rect 1021 85 1036 101
rect 853 67 1036 85
rect 1070 67 1082 101
rect 853 51 1082 67
rect 1116 93 1159 109
rect 1116 59 1125 93
rect 1116 17 1159 59
rect 1193 93 1259 127
rect 1193 59 1209 93
rect 1243 59 1259 93
rect 1193 51 1259 59
rect 1317 169 1555 177
rect 1317 161 1506 169
rect 1317 127 1333 161
rect 1367 143 1506 161
rect 1367 127 1383 143
rect 1317 93 1383 127
rect 1494 135 1506 143
rect 1540 135 1555 169
rect 1317 59 1333 93
rect 1367 59 1383 93
rect 1317 51 1383 59
rect 1417 93 1460 109
rect 1451 59 1460 93
rect 1417 17 1460 59
rect 1494 101 1555 135
rect 1589 153 1655 177
rect 1589 119 1605 153
rect 1639 119 1655 153
rect 1689 138 1723 154
rect 1494 67 1506 101
rect 1540 85 1555 101
rect 1757 151 1791 241
rect 1846 249 1913 259
rect 1846 215 1862 249
rect 1896 215 1913 249
rect 1846 205 1913 215
rect 1951 249 2018 259
rect 1951 215 1968 249
rect 2002 215 2018 249
rect 1951 205 2018 215
rect 2073 251 2106 261
rect 2140 251 2156 285
rect 2073 241 2156 251
rect 2073 151 2107 241
rect 2225 177 2259 351
rect 2397 485 2457 527
rect 2397 451 2413 485
rect 2447 451 2457 485
rect 2397 421 2457 451
rect 2491 485 2557 493
rect 2491 451 2507 485
rect 2541 451 2557 485
rect 2491 442 2557 451
rect 2397 405 2463 421
rect 2397 371 2413 405
rect 2447 371 2463 405
rect 2397 367 2463 371
rect 2497 417 2557 442
rect 2497 383 2507 417
rect 2541 383 2557 417
rect 2319 333 2353 339
rect 2497 349 2557 383
rect 2497 333 2507 349
rect 2319 315 2507 333
rect 2541 315 2557 349
rect 2319 299 2557 315
rect 2595 485 2661 493
rect 2595 451 2611 485
rect 2645 451 2661 485
rect 2595 442 2661 451
rect 2695 485 2755 527
rect 2695 451 2705 485
rect 2739 451 2755 485
rect 2595 417 2655 442
rect 2695 421 2755 451
rect 2595 383 2611 417
rect 2645 383 2655 417
rect 2595 349 2655 383
rect 2689 405 2755 421
rect 2689 371 2705 405
rect 2739 371 2755 405
rect 2689 367 2755 371
rect 2799 477 3032 493
rect 2833 459 2998 477
rect 2799 373 2833 443
rect 2595 315 2611 349
rect 2645 333 2655 349
rect 2869 421 2955 425
rect 2869 391 2904 421
rect 2869 357 2881 391
rect 2938 387 2955 421
rect 2915 357 2955 387
rect 2869 351 2955 357
rect 2998 379 3032 443
rect 2799 333 2833 339
rect 2645 315 2833 333
rect 2595 299 2833 315
rect 2393 249 2557 265
rect 2393 215 2409 249
rect 2443 215 2477 249
rect 2511 215 2557 249
rect 2393 211 2557 215
rect 2595 249 2759 265
rect 2595 215 2641 249
rect 2675 215 2709 249
rect 2743 215 2759 249
rect 2595 211 2759 215
rect 2309 177 2370 185
rect 2782 177 2843 185
rect 2893 177 2927 351
rect 2998 329 3032 345
rect 3086 479 3152 493
rect 3086 445 3102 479
rect 3136 445 3152 479
rect 3086 411 3152 445
rect 3086 377 3102 411
rect 3136 377 3152 411
rect 3086 343 3152 377
rect 3086 327 3102 343
rect 3066 309 3102 327
rect 3136 309 3152 343
rect 3066 295 3152 309
rect 2996 293 3152 295
rect 3187 479 3253 527
rect 3187 445 3203 479
rect 3237 445 3253 479
rect 3187 411 3253 445
rect 3187 377 3203 411
rect 3237 377 3253 411
rect 3187 343 3253 377
rect 3187 309 3203 343
rect 3237 309 3253 343
rect 3187 293 3253 309
rect 3288 479 3354 493
rect 3288 445 3304 479
rect 3338 445 3354 479
rect 3288 411 3354 445
rect 3288 377 3304 411
rect 3338 377 3354 411
rect 3288 343 3354 377
rect 3288 309 3304 343
rect 3338 327 3354 343
rect 3408 477 3641 493
rect 3442 459 3607 477
rect 3408 379 3442 443
rect 3485 421 3571 425
rect 3485 387 3502 421
rect 3536 391 3571 421
rect 3485 357 3525 387
rect 3559 357 3571 391
rect 3485 351 3571 357
rect 3607 373 3641 443
rect 3408 329 3442 345
rect 3338 309 3374 327
rect 3288 295 3374 309
rect 3288 293 3444 295
rect 2996 285 3100 293
rect 2996 251 3012 285
rect 3046 261 3100 285
rect 3340 285 3444 293
rect 3340 261 3394 285
rect 3046 251 3079 261
rect 2996 241 3079 251
rect 1757 117 1873 151
rect 1689 85 1723 104
rect 1540 67 1723 85
rect 1494 51 1723 67
rect 1823 116 1873 117
rect 1823 82 1831 116
rect 1865 82 1873 116
rect 1823 66 1873 82
rect 1907 116 1957 132
rect 1907 82 1915 116
rect 1949 82 1957 116
rect 1907 17 1957 82
rect 1991 117 2107 151
rect 2141 138 2175 154
rect 1991 116 2041 117
rect 1991 82 1999 116
rect 2033 82 2041 116
rect 1991 66 2041 82
rect 2209 153 2275 177
rect 2209 119 2225 153
rect 2259 119 2275 153
rect 2309 169 2547 177
rect 2309 135 2324 169
rect 2358 161 2547 169
rect 2358 143 2497 161
rect 2358 135 2370 143
rect 2141 85 2175 104
rect 2309 101 2370 135
rect 2481 127 2497 143
rect 2531 127 2547 161
rect 2309 85 2324 101
rect 2141 67 2324 85
rect 2358 67 2370 101
rect 2141 51 2370 67
rect 2404 93 2447 109
rect 2404 59 2413 93
rect 2404 17 2447 59
rect 2481 93 2547 127
rect 2481 59 2497 93
rect 2531 59 2547 93
rect 2481 51 2547 59
rect 2605 169 2843 177
rect 2605 161 2794 169
rect 2605 127 2621 161
rect 2655 143 2794 161
rect 2655 127 2671 143
rect 2605 93 2671 127
rect 2782 135 2794 143
rect 2828 135 2843 169
rect 2605 59 2621 93
rect 2655 59 2671 93
rect 2605 51 2671 59
rect 2705 93 2748 109
rect 2739 59 2748 93
rect 2705 17 2748 59
rect 2782 101 2843 135
rect 2877 153 2943 177
rect 2877 119 2893 153
rect 2927 119 2943 153
rect 2977 138 3011 154
rect 2782 67 2794 101
rect 2828 85 2843 101
rect 3045 151 3079 241
rect 3134 249 3201 259
rect 3134 215 3150 249
rect 3184 215 3201 249
rect 3134 205 3201 215
rect 3239 249 3306 259
rect 3239 215 3256 249
rect 3290 215 3306 249
rect 3239 205 3306 215
rect 3361 251 3394 261
rect 3428 251 3444 285
rect 3361 241 3444 251
rect 3361 151 3395 241
rect 3513 177 3547 351
rect 3685 485 3745 527
rect 3685 451 3701 485
rect 3735 451 3745 485
rect 3685 421 3745 451
rect 3779 485 3845 493
rect 3779 451 3795 485
rect 3829 451 3845 485
rect 3779 442 3845 451
rect 3685 405 3751 421
rect 3685 371 3701 405
rect 3735 371 3751 405
rect 3685 367 3751 371
rect 3785 417 3845 442
rect 3785 383 3795 417
rect 3829 383 3845 417
rect 3607 333 3641 339
rect 3785 349 3845 383
rect 3785 333 3795 349
rect 3607 315 3795 333
rect 3829 315 3845 349
rect 3607 299 3845 315
rect 3883 485 3949 493
rect 3883 451 3899 485
rect 3933 451 3949 485
rect 3883 442 3949 451
rect 3983 485 4043 527
rect 3983 451 3993 485
rect 4027 451 4043 485
rect 3883 417 3943 442
rect 3983 421 4043 451
rect 3883 383 3899 417
rect 3933 383 3943 417
rect 3883 349 3943 383
rect 3977 405 4043 421
rect 3977 371 3993 405
rect 4027 371 4043 405
rect 3977 367 4043 371
rect 4087 477 4320 493
rect 4121 459 4286 477
rect 4087 373 4121 443
rect 3883 315 3899 349
rect 3933 333 3943 349
rect 4157 421 4243 425
rect 4157 391 4192 421
rect 4157 357 4169 391
rect 4226 387 4243 421
rect 4203 357 4243 387
rect 4157 351 4243 357
rect 4286 379 4320 443
rect 4087 333 4121 339
rect 3933 315 4121 333
rect 3883 299 4121 315
rect 3681 249 3845 265
rect 3681 215 3697 249
rect 3731 215 3765 249
rect 3799 215 3845 249
rect 3681 211 3845 215
rect 3883 249 4047 265
rect 3883 215 3929 249
rect 3963 215 3997 249
rect 4031 215 4047 249
rect 3883 211 4047 215
rect 3597 177 3658 185
rect 4070 177 4131 185
rect 4181 177 4215 351
rect 4286 329 4320 345
rect 4374 479 4440 493
rect 4374 445 4390 479
rect 4424 445 4440 479
rect 4374 411 4440 445
rect 4374 377 4390 411
rect 4424 377 4440 411
rect 4374 343 4440 377
rect 4374 327 4390 343
rect 4354 309 4390 327
rect 4424 309 4440 343
rect 4354 295 4440 309
rect 4284 293 4440 295
rect 4475 479 4541 527
rect 4475 445 4491 479
rect 4525 445 4541 479
rect 4475 411 4541 445
rect 4475 377 4491 411
rect 4525 377 4541 411
rect 4475 343 4541 377
rect 4475 309 4491 343
rect 4525 309 4541 343
rect 4475 293 4541 309
rect 4576 479 4642 493
rect 4576 445 4592 479
rect 4626 445 4642 479
rect 4576 411 4642 445
rect 4576 377 4592 411
rect 4626 377 4642 411
rect 4576 343 4642 377
rect 4576 309 4592 343
rect 4626 327 4642 343
rect 4696 477 4929 493
rect 4730 459 4895 477
rect 4696 379 4730 443
rect 4773 421 4859 425
rect 4773 387 4790 421
rect 4824 391 4859 421
rect 4773 357 4813 387
rect 4847 357 4859 391
rect 4773 351 4859 357
rect 4895 373 4929 443
rect 4696 329 4730 345
rect 4626 309 4662 327
rect 4576 295 4662 309
rect 4576 293 4732 295
rect 4284 285 4388 293
rect 4284 251 4300 285
rect 4334 261 4388 285
rect 4628 285 4732 293
rect 4628 261 4682 285
rect 4334 251 4367 261
rect 4284 241 4367 251
rect 3045 117 3161 151
rect 2977 85 3011 104
rect 2828 67 3011 85
rect 2782 51 3011 67
rect 3111 116 3161 117
rect 3111 82 3119 116
rect 3153 82 3161 116
rect 3111 66 3161 82
rect 3195 116 3245 132
rect 3195 82 3203 116
rect 3237 82 3245 116
rect 3195 17 3245 82
rect 3279 117 3395 151
rect 3429 138 3463 154
rect 3279 116 3329 117
rect 3279 82 3287 116
rect 3321 82 3329 116
rect 3279 66 3329 82
rect 3497 153 3563 177
rect 3497 119 3513 153
rect 3547 119 3563 153
rect 3597 169 3835 177
rect 3597 135 3612 169
rect 3646 161 3835 169
rect 3646 143 3785 161
rect 3646 135 3658 143
rect 3429 85 3463 104
rect 3597 101 3658 135
rect 3769 127 3785 143
rect 3819 127 3835 161
rect 3597 85 3612 101
rect 3429 67 3612 85
rect 3646 67 3658 101
rect 3429 51 3658 67
rect 3692 93 3735 109
rect 3692 59 3701 93
rect 3692 17 3735 59
rect 3769 93 3835 127
rect 3769 59 3785 93
rect 3819 59 3835 93
rect 3769 51 3835 59
rect 3893 169 4131 177
rect 3893 161 4082 169
rect 3893 127 3909 161
rect 3943 143 4082 161
rect 3943 127 3959 143
rect 3893 93 3959 127
rect 4070 135 4082 143
rect 4116 135 4131 169
rect 3893 59 3909 93
rect 3943 59 3959 93
rect 3893 51 3959 59
rect 3993 93 4036 109
rect 4027 59 4036 93
rect 3993 17 4036 59
rect 4070 101 4131 135
rect 4165 153 4231 177
rect 4165 119 4181 153
rect 4215 119 4231 153
rect 4265 138 4299 154
rect 4070 67 4082 101
rect 4116 85 4131 101
rect 4333 151 4367 241
rect 4422 249 4489 259
rect 4422 215 4438 249
rect 4472 215 4489 249
rect 4422 205 4489 215
rect 4527 249 4594 259
rect 4527 215 4544 249
rect 4578 215 4594 249
rect 4527 205 4594 215
rect 4649 251 4682 261
rect 4716 251 4732 285
rect 4649 241 4732 251
rect 4649 151 4683 241
rect 4801 177 4835 351
rect 4973 485 5033 527
rect 4973 451 4989 485
rect 5023 451 5033 485
rect 4973 421 5033 451
rect 5067 485 5133 493
rect 5067 451 5083 485
rect 5117 451 5133 485
rect 5067 442 5133 451
rect 4973 405 5039 421
rect 4973 371 4989 405
rect 5023 371 5039 405
rect 4973 367 5039 371
rect 5073 417 5133 442
rect 5073 383 5083 417
rect 5117 383 5133 417
rect 4895 333 4929 339
rect 5073 349 5133 383
rect 5073 333 5083 349
rect 4895 315 5083 333
rect 5117 315 5133 349
rect 4895 299 5133 315
rect 4969 249 5133 265
rect 4969 215 4985 249
rect 5019 215 5053 249
rect 5087 215 5133 249
rect 4969 211 5133 215
rect 4885 177 4946 185
rect 4333 117 4449 151
rect 4265 85 4299 104
rect 4116 67 4299 85
rect 4070 51 4299 67
rect 4399 116 4449 117
rect 4399 82 4407 116
rect 4441 82 4449 116
rect 4399 66 4449 82
rect 4483 116 4533 132
rect 4483 82 4491 116
rect 4525 82 4533 116
rect 4483 17 4533 82
rect 4567 117 4683 151
rect 4717 138 4751 154
rect 4567 116 4617 117
rect 4567 82 4575 116
rect 4609 82 4617 116
rect 4567 66 4617 82
rect 4785 153 4851 177
rect 4785 119 4801 153
rect 4835 119 4851 153
rect 4885 169 5123 177
rect 4885 135 4900 169
rect 4934 161 5123 169
rect 4934 143 5073 161
rect 4934 135 4946 143
rect 4717 85 4751 104
rect 4885 101 4946 135
rect 5057 127 5073 143
rect 5107 127 5123 161
rect 4885 85 4900 101
rect 4717 67 4900 85
rect 4934 67 4946 101
rect 4717 51 4946 67
rect 4980 93 5023 109
rect 4980 59 4989 93
rect 4980 17 5023 59
rect 5057 93 5123 127
rect 5057 59 5073 93
rect 5107 59 5123 93
rect 5057 51 5123 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3341 17
rect 3375 -17 3433 17
rect 3467 -17 3525 17
rect 3559 -17 3617 17
rect 3651 -17 3709 17
rect 3743 -17 3801 17
rect 3835 -17 3893 17
rect 3927 -17 3985 17
rect 4019 -17 4077 17
rect 4111 -17 4169 17
rect 4203 -17 4261 17
rect 4295 -17 4353 17
rect 4387 -17 4445 17
rect 4479 -17 4537 17
rect 4571 -17 4629 17
rect 4663 -17 4721 17
rect 4755 -17 4813 17
rect 4847 -17 4905 17
rect 4939 -17 4997 17
rect 5031 -17 5089 17
rect 5123 -17 5152 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 2881 527 2915 561
rect 2973 527 3007 561
rect 3065 527 3099 561
rect 3157 527 3191 561
rect 3249 527 3283 561
rect 3341 527 3375 561
rect 3433 527 3467 561
rect 3525 527 3559 561
rect 3617 527 3651 561
rect 3709 527 3743 561
rect 3801 527 3835 561
rect 3893 527 3927 561
rect 3985 527 4019 561
rect 4077 527 4111 561
rect 4169 527 4203 561
rect 4261 527 4295 561
rect 4353 527 4387 561
rect 4445 527 4479 561
rect 4537 527 4571 561
rect 4629 527 4663 561
rect 4721 527 4755 561
rect 4813 527 4847 561
rect 4905 527 4939 561
rect 4997 527 5031 561
rect 5089 527 5123 561
rect 305 387 328 391
rect 328 387 339 391
rect 305 357 339 387
rect 949 387 960 391
rect 960 387 983 391
rect 949 357 983 387
rect 1593 387 1616 391
rect 1616 387 1627 391
rect 1593 357 1627 387
rect 2237 387 2248 391
rect 2248 387 2271 391
rect 2237 357 2271 387
rect 2881 387 2904 391
rect 2904 387 2915 391
rect 2881 357 2915 387
rect 3525 387 3536 391
rect 3536 387 3559 391
rect 3525 357 3559 387
rect 4169 387 4192 391
rect 4192 387 4203 391
rect 4169 357 4203 387
rect 4813 387 4824 391
rect 4824 387 4847 391
rect 4813 357 4847 387
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
rect 2881 -17 2915 17
rect 2973 -17 3007 17
rect 3065 -17 3099 17
rect 3157 -17 3191 17
rect 3249 -17 3283 17
rect 3341 -17 3375 17
rect 3433 -17 3467 17
rect 3525 -17 3559 17
rect 3617 -17 3651 17
rect 3709 -17 3743 17
rect 3801 -17 3835 17
rect 3893 -17 3927 17
rect 3985 -17 4019 17
rect 4077 -17 4111 17
rect 4169 -17 4203 17
rect 4261 -17 4295 17
rect 4353 -17 4387 17
rect 4445 -17 4479 17
rect 4537 -17 4571 17
rect 4629 -17 4663 17
rect 4721 -17 4755 17
rect 4813 -17 4847 17
rect 4905 -17 4939 17
rect 4997 -17 5031 17
rect 5089 -17 5123 17
<< metal1 >>
rect 0 561 5152 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3157 561
rect 3191 527 3249 561
rect 3283 527 3341 561
rect 3375 527 3433 561
rect 3467 527 3525 561
rect 3559 527 3617 561
rect 3651 527 3709 561
rect 3743 527 3801 561
rect 3835 527 3893 561
rect 3927 527 3985 561
rect 4019 527 4077 561
rect 4111 527 4169 561
rect 4203 527 4261 561
rect 4295 527 4353 561
rect 4387 527 4445 561
rect 4479 527 4537 561
rect 4571 527 4629 561
rect 4663 527 4721 561
rect 4755 527 4813 561
rect 4847 527 4905 561
rect 4939 527 4997 561
rect 5031 527 5089 561
rect 5123 527 5152 561
rect 0 496 5152 527
rect 293 391 351 397
rect 293 357 305 391
rect 339 388 351 391
rect 937 391 995 397
rect 937 388 949 391
rect 339 360 949 388
rect 339 357 351 360
rect 293 351 351 357
rect 937 357 949 360
rect 983 388 995 391
rect 1581 391 1639 397
rect 1581 388 1593 391
rect 983 360 1593 388
rect 983 357 995 360
rect 937 351 995 357
rect 1581 357 1593 360
rect 1627 388 1639 391
rect 2225 391 2283 397
rect 2225 388 2237 391
rect 1627 360 2237 388
rect 1627 357 1639 360
rect 1581 351 1639 357
rect 2225 357 2237 360
rect 2271 388 2283 391
rect 2869 391 2927 397
rect 2869 388 2881 391
rect 2271 360 2881 388
rect 2271 357 2283 360
rect 2225 351 2283 357
rect 2869 357 2881 360
rect 2915 388 2927 391
rect 3513 391 3571 397
rect 3513 388 3525 391
rect 2915 360 3525 388
rect 2915 357 2927 360
rect 2869 351 2927 357
rect 3513 357 3525 360
rect 3559 388 3571 391
rect 4157 391 4215 397
rect 4157 388 4169 391
rect 3559 360 4169 388
rect 3559 357 3571 360
rect 3513 351 3571 357
rect 4157 357 4169 360
rect 4203 388 4215 391
rect 4801 391 4859 397
rect 4801 388 4813 391
rect 4203 360 4813 388
rect 4203 357 4215 360
rect 4157 351 4215 357
rect 4801 357 4813 360
rect 4847 357 4859 391
rect 4801 351 4859 357
rect 0 17 5152 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3341 17
rect 3375 -17 3433 17
rect 3467 -17 3525 17
rect 3559 -17 3617 17
rect 3651 -17 3709 17
rect 3743 -17 3801 17
rect 3835 -17 3893 17
rect 3927 -17 3985 17
rect 4019 -17 4077 17
rect 4111 -17 4169 17
rect 4203 -17 4261 17
rect 4295 -17 4353 17
rect 4387 -17 4445 17
rect 4479 -17 4537 17
rect 4571 -17 4629 17
rect 4663 -17 4721 17
rect 4755 -17 4813 17
rect 4847 -17 4905 17
rect 4939 -17 4997 17
rect 5031 -17 5089 17
rect 5123 -17 5152 17
rect 0 -48 5152 -17
<< labels >>
rlabel comment s 0 0 0 0 4 muxb8to1_2
flabel metal1 s 305 357 339 391 0 FreeSans 200 0 0 0 Z
port 21 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 17 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 20 nsew
flabel metal1 s 2605 -17 2639 17 0 FreeSans 200 0 0 0 VGND
port 17 nsew
flabel metal1 s 2605 527 2639 561 0 FreeSans 200 0 0 0 VPWR
port 20 nsew
flabel metal1 s 2513 -17 2547 17 0 FreeSans 200 180 0 0 VGND
port 17 nsew
flabel metal1 s 2513 527 2547 561 0 FreeSans 200 180 0 0 VPWR
port 20 nsew
flabel metal1 s 1317 -17 1351 17 0 FreeSans 200 0 0 0 VGND
port 17 nsew
flabel metal1 s 1317 527 1351 561 0 FreeSans 200 0 0 0 VPWR
port 20 nsew
flabel metal1 s 1225 -17 1259 17 0 FreeSans 200 180 0 0 VGND
port 17 nsew
flabel metal1 s 1225 527 1259 561 0 FreeSans 200 180 0 0 VPWR
port 20 nsew
flabel metal1 s 46 0 46 0 0 FreeSans 200 0 0 0 VGND
port 17 nsew
flabel metal1 s 46 544 46 544 0 FreeSans 200 0 0 0 VPWR
port 20 nsew
flabel metal1 s 3801 527 3835 561 0 FreeSans 200 180 0 0 VPWR
port 20 nsew
flabel metal1 s 3801 -17 3835 17 0 FreeSans 200 180 0 0 VGND
port 17 nsew
flabel metal1 s 3893 527 3927 561 0 FreeSans 200 0 0 0 VPWR
port 20 nsew
flabel metal1 s 3893 -17 3927 17 0 FreeSans 200 0 0 0 VGND
port 17 nsew
flabel metal1 s 5089 527 5123 561 0 FreeSans 200 180 0 0 VPWR
port 20 nsew
flabel metal1 s 5089 -17 5123 17 0 FreeSans 200 180 0 0 VGND
port 17 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 18 nsew
flabel pwell s 2605 -17 2639 17 0 FreeSans 200 0 0 0 VNB
port 18 nsew
flabel pwell s 2513 -17 2547 17 0 FreeSans 200 180 0 0 VNB
port 18 nsew
flabel pwell s 1317 -17 1351 17 0 FreeSans 200 0 0 0 VNB
port 18 nsew
flabel pwell s 1225 -17 1259 17 0 FreeSans 200 180 0 0 VNB
port 18 nsew
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
port 18 nsew
flabel pwell s 3801 -17 3835 17 0 FreeSans 200 180 0 0 VNB
port 18 nsew
flabel pwell s 3893 -17 3927 17 0 FreeSans 200 0 0 0 VNB
port 18 nsew
flabel pwell s 5089 -17 5123 17 0 FreeSans 200 180 0 0 VNB
port 18 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 19 nsew
flabel nbase s 2605 527 2639 561 0 FreeSans 200 0 0 0 VPB
port 19 nsew
flabel nbase s 2513 527 2547 561 0 FreeSans 200 180 0 0 VPB
port 19 nsew
flabel nbase s 1317 527 1351 561 0 FreeSans 200 0 0 0 VPB
port 19 nsew
flabel nbase s 1225 527 1259 561 0 FreeSans 200 180 0 0 VPB
port 19 nsew
flabel nbase s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
port 19 nsew
flabel nbase s 3801 527 3835 561 0 FreeSans 200 180 0 0 VPB
port 19 nsew
flabel nbase s 3893 527 3927 561 0 FreeSans 200 0 0 0 VPB
port 19 nsew
flabel nbase s 5089 527 5123 561 0 FreeSans 200 180 0 0 VPB
port 19 nsew
flabel corelocali s 1317 221 1351 255 0 FreeSans 200 0 0 0 D[2]
port 6 nsew
flabel corelocali s 1225 221 1259 255 0 FreeSans 200 0 0 0 D[1]
port 7 nsew
flabel corelocali s 4537 221 4571 255 0 FreeSans 200 0 0 0 S[7]
port 9 nsew
flabel corelocali s 4445 221 4479 255 0 FreeSans 200 0 0 0 S[6]
port 10 nsew
flabel corelocali s 3249 221 3283 255 0 FreeSans 200 0 0 0 S[5]
port 11 nsew
flabel corelocali s 3157 221 3191 255 0 FreeSans 200 0 0 0 S[4]
port 12 nsew
flabel corelocali s 1961 221 1995 255 0 FreeSans 200 0 0 0 S[3]
port 13 nsew
flabel corelocali s 1869 221 1903 255 0 FreeSans 200 0 0 0 S[2]
port 14 nsew
flabel corelocali s 673 221 707 255 0 FreeSans 200 0 0 0 S[1]
port 15 nsew
flabel corelocali s 581 221 615 255 0 FreeSans 200 0 0 0 S[0]
port 16 nsew
flabel corelocali s 5089 221 5123 255 0 FreeSans 200 0 0 0 D[7]
port 1 nsew
flabel corelocali s 3893 221 3927 255 0 FreeSans 200 0 0 0 D[6]
port 2 nsew
flabel corelocali s 3801 221 3835 255 0 FreeSans 200 0 0 0 D[5]
port 3 nsew
flabel corelocali s 2605 221 2639 255 0 FreeSans 200 0 0 0 D[4]
port 4 nsew
flabel corelocali s 2513 221 2547 255 0 FreeSans 200 0 0 0 D[3]
port 5 nsew
flabel corelocali s 29 221 63 255 0 FreeSans 200 0 0 0 D[0]
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 5152 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2893436
string GDS_START 2834862
<< end >>
