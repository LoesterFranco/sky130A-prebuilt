magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 1359 424 1393 547
rect 1539 424 1579 547
rect 1359 390 1579 424
rect 25 270 455 356
rect 501 270 771 356
rect 889 260 1223 356
rect 1273 270 1511 356
rect 1545 236 1703 390
rect 1264 226 1703 236
rect 514 202 1703 226
rect 514 192 1298 202
rect 514 157 752 192
rect 1076 70 1126 192
rect 1264 70 1298 192
rect 1436 70 1703 202
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 69 424 135 596
rect 175 458 209 649
rect 249 424 299 596
rect 339 458 405 649
rect 445 424 479 596
rect 519 458 585 649
rect 625 424 659 596
rect 699 458 765 649
rect 805 424 855 596
rect 893 581 1679 615
rect 893 458 959 581
rect 999 424 1033 547
rect 1073 458 1139 581
rect 1179 424 1229 547
rect 69 390 1229 424
rect 1263 390 1319 581
rect 1433 458 1499 581
rect 1613 424 1679 581
rect 805 364 855 390
rect 84 202 478 236
rect 84 70 134 202
rect 170 17 236 168
rect 272 70 306 202
rect 342 17 408 168
rect 444 123 478 202
rect 444 70 838 123
rect 1162 17 1228 158
rect 1334 17 1400 168
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
<< metal1 >>
rect 0 683 1728 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 0 617 1728 649
rect 0 17 1728 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
rect 0 -49 1728 -17
<< labels >>
rlabel locali s 501 270 771 356 6 A1
port 1 nsew signal input
rlabel locali s 25 270 455 356 6 A2
port 2 nsew signal input
rlabel locali s 889 260 1223 356 6 B1
port 3 nsew signal input
rlabel locali s 1273 270 1511 356 6 C1
port 4 nsew signal input
rlabel locali s 1545 236 1703 390 6 Y
port 5 nsew signal output
rlabel locali s 1539 424 1579 547 6 Y
port 5 nsew signal output
rlabel locali s 1436 70 1703 202 6 Y
port 5 nsew signal output
rlabel locali s 1359 424 1393 547 6 Y
port 5 nsew signal output
rlabel locali s 1359 390 1579 424 6 Y
port 5 nsew signal output
rlabel locali s 1264 226 1703 236 6 Y
port 5 nsew signal output
rlabel locali s 1264 70 1298 192 6 Y
port 5 nsew signal output
rlabel locali s 1076 70 1126 192 6 Y
port 5 nsew signal output
rlabel locali s 514 202 1703 226 6 Y
port 5 nsew signal output
rlabel locali s 514 192 1298 202 6 Y
port 5 nsew signal output
rlabel locali s 514 157 752 192 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -49 1728 49 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1728 715 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1728 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 4071700
string GDS_START 4057012
<< end >>
