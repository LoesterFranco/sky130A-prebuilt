magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1012 561
rect 19 305 78 493
rect 198 305 250 493
rect 284 347 336 492
rect 370 381 422 493
rect 456 347 508 492
rect 542 381 594 493
rect 628 347 680 492
rect 714 381 766 493
rect 800 347 852 492
rect 886 381 945 493
rect 284 299 946 347
rect 17 143 80 265
rect 29 17 78 109
rect 752 181 946 299
rect 284 147 946 181
rect 198 17 250 122
rect 284 56 336 147
rect 370 17 422 113
rect 456 56 508 147
rect 542 17 594 113
rect 628 56 680 147
rect 714 17 766 113
rect 800 56 852 147
rect 886 17 946 113
rect 0 -17 1012 17
<< obsli1 >>
rect 114 265 164 492
rect 114 215 718 265
rect 114 53 164 215
<< metal1 >>
rect 0 496 1012 592
rect 14 428 998 468
rect 23 416 81 428
rect 195 416 253 428
rect 366 416 424 428
rect 536 416 594 428
rect 712 416 770 428
rect 884 416 942 428
rect 0 -48 1012 48
<< labels >>
rlabel locali s 17 143 80 265 6 A
port 1 nsew signal input
rlabel locali s 800 347 852 492 6 X
port 2 nsew signal output
rlabel locali s 800 56 852 147 6 X
port 2 nsew signal output
rlabel locali s 752 181 946 299 6 X
port 2 nsew signal output
rlabel locali s 628 347 680 492 6 X
port 2 nsew signal output
rlabel locali s 628 56 680 147 6 X
port 2 nsew signal output
rlabel locali s 456 347 508 492 6 X
port 2 nsew signal output
rlabel locali s 456 56 508 147 6 X
port 2 nsew signal output
rlabel locali s 284 347 336 492 6 X
port 2 nsew signal output
rlabel locali s 284 299 946 347 6 X
port 2 nsew signal output
rlabel locali s 284 147 946 181 6 X
port 2 nsew signal output
rlabel locali s 284 56 336 147 6 X
port 2 nsew signal output
rlabel locali s 19 305 78 493 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 198 305 250 493 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 370 381 422 493 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 542 381 594 493 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 714 381 766 493 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 886 381 945 493 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 884 416 942 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 712 416 770 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 536 416 594 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 366 416 424 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 195 416 253 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 23 416 81 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 14 428 998 468 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel locali s 886 17 946 113 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 714 17 766 113 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 542 17 594 113 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 370 17 422 113 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 198 17 250 122 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 29 17 78 109 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 1012 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1012 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 527 1012 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 1012 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1012 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2183900
string GDS_START 2175056
<< end >>
