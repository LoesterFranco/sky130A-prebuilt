magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1472 561
rect 27 149 70 325
rect 459 451 525 527
rect 627 451 693 527
rect 795 451 861 527
rect 963 451 1035 527
rect 1143 451 1209 527
rect 1387 359 1454 527
rect 212 257 251 325
rect 543 309 777 343
rect 212 215 301 257
rect 582 177 621 309
rect 903 215 989 257
rect 1051 215 1208 257
rect 459 143 661 177
rect 19 17 69 113
rect 203 17 237 109
rect 371 17 405 109
rect 459 93 493 143
rect 439 59 509 93
rect 543 17 577 109
rect 627 93 661 143
rect 611 59 677 93
rect 711 17 813 109
rect 955 17 989 109
rect 1389 215 1455 323
rect 0 -17 1472 17
<< obsli1 >>
rect 35 459 405 493
rect 35 359 69 459
rect 103 391 169 425
rect 119 177 153 391
rect 203 359 237 459
rect 287 325 321 425
rect 371 359 405 459
rect 895 417 929 493
rect 1075 417 1109 493
rect 1319 417 1353 493
rect 439 383 1353 417
rect 439 325 477 383
rect 895 359 929 383
rect 1075 359 1109 383
rect 1319 359 1353 383
rect 287 291 477 325
rect 371 215 541 249
rect 371 177 405 215
rect 830 291 1337 325
rect 830 249 864 291
rect 655 215 864 249
rect 119 143 405 177
rect 119 93 153 143
rect 103 59 169 93
rect 287 93 321 143
rect 271 59 337 93
rect 871 143 1201 177
rect 871 93 905 143
rect 1135 129 1201 143
rect 855 59 921 93
rect 1235 93 1269 177
rect 1303 165 1337 291
rect 1303 129 1369 165
rect 1403 100 1454 181
rect 1051 85 1269 93
rect 1387 85 1454 100
rect 1051 51 1454 85
<< metal1 >>
rect 0 496 1472 592
rect 0 -48 1472 48
<< labels >>
rlabel locali s 1389 215 1455 323 6 A1
port 1 nsew signal input
rlabel locali s 1051 215 1208 257 6 A2
port 2 nsew signal input
rlabel locali s 903 215 989 257 6 A3
port 3 nsew signal input
rlabel locali s 212 257 251 325 6 B1
port 4 nsew signal input
rlabel locali s 212 215 301 257 6 B1
port 4 nsew signal input
rlabel locali s 27 149 70 325 6 C1
port 5 nsew signal input
rlabel locali s 627 93 661 143 6 X
port 6 nsew signal output
rlabel locali s 611 59 677 93 6 X
port 6 nsew signal output
rlabel locali s 582 177 621 309 6 X
port 6 nsew signal output
rlabel locali s 543 309 777 343 6 X
port 6 nsew signal output
rlabel locali s 459 143 661 177 6 X
port 6 nsew signal output
rlabel locali s 459 93 493 143 6 X
port 6 nsew signal output
rlabel locali s 439 59 509 93 6 X
port 6 nsew signal output
rlabel locali s 955 17 989 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 711 17 813 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 543 17 577 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 371 17 405 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 203 17 237 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 19 17 69 113 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 1472 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1472 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1387 359 1454 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1143 451 1209 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 963 451 1035 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 795 451 861 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 627 451 693 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 459 451 525 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 1472 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 1472 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1472 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3613270
string GDS_START 3601548
<< end >>
