magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 828 561
rect 150 370 198 527
rect 17 195 69 265
rect 300 255 358 341
rect 177 215 246 255
rect 280 215 358 255
rect 396 257 457 341
rect 559 359 625 527
rect 659 409 709 493
rect 743 443 811 527
rect 659 375 811 409
rect 396 215 493 257
rect 527 215 615 257
rect 749 181 811 375
rect 423 17 457 111
rect 591 17 625 181
rect 659 147 811 181
rect 659 53 725 147
rect 759 17 793 113
rect 0 -17 828 17
<< obsli1 >>
rect 50 334 116 493
rect 310 409 461 493
rect 232 375 525 409
rect 232 334 266 375
rect 50 299 266 334
rect 109 289 266 299
rect 109 161 143 289
rect 491 325 525 375
rect 491 291 683 325
rect 649 257 683 291
rect 649 215 715 257
rect 34 127 143 161
rect 217 147 557 181
rect 217 129 294 147
rect 34 51 100 127
rect 134 59 371 93
rect 491 54 557 147
<< metal1 >>
rect 0 496 828 592
rect 0 -48 828 48
<< labels >>
rlabel locali s 527 215 615 257 6 A1
port 1 nsew signal input
rlabel locali s 396 257 457 341 6 A2
port 2 nsew signal input
rlabel locali s 396 215 493 257 6 A2
port 2 nsew signal input
rlabel locali s 177 215 246 255 6 B1
port 3 nsew signal input
rlabel locali s 300 255 358 341 6 B2
port 4 nsew signal input
rlabel locali s 280 215 358 255 6 B2
port 4 nsew signal input
rlabel locali s 17 195 69 265 6 C1
port 5 nsew signal input
rlabel locali s 749 181 811 375 6 X
port 6 nsew signal output
rlabel locali s 659 409 709 493 6 X
port 6 nsew signal output
rlabel locali s 659 375 811 409 6 X
port 6 nsew signal output
rlabel locali s 659 147 811 181 6 X
port 6 nsew signal output
rlabel locali s 659 53 725 147 6 X
port 6 nsew signal output
rlabel locali s 759 17 793 113 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 591 17 625 181 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 423 17 457 111 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 828 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 828 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 743 443 811 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 559 359 625 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 150 370 198 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 828 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 828 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1427202
string GDS_START 1419732
<< end >>
