magic
tech sky130A
magscale 1 2
timestamp 1604502705
<< nwell >>
rect -38 332 2918 704
<< pwell >>
rect 0 0 2880 49
<< scnmos >>
rect 84 74 114 222
rect 170 74 200 222
rect 368 119 398 203
rect 499 119 529 203
rect 571 119 601 203
rect 657 119 687 203
rect 924 125 954 235
rect 1010 125 1040 235
rect 1110 125 1140 235
rect 1210 125 1240 235
rect 1305 112 1335 222
rect 1610 138 1640 222
rect 1688 138 1718 222
rect 1802 74 1832 222
rect 1888 74 1918 222
rect 1982 74 2012 222
rect 2193 164 2223 248
rect 2301 100 2331 248
rect 2387 100 2417 248
rect 2588 74 2618 202
rect 2683 74 2713 222
rect 2769 74 2799 222
<< pmoshvt >>
rect 84 368 114 592
rect 174 368 204 592
rect 387 503 417 587
rect 506 503 536 587
rect 590 503 620 587
rect 692 503 722 587
rect 900 424 930 592
rect 984 424 1014 592
rect 1086 424 1116 592
rect 1282 424 1312 592
rect 1366 424 1396 592
rect 1474 508 1504 592
rect 1558 508 1588 592
rect 1777 392 1807 592
rect 1901 392 1931 592
rect 1985 392 2015 592
rect 2181 368 2211 496
rect 2286 368 2316 592
rect 2376 368 2406 592
rect 2572 368 2602 568
rect 2676 368 2706 592
rect 2766 368 2796 592
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 142 170 222
rect 114 108 125 142
rect 159 108 170 142
rect 114 74 170 108
rect 200 210 257 222
rect 200 176 211 210
rect 245 176 257 210
rect 200 120 257 176
rect 200 86 211 120
rect 245 86 257 120
rect 311 175 368 203
rect 311 141 323 175
rect 357 141 368 175
rect 311 119 368 141
rect 398 134 499 203
rect 398 119 431 134
rect 413 100 431 119
rect 465 119 499 134
rect 529 119 571 203
rect 601 172 657 203
rect 601 138 612 172
rect 646 138 657 172
rect 601 119 657 138
rect 687 123 813 203
rect 867 173 924 235
rect 867 139 879 173
rect 913 139 924 173
rect 867 125 924 139
rect 954 189 1010 235
rect 954 155 965 189
rect 999 155 1010 189
rect 954 125 1010 155
rect 1040 189 1110 235
rect 1040 155 1065 189
rect 1099 155 1110 189
rect 1040 125 1110 155
rect 1140 189 1210 235
rect 1140 155 1165 189
rect 1199 155 1210 189
rect 1140 125 1210 155
rect 1240 222 1290 235
rect 2137 236 2193 248
rect 1240 125 1305 222
rect 687 119 740 123
rect 465 100 484 119
rect 413 88 484 100
rect 200 74 257 86
rect 702 89 740 119
rect 774 89 813 123
rect 1255 112 1305 125
rect 1335 186 1610 222
rect 1335 152 1346 186
rect 1380 152 1419 186
rect 1453 152 1492 186
rect 1526 152 1565 186
rect 1599 152 1610 186
rect 1335 138 1610 152
rect 1640 138 1688 222
rect 1718 138 1802 222
rect 1335 112 1385 138
rect 1745 136 1802 138
rect 702 77 813 89
rect 1745 102 1757 136
rect 1791 102 1802 136
rect 1745 74 1802 102
rect 1832 136 1888 222
rect 1832 102 1843 136
rect 1877 102 1888 136
rect 1832 74 1888 102
rect 1918 160 1982 222
rect 1918 126 1937 160
rect 1971 126 1982 160
rect 1918 74 1982 126
rect 2012 100 2083 222
rect 2137 202 2148 236
rect 2182 202 2193 236
rect 2137 164 2193 202
rect 2223 164 2301 248
rect 2251 100 2301 164
rect 2331 220 2387 248
rect 2331 186 2342 220
rect 2376 186 2387 220
rect 2331 146 2387 186
rect 2331 112 2342 146
rect 2376 112 2387 146
rect 2331 100 2387 112
rect 2417 236 2477 248
rect 2417 202 2431 236
rect 2465 202 2477 236
rect 2633 202 2683 222
rect 2417 146 2477 202
rect 2417 112 2431 146
rect 2465 112 2477 146
rect 2417 100 2477 112
rect 2531 194 2588 202
rect 2531 160 2543 194
rect 2577 160 2588 194
rect 2531 120 2588 160
rect 2012 74 2038 100
rect 2027 66 2038 74
rect 2072 66 2083 100
rect 2027 54 2083 66
rect 2137 84 2286 100
rect 2137 50 2149 84
rect 2183 50 2240 84
rect 2274 50 2286 84
rect 2531 86 2543 120
rect 2577 86 2588 120
rect 2531 74 2588 86
rect 2618 194 2683 202
rect 2618 160 2635 194
rect 2669 160 2683 194
rect 2618 116 2683 160
rect 2618 82 2635 116
rect 2669 82 2683 116
rect 2618 74 2683 82
rect 2713 204 2769 222
rect 2713 170 2724 204
rect 2758 170 2769 204
rect 2713 120 2769 170
rect 2713 86 2724 120
rect 2758 86 2769 120
rect 2713 74 2769 86
rect 2799 120 2853 222
rect 2799 86 2810 120
rect 2844 86 2853 120
rect 2799 74 2853 86
rect 2137 38 2286 50
<< pdiff >>
rect 1606 628 1664 639
rect 27 580 84 592
rect 27 546 37 580
rect 71 546 84 580
rect 27 510 84 546
rect 27 476 37 510
rect 71 476 84 510
rect 27 440 84 476
rect 27 406 37 440
rect 71 406 84 440
rect 27 368 84 406
rect 114 580 174 592
rect 114 546 127 580
rect 161 546 174 580
rect 114 508 174 546
rect 114 474 127 508
rect 161 474 174 508
rect 114 368 174 474
rect 204 580 260 592
rect 1606 594 1618 628
rect 1652 594 1664 628
rect 1825 628 1883 639
rect 1606 592 1664 594
rect 1825 594 1837 628
rect 1871 594 1883 628
rect 1825 592 1883 594
rect 204 546 217 580
rect 251 546 260 580
rect 204 497 260 546
rect 204 463 217 497
rect 251 463 260 497
rect 314 531 387 587
rect 314 497 323 531
rect 357 503 387 531
rect 417 565 506 587
rect 417 531 459 565
rect 493 531 506 565
rect 417 503 506 531
rect 536 503 590 587
rect 620 547 692 587
rect 620 513 639 547
rect 673 513 692 547
rect 620 503 692 513
rect 722 531 790 587
rect 722 503 748 531
rect 357 497 369 503
rect 314 485 369 497
rect 740 497 748 503
rect 782 497 790 531
rect 204 414 260 463
rect 204 380 217 414
rect 251 380 260 414
rect 204 368 260 380
rect 740 485 790 497
rect 844 580 900 592
rect 844 546 853 580
rect 887 546 900 580
rect 844 495 900 546
rect 844 461 853 495
rect 887 461 900 495
rect 844 424 900 461
rect 930 424 984 592
rect 1014 573 1086 592
rect 1014 539 1027 573
rect 1061 539 1086 573
rect 1014 424 1086 539
rect 1116 580 1172 592
rect 1116 546 1129 580
rect 1163 546 1172 580
rect 1116 498 1172 546
rect 1116 464 1129 498
rect 1163 464 1172 498
rect 1116 424 1172 464
rect 1226 573 1282 592
rect 1226 539 1235 573
rect 1269 539 1282 573
rect 1226 424 1282 539
rect 1312 424 1366 592
rect 1396 580 1474 592
rect 1396 546 1409 580
rect 1443 546 1474 580
rect 1396 508 1474 546
rect 1504 508 1558 592
rect 1588 508 1664 592
rect 1718 578 1777 592
rect 1718 544 1730 578
rect 1764 544 1777 578
rect 1396 470 1455 508
rect 1396 436 1409 470
rect 1443 436 1455 470
rect 1396 424 1455 436
rect 1718 392 1777 544
rect 1807 392 1901 592
rect 1931 392 1985 592
rect 2015 580 2071 592
rect 2015 546 2028 580
rect 2062 546 2071 580
rect 2015 508 2071 546
rect 2229 578 2286 592
rect 2229 544 2239 578
rect 2273 544 2286 578
rect 2015 474 2028 508
rect 2062 474 2071 508
rect 2229 496 2286 544
rect 2015 392 2071 474
rect 2125 424 2181 496
rect 2125 390 2134 424
rect 2168 390 2181 424
rect 2125 368 2181 390
rect 2211 368 2286 496
rect 2316 580 2376 592
rect 2316 546 2329 580
rect 2363 546 2376 580
rect 2316 500 2376 546
rect 2316 466 2329 500
rect 2363 466 2376 500
rect 2316 420 2376 466
rect 2316 386 2329 420
rect 2363 386 2376 420
rect 2316 368 2376 386
rect 2406 580 2462 592
rect 2406 546 2419 580
rect 2453 546 2462 580
rect 2620 568 2676 592
rect 2406 488 2462 546
rect 2406 454 2419 488
rect 2453 454 2462 488
rect 2406 368 2462 454
rect 2516 556 2572 568
rect 2516 522 2525 556
rect 2559 522 2572 556
rect 2516 485 2572 522
rect 2516 451 2525 485
rect 2559 451 2572 485
rect 2516 414 2572 451
rect 2516 380 2525 414
rect 2559 380 2572 414
rect 2516 368 2572 380
rect 2602 556 2676 568
rect 2602 522 2629 556
rect 2663 522 2676 556
rect 2602 485 2676 522
rect 2602 451 2629 485
rect 2663 451 2676 485
rect 2602 414 2676 451
rect 2602 380 2629 414
rect 2663 380 2676 414
rect 2602 368 2676 380
rect 2706 580 2766 592
rect 2706 546 2719 580
rect 2753 546 2766 580
rect 2706 497 2766 546
rect 2706 463 2719 497
rect 2753 463 2766 497
rect 2706 414 2766 463
rect 2706 380 2719 414
rect 2753 380 2766 414
rect 2706 368 2766 380
rect 2796 580 2853 592
rect 2796 546 2809 580
rect 2843 546 2853 580
rect 2796 472 2853 546
rect 2796 438 2809 472
rect 2843 438 2853 472
rect 2796 368 2853 438
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 125 108 159 142
rect 211 176 245 210
rect 211 86 245 120
rect 323 141 357 175
rect 431 100 465 134
rect 612 138 646 172
rect 879 139 913 173
rect 965 155 999 189
rect 1065 155 1099 189
rect 1165 155 1199 189
rect 740 89 774 123
rect 1346 152 1380 186
rect 1419 152 1453 186
rect 1492 152 1526 186
rect 1565 152 1599 186
rect 1757 102 1791 136
rect 1843 102 1877 136
rect 1937 126 1971 160
rect 2148 202 2182 236
rect 2342 186 2376 220
rect 2342 112 2376 146
rect 2431 202 2465 236
rect 2431 112 2465 146
rect 2543 160 2577 194
rect 2038 66 2072 100
rect 2149 50 2183 84
rect 2240 50 2274 84
rect 2543 86 2577 120
rect 2635 160 2669 194
rect 2635 82 2669 116
rect 2724 170 2758 204
rect 2724 86 2758 120
rect 2810 86 2844 120
<< pdiffc >>
rect 37 546 71 580
rect 37 476 71 510
rect 37 406 71 440
rect 127 546 161 580
rect 127 474 161 508
rect 1618 594 1652 628
rect 1837 594 1871 628
rect 217 546 251 580
rect 217 463 251 497
rect 323 497 357 531
rect 459 531 493 565
rect 639 513 673 547
rect 748 497 782 531
rect 217 380 251 414
rect 853 546 887 580
rect 853 461 887 495
rect 1027 539 1061 573
rect 1129 546 1163 580
rect 1129 464 1163 498
rect 1235 539 1269 573
rect 1409 546 1443 580
rect 1730 544 1764 578
rect 1409 436 1443 470
rect 2028 546 2062 580
rect 2239 544 2273 578
rect 2028 474 2062 508
rect 2134 390 2168 424
rect 2329 546 2363 580
rect 2329 466 2363 500
rect 2329 386 2363 420
rect 2419 546 2453 580
rect 2419 454 2453 488
rect 2525 522 2559 556
rect 2525 451 2559 485
rect 2525 380 2559 414
rect 2629 522 2663 556
rect 2629 451 2663 485
rect 2629 380 2663 414
rect 2719 546 2753 580
rect 2719 463 2753 497
rect 2719 380 2753 414
rect 2809 546 2843 580
rect 2809 438 2843 472
<< poly >>
rect 84 592 114 618
rect 174 592 204 618
rect 387 587 417 613
rect 506 587 536 613
rect 590 587 620 613
rect 692 587 722 613
rect 900 592 930 618
rect 984 592 1014 618
rect 1086 592 1116 618
rect 1282 592 1312 618
rect 1366 592 1396 618
rect 1474 592 1504 618
rect 1558 592 1588 618
rect 1777 592 1807 618
rect 1901 592 1931 618
rect 1985 592 2015 618
rect 2286 592 2316 618
rect 2376 592 2406 618
rect 387 488 417 503
rect 506 488 536 503
rect 590 488 620 503
rect 692 488 722 503
rect 84 353 114 368
rect 174 353 204 368
rect 81 326 117 353
rect 171 326 207 353
rect 33 310 117 326
rect 33 276 49 310
rect 83 276 117 310
rect 33 260 117 276
rect 159 310 225 326
rect 159 276 175 310
rect 209 276 225 310
rect 384 302 420 488
rect 503 471 539 488
rect 587 471 623 488
rect 473 455 539 471
rect 473 421 489 455
rect 523 421 539 455
rect 473 405 539 421
rect 581 455 647 471
rect 581 421 597 455
rect 631 421 647 455
rect 581 405 647 421
rect 159 260 225 276
rect 368 286 457 302
rect 84 222 114 260
rect 170 222 200 260
rect 368 252 407 286
rect 441 252 457 286
rect 368 236 457 252
rect 368 203 398 236
rect 499 203 529 405
rect 689 363 725 488
rect 1474 493 1504 508
rect 1558 493 1588 508
rect 900 409 930 424
rect 984 409 1014 424
rect 1086 409 1116 424
rect 1282 409 1312 424
rect 1366 409 1396 424
rect 571 333 725 363
rect 897 359 933 409
rect 981 388 1017 409
rect 1083 392 1119 409
rect 1279 392 1315 409
rect 767 343 933 359
rect 571 203 601 333
rect 767 309 783 343
rect 817 309 933 343
rect 975 372 1041 388
rect 975 338 991 372
rect 1025 338 1041 372
rect 975 322 1041 338
rect 1083 376 1149 392
rect 1083 342 1099 376
rect 1133 342 1149 376
rect 1083 326 1149 342
rect 1210 376 1315 392
rect 1363 382 1399 409
rect 1471 388 1507 493
rect 1555 476 1591 493
rect 1555 460 1681 476
rect 1555 426 1601 460
rect 1635 426 1681 460
rect 1555 410 1681 426
rect 1210 342 1226 376
rect 1260 342 1315 376
rect 1210 326 1315 342
rect 1357 366 1423 382
rect 1357 332 1373 366
rect 1407 332 1423 366
rect 767 293 933 309
rect 643 275 709 291
rect 643 241 659 275
rect 693 241 709 275
rect 903 280 933 293
rect 903 250 954 280
rect 643 225 709 241
rect 924 235 954 250
rect 1010 235 1040 322
rect 1110 235 1140 326
rect 1210 235 1240 326
rect 1357 316 1423 332
rect 1465 358 1507 388
rect 1651 377 1681 410
rect 2181 496 2211 522
rect 1777 377 1807 392
rect 1901 377 1931 392
rect 1985 377 2015 392
rect 1465 267 1495 358
rect 1651 347 1718 377
rect 1774 356 1810 377
rect 1305 237 1495 267
rect 1537 294 1603 310
rect 1537 260 1553 294
rect 1587 274 1603 294
rect 1587 260 1640 274
rect 1537 244 1640 260
rect 657 203 687 225
rect 368 93 398 119
rect 1305 222 1335 237
rect 1610 222 1640 244
rect 1688 222 1718 347
rect 1766 340 1832 356
rect 1766 306 1782 340
rect 1816 306 1832 340
rect 1898 310 1934 377
rect 1982 360 2018 377
rect 2572 568 2602 594
rect 2676 592 2706 618
rect 2766 592 2796 618
rect 1982 344 2048 360
rect 2181 353 2211 368
rect 2286 353 2316 368
rect 2376 353 2406 368
rect 2572 353 2602 368
rect 2676 353 2706 368
rect 2766 353 2796 368
rect 1982 310 1998 344
rect 2032 310 2048 344
rect 2178 336 2214 353
rect 2283 336 2319 353
rect 2373 336 2409 353
rect 2569 336 2605 353
rect 1766 290 1832 306
rect 1802 222 1832 290
rect 1874 294 1940 310
rect 1874 260 1890 294
rect 1924 260 1940 294
rect 1874 244 1940 260
rect 1982 294 2048 310
rect 2157 320 2223 336
rect 1888 222 1918 244
rect 1982 222 2012 294
rect 2157 286 2173 320
rect 2207 286 2223 320
rect 2157 270 2223 286
rect 2265 320 2605 336
rect 2265 286 2281 320
rect 2315 300 2605 320
rect 2673 320 2709 353
rect 2763 320 2799 353
rect 2673 304 2799 320
rect 2315 286 2618 300
rect 2265 270 2618 286
rect 2193 248 2223 270
rect 2301 248 2331 270
rect 2387 248 2417 270
rect 499 93 529 119
rect 84 48 114 74
rect 170 51 200 74
rect 571 51 601 119
rect 657 93 687 119
rect 924 99 954 125
rect 1010 99 1040 125
rect 1110 99 1140 125
rect 1210 99 1240 125
rect 1610 112 1640 138
rect 1688 112 1718 138
rect 1305 51 1335 112
rect 2193 138 2223 164
rect 2588 202 2618 270
rect 2673 270 2689 304
rect 2723 270 2799 304
rect 2673 254 2799 270
rect 2683 222 2713 254
rect 2769 222 2799 254
rect 170 21 1335 51
rect 1802 48 1832 74
rect 1888 48 1918 74
rect 1982 48 2012 74
rect 2301 74 2331 100
rect 2387 74 2417 100
rect 2588 48 2618 74
rect 2683 48 2713 74
rect 2769 48 2799 74
<< polycont >>
rect 49 276 83 310
rect 175 276 209 310
rect 489 421 523 455
rect 597 421 631 455
rect 407 252 441 286
rect 783 309 817 343
rect 991 338 1025 372
rect 1099 342 1133 376
rect 1601 426 1635 460
rect 1226 342 1260 376
rect 1373 332 1407 366
rect 659 241 693 275
rect 1553 260 1587 294
rect 1782 306 1816 340
rect 1998 310 2032 344
rect 1890 260 1924 294
rect 2173 286 2207 320
rect 2281 286 2315 320
rect 2689 270 2723 304
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2880 683
rect 21 580 87 596
rect 21 546 37 580
rect 71 546 87 580
rect 21 510 87 546
rect 21 476 37 510
rect 71 476 87 510
rect 21 440 87 476
rect 127 580 161 649
rect 127 508 161 546
rect 127 458 161 474
rect 201 581 425 615
rect 201 580 289 581
rect 201 546 217 580
rect 251 546 289 580
rect 201 497 289 546
rect 201 463 217 497
rect 251 463 289 497
rect 21 406 37 440
rect 71 424 87 440
rect 71 406 167 424
rect 21 390 167 406
rect 25 310 99 356
rect 25 276 49 310
rect 83 276 99 310
rect 25 260 99 276
rect 133 326 167 390
rect 201 414 289 463
rect 201 380 217 414
rect 251 380 289 414
rect 201 364 289 380
rect 133 310 221 326
rect 133 276 175 310
rect 209 276 221 310
rect 133 260 221 276
rect 133 226 167 260
rect 255 226 289 364
rect 23 210 167 226
rect 23 176 39 210
rect 73 192 167 210
rect 211 210 289 226
rect 23 120 73 176
rect 245 176 289 210
rect 23 86 39 120
rect 23 70 73 86
rect 109 142 175 158
rect 109 108 125 142
rect 159 108 175 142
rect 109 17 175 108
rect 211 120 289 176
rect 245 86 289 120
rect 323 531 357 547
rect 323 202 357 497
rect 391 371 425 581
rect 459 565 493 649
rect 459 505 493 531
rect 527 581 921 615
rect 527 471 561 581
rect 837 580 921 581
rect 617 513 639 547
rect 673 513 714 547
rect 473 455 561 471
rect 473 421 489 455
rect 523 421 561 455
rect 473 405 561 421
rect 595 455 646 471
rect 595 421 597 455
rect 631 421 646 455
rect 595 371 646 421
rect 391 337 646 371
rect 391 286 551 302
rect 391 252 407 286
rect 441 252 551 286
rect 391 236 551 252
rect 601 291 646 337
rect 680 359 714 513
rect 748 531 798 547
rect 782 497 798 531
rect 748 427 798 497
rect 837 546 853 580
rect 887 546 921 580
rect 837 498 921 546
rect 1011 573 1077 649
rect 1011 539 1027 573
rect 1061 539 1077 573
rect 1011 532 1077 539
rect 1113 580 1179 596
rect 1113 546 1129 580
rect 1163 546 1179 580
rect 1113 498 1179 546
rect 1219 573 1285 649
rect 1602 628 1668 649
rect 1219 539 1235 573
rect 1269 539 1285 573
rect 1219 532 1285 539
rect 1393 580 1491 596
rect 1602 594 1618 628
rect 1652 594 1668 628
rect 1821 628 1887 649
rect 1393 546 1409 580
rect 1443 546 1491 580
rect 1714 578 1780 596
rect 1821 594 1837 628
rect 1871 594 1887 628
rect 1714 560 1730 578
rect 837 495 1129 498
rect 837 461 853 495
rect 887 464 1129 495
rect 1163 464 1276 498
rect 887 461 955 464
rect 748 393 887 427
rect 680 343 819 359
rect 680 325 783 343
rect 743 309 783 325
rect 817 309 819 343
rect 743 293 819 309
rect 601 276 709 291
rect 601 242 607 276
rect 641 275 709 276
rect 641 242 659 275
rect 601 241 659 242
rect 693 241 709 275
rect 601 225 709 241
rect 323 175 556 202
rect 743 191 777 293
rect 853 259 887 393
rect 357 168 556 175
rect 357 141 373 168
rect 323 115 373 141
rect 211 70 289 86
rect 409 100 431 134
rect 465 100 488 134
rect 409 17 488 100
rect 522 85 556 168
rect 596 172 777 191
rect 596 138 612 172
rect 646 157 777 172
rect 811 225 887 259
rect 921 259 955 461
rect 1083 424 1149 430
rect 1083 390 1087 424
rect 1121 390 1149 424
rect 989 372 1049 388
rect 989 338 991 372
rect 1025 338 1049 372
rect 989 322 1049 338
rect 1083 376 1149 390
rect 1083 342 1099 376
rect 1133 342 1149 376
rect 1083 326 1149 342
rect 1210 376 1276 464
rect 1393 470 1491 546
rect 1393 436 1409 470
rect 1443 436 1491 470
rect 1393 420 1491 436
rect 1210 342 1226 376
rect 1260 342 1276 376
rect 1210 326 1276 342
rect 1357 366 1423 382
rect 1357 332 1373 366
rect 1407 332 1423 366
rect 1457 378 1491 420
rect 1585 544 1730 560
rect 1764 560 1780 578
rect 2012 580 2078 596
rect 2012 560 2028 580
rect 1764 546 2028 560
rect 2062 546 2078 580
rect 1764 544 2078 546
rect 1585 526 2078 544
rect 2223 578 2289 649
rect 2223 544 2239 578
rect 2273 544 2289 578
rect 2223 526 2289 544
rect 2329 580 2363 596
rect 1585 460 1651 526
rect 2012 508 2078 526
rect 1585 426 1601 460
rect 1635 426 1651 460
rect 1585 412 1651 426
rect 1685 458 1978 492
rect 2012 474 2028 508
rect 2062 492 2078 508
rect 2329 500 2363 546
rect 2062 474 2292 492
rect 2012 458 2292 474
rect 1685 378 1719 458
rect 1457 344 1719 378
rect 1753 390 1759 424
rect 1793 390 1799 424
rect 1753 356 1799 390
rect 1944 378 1978 458
rect 2075 390 2134 424
rect 2168 390 2184 424
rect 1015 292 1049 322
rect 921 225 981 259
rect 1015 258 1283 292
rect 646 138 662 157
rect 596 119 662 138
rect 811 123 845 225
rect 947 224 981 225
rect 698 89 740 123
rect 774 89 845 123
rect 698 85 845 89
rect 522 51 845 85
rect 879 173 913 191
rect 879 87 913 139
rect 947 189 1015 224
rect 947 155 965 189
rect 999 155 1015 189
rect 947 121 1015 155
rect 1049 189 1115 205
rect 1049 155 1065 189
rect 1099 155 1115 189
rect 1049 87 1115 155
rect 879 53 1115 87
rect 1149 189 1215 205
rect 1149 155 1165 189
rect 1199 155 1215 189
rect 1149 17 1215 155
rect 1249 102 1283 258
rect 1357 282 1423 332
rect 1537 294 1587 310
rect 1537 282 1553 294
rect 1357 276 1553 282
rect 1357 242 1375 276
rect 1409 260 1553 276
rect 1409 242 1587 260
rect 1357 236 1587 242
rect 1621 202 1655 344
rect 1753 340 1832 356
rect 1944 344 2041 378
rect 1753 306 1782 340
rect 1816 306 1832 340
rect 1982 310 1998 344
rect 2032 310 2041 344
rect 1753 290 1832 306
rect 1874 294 1940 310
rect 1982 294 2041 310
rect 1874 260 1890 294
rect 1924 260 1940 294
rect 1874 236 1940 260
rect 2075 236 2109 390
rect 2143 320 2223 356
rect 2143 286 2173 320
rect 2207 286 2223 320
rect 2143 270 2223 286
rect 2258 336 2292 458
rect 2329 420 2363 466
rect 2403 580 2469 649
rect 2403 546 2419 580
rect 2453 546 2469 580
rect 2403 488 2469 546
rect 2403 454 2419 488
rect 2453 454 2469 488
rect 2403 438 2469 454
rect 2509 556 2575 572
rect 2509 522 2525 556
rect 2559 522 2575 556
rect 2509 485 2575 522
rect 2509 451 2525 485
rect 2559 451 2575 485
rect 2509 414 2575 451
rect 2363 386 2397 404
rect 2329 370 2397 386
rect 2258 320 2329 336
rect 2258 286 2281 320
rect 2315 286 2329 320
rect 2258 270 2329 286
rect 1330 186 1655 202
rect 1330 152 1346 186
rect 1380 152 1419 186
rect 1453 152 1492 186
rect 1526 152 1565 186
rect 1599 152 1655 186
rect 1330 136 1655 152
rect 1689 202 2148 236
rect 2182 202 2198 236
rect 1689 102 1723 202
rect 2258 168 2292 270
rect 2363 236 2397 370
rect 2509 380 2525 414
rect 2559 380 2575 414
rect 2509 364 2575 380
rect 2613 556 2663 649
rect 2613 522 2629 556
rect 2613 485 2663 522
rect 2613 451 2629 485
rect 2613 414 2663 451
rect 2613 380 2629 414
rect 2613 364 2663 380
rect 2703 580 2769 596
rect 2703 546 2719 580
rect 2753 546 2769 580
rect 2703 497 2769 546
rect 2703 463 2719 497
rect 2753 463 2769 497
rect 2703 414 2769 463
rect 2809 580 2859 649
rect 2843 546 2859 580
rect 2809 472 2859 546
rect 2843 438 2859 472
rect 2809 422 2859 438
rect 2703 380 2719 414
rect 2753 388 2769 414
rect 2753 380 2807 388
rect 2527 320 2575 364
rect 2703 354 2807 380
rect 2527 304 2739 320
rect 2527 270 2689 304
rect 2723 270 2739 304
rect 2527 254 2739 270
rect 1249 68 1723 102
rect 1757 136 1791 168
rect 1757 17 1791 102
rect 1827 136 1877 168
rect 1827 102 1843 136
rect 1921 160 2292 168
rect 1921 126 1937 160
rect 1971 134 2292 160
rect 2326 220 2397 236
rect 2326 186 2342 220
rect 2376 186 2397 220
rect 2326 146 2397 186
rect 1971 126 1987 134
rect 1921 119 1987 126
rect 1827 85 1877 102
rect 2326 112 2342 146
rect 2376 112 2397 146
rect 2022 85 2038 100
rect 1827 66 2038 85
rect 2072 66 2088 100
rect 1827 51 2088 66
rect 2133 84 2290 100
rect 2326 88 2397 112
rect 2431 236 2481 252
rect 2465 202 2481 236
rect 2431 146 2481 202
rect 2465 112 2481 146
rect 2133 50 2149 84
rect 2183 50 2240 84
rect 2274 50 2290 84
rect 2133 17 2290 50
rect 2431 17 2481 112
rect 2527 194 2577 254
rect 2773 220 2807 354
rect 2527 160 2543 194
rect 2527 120 2577 160
rect 2527 86 2543 120
rect 2527 70 2577 86
rect 2619 194 2674 210
rect 2619 160 2635 194
rect 2669 160 2674 194
rect 2619 116 2674 160
rect 2619 82 2635 116
rect 2669 82 2674 116
rect 2619 17 2674 82
rect 2708 204 2807 220
rect 2708 170 2724 204
rect 2758 170 2807 204
rect 2708 120 2760 170
rect 2708 86 2724 120
rect 2758 86 2760 120
rect 2708 70 2760 86
rect 2794 120 2860 136
rect 2794 86 2810 120
rect 2844 86 2860 120
rect 2794 17 2860 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2880 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 607 242 641 276
rect 1087 390 1121 424
rect 1759 390 1793 424
rect 1375 242 1409 276
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
<< metal1 >>
rect 0 683 2880 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2880 683
rect 0 617 2880 649
rect 1075 424 1133 430
rect 1075 390 1087 424
rect 1121 421 1133 424
rect 1747 424 1805 430
rect 1747 421 1759 424
rect 1121 393 1759 421
rect 1121 390 1133 393
rect 1075 384 1133 390
rect 1747 390 1759 393
rect 1793 390 1805 424
rect 1747 384 1805 390
rect 595 276 653 282
rect 595 242 607 276
rect 641 273 653 276
rect 1363 276 1421 282
rect 1363 273 1375 276
rect 641 245 1375 273
rect 641 242 653 245
rect 595 236 653 242
rect 1363 242 1375 245
rect 1409 242 1421 276
rect 1363 236 1421 242
rect 0 17 2880 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2880 17
rect 0 -49 2880 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dfbbn_2
flabel pwell s 0 0 2880 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 2880 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 1759 390 1793 424 0 FreeSans 340 0 0 0 SET_B
port 4 nsew
flabel metal1 s 0 617 2880 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 2880 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 2143 316 2177 350 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew
flabel corelocali s 415 242 449 276 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 511 242 545 276 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 CLK_N
port 1 nsew
flabel corelocali s 2335 94 2369 128 0 FreeSans 340 0 0 0 Q_N
port 10 nsew
flabel corelocali s 2335 168 2369 202 0 FreeSans 340 0 0 0 Q_N
port 10 nsew
flabel corelocali s 2719 390 2753 424 0 FreeSans 340 0 0 0 Q
port 9 nsew
flabel corelocali s 2719 464 2753 498 0 FreeSans 340 0 0 0 Q
port 9 nsew
flabel corelocali s 2719 538 2753 572 0 FreeSans 340 0 0 0 Q
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 2880 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2510456
string GDS_START 2489068
<< end >>
