magic
tech sky130A
magscale 1 2
timestamp 1599588238
<< locali >>
rect 181 458 237 596
rect 181 378 215 458
rect 106 344 215 378
rect 106 70 172 344
rect 317 270 381 356
rect 415 270 499 356
rect 541 270 647 356
rect 681 270 747 356
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 97 412 147 649
rect 277 458 343 649
rect 385 581 645 615
rect 385 458 451 581
rect 491 424 541 547
rect 249 390 541 424
rect 575 390 645 581
rect 679 390 745 649
rect 20 17 70 226
rect 249 310 283 390
rect 217 236 283 310
rect 217 202 466 236
rect 208 17 258 168
rect 300 85 366 168
rect 400 119 466 202
rect 500 202 740 236
rect 500 85 534 202
rect 300 51 534 85
rect 574 17 640 168
rect 674 70 740 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel locali s 317 270 381 356 6 A1
port 1 nsew signal input
rlabel locali s 681 270 747 356 6 A2
port 2 nsew signal input
rlabel locali s 415 270 499 356 6 B1
port 3 nsew signal input
rlabel locali s 541 270 647 356 6 B2
port 4 nsew signal input
rlabel locali s 181 458 237 596 6 X
port 5 nsew signal output
rlabel locali s 181 378 215 458 6 X
port 5 nsew signal output
rlabel locali s 106 344 215 378 6 X
port 5 nsew signal output
rlabel locali s 106 70 172 344 6 X
port 5 nsew signal output
rlabel metal1 s 0 -49 768 49 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 617 768 715 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3456310
string GDS_START 3449082
<< end >>
