magic
tech sky130A
magscale 1 2
timestamp 1601050056
<< nwell >>
rect -38 332 998 704
<< pwell >>
rect 0 0 960 49
<< scpmos >>
rect 83 368 119 592
rect 167 368 203 592
rect 281 368 317 592
rect 395 368 431 592
rect 509 368 545 568
rect 751 368 787 592
rect 841 368 877 592
<< nmoslvt >>
rect 84 74 114 222
rect 198 74 228 222
rect 284 74 314 222
rect 431 74 461 222
rect 520 74 550 222
rect 746 74 776 222
rect 832 74 862 222
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 136 198 222
rect 114 102 139 136
rect 173 102 198 136
rect 114 74 198 102
rect 228 210 284 222
rect 228 176 239 210
rect 273 176 284 210
rect 228 120 284 176
rect 228 86 239 120
rect 273 86 284 120
rect 228 74 284 86
rect 314 140 431 222
rect 314 106 357 140
rect 391 106 431 140
rect 314 74 431 106
rect 461 210 520 222
rect 461 176 475 210
rect 509 176 520 210
rect 461 120 520 176
rect 461 86 475 120
rect 509 86 520 120
rect 461 74 520 86
rect 550 210 621 222
rect 550 176 561 210
rect 595 176 621 210
rect 550 120 621 176
rect 550 86 561 120
rect 595 86 621 120
rect 550 74 621 86
rect 675 148 746 222
rect 675 114 701 148
rect 735 114 746 148
rect 675 74 746 114
rect 776 210 832 222
rect 776 176 787 210
rect 821 176 832 210
rect 776 120 832 176
rect 776 86 787 120
rect 821 86 832 120
rect 776 74 832 86
rect 862 186 933 222
rect 862 152 873 186
rect 907 152 933 186
rect 862 116 933 152
rect 862 82 873 116
rect 907 82 933 116
rect 862 74 933 82
<< pdiff >>
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 510 83 546
rect 27 476 39 510
rect 73 476 83 510
rect 27 440 83 476
rect 27 406 39 440
rect 73 406 83 440
rect 27 368 83 406
rect 119 368 167 592
rect 203 368 281 592
rect 317 368 395 592
rect 431 580 487 592
rect 431 546 441 580
rect 475 568 487 580
rect 701 568 751 592
rect 475 546 509 568
rect 431 510 509 546
rect 431 476 441 510
rect 475 476 509 510
rect 431 440 509 476
rect 431 406 441 440
rect 475 406 509 440
rect 431 368 509 406
rect 545 560 751 568
rect 545 526 555 560
rect 589 526 626 560
rect 660 526 706 560
rect 740 526 751 560
rect 545 492 751 526
rect 545 458 555 492
rect 589 458 626 492
rect 660 458 706 492
rect 740 458 751 492
rect 545 368 751 458
rect 787 580 841 592
rect 787 546 797 580
rect 831 546 841 580
rect 787 497 841 546
rect 787 463 797 497
rect 831 463 841 497
rect 787 414 841 463
rect 787 380 797 414
rect 831 380 841 414
rect 787 368 841 380
rect 877 580 933 592
rect 877 546 887 580
rect 921 546 933 580
rect 877 497 933 546
rect 877 463 887 497
rect 921 463 933 497
rect 877 414 933 463
rect 877 380 887 414
rect 921 380 933 414
rect 877 368 933 380
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 139 102 173 136
rect 239 176 273 210
rect 239 86 273 120
rect 357 106 391 140
rect 475 176 509 210
rect 475 86 509 120
rect 561 176 595 210
rect 561 86 595 120
rect 701 114 735 148
rect 787 176 821 210
rect 787 86 821 120
rect 873 152 907 186
rect 873 82 907 116
<< pdiffc >>
rect 39 546 73 580
rect 39 476 73 510
rect 39 406 73 440
rect 441 546 475 580
rect 441 476 475 510
rect 441 406 475 440
rect 555 526 589 560
rect 626 526 660 560
rect 706 526 740 560
rect 555 458 589 492
rect 626 458 660 492
rect 706 458 740 492
rect 797 546 831 580
rect 797 463 831 497
rect 797 380 831 414
rect 887 546 921 580
rect 887 463 921 497
rect 887 380 921 414
<< poly >>
rect 83 592 119 618
rect 167 592 203 618
rect 281 592 317 618
rect 395 592 431 618
rect 509 568 545 594
rect 751 592 787 618
rect 841 592 877 618
rect 83 336 119 368
rect 53 320 119 336
rect 53 286 69 320
rect 103 286 119 320
rect 53 270 119 286
rect 167 336 203 368
rect 281 336 317 368
rect 395 336 431 368
rect 509 336 545 368
rect 167 320 233 336
rect 167 286 183 320
rect 217 286 233 320
rect 167 270 233 286
rect 281 320 347 336
rect 281 286 297 320
rect 331 286 347 320
rect 281 270 347 286
rect 395 320 461 336
rect 395 286 411 320
rect 445 286 461 320
rect 395 270 461 286
rect 509 320 575 336
rect 751 326 787 368
rect 841 326 877 368
rect 509 286 525 320
rect 559 286 575 320
rect 509 270 575 286
rect 681 310 877 326
rect 681 276 697 310
rect 731 296 877 310
rect 731 276 862 296
rect 84 222 114 270
rect 198 222 228 270
rect 284 222 314 270
rect 431 222 461 270
rect 520 222 550 270
rect 681 260 862 276
rect 746 222 776 260
rect 832 222 862 260
rect 84 48 114 74
rect 198 48 228 74
rect 284 48 314 74
rect 431 48 461 74
rect 520 48 550 74
rect 746 48 776 74
rect 832 48 862 74
<< polycont >>
rect 69 286 103 320
rect 183 286 217 320
rect 297 286 331 320
rect 411 286 445 320
rect 525 286 559 320
rect 697 276 731 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 23 580 89 649
rect 23 546 39 580
rect 73 546 89 580
rect 425 580 491 596
rect 23 510 89 546
rect 23 476 39 510
rect 73 476 89 510
rect 23 440 89 476
rect 23 406 39 440
rect 73 406 89 440
rect 23 390 89 406
rect 167 384 263 578
rect 25 320 119 356
rect 25 286 69 320
rect 103 286 119 320
rect 25 270 119 286
rect 167 320 233 384
rect 313 336 359 578
rect 425 546 441 580
rect 475 546 491 580
rect 425 510 491 546
rect 425 476 441 510
rect 475 476 491 510
rect 425 440 491 476
rect 539 560 756 649
rect 539 526 555 560
rect 589 526 626 560
rect 660 526 706 560
rect 740 526 756 560
rect 539 492 756 526
rect 539 458 555 492
rect 589 458 626 492
rect 660 458 706 492
rect 740 458 756 492
rect 790 580 831 596
rect 790 546 797 580
rect 790 497 831 546
rect 790 463 797 497
rect 425 406 441 440
rect 475 424 491 440
rect 475 406 747 424
rect 425 390 747 406
rect 167 286 183 320
rect 217 286 233 320
rect 167 270 233 286
rect 281 320 359 336
rect 281 286 297 320
rect 331 286 359 320
rect 281 270 359 286
rect 395 320 461 356
rect 395 286 411 320
rect 445 286 461 320
rect 395 270 461 286
rect 505 320 647 356
rect 505 286 525 320
rect 559 286 647 320
rect 505 270 647 286
rect 681 310 747 390
rect 681 276 697 310
rect 731 276 747 310
rect 681 260 747 276
rect 790 414 831 463
rect 790 380 797 414
rect 790 282 831 380
rect 871 580 937 649
rect 871 546 887 580
rect 921 546 937 580
rect 871 497 937 546
rect 871 463 887 497
rect 921 463 937 497
rect 871 414 937 463
rect 871 380 887 414
rect 921 380 937 414
rect 871 364 937 380
rect 681 236 715 260
rect 23 210 525 236
rect 23 176 39 210
rect 73 202 239 210
rect 73 176 89 202
rect 23 120 89 176
rect 223 176 239 202
rect 273 202 475 210
rect 273 176 289 202
rect 23 86 39 120
rect 73 86 89 120
rect 23 70 89 86
rect 123 136 189 168
rect 123 102 139 136
rect 173 102 189 136
rect 123 17 189 102
rect 223 120 289 176
rect 459 176 475 202
rect 509 176 525 210
rect 223 86 239 120
rect 273 86 289 120
rect 223 70 289 86
rect 323 140 425 163
rect 323 106 357 140
rect 391 106 425 140
rect 323 17 425 106
rect 459 120 525 176
rect 459 86 475 120
rect 509 86 525 120
rect 459 70 525 86
rect 559 210 715 236
rect 790 236 839 282
rect 790 226 837 236
rect 559 176 561 210
rect 595 202 715 210
rect 771 210 837 226
rect 595 176 625 202
rect 559 120 625 176
rect 771 176 787 210
rect 821 176 837 210
rect 559 86 561 120
rect 595 86 625 120
rect 559 70 625 86
rect 671 148 737 164
rect 671 114 701 148
rect 735 114 737 148
rect 671 17 737 114
rect 771 120 837 176
rect 771 86 787 120
rect 821 86 837 120
rect 771 70 837 86
rect 871 186 923 202
rect 871 152 873 186
rect 907 152 923 186
rect 871 116 923 152
rect 871 82 873 116
rect 907 82 923 116
rect 871 17 923 82
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
rlabel comment s 0 0 0 0 4 o41a_2
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 223 390 257 424 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 223 464 257 498 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 223 538 257 572 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 319 390 353 424 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 319 464 353 498 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 319 538 353 572 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A4
port 4 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 B1
port 5 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 5 nsew
flabel corelocali s 799 242 833 276 0 FreeSans 340 0 0 0 X
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 960 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 709074
string GDS_START 700574
<< end >>
