magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 335 2246 704
rect -38 332 278 335
rect 1064 332 2246 335
rect 1064 311 1280 332
<< pwell >>
rect 0 0 2208 49
<< scnmos >>
rect 87 78 117 162
rect 165 78 195 162
rect 375 119 405 267
rect 485 119 515 267
rect 686 138 716 222
rect 786 138 816 222
rect 864 138 894 222
rect 942 138 972 222
rect 1073 74 1103 222
rect 1236 74 1266 222
rect 1446 81 1476 165
rect 1524 81 1554 165
rect 1626 81 1656 165
rect 1698 81 1728 165
rect 1896 74 1926 184
rect 2094 74 2124 222
<< pmoshvt >>
rect 84 508 114 592
rect 171 508 201 592
rect 370 390 400 590
rect 460 390 490 590
rect 665 457 695 541
rect 755 457 785 541
rect 833 457 863 541
rect 957 457 987 541
rect 1161 347 1191 547
rect 1262 377 1292 577
rect 1438 493 1468 577
rect 1522 493 1552 577
rect 1637 493 1667 577
rect 1727 493 1757 577
rect 1834 409 1864 577
rect 2091 368 2121 592
<< ndiff >>
rect 316 210 375 267
rect 316 180 330 210
rect 306 176 330 180
rect 364 176 375 210
rect 30 137 87 162
rect 30 103 42 137
rect 76 103 87 137
rect 30 78 87 103
rect 117 78 165 162
rect 195 137 252 162
rect 195 103 206 137
rect 240 103 252 137
rect 195 78 252 103
rect 306 142 375 176
rect 306 108 318 142
rect 352 119 375 142
rect 405 160 485 267
rect 405 126 428 160
rect 462 126 485 160
rect 405 119 485 126
rect 515 161 574 267
rect 515 127 528 161
rect 562 127 574 161
rect 629 193 686 222
rect 629 159 641 193
rect 675 159 686 193
rect 629 138 686 159
rect 716 189 786 222
rect 716 155 741 189
rect 775 155 786 189
rect 716 138 786 155
rect 816 138 864 222
rect 894 138 942 222
rect 972 138 1073 222
rect 515 119 574 127
rect 352 108 360 119
rect 306 96 360 108
rect 420 96 470 119
rect 987 79 1073 138
rect 987 45 1005 79
rect 1039 74 1073 79
rect 1103 188 1236 222
rect 1103 154 1180 188
rect 1214 154 1236 188
rect 1103 74 1236 154
rect 1266 165 1316 222
rect 2037 210 2094 222
rect 1266 153 1446 165
rect 1266 119 1280 153
rect 1314 119 1366 153
rect 1400 119 1446 153
rect 1266 81 1446 119
rect 1476 81 1524 165
rect 1554 140 1626 165
rect 1554 106 1565 140
rect 1599 106 1626 140
rect 1554 81 1626 106
rect 1656 81 1698 165
rect 1728 140 1785 165
rect 1728 106 1739 140
rect 1773 106 1785 140
rect 1728 81 1785 106
rect 1839 136 1896 184
rect 1839 102 1851 136
rect 1885 102 1896 136
rect 1266 74 1316 81
rect 1039 45 1058 74
rect 1839 74 1896 102
rect 1926 146 1983 184
rect 1926 112 1937 146
rect 1971 112 1983 146
rect 1926 74 1983 112
rect 2037 176 2049 210
rect 2083 176 2094 210
rect 2037 120 2094 176
rect 2037 86 2049 120
rect 2083 86 2094 120
rect 2037 74 2094 86
rect 2124 210 2181 222
rect 2124 176 2135 210
rect 2169 176 2181 210
rect 2124 120 2181 176
rect 2124 86 2135 120
rect 2169 86 2181 120
rect 2124 74 2181 86
rect 987 33 1058 45
<< pdiff >>
rect 27 567 84 592
rect 27 533 37 567
rect 71 533 84 567
rect 27 508 84 533
rect 114 567 171 592
rect 114 533 126 567
rect 160 533 171 567
rect 114 508 171 533
rect 201 580 254 592
rect 201 546 212 580
rect 246 546 254 580
rect 201 508 254 546
rect 308 432 370 590
rect 308 398 323 432
rect 357 398 370 432
rect 308 390 370 398
rect 400 582 460 590
rect 400 548 413 582
rect 447 548 460 582
rect 400 390 460 548
rect 490 441 547 590
rect 490 407 505 441
rect 539 407 547 441
rect 490 390 547 407
rect 881 582 939 594
rect 881 548 893 582
rect 927 548 939 582
rect 2023 580 2091 592
rect 881 541 939 548
rect 1209 547 1262 577
rect 607 516 665 541
rect 607 482 618 516
rect 652 482 665 516
rect 607 457 665 482
rect 695 533 755 541
rect 695 499 708 533
rect 742 499 755 533
rect 695 457 755 499
rect 785 457 833 541
rect 863 457 957 541
rect 987 514 1046 541
rect 987 480 1000 514
rect 1034 480 1046 514
rect 987 457 1046 480
rect 1100 535 1161 547
rect 1100 501 1112 535
rect 1146 501 1161 535
rect 1100 467 1161 501
rect 1100 433 1112 467
rect 1146 433 1161 467
rect 1100 399 1161 433
rect 1100 365 1112 399
rect 1146 365 1161 399
rect 1100 347 1161 365
rect 1191 535 1262 547
rect 1191 501 1212 535
rect 1246 501 1262 535
rect 1191 423 1262 501
rect 1191 389 1212 423
rect 1246 389 1262 423
rect 1191 377 1262 389
rect 1292 545 1438 577
rect 1292 511 1312 545
rect 1346 511 1391 545
rect 1425 511 1438 545
rect 1292 493 1438 511
rect 1468 493 1522 577
rect 1552 552 1637 577
rect 1552 518 1577 552
rect 1611 518 1637 552
rect 1552 493 1637 518
rect 1667 552 1727 577
rect 1667 518 1680 552
rect 1714 518 1727 552
rect 1667 493 1727 518
rect 1757 565 1834 577
rect 1757 531 1787 565
rect 1821 531 1834 565
rect 1757 493 1834 531
rect 1292 377 1345 493
rect 1775 489 1834 493
rect 1191 347 1244 377
rect 1775 455 1787 489
rect 1821 455 1834 489
rect 1775 409 1834 455
rect 1864 565 1923 577
rect 1864 531 1877 565
rect 1911 531 1923 565
rect 1864 455 1923 531
rect 1864 421 1877 455
rect 1911 421 1923 455
rect 1864 409 1923 421
rect 2023 546 2035 580
rect 2069 546 2091 580
rect 2023 503 2091 546
rect 2023 469 2035 503
rect 2069 469 2091 503
rect 2023 427 2091 469
rect 2023 393 2035 427
rect 2069 393 2091 427
rect 2023 368 2091 393
rect 2121 580 2181 592
rect 2121 546 2135 580
rect 2169 546 2181 580
rect 2121 497 2181 546
rect 2121 463 2135 497
rect 2169 463 2181 497
rect 2121 414 2181 463
rect 2121 380 2135 414
rect 2169 380 2181 414
rect 2121 368 2181 380
<< ndiffc >>
rect 330 176 364 210
rect 42 103 76 137
rect 206 103 240 137
rect 318 108 352 142
rect 428 126 462 160
rect 528 127 562 161
rect 641 159 675 193
rect 741 155 775 189
rect 1005 45 1039 79
rect 1180 154 1214 188
rect 1280 119 1314 153
rect 1366 119 1400 153
rect 1565 106 1599 140
rect 1739 106 1773 140
rect 1851 102 1885 136
rect 1937 112 1971 146
rect 2049 176 2083 210
rect 2049 86 2083 120
rect 2135 176 2169 210
rect 2135 86 2169 120
<< pdiffc >>
rect 37 533 71 567
rect 126 533 160 567
rect 212 546 246 580
rect 323 398 357 432
rect 413 548 447 582
rect 505 407 539 441
rect 893 548 927 582
rect 618 482 652 516
rect 708 499 742 533
rect 1000 480 1034 514
rect 1112 501 1146 535
rect 1112 433 1146 467
rect 1112 365 1146 399
rect 1212 501 1246 535
rect 1212 389 1246 423
rect 1312 511 1346 545
rect 1391 511 1425 545
rect 1577 518 1611 552
rect 1680 518 1714 552
rect 1787 531 1821 565
rect 1787 455 1821 489
rect 1877 531 1911 565
rect 1877 421 1911 455
rect 2035 546 2069 580
rect 2035 469 2069 503
rect 2035 393 2069 427
rect 2135 546 2169 580
rect 2135 463 2169 497
rect 2135 380 2169 414
<< poly >>
rect 84 592 114 618
rect 171 592 201 618
rect 370 590 400 616
rect 460 590 490 616
rect 562 615 1295 645
rect 84 493 114 508
rect 171 493 201 508
rect 81 402 117 493
rect 171 428 207 493
rect 44 386 117 402
rect 44 352 60 386
rect 94 352 117 386
rect 44 318 117 352
rect 44 284 60 318
rect 94 284 117 318
rect 44 250 117 284
rect 44 216 60 250
rect 94 216 117 250
rect 44 200 117 216
rect 87 162 117 200
rect 165 412 264 428
rect 165 378 214 412
rect 248 378 264 412
rect 165 344 264 378
rect 370 355 400 390
rect 460 355 490 390
rect 562 355 592 615
rect 665 541 695 567
rect 755 541 785 615
rect 1259 592 1295 615
rect 833 541 863 567
rect 1262 577 1292 592
rect 1438 577 1468 603
rect 1522 577 1552 603
rect 1637 577 1667 603
rect 1727 577 1757 603
rect 1834 577 1864 603
rect 2091 592 2121 618
rect 957 541 987 567
rect 1161 547 1191 573
rect 665 442 695 457
rect 665 397 700 442
rect 755 431 785 457
rect 833 442 863 457
rect 957 442 987 457
rect 165 310 214 344
rect 248 310 264 344
rect 165 276 264 310
rect 349 339 415 355
rect 349 305 365 339
rect 399 305 415 339
rect 349 287 415 305
rect 460 339 592 355
rect 634 381 700 397
rect 634 347 650 381
rect 684 347 700 381
rect 830 425 866 442
rect 954 425 990 442
rect 830 409 904 425
rect 830 375 854 409
rect 888 375 904 409
rect 830 359 904 375
rect 954 409 1057 425
rect 954 375 1007 409
rect 1041 375 1057 409
rect 954 359 1057 375
rect 634 342 700 347
rect 634 339 788 342
rect 460 305 505 339
rect 539 314 592 339
rect 636 335 788 339
rect 638 333 788 335
rect 642 331 788 333
rect 649 324 788 331
rect 539 310 596 314
rect 657 312 788 324
rect 758 311 788 312
rect 539 306 601 310
rect 539 305 603 306
rect 460 304 603 305
rect 460 302 607 304
rect 460 300 609 302
rect 460 297 611 300
rect 460 294 614 297
rect 165 242 214 276
rect 248 242 264 276
rect 375 267 405 287
rect 460 282 619 294
rect 485 267 515 282
rect 582 280 619 282
rect 758 281 816 311
rect 585 278 619 280
rect 587 276 619 278
rect 589 270 619 276
rect 165 226 264 242
rect 165 162 195 226
rect 589 240 716 270
rect 686 222 716 240
rect 786 222 816 281
rect 864 222 894 359
rect 960 267 990 359
rect 1438 478 1468 493
rect 1522 478 1552 493
rect 1637 478 1667 493
rect 1727 478 1757 493
rect 1435 461 1471 478
rect 1393 445 1471 461
rect 1393 411 1409 445
rect 1443 411 1471 445
rect 1393 395 1471 411
rect 1262 362 1292 377
rect 1259 347 1295 362
rect 1519 349 1555 478
rect 1634 451 1670 478
rect 1603 435 1670 451
rect 1603 401 1619 435
rect 1653 401 1670 435
rect 1603 385 1670 401
rect 1161 332 1191 347
rect 1158 315 1194 332
rect 1259 317 1476 347
rect 942 237 990 267
rect 1064 299 1194 315
rect 1064 265 1080 299
rect 1114 285 1194 299
rect 1114 265 1130 285
rect 1064 249 1130 265
rect 1236 253 1404 269
rect 942 222 972 237
rect 1073 222 1103 249
rect 1236 239 1354 253
rect 1236 222 1266 239
rect 375 93 405 119
rect 485 93 515 119
rect 686 112 716 138
rect 786 112 816 138
rect 864 112 894 138
rect 87 52 117 78
rect 165 51 195 78
rect 942 51 972 138
rect 165 21 972 51
rect 1338 219 1354 239
rect 1388 219 1404 253
rect 1338 203 1404 219
rect 1446 165 1476 317
rect 1519 269 1549 349
rect 1518 253 1584 269
rect 1518 219 1534 253
rect 1568 219 1584 253
rect 1518 203 1584 219
rect 1524 165 1554 203
rect 1626 165 1656 385
rect 1724 337 1760 478
rect 1834 394 1864 409
rect 1831 337 1867 394
rect 2091 353 2121 368
rect 2088 343 2124 353
rect 1704 321 1867 337
rect 1704 301 1720 321
rect 1698 287 1720 301
rect 1754 287 1867 321
rect 1698 271 1867 287
rect 1921 327 2124 343
rect 1921 293 1937 327
rect 1971 293 2124 327
rect 1921 277 2124 293
rect 1698 165 1728 271
rect 1831 229 1861 271
rect 1831 199 1926 229
rect 2094 222 2124 277
rect 1896 184 1926 199
rect 1073 48 1103 74
rect 1236 48 1266 74
rect 1446 55 1476 81
rect 1524 55 1554 81
rect 1626 55 1656 81
rect 1698 55 1728 81
rect 1896 48 1926 74
rect 2094 48 2124 74
<< polycont >>
rect 60 352 94 386
rect 60 284 94 318
rect 60 216 94 250
rect 214 378 248 412
rect 214 310 248 344
rect 365 305 399 339
rect 650 347 684 381
rect 854 375 888 409
rect 1007 375 1041 409
rect 505 305 539 339
rect 214 242 248 276
rect 1409 411 1443 445
rect 1619 401 1653 435
rect 1080 265 1114 299
rect 1354 219 1388 253
rect 1534 219 1568 253
rect 1720 287 1754 321
rect 1937 293 1971 327
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 21 567 71 649
rect 21 533 37 567
rect 21 504 71 533
rect 111 567 162 596
rect 111 533 126 567
rect 160 533 162 567
rect 196 580 262 649
rect 196 546 212 580
rect 246 546 262 580
rect 397 582 463 649
rect 397 548 413 582
rect 447 548 463 582
rect 877 582 943 649
rect 877 548 893 582
rect 927 548 943 582
rect 111 528 162 533
rect 111 521 167 528
rect 111 512 172 521
rect 287 518 372 522
rect 287 517 378 518
rect 281 516 378 517
rect 602 516 658 545
rect 281 515 382 516
rect 281 514 385 515
rect 602 514 618 516
rect 281 512 618 514
rect 111 504 618 512
rect 137 482 618 504
rect 652 482 658 516
rect 692 533 843 545
rect 692 499 708 533
rect 742 514 843 533
rect 1096 535 1162 649
rect 742 499 1000 514
rect 137 478 306 482
rect 367 481 658 482
rect 370 480 658 481
rect 374 478 658 480
rect 137 475 302 478
rect 379 475 658 478
rect 137 472 298 475
rect 602 474 658 475
rect 786 480 1000 499
rect 1034 480 1050 514
rect 137 467 293 472
rect 137 462 287 467
rect 602 465 667 474
rect 25 386 103 434
rect 25 352 60 386
rect 94 352 103 386
rect 25 318 103 352
rect 25 284 60 318
rect 94 284 103 318
rect 25 250 103 284
rect 25 216 60 250
rect 94 216 103 250
rect 25 200 103 216
rect 137 166 171 462
rect 323 441 357 448
rect 602 441 752 465
rect 323 432 373 441
rect 205 424 257 428
rect 205 412 223 424
rect 205 378 214 412
rect 248 378 257 390
rect 205 344 257 378
rect 205 310 214 344
rect 248 310 257 344
rect 205 276 257 310
rect 205 242 214 276
rect 248 242 257 276
rect 205 226 257 242
rect 291 398 323 428
rect 357 398 373 432
rect 291 389 373 398
rect 489 407 505 441
rect 539 407 555 441
rect 637 431 752 441
rect 489 397 612 407
rect 291 228 325 389
rect 489 381 684 397
rect 489 373 650 381
rect 580 364 650 373
rect 409 355 455 356
rect 359 339 455 355
rect 589 347 650 364
rect 359 305 365 339
rect 399 305 455 339
rect 359 262 455 305
rect 489 305 505 339
rect 539 305 555 339
rect 489 298 555 305
rect 589 312 684 347
rect 489 228 539 298
rect 589 269 623 312
rect 718 278 752 431
rect 291 210 539 228
rect 291 176 330 210
rect 364 195 539 210
rect 573 239 623 269
rect 657 244 752 278
rect 364 194 501 195
rect 364 176 368 194
rect 26 137 171 166
rect 26 103 42 137
rect 76 132 171 137
rect 206 137 256 166
rect 76 103 92 132
rect 26 74 92 103
rect 240 103 256 137
rect 206 17 256 103
rect 291 142 368 176
rect 573 161 607 239
rect 657 209 691 244
rect 786 210 820 480
rect 923 464 1050 480
rect 1096 501 1112 535
rect 1146 501 1162 535
rect 1096 467 1162 501
rect 291 108 318 142
rect 352 108 368 142
rect 291 70 368 108
rect 412 126 428 160
rect 462 126 478 160
rect 412 17 478 126
rect 512 127 528 161
rect 562 127 607 161
rect 641 193 691 209
rect 675 159 691 193
rect 641 134 691 159
rect 725 189 820 210
rect 725 155 741 189
rect 775 155 820 189
rect 854 409 889 425
rect 888 375 889 409
rect 854 215 889 375
rect 923 315 957 464
rect 1096 433 1112 467
rect 1146 433 1162 467
rect 991 424 1057 430
rect 1025 409 1057 424
rect 991 375 1007 390
rect 1041 375 1057 409
rect 991 359 1057 375
rect 1096 399 1162 433
rect 1096 365 1112 399
rect 1146 365 1162 399
rect 1096 349 1162 365
rect 1196 535 1262 551
rect 1196 501 1212 535
rect 1246 501 1262 535
rect 1196 423 1262 501
rect 1196 389 1212 423
rect 1246 389 1262 423
rect 1196 373 1262 389
rect 1296 545 1527 561
rect 1296 511 1312 545
rect 1346 511 1391 545
rect 1425 511 1527 545
rect 1296 495 1527 511
rect 923 299 1130 315
rect 923 265 1080 299
rect 1114 265 1130 299
rect 923 249 1130 265
rect 1196 226 1230 373
rect 1296 337 1330 495
rect 1164 215 1230 226
rect 854 188 1230 215
rect 854 181 1180 188
rect 725 134 820 155
rect 1164 154 1180 181
rect 1214 154 1230 188
rect 512 100 607 127
rect 854 113 1130 147
rect 1164 133 1230 154
rect 1264 303 1330 337
rect 1393 445 1459 461
rect 1393 411 1409 445
rect 1443 411 1459 445
rect 1264 169 1298 303
rect 1393 269 1459 411
rect 1493 337 1527 495
rect 1561 552 1627 649
rect 1561 518 1577 552
rect 1611 518 1627 552
rect 1561 489 1627 518
rect 1664 552 1737 581
rect 1664 518 1680 552
rect 1714 518 1737 552
rect 1664 489 1737 518
rect 1561 435 1669 451
rect 1561 424 1619 435
rect 1561 390 1567 424
rect 1601 401 1619 424
rect 1653 401 1669 435
rect 1601 390 1669 401
rect 1561 384 1669 390
rect 1703 405 1737 489
rect 1771 565 1837 649
rect 1771 531 1787 565
rect 1821 531 1837 565
rect 1771 489 1837 531
rect 1771 455 1787 489
rect 1821 455 1837 489
rect 1771 439 1837 455
rect 1877 565 1911 581
rect 1877 455 1911 531
rect 1703 371 1838 405
rect 1493 321 1770 337
rect 1493 303 1720 321
rect 1704 287 1720 303
rect 1754 287 1770 321
rect 1704 271 1770 287
rect 1338 253 1484 269
rect 1338 219 1354 253
rect 1388 219 1484 253
rect 1338 203 1484 219
rect 1518 253 1584 269
rect 1518 219 1534 253
rect 1568 237 1584 253
rect 1804 237 1838 371
rect 1877 343 1911 421
rect 1945 580 2085 596
rect 1945 546 2035 580
rect 2069 546 2085 580
rect 1945 503 2085 546
rect 1945 469 2035 503
rect 2069 469 2085 503
rect 1945 427 2085 469
rect 1945 393 2035 427
rect 2069 393 2085 427
rect 1945 377 2085 393
rect 1877 327 1987 343
rect 1877 293 1937 327
rect 1971 293 1987 327
rect 1877 277 1987 293
rect 1568 219 1838 237
rect 1518 203 1838 219
rect 1264 153 1416 169
rect 1264 119 1280 153
rect 1314 119 1366 153
rect 1400 119 1416 153
rect 854 100 888 113
rect 512 66 888 100
rect 1096 85 1130 113
rect 1450 85 1484 203
rect 983 45 1005 79
rect 1039 45 1062 79
rect 1096 51 1484 85
rect 1549 140 1615 169
rect 1549 106 1565 140
rect 1599 106 1615 140
rect 983 17 1062 45
rect 1549 17 1615 106
rect 1723 140 1789 203
rect 1723 106 1739 140
rect 1773 106 1789 140
rect 1723 77 1789 106
rect 1835 136 1885 169
rect 1835 102 1851 136
rect 1835 17 1885 102
rect 1921 146 1987 277
rect 1921 112 1937 146
rect 1971 112 1987 146
rect 1921 70 1987 112
rect 2033 226 2085 377
rect 2119 580 2185 649
rect 2119 546 2135 580
rect 2169 546 2185 580
rect 2119 497 2185 546
rect 2119 463 2135 497
rect 2169 463 2185 497
rect 2119 414 2185 463
rect 2119 380 2135 414
rect 2169 380 2185 414
rect 2119 364 2185 380
rect 2033 210 2099 226
rect 2033 176 2049 210
rect 2083 176 2099 210
rect 2033 120 2099 176
rect 2033 86 2049 120
rect 2083 86 2099 120
rect 2033 70 2099 86
rect 2135 210 2185 226
rect 2169 176 2185 210
rect 2135 120 2185 176
rect 2169 86 2185 120
rect 2135 17 2185 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 223 412 257 424
rect 223 390 248 412
rect 248 390 257 412
rect 991 409 1025 424
rect 991 390 1007 409
rect 1007 390 1025 409
rect 1567 390 1601 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
<< metal1 >>
rect 0 683 2208 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 0 617 2208 649
rect 211 424 269 430
rect 211 390 223 424
rect 257 421 269 424
rect 979 424 1037 430
rect 979 421 991 424
rect 257 393 991 421
rect 257 390 269 393
rect 211 384 269 390
rect 979 390 991 393
rect 1025 421 1037 424
rect 1555 424 1613 430
rect 1555 421 1567 424
rect 1025 393 1567 421
rect 1025 390 1037 393
rect 979 384 1037 390
rect 1555 390 1567 393
rect 1601 390 1613 424
rect 1555 384 1613 390
rect 0 17 2208 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
rect 0 -49 2208 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dfrtp_1
flabel comment s 927 630 927 630 0 FreeSans 300 0 0 0 no_jumper_check
flabel comment s 565 36 565 36 0 FreeSans 300 0 0 0 no_jumper_check
flabel pwell s 0 0 2208 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 2208 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 223 390 257 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew
flabel metal1 s 0 617 2208 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 2208 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 1951 390 1985 424 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 1951 464 1985 498 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 1951 538 1985 572 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 31 390 65 424 0 FreeSans 340 0 0 0 D
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 2208 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2604976
string GDS_START 2586002
<< end >>
