magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 89 47 119 131
rect 173 47 203 131
rect 269 47 299 131
rect 367 47 397 131
rect 487 47 517 177
<< pmoshvt >>
rect 81 413 117 497
rect 175 413 211 497
rect 271 413 307 497
rect 369 413 405 497
rect 479 297 515 497
<< ndiff >>
rect 412 131 487 177
rect 27 101 89 131
rect 27 67 35 101
rect 69 67 89 101
rect 27 47 89 67
rect 119 47 173 131
rect 203 47 269 131
rect 299 47 367 131
rect 397 93 487 131
rect 397 59 418 93
rect 452 59 487 93
rect 397 47 487 59
rect 517 161 607 177
rect 517 127 565 161
rect 599 127 607 161
rect 517 93 607 127
rect 517 59 565 93
rect 599 59 607 93
rect 517 47 607 59
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 413 81 451
rect 117 477 175 497
rect 117 443 129 477
rect 163 443 175 477
rect 117 413 175 443
rect 211 485 271 497
rect 211 451 223 485
rect 257 451 271 485
rect 211 413 271 451
rect 307 477 369 497
rect 307 443 320 477
rect 354 443 369 477
rect 307 413 369 443
rect 405 485 479 497
rect 405 451 433 485
rect 467 451 479 485
rect 405 417 479 451
rect 405 413 433 417
rect 422 383 433 413
rect 467 383 479 417
rect 422 297 479 383
rect 515 485 607 497
rect 515 451 565 485
rect 599 451 607 485
rect 515 417 607 451
rect 515 383 565 417
rect 599 383 607 417
rect 515 349 607 383
rect 515 315 565 349
rect 599 315 607 349
rect 515 297 607 315
<< ndiffc >>
rect 35 67 69 101
rect 418 59 452 93
rect 565 127 599 161
rect 565 59 599 93
<< pdiffc >>
rect 35 451 69 485
rect 129 443 163 477
rect 223 451 257 485
rect 320 443 354 477
rect 433 451 467 485
rect 433 383 467 417
rect 565 451 599 485
rect 565 383 599 417
rect 565 315 599 349
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 271 497 307 523
rect 369 497 405 523
rect 479 497 515 523
rect 81 398 117 413
rect 175 398 211 413
rect 271 398 307 413
rect 369 398 405 413
rect 79 265 119 398
rect 21 249 119 265
rect 21 215 31 249
rect 65 215 119 249
rect 21 199 119 215
rect 89 131 119 199
rect 173 265 213 398
rect 269 265 309 398
rect 367 265 407 398
rect 479 282 515 297
rect 477 265 517 282
rect 173 249 227 265
rect 173 215 183 249
rect 217 215 227 249
rect 173 199 227 215
rect 269 249 325 265
rect 269 215 281 249
rect 315 215 325 249
rect 269 199 325 215
rect 367 249 421 265
rect 367 215 377 249
rect 411 215 421 249
rect 367 199 421 215
rect 463 249 517 265
rect 463 215 473 249
rect 507 215 517 249
rect 463 199 517 215
rect 173 131 203 199
rect 269 131 299 199
rect 367 131 397 199
rect 487 177 517 199
rect 89 21 119 47
rect 173 21 203 47
rect 269 21 299 47
rect 367 21 397 47
rect 487 21 517 47
<< polycont >>
rect 31 215 65 249
rect 183 215 217 249
rect 281 215 315 249
rect 377 215 411 249
rect 473 215 507 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 18 485 85 527
rect 18 451 35 485
rect 69 451 85 485
rect 121 477 171 493
rect 121 443 129 477
rect 163 443 171 477
rect 17 249 65 415
rect 121 333 171 443
rect 207 485 273 527
rect 207 451 223 485
rect 257 451 273 485
rect 207 383 273 451
rect 312 477 362 493
rect 312 443 320 477
rect 354 443 362 477
rect 312 333 362 443
rect 401 485 475 527
rect 401 451 433 485
rect 467 451 475 485
rect 401 417 475 451
rect 539 485 617 493
rect 539 451 565 485
rect 599 451 617 485
rect 539 441 617 451
rect 401 383 433 417
rect 467 383 475 417
rect 401 367 475 383
rect 565 417 617 441
rect 599 383 617 417
rect 565 349 617 383
rect 17 215 31 249
rect 17 153 65 215
rect 99 299 507 333
rect 99 117 137 299
rect 34 101 137 117
rect 34 67 35 101
rect 69 67 137 101
rect 171 249 247 265
rect 171 215 183 249
rect 217 215 247 249
rect 171 72 247 215
rect 281 249 339 265
rect 315 215 339 249
rect 281 71 339 215
rect 377 249 433 265
rect 411 215 433 249
rect 377 143 433 215
rect 467 249 507 299
rect 467 215 473 249
rect 467 199 507 215
rect 599 315 617 349
rect 565 161 617 315
rect 539 127 565 161
rect 599 127 617 161
rect 413 93 467 109
rect 34 51 137 67
rect 413 59 418 93
rect 452 59 467 93
rect 539 93 617 127
rect 539 59 565 93
rect 599 59 617 93
rect 413 17 467 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel corelocali s 571 425 605 459 0 FreeSans 200 0 0 0 X
port 9 nsew
flabel corelocali s 288 102 288 102 0 FreeSans 200 0 0 0 C
port 3 nsew
flabel corelocali s 288 170 288 170 0 FreeSans 200 0 0 0 C
port 3 nsew
flabel corelocali s 29 221 63 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 288 238 288 238 0 FreeSans 200 0 0 0 C
port 3 nsew
flabel corelocali s 193 102 193 102 0 FreeSans 200 0 0 0 B
port 2 nsew
flabel corelocali s 193 170 193 170 0 FreeSans 200 0 0 0 B
port 2 nsew
flabel corelocali s 382 238 382 238 0 FreeSans 200 0 0 0 D
port 4 nsew
flabel corelocali s 571 85 605 119 0 FreeSans 200 0 0 0 X
port 9 nsew
flabel corelocali s 571 153 605 187 0 FreeSans 200 0 0 0 X
port 9 nsew
flabel corelocali s 571 221 605 255 0 FreeSans 200 0 0 0 X
port 9 nsew
flabel corelocali s 571 289 605 323 0 FreeSans 200 0 0 0 X
port 9 nsew
flabel corelocali s 571 357 605 391 0 FreeSans 200 0 0 0 X
port 9 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
rlabel comment s 0 0 0 0 4 and4_1
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1558150
string GDS_START 1551716
<< end >>
