magic
tech sky130A
magscale 1 2
timestamp 1601050047
<< nwell >>
rect -38 332 806 704
<< pwell >>
rect 0 0 768 49
<< scpmos >>
rect 100 368 130 592
rect 190 368 220 592
rect 332 368 362 568
rect 422 368 452 568
rect 550 368 580 568
rect 650 368 680 568
<< nmoslvt >>
rect 98 74 128 222
rect 184 74 214 222
rect 341 74 371 222
rect 419 74 449 222
rect 533 74 563 222
rect 647 74 677 222
<< ndiff >>
rect 27 210 98 222
rect 27 176 39 210
rect 73 176 98 210
rect 27 120 98 176
rect 27 86 39 120
rect 73 86 98 120
rect 27 74 98 86
rect 128 210 184 222
rect 128 176 139 210
rect 173 176 184 210
rect 128 120 184 176
rect 128 86 139 120
rect 173 86 184 120
rect 128 74 184 86
rect 214 120 341 222
rect 214 86 228 120
rect 262 86 296 120
rect 330 86 341 120
rect 214 74 341 86
rect 371 74 419 222
rect 449 74 533 222
rect 563 202 647 222
rect 563 168 586 202
rect 620 168 647 202
rect 563 116 647 168
rect 563 82 586 116
rect 620 82 647 116
rect 563 74 647 82
rect 677 188 734 222
rect 677 154 688 188
rect 722 154 734 188
rect 677 120 734 154
rect 677 86 688 120
rect 722 86 734 120
rect 677 74 734 86
<< pdiff >>
rect 41 580 100 592
rect 41 546 53 580
rect 87 546 100 580
rect 41 497 100 546
rect 41 463 53 497
rect 87 463 100 497
rect 41 414 100 463
rect 41 380 53 414
rect 87 380 100 414
rect 41 368 100 380
rect 130 580 190 592
rect 130 546 143 580
rect 177 546 190 580
rect 130 497 190 546
rect 130 463 143 497
rect 177 463 190 497
rect 130 414 190 463
rect 130 380 143 414
rect 177 380 190 414
rect 130 368 190 380
rect 220 584 308 592
rect 220 550 234 584
rect 268 568 308 584
rect 268 550 332 568
rect 220 516 332 550
rect 220 482 284 516
rect 318 482 332 516
rect 220 446 332 482
rect 220 412 234 446
rect 268 412 332 446
rect 220 368 332 412
rect 362 556 422 568
rect 362 522 375 556
rect 409 522 422 556
rect 362 449 422 522
rect 362 415 375 449
rect 409 415 422 449
rect 362 368 422 415
rect 452 530 550 568
rect 452 496 486 530
rect 520 496 550 530
rect 452 368 550 496
rect 580 556 650 568
rect 580 522 593 556
rect 627 522 650 556
rect 580 451 650 522
rect 580 417 593 451
rect 627 417 650 451
rect 580 368 650 417
rect 680 556 741 568
rect 680 522 694 556
rect 728 522 741 556
rect 680 485 741 522
rect 680 451 694 485
rect 728 451 741 485
rect 680 414 741 451
rect 680 380 694 414
rect 728 380 741 414
rect 680 368 741 380
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 139 176 173 210
rect 139 86 173 120
rect 228 86 262 120
rect 296 86 330 120
rect 586 168 620 202
rect 586 82 620 116
rect 688 154 722 188
rect 688 86 722 120
<< pdiffc >>
rect 53 546 87 580
rect 53 463 87 497
rect 53 380 87 414
rect 143 546 177 580
rect 143 463 177 497
rect 143 380 177 414
rect 234 550 268 584
rect 284 482 318 516
rect 234 412 268 446
rect 375 522 409 556
rect 375 415 409 449
rect 486 496 520 530
rect 593 522 627 556
rect 593 417 627 451
rect 694 522 728 556
rect 694 451 728 485
rect 694 380 728 414
<< poly >>
rect 100 592 130 618
rect 190 592 220 618
rect 332 568 362 594
rect 422 568 452 594
rect 550 568 580 594
rect 650 568 680 594
rect 100 353 130 368
rect 190 353 220 368
rect 332 353 362 368
rect 422 353 452 368
rect 550 353 580 368
rect 650 353 680 368
rect 97 326 133 353
rect 187 326 223 353
rect 97 310 257 326
rect 329 310 365 353
rect 419 310 455 353
rect 547 310 583 353
rect 647 310 683 353
rect 97 296 207 310
rect 98 276 207 296
rect 241 276 257 310
rect 98 260 257 276
rect 305 294 371 310
rect 305 260 321 294
rect 355 260 371 294
rect 98 222 128 260
rect 184 222 214 260
rect 305 244 371 260
rect 341 222 371 244
rect 419 294 485 310
rect 419 260 435 294
rect 469 260 485 294
rect 419 244 485 260
rect 533 294 599 310
rect 533 260 549 294
rect 583 260 599 294
rect 533 244 599 260
rect 647 294 747 310
rect 647 260 697 294
rect 731 260 747 294
rect 647 244 747 260
rect 419 222 449 244
rect 533 222 563 244
rect 647 222 677 244
rect 98 48 128 74
rect 184 48 214 74
rect 341 48 371 74
rect 419 48 449 74
rect 533 48 563 74
rect 647 48 677 74
<< polycont >>
rect 207 276 241 310
rect 321 260 355 294
rect 435 260 469 294
rect 549 260 583 294
rect 697 260 731 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 37 580 87 649
rect 37 546 53 580
rect 37 497 87 546
rect 37 463 53 497
rect 37 414 87 463
rect 37 380 53 414
rect 37 364 87 380
rect 121 580 184 596
rect 121 546 143 580
rect 177 546 184 580
rect 121 497 184 546
rect 121 463 143 497
rect 177 463 184 497
rect 121 414 184 463
rect 121 380 143 414
rect 177 380 184 414
rect 218 584 325 649
rect 218 550 234 584
rect 268 550 325 584
rect 218 516 325 550
rect 218 482 284 516
rect 318 482 325 516
rect 218 446 325 482
rect 218 412 234 446
rect 268 412 325 446
rect 359 556 425 572
rect 359 522 375 556
rect 409 522 425 556
rect 359 449 425 522
rect 470 530 536 649
rect 470 496 486 530
rect 520 496 536 530
rect 470 480 536 496
rect 577 556 643 572
rect 577 522 593 556
rect 627 522 643 556
rect 359 415 375 449
rect 409 446 425 449
rect 577 451 643 522
rect 577 446 593 451
rect 409 417 593 446
rect 627 417 643 451
rect 409 415 643 417
rect 359 412 643 415
rect 677 556 745 572
rect 677 522 694 556
rect 728 522 745 556
rect 677 485 745 522
rect 677 451 694 485
rect 728 451 745 485
rect 677 414 745 451
rect 121 364 184 380
rect 677 380 694 414
rect 728 380 745 414
rect 677 378 745 380
rect 123 226 157 364
rect 227 344 745 378
rect 227 326 261 344
rect 191 310 261 326
rect 191 276 207 310
rect 241 276 261 310
rect 191 260 261 276
rect 23 210 89 226
rect 23 176 39 210
rect 73 176 89 210
rect 23 120 89 176
rect 23 86 39 120
rect 73 86 89 120
rect 23 17 89 86
rect 123 210 178 226
rect 123 176 139 210
rect 173 176 178 210
rect 123 120 178 176
rect 227 202 261 260
rect 305 294 371 310
rect 305 260 321 294
rect 355 260 371 294
rect 305 236 371 260
rect 409 294 485 310
rect 409 260 435 294
rect 469 260 485 294
rect 409 236 485 260
rect 533 294 647 310
rect 533 260 549 294
rect 583 260 647 294
rect 533 236 647 260
rect 681 294 747 310
rect 681 260 697 294
rect 731 260 747 294
rect 681 236 747 260
rect 227 168 586 202
rect 620 168 636 202
rect 123 86 139 120
rect 173 86 178 120
rect 123 70 178 86
rect 212 86 228 120
rect 262 86 296 120
rect 330 86 346 120
rect 212 17 346 86
rect 570 116 636 168
rect 570 82 586 116
rect 620 82 636 116
rect 570 70 636 82
rect 672 188 738 202
rect 672 154 688 188
rect 722 154 738 188
rect 672 120 738 154
rect 672 86 688 120
rect 722 86 738 120
rect 672 17 738 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a31o_2
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 607 242 641 276 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 415 242 449 276 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 319 242 353 276 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 703 242 737 276 0 FreeSans 340 0 0 0 B1
port 4 nsew
flabel corelocali s 127 390 161 424 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 127 464 161 498 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 127 538 161 572 0 FreeSans 340 0 0 0 X
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 768 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3809844
string GDS_START 3802838
<< end >>
