magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 902 704
<< pwell >>
rect 0 0 864 49
<< scnmos >>
rect 84 112 114 222
rect 186 74 216 222
rect 272 74 302 222
rect 429 74 459 222
rect 507 74 537 222
rect 615 74 645 222
rect 723 74 753 222
<< pmoshvt >>
rect 86 368 116 536
rect 195 368 225 592
rect 285 368 315 592
rect 409 368 439 568
rect 504 368 534 568
rect 628 368 658 568
rect 726 368 756 568
<< ndiff >>
rect 27 184 84 222
rect 27 150 39 184
rect 73 150 84 184
rect 27 112 84 150
rect 114 142 186 222
rect 114 112 141 142
rect 129 108 141 112
rect 175 108 186 142
rect 129 74 186 108
rect 216 210 272 222
rect 216 176 227 210
rect 261 176 272 210
rect 216 120 272 176
rect 216 86 227 120
rect 261 86 272 120
rect 216 74 272 86
rect 302 142 429 222
rect 302 108 313 142
rect 347 108 384 142
rect 418 108 429 142
rect 302 74 429 108
rect 459 74 507 222
rect 537 74 615 222
rect 645 74 723 222
rect 753 210 810 222
rect 753 176 764 210
rect 798 176 810 210
rect 753 120 810 176
rect 753 86 764 120
rect 798 86 810 120
rect 753 74 810 86
<< pdiff >>
rect 134 578 195 592
rect 134 544 146 578
rect 180 544 195 578
rect 134 536 195 544
rect 27 524 86 536
rect 27 490 39 524
rect 73 490 86 524
rect 27 440 86 490
rect 27 406 39 440
rect 73 406 86 440
rect 27 368 86 406
rect 116 368 195 536
rect 225 419 285 592
rect 225 385 238 419
rect 272 385 285 419
rect 225 368 285 385
rect 315 578 391 592
rect 315 544 345 578
rect 379 568 391 578
rect 552 578 610 586
rect 552 568 564 578
rect 379 544 409 568
rect 315 368 409 544
rect 439 424 504 568
rect 439 390 454 424
rect 488 390 504 424
rect 439 368 504 390
rect 534 544 564 568
rect 598 568 610 578
rect 774 578 837 586
rect 774 568 788 578
rect 598 544 628 568
rect 534 368 628 544
rect 658 424 726 568
rect 658 390 675 424
rect 709 390 726 424
rect 658 368 726 390
rect 756 544 788 568
rect 822 544 837 578
rect 756 368 837 544
<< ndiffc >>
rect 39 150 73 184
rect 141 108 175 142
rect 227 176 261 210
rect 227 86 261 120
rect 313 108 347 142
rect 384 108 418 142
rect 764 176 798 210
rect 764 86 798 120
<< pdiffc >>
rect 146 544 180 578
rect 39 490 73 524
rect 39 406 73 440
rect 238 385 272 419
rect 345 544 379 578
rect 454 390 488 424
rect 564 544 598 578
rect 675 390 709 424
rect 788 544 822 578
<< poly >>
rect 195 592 225 618
rect 285 592 315 618
rect 86 536 116 562
rect 409 568 439 594
rect 504 568 534 594
rect 628 568 658 594
rect 726 568 756 594
rect 86 353 116 368
rect 195 353 225 368
rect 285 353 315 368
rect 409 353 439 368
rect 504 353 534 368
rect 628 353 658 368
rect 726 353 756 368
rect 83 326 119 353
rect 25 310 119 326
rect 25 276 41 310
rect 75 276 119 310
rect 192 326 228 353
rect 282 326 318 353
rect 406 336 442 353
rect 501 336 537 353
rect 625 336 661 353
rect 723 336 759 353
rect 192 310 345 326
rect 192 290 295 310
rect 25 260 119 276
rect 186 276 295 290
rect 329 276 345 310
rect 186 260 345 276
rect 393 320 459 336
rect 393 286 409 320
rect 443 286 459 320
rect 393 270 459 286
rect 501 320 567 336
rect 501 286 517 320
rect 551 286 567 320
rect 501 270 567 286
rect 615 320 681 336
rect 615 286 631 320
rect 665 286 681 320
rect 615 270 681 286
rect 723 320 789 336
rect 723 286 739 320
rect 773 286 789 320
rect 723 270 789 286
rect 84 222 114 260
rect 186 222 216 260
rect 272 222 302 260
rect 429 222 459 270
rect 507 222 537 270
rect 615 222 645 270
rect 723 222 753 270
rect 84 86 114 112
rect 186 48 216 74
rect 272 48 302 74
rect 429 48 459 74
rect 507 48 537 74
rect 615 48 645 74
rect 723 48 753 74
<< polycont >>
rect 41 276 75 310
rect 295 276 329 310
rect 409 286 443 320
rect 517 286 551 320
rect 631 286 665 320
rect 739 286 773 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 130 578 196 649
rect 130 544 146 578
rect 180 544 196 578
rect 130 542 196 544
rect 329 578 395 649
rect 329 544 345 578
rect 379 544 395 578
rect 329 542 395 544
rect 548 578 614 649
rect 548 544 564 578
rect 598 544 614 578
rect 548 542 614 544
rect 770 578 841 649
rect 770 544 788 578
rect 822 544 841 578
rect 770 542 841 544
rect 23 524 89 540
rect 23 490 39 524
rect 73 508 89 524
rect 73 490 797 508
rect 23 474 797 490
rect 23 440 159 474
rect 23 406 39 440
rect 73 406 159 440
rect 23 390 159 406
rect 25 310 91 356
rect 25 276 41 310
rect 75 276 91 310
rect 25 260 91 276
rect 125 226 159 390
rect 23 192 159 226
rect 211 419 288 440
rect 211 385 238 419
rect 272 385 288 419
rect 211 364 288 385
rect 322 424 729 440
rect 322 390 454 424
rect 488 390 675 424
rect 709 390 729 424
rect 211 226 245 364
rect 322 326 356 390
rect 279 310 356 326
rect 279 276 295 310
rect 329 276 356 310
rect 279 260 356 276
rect 393 320 459 356
rect 393 286 409 320
rect 443 286 459 320
rect 393 270 459 286
rect 501 320 567 356
rect 501 286 517 320
rect 551 286 567 320
rect 501 270 567 286
rect 601 320 681 356
rect 763 336 797 474
rect 601 286 631 320
rect 665 286 681 320
rect 601 270 681 286
rect 723 320 797 336
rect 723 286 739 320
rect 773 286 797 320
rect 723 270 797 286
rect 322 226 356 260
rect 211 210 277 226
rect 23 184 89 192
rect 23 150 39 184
rect 73 150 89 184
rect 211 176 227 210
rect 261 176 277 210
rect 322 210 814 226
rect 322 192 764 210
rect 23 108 89 150
rect 125 142 175 158
rect 125 108 141 142
rect 125 17 175 108
rect 211 120 277 176
rect 748 176 764 192
rect 798 176 814 210
rect 211 86 227 120
rect 261 86 277 120
rect 211 70 277 86
rect 311 142 433 158
rect 311 108 313 142
rect 347 108 384 142
rect 418 108 433 142
rect 311 17 433 108
rect 748 120 814 176
rect 748 86 764 120
rect 798 86 814 120
rect 748 70 814 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel comment s 0 0 0 0 4 and4b_2
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 223 390 257 424 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 D
port 4 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 B
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 864 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3194862
string GDS_START 3188264
<< end >>
