magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 828 561
rect 103 441 169 527
rect 85 199 155 339
rect 189 199 247 265
rect 496 425 624 491
rect 658 367 714 527
rect 756 299 811 493
rect 523 199 654 265
rect 131 17 165 165
rect 777 152 811 299
rect 294 17 369 97
rect 474 17 540 97
rect 642 17 718 97
rect 756 83 811 152
rect 0 -17 828 17
<< obsli1 >>
rect 17 407 69 491
rect 302 441 451 475
rect 17 373 383 407
rect 17 165 51 373
rect 198 305 315 339
rect 281 249 315 305
rect 349 317 383 373
rect 417 391 451 441
rect 417 357 624 391
rect 590 333 624 357
rect 349 283 479 317
rect 590 299 722 333
rect 281 215 366 249
rect 281 165 315 215
rect 445 199 479 283
rect 688 265 722 299
rect 688 199 743 265
rect 688 165 722 199
rect 17 90 80 165
rect 215 131 315 165
rect 403 131 722 165
rect 215 90 249 131
rect 403 61 437 131
rect 574 61 608 131
<< metal1 >>
rect 0 496 828 592
rect 0 -48 828 48
<< labels >>
rlabel locali s 523 199 654 265 6 A
port 1 nsew signal input
rlabel locali s 496 425 624 491 6 B
port 2 nsew signal input
rlabel locali s 85 199 155 339 6 C_N
port 3 nsew signal input
rlabel locali s 189 199 247 265 6 D_N
port 4 nsew signal input
rlabel locali s 777 152 811 299 6 X
port 5 nsew signal output
rlabel locali s 756 299 811 493 6 X
port 5 nsew signal output
rlabel locali s 756 83 811 152 6 X
port 5 nsew signal output
rlabel locali s 642 17 718 97 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 474 17 540 97 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 294 17 369 97 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 131 17 165 165 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 828 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 828 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 658 367 714 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 103 441 169 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 828 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 828 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1112386
string GDS_START 1105338
<< end >>
