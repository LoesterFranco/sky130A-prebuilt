magic
tech sky130A
magscale 1 2
timestamp 1604502697
<< nwell >>
rect -38 261 2154 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 93 47 123 177
rect 187 47 217 177
rect 281 47 311 177
rect 375 47 405 177
rect 473 47 503 177
rect 567 47 597 177
rect 661 47 691 177
rect 855 47 885 177
rect 949 47 979 177
rect 1043 47 1073 177
rect 1147 47 1177 177
rect 1241 47 1271 177
rect 1345 47 1375 177
rect 1429 47 1459 177
rect 1523 47 1553 177
rect 1617 47 1647 177
rect 1721 47 1751 177
rect 1805 47 1835 177
rect 1899 47 1929 177
rect 1993 47 2023 177
<< pmoshvt >>
rect 85 297 121 497
rect 179 297 215 497
rect 273 297 309 497
rect 367 297 403 497
rect 575 297 611 497
rect 669 297 705 497
rect 763 297 799 497
rect 857 297 893 497
rect 951 297 987 497
rect 1045 297 1081 497
rect 1139 297 1175 497
rect 1233 297 1269 497
rect 1337 297 1373 497
rect 1431 297 1467 497
rect 1525 297 1561 497
rect 1619 297 1655 497
rect 1713 297 1749 497
rect 1807 297 1843 497
rect 1901 297 1937 497
rect 1995 297 2031 497
<< ndiff >>
rect 27 163 93 177
rect 27 129 39 163
rect 73 129 93 163
rect 27 95 93 129
rect 27 61 39 95
rect 73 61 93 95
rect 27 47 93 61
rect 123 163 187 177
rect 123 129 133 163
rect 167 129 187 163
rect 123 95 187 129
rect 123 61 133 95
rect 167 61 187 95
rect 123 47 187 61
rect 217 95 281 177
rect 217 61 227 95
rect 261 61 281 95
rect 217 47 281 61
rect 311 163 375 177
rect 311 129 321 163
rect 355 129 375 163
rect 311 95 375 129
rect 311 61 321 95
rect 355 61 375 95
rect 311 47 375 61
rect 405 95 473 177
rect 405 61 415 95
rect 449 61 473 95
rect 405 47 473 61
rect 503 95 567 177
rect 503 61 513 95
rect 547 61 567 95
rect 503 47 567 61
rect 597 169 661 177
rect 597 135 607 169
rect 641 135 661 169
rect 597 47 661 135
rect 691 95 855 177
rect 691 61 701 95
rect 735 61 811 95
rect 845 61 855 95
rect 691 47 855 61
rect 885 163 949 177
rect 885 129 905 163
rect 939 129 949 163
rect 885 47 949 129
rect 979 95 1043 177
rect 979 61 999 95
rect 1033 61 1043 95
rect 979 47 1043 61
rect 1073 163 1147 177
rect 1073 129 1093 163
rect 1127 129 1147 163
rect 1073 47 1147 129
rect 1177 95 1241 177
rect 1177 61 1187 95
rect 1221 61 1241 95
rect 1177 47 1241 61
rect 1271 95 1345 177
rect 1271 61 1291 95
rect 1325 61 1345 95
rect 1271 47 1345 61
rect 1375 95 1429 177
rect 1375 61 1385 95
rect 1419 61 1429 95
rect 1375 47 1429 61
rect 1459 163 1523 177
rect 1459 129 1479 163
rect 1513 129 1523 163
rect 1459 47 1523 129
rect 1553 95 1617 177
rect 1553 61 1573 95
rect 1607 61 1617 95
rect 1553 47 1617 61
rect 1647 163 1721 177
rect 1647 129 1667 163
rect 1701 129 1721 163
rect 1647 47 1721 129
rect 1751 163 1805 177
rect 1751 129 1761 163
rect 1795 129 1805 163
rect 1751 95 1805 129
rect 1751 61 1761 95
rect 1795 61 1805 95
rect 1751 47 1805 61
rect 1835 95 1899 177
rect 1835 61 1855 95
rect 1889 61 1899 95
rect 1835 47 1899 61
rect 1929 163 1993 177
rect 1929 129 1949 163
rect 1983 129 1993 163
rect 1929 95 1993 129
rect 1929 61 1949 95
rect 1983 61 1993 95
rect 1929 47 1993 61
rect 2023 163 2080 177
rect 2023 129 2033 163
rect 2067 129 2080 163
rect 2023 95 2080 129
rect 2023 61 2033 95
rect 2067 61 2080 95
rect 2023 47 2080 61
<< pdiff >>
rect 27 477 85 497
rect 27 443 39 477
rect 73 443 85 477
rect 27 409 85 443
rect 27 375 39 409
rect 73 375 85 409
rect 27 341 85 375
rect 27 307 39 341
rect 73 307 85 341
rect 27 297 85 307
rect 121 409 179 497
rect 121 375 133 409
rect 167 375 179 409
rect 121 341 179 375
rect 121 307 133 341
rect 167 307 179 341
rect 121 297 179 307
rect 215 477 273 497
rect 215 443 227 477
rect 261 443 273 477
rect 215 409 273 443
rect 215 375 227 409
rect 261 375 273 409
rect 215 297 273 375
rect 309 409 367 497
rect 309 375 321 409
rect 355 375 367 409
rect 309 341 367 375
rect 309 307 321 341
rect 355 307 367 341
rect 309 297 367 307
rect 403 479 457 497
rect 403 445 415 479
rect 449 445 457 479
rect 403 411 457 445
rect 403 377 415 411
rect 449 377 457 411
rect 403 343 457 377
rect 403 309 415 343
rect 449 309 457 343
rect 403 297 457 309
rect 511 477 575 497
rect 511 443 529 477
rect 563 443 575 477
rect 511 409 575 443
rect 511 375 529 409
rect 563 375 575 409
rect 511 297 575 375
rect 611 409 669 497
rect 611 375 623 409
rect 657 375 669 409
rect 611 341 669 375
rect 611 307 623 341
rect 657 307 669 341
rect 611 297 669 307
rect 705 477 763 497
rect 705 443 717 477
rect 751 443 763 477
rect 705 297 763 443
rect 799 409 857 497
rect 799 375 811 409
rect 845 375 857 409
rect 799 297 857 375
rect 893 477 951 497
rect 893 443 905 477
rect 939 443 951 477
rect 893 297 951 443
rect 987 409 1045 497
rect 987 375 999 409
rect 1033 375 1045 409
rect 987 297 1045 375
rect 1081 477 1139 497
rect 1081 443 1093 477
rect 1127 443 1139 477
rect 1081 297 1139 443
rect 1175 409 1233 497
rect 1175 375 1187 409
rect 1221 375 1233 409
rect 1175 297 1233 375
rect 1269 477 1337 497
rect 1269 443 1289 477
rect 1323 443 1337 477
rect 1269 409 1337 443
rect 1269 375 1289 409
rect 1323 375 1337 409
rect 1269 297 1337 375
rect 1373 477 1431 497
rect 1373 443 1385 477
rect 1419 443 1431 477
rect 1373 297 1431 443
rect 1467 409 1525 497
rect 1467 375 1479 409
rect 1513 375 1525 409
rect 1467 297 1525 375
rect 1561 477 1619 497
rect 1561 443 1573 477
rect 1607 443 1619 477
rect 1561 297 1619 443
rect 1655 409 1713 497
rect 1655 375 1667 409
rect 1701 375 1713 409
rect 1655 297 1713 375
rect 1749 477 1807 497
rect 1749 443 1761 477
rect 1795 443 1807 477
rect 1749 297 1807 443
rect 1843 477 1901 497
rect 1843 443 1855 477
rect 1889 443 1901 477
rect 1843 409 1901 443
rect 1843 375 1855 409
rect 1889 375 1901 409
rect 1843 297 1901 375
rect 1937 477 1995 497
rect 1937 443 1949 477
rect 1983 443 1995 477
rect 1937 409 1995 443
rect 1937 375 1949 409
rect 1983 375 1995 409
rect 1937 297 1995 375
rect 2031 449 2089 497
rect 2031 415 2043 449
rect 2077 415 2089 449
rect 2031 381 2089 415
rect 2031 347 2043 381
rect 2077 347 2089 381
rect 2031 297 2089 347
<< ndiffc >>
rect 39 129 73 163
rect 39 61 73 95
rect 133 129 167 163
rect 133 61 167 95
rect 227 61 261 95
rect 321 129 355 163
rect 321 61 355 95
rect 415 61 449 95
rect 513 61 547 95
rect 607 135 641 169
rect 701 61 735 95
rect 811 61 845 95
rect 905 129 939 163
rect 999 61 1033 95
rect 1093 129 1127 163
rect 1187 61 1221 95
rect 1291 61 1325 95
rect 1385 61 1419 95
rect 1479 129 1513 163
rect 1573 61 1607 95
rect 1667 129 1701 163
rect 1761 129 1795 163
rect 1761 61 1795 95
rect 1855 61 1889 95
rect 1949 129 1983 163
rect 1949 61 1983 95
rect 2033 129 2067 163
rect 2033 61 2067 95
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 133 375 167 409
rect 133 307 167 341
rect 227 443 261 477
rect 227 375 261 409
rect 321 375 355 409
rect 321 307 355 341
rect 415 445 449 479
rect 415 377 449 411
rect 415 309 449 343
rect 529 443 563 477
rect 529 375 563 409
rect 623 375 657 409
rect 623 307 657 341
rect 717 443 751 477
rect 811 375 845 409
rect 905 443 939 477
rect 999 375 1033 409
rect 1093 443 1127 477
rect 1187 375 1221 409
rect 1289 443 1323 477
rect 1289 375 1323 409
rect 1385 443 1419 477
rect 1479 375 1513 409
rect 1573 443 1607 477
rect 1667 375 1701 409
rect 1761 443 1795 477
rect 1855 443 1889 477
rect 1855 375 1889 409
rect 1949 443 1983 477
rect 1949 375 1983 409
rect 2043 415 2077 449
rect 2043 347 2077 381
<< poly >>
rect 85 497 121 523
rect 179 497 215 523
rect 273 497 309 523
rect 367 497 403 523
rect 575 497 611 523
rect 669 497 705 523
rect 763 497 799 523
rect 857 497 893 523
rect 951 497 987 523
rect 1045 497 1081 523
rect 1139 497 1175 523
rect 1233 497 1269 523
rect 1337 497 1373 523
rect 1431 497 1467 523
rect 1525 497 1561 523
rect 1619 497 1655 523
rect 1713 497 1749 523
rect 1807 497 1843 523
rect 1901 497 1937 523
rect 1995 497 2031 523
rect 85 282 121 297
rect 179 282 215 297
rect 273 282 309 297
rect 367 282 403 297
rect 575 282 611 297
rect 669 282 705 297
rect 763 282 799 297
rect 857 282 893 297
rect 951 282 987 297
rect 1045 282 1081 297
rect 1139 282 1175 297
rect 1233 282 1269 297
rect 1337 282 1373 297
rect 1431 282 1467 297
rect 1525 282 1561 297
rect 1619 282 1655 297
rect 1713 282 1749 297
rect 1807 282 1843 297
rect 1901 282 1937 297
rect 1995 282 2031 297
rect 83 265 123 282
rect 177 265 217 282
rect 271 265 311 282
rect 365 265 405 282
rect 573 265 613 282
rect 667 265 707 282
rect 761 265 801 282
rect 855 265 895 282
rect 949 265 989 282
rect 1043 265 1083 282
rect 1137 265 1177 282
rect 1231 265 1271 282
rect 1335 265 1375 282
rect 1429 265 1469 282
rect 1523 265 1563 282
rect 1617 265 1657 282
rect 1711 265 1751 282
rect 65 249 405 265
rect 65 215 81 249
rect 115 215 159 249
rect 193 215 237 249
rect 271 215 405 249
rect 65 199 405 215
rect 93 177 123 199
rect 187 177 217 199
rect 281 177 311 199
rect 375 177 405 199
rect 473 249 807 265
rect 473 215 753 249
rect 787 215 807 249
rect 473 199 807 215
rect 855 249 1177 265
rect 855 215 883 249
rect 917 215 961 249
rect 995 215 1039 249
rect 1073 215 1117 249
rect 1151 215 1177 249
rect 855 199 1177 215
rect 1219 249 1281 265
rect 1219 215 1229 249
rect 1263 215 1281 249
rect 1219 199 1281 215
rect 1323 249 1387 265
rect 1323 215 1333 249
rect 1367 215 1387 249
rect 1323 199 1387 215
rect 1429 249 1751 265
rect 1429 215 1445 249
rect 1479 215 1523 249
rect 1557 215 1601 249
rect 1635 215 1751 249
rect 1429 199 1751 215
rect 473 177 503 199
rect 567 177 597 199
rect 661 177 691 199
rect 855 177 885 199
rect 949 177 979 199
rect 1043 177 1073 199
rect 1147 177 1177 199
rect 1241 177 1271 199
rect 1345 177 1375 199
rect 1429 177 1459 199
rect 1523 177 1553 199
rect 1617 177 1647 199
rect 1721 177 1751 199
rect 1805 265 1845 282
rect 1899 265 1939 282
rect 1993 265 2033 282
rect 1805 249 2042 265
rect 1805 215 1821 249
rect 1855 215 1899 249
rect 1933 215 1977 249
rect 2011 215 2042 249
rect 1805 199 2042 215
rect 1805 177 1835 199
rect 1899 177 1929 199
rect 1993 177 2023 199
rect 93 21 123 47
rect 187 21 217 47
rect 281 21 311 47
rect 375 21 405 47
rect 473 21 503 47
rect 567 21 597 47
rect 661 21 691 47
rect 855 21 885 47
rect 949 21 979 47
rect 1043 21 1073 47
rect 1147 21 1177 47
rect 1241 21 1271 47
rect 1345 21 1375 47
rect 1429 21 1459 47
rect 1523 21 1553 47
rect 1617 21 1647 47
rect 1721 21 1751 47
rect 1805 21 1835 47
rect 1899 21 1929 47
rect 1993 21 2023 47
<< polycont >>
rect 81 215 115 249
rect 159 215 193 249
rect 237 215 271 249
rect 753 215 787 249
rect 883 215 917 249
rect 961 215 995 249
rect 1039 215 1073 249
rect 1117 215 1151 249
rect 1229 215 1263 249
rect 1333 215 1367 249
rect 1445 215 1479 249
rect 1523 215 1557 249
rect 1601 215 1635 249
rect 1821 215 1855 249
rect 1899 215 1933 249
rect 1977 215 2011 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 18 479 465 493
rect 18 477 415 479
rect 18 443 39 477
rect 73 459 227 477
rect 73 443 81 459
rect 18 409 81 443
rect 219 443 227 459
rect 261 459 415 477
rect 261 443 269 459
rect 18 375 39 409
rect 73 375 81 409
rect 18 341 81 375
rect 18 307 39 341
rect 73 307 81 341
rect 18 289 81 307
rect 125 409 175 425
rect 125 375 133 409
rect 167 375 175 409
rect 125 341 175 375
rect 219 409 269 443
rect 449 445 465 479
rect 219 375 227 409
rect 261 375 269 409
rect 219 357 269 375
rect 313 409 363 425
rect 313 375 321 409
rect 355 375 363 409
rect 125 307 133 341
rect 167 323 175 341
rect 313 341 363 375
rect 313 323 321 341
rect 167 307 321 323
rect 355 323 363 341
rect 415 411 465 445
rect 449 377 465 411
rect 415 343 465 377
rect 513 477 1331 493
rect 513 443 529 477
rect 563 443 717 477
rect 751 443 905 477
rect 939 443 1093 477
rect 1127 443 1289 477
rect 1323 443 1331 477
rect 1365 477 1817 527
rect 1365 443 1385 477
rect 1419 443 1573 477
rect 1607 443 1761 477
rect 1795 443 1817 477
rect 1855 477 1889 493
rect 513 409 563 443
rect 1281 409 1331 443
rect 1855 409 1889 443
rect 1949 477 1983 527
rect 1949 409 1983 443
rect 513 375 529 409
rect 513 359 563 375
rect 607 375 623 409
rect 657 375 811 409
rect 845 375 999 409
rect 1033 375 1187 409
rect 1221 375 1237 409
rect 607 367 1237 375
rect 1281 375 1289 409
rect 1323 375 1479 409
rect 1513 375 1667 409
rect 1701 375 1855 409
rect 1889 375 1905 409
rect 355 307 371 323
rect 125 289 371 307
rect 449 323 465 343
rect 607 341 666 367
rect 1281 357 1905 375
rect 1949 359 1983 375
rect 2035 449 2085 493
rect 2035 415 2043 449
rect 2077 415 2085 449
rect 2035 381 2085 415
rect 607 323 623 341
rect 449 309 623 323
rect 415 307 623 309
rect 657 307 666 341
rect 1871 323 1905 357
rect 2035 347 2043 381
rect 2077 347 2085 381
rect 2035 323 2085 347
rect 415 289 666 307
rect 789 289 1282 323
rect 331 255 371 289
rect 789 265 833 289
rect 18 249 287 255
rect 18 215 81 249
rect 115 215 159 249
rect 193 215 237 249
rect 271 215 287 249
rect 331 219 719 255
rect 331 181 371 219
rect 23 163 73 179
rect 23 129 39 163
rect 23 95 73 129
rect 23 61 39 95
rect 23 17 73 61
rect 107 163 371 181
rect 107 129 133 163
rect 167 145 321 163
rect 167 129 183 145
rect 107 95 183 129
rect 295 129 321 145
rect 355 129 371 163
rect 107 61 133 95
rect 167 61 183 95
rect 107 51 183 61
rect 227 95 261 111
rect 227 17 261 61
rect 295 95 371 129
rect 295 61 321 95
rect 355 61 371 95
rect 295 51 371 61
rect 415 169 641 185
rect 415 135 607 169
rect 415 129 641 135
rect 675 164 719 219
rect 753 249 833 265
rect 787 215 833 249
rect 753 199 833 215
rect 867 249 1177 255
rect 867 215 883 249
rect 917 215 961 249
rect 995 215 1039 249
rect 1073 215 1117 249
rect 1151 215 1177 249
rect 1213 249 1282 289
rect 1213 215 1229 249
rect 1263 215 1282 249
rect 1317 289 1827 323
rect 1871 289 2085 323
rect 1317 249 1393 289
rect 1793 255 1827 289
rect 1317 215 1333 249
rect 1367 215 1393 249
rect 1429 249 1751 255
rect 1429 215 1445 249
rect 1479 215 1523 249
rect 1557 215 1601 249
rect 1635 215 1751 249
rect 1793 249 2080 255
rect 1793 215 1821 249
rect 1855 215 1899 249
rect 1933 215 1977 249
rect 2011 215 2080 249
rect 867 199 1177 215
rect 1222 164 1426 181
rect 675 163 1717 164
rect 675 129 905 163
rect 939 129 1093 163
rect 1127 147 1479 163
rect 1127 129 1256 147
rect 1392 129 1479 147
rect 1513 129 1667 163
rect 1701 129 1717 163
rect 1761 163 1999 181
rect 1795 145 1949 163
rect 1795 129 1811 145
rect 415 95 449 129
rect 607 119 641 129
rect 1291 95 1325 111
rect 1761 95 1811 129
rect 1923 129 1949 145
rect 1983 129 1999 163
rect 415 17 449 61
rect 487 61 513 95
rect 547 85 572 95
rect 667 85 701 95
rect 547 61 701 85
rect 735 61 811 95
rect 845 61 999 95
rect 1033 61 1187 95
rect 1221 61 1237 95
rect 487 51 1237 61
rect 1291 17 1325 61
rect 1359 61 1385 95
rect 1419 61 1573 95
rect 1607 61 1761 95
rect 1795 61 1811 95
rect 1359 51 1811 61
rect 1855 95 1889 111
rect 1855 17 1889 61
rect 1923 95 1999 129
rect 1923 61 1949 95
rect 1983 61 1999 95
rect 1923 51 1999 61
rect 2033 163 2067 181
rect 2033 95 2067 129
rect 2033 17 2067 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
<< metal1 >>
rect 0 561 2116 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 0 496 2116 527
rect 0 17 2116 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
rect 0 -48 2116 -17
<< labels >>
flabel corelocali s 1860 238 1860 238 0 FreeSans 400 180 0 0 A2
port 2 nsew
flabel corelocali s 336 221 370 255 0 FreeSans 400 180 0 0 Y
port 10 nsew
flabel corelocali s 214 221 248 255 0 FreeSans 400 0 0 0 C1
port 5 nsew
flabel corelocali s 1502 221 1536 255 0 FreeSans 400 180 0 0 A1
port 1 nsew
flabel corelocali s 850 289 884 323 0 FreeSans 400 0 0 0 B2
port 4 nsew
flabel corelocali s 952 221 986 255 0 FreeSans 400 0 0 0 B1
port 3 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 2116 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1245370
string GDS_START 1231422
<< end >>
