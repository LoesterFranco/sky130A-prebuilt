magic
tech sky130A
magscale 1 2
timestamp 1599588244
<< locali >>
rect 25 270 114 356
rect 713 394 766 596
rect 899 394 949 596
rect 1077 394 1131 596
rect 1257 394 1311 596
rect 713 360 1311 394
rect 1251 356 1311 360
rect 1251 254 1415 356
rect 1251 226 1317 254
rect 695 176 1317 226
rect 695 70 761 176
rect 1251 70 1317 176
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 23 440 76 540
rect 113 474 184 649
rect 23 390 184 440
rect 150 326 184 390
rect 218 364 296 596
rect 330 398 396 596
rect 430 432 476 649
rect 510 398 576 596
rect 330 364 576 398
rect 610 364 676 649
rect 807 428 858 649
rect 986 428 1041 649
rect 1167 428 1221 649
rect 262 326 296 364
rect 534 326 576 364
rect 1347 390 1408 649
rect 150 260 228 326
rect 262 260 500 326
rect 534 260 1204 326
rect 150 236 184 260
rect 23 202 184 236
rect 262 226 296 260
rect 534 226 625 260
rect 23 108 89 202
rect 125 17 191 168
rect 225 70 296 226
rect 337 176 625 226
rect 337 70 387 176
rect 423 17 489 142
rect 595 17 661 142
rect 795 17 861 142
rect 967 17 1033 142
rect 1151 17 1217 142
rect 1351 17 1417 220
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 683 1440 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 0 617 1440 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 1440 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -49 1440 -17
<< labels >>
rlabel locali s 25 270 114 356 6 A
port 1 nsew signal input
rlabel locali s 1257 394 1311 596 6 X
port 2 nsew signal output
rlabel locali s 1251 356 1311 360 6 X
port 2 nsew signal output
rlabel locali s 1251 254 1415 356 6 X
port 2 nsew signal output
rlabel locali s 1251 226 1317 254 6 X
port 2 nsew signal output
rlabel locali s 1251 70 1317 176 6 X
port 2 nsew signal output
rlabel locali s 1077 394 1131 596 6 X
port 2 nsew signal output
rlabel locali s 899 394 949 596 6 X
port 2 nsew signal output
rlabel locali s 713 394 766 596 6 X
port 2 nsew signal output
rlabel locali s 713 360 1311 394 6 X
port 2 nsew signal output
rlabel locali s 695 176 1317 226 6 X
port 2 nsew signal output
rlabel locali s 695 70 761 176 6 X
port 2 nsew signal output
rlabel metal1 s 0 -49 1440 49 8 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 4 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 617 1440 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1440 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3321776
string GDS_START 3311222
<< end >>
