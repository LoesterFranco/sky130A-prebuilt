magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 1671 378 1705 547
rect 1851 378 1885 547
rect 105 270 375 356
rect 409 270 743 356
rect 927 270 1223 356
rect 1671 344 1885 378
rect 1355 264 1557 330
rect 1355 236 1511 264
rect 1613 244 1815 310
rect 1657 236 1815 244
rect 866 202 1276 226
rect 1552 202 1602 210
rect 1851 202 1885 344
rect 866 170 1885 202
rect 866 154 932 170
rect 1226 168 1885 170
rect 1226 70 1276 168
rect 1552 70 1602 168
rect 1740 134 1885 168
rect 1740 70 1991 134
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 21 364 71 649
rect 111 424 161 596
rect 201 458 267 649
rect 307 424 341 596
rect 381 458 447 649
rect 487 424 521 596
rect 561 458 627 649
rect 667 424 701 596
rect 741 458 807 649
rect 847 424 881 596
rect 921 458 971 649
rect 1011 424 1061 596
rect 1101 458 1167 649
rect 1205 581 1991 615
rect 1205 464 1271 581
rect 1305 430 1351 547
rect 1385 464 1451 581
rect 1485 430 1531 547
rect 1295 424 1531 430
rect 111 390 1531 424
rect 847 364 881 390
rect 1295 364 1531 390
rect 1565 364 1631 581
rect 1745 412 1811 581
rect 1925 364 1991 581
rect 30 202 784 236
rect 30 70 80 202
rect 116 17 166 168
rect 202 70 252 202
rect 390 195 784 202
rect 288 17 354 168
rect 390 70 424 195
rect 546 154 612 195
rect 718 154 784 195
rect 460 120 512 136
rect 646 120 684 136
rect 1124 120 1190 136
rect 460 70 1190 120
rect 1310 17 1518 134
rect 1638 17 1704 134
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
rlabel locali s 927 270 1223 356 6 A1
port 1 nsew signal input
rlabel locali s 409 270 743 356 6 A2
port 2 nsew signal input
rlabel locali s 105 270 375 356 6 A3
port 3 nsew signal input
rlabel locali s 1355 264 1557 330 6 B1
port 4 nsew signal input
rlabel locali s 1355 236 1511 264 6 B1
port 4 nsew signal input
rlabel locali s 1657 236 1815 244 6 C1
port 5 nsew signal input
rlabel locali s 1613 244 1815 310 6 C1
port 5 nsew signal input
rlabel locali s 1851 378 1885 547 6 Y
port 6 nsew signal output
rlabel locali s 1851 202 1885 344 6 Y
port 6 nsew signal output
rlabel locali s 1740 134 1885 168 6 Y
port 6 nsew signal output
rlabel locali s 1740 70 1991 134 6 Y
port 6 nsew signal output
rlabel locali s 1671 378 1705 547 6 Y
port 6 nsew signal output
rlabel locali s 1671 344 1885 378 6 Y
port 6 nsew signal output
rlabel locali s 1552 202 1602 210 6 Y
port 6 nsew signal output
rlabel locali s 1552 70 1602 168 6 Y
port 6 nsew signal output
rlabel locali s 1226 168 1885 170 6 Y
port 6 nsew signal output
rlabel locali s 1226 70 1276 168 6 Y
port 6 nsew signal output
rlabel locali s 866 202 1276 226 6 Y
port 6 nsew signal output
rlabel locali s 866 170 1885 202 6 Y
port 6 nsew signal output
rlabel locali s 866 154 932 170 6 Y
port 6 nsew signal output
rlabel metal1 s 0 -49 2016 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 617 2016 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2016 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3689342
string GDS_START 3672944
<< end >>
