magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 22 215 89 273
rect 201 215 279 265
rect 388 283 687 341
rect 653 181 687 283
rect 1130 215 1561 257
rect 1615 215 2002 257
rect 407 145 1903 181
rect 407 51 483 145
rect 595 51 671 145
rect 783 51 859 145
rect 971 51 1047 145
rect 1263 51 1339 145
rect 1451 51 1527 145
rect 1639 51 1715 145
rect 1827 51 1903 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 17 409 73 493
rect 107 443 183 527
rect 323 459 1139 493
rect 323 443 765 459
rect 17 375 765 409
rect 17 307 167 375
rect 201 307 347 341
rect 133 179 167 307
rect 313 249 347 307
rect 313 215 619 249
rect 313 181 347 215
rect 731 257 765 375
rect 809 325 851 425
rect 895 359 945 459
rect 989 325 1039 425
rect 1083 359 1139 459
rect 1176 459 1613 493
rect 1176 359 1237 459
rect 1281 325 1331 425
rect 1375 359 1425 459
rect 1469 325 1519 425
rect 809 291 1519 325
rect 1563 325 1613 459
rect 1657 359 1707 527
rect 1751 325 1801 493
rect 1845 359 1895 527
rect 1939 325 2002 493
rect 1563 291 2002 325
rect 731 215 1081 257
rect 17 145 167 179
rect 201 147 347 181
rect 17 51 89 145
rect 133 17 167 111
rect 201 51 277 147
rect 339 17 373 111
rect 527 17 561 111
rect 715 17 749 111
rect 903 17 937 111
rect 1091 17 1229 111
rect 1383 17 1417 111
rect 1571 17 1605 111
rect 1759 17 1793 111
rect 1947 17 2002 181
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
<< metal1 >>
rect 0 561 2024 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 0 496 2024 527
rect 0 17 2024 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
rect 0 -48 2024 -17
<< labels >>
rlabel locali s 1615 215 2002 257 6 A
port 1 nsew signal input
rlabel locali s 1130 215 1561 257 6 B
port 2 nsew signal input
rlabel locali s 22 215 89 273 6 C_N
port 3 nsew signal input
rlabel locali s 201 215 279 265 6 D_N
port 4 nsew signal input
rlabel locali s 1827 51 1903 145 6 Y
port 5 nsew signal output
rlabel locali s 1639 51 1715 145 6 Y
port 5 nsew signal output
rlabel locali s 1451 51 1527 145 6 Y
port 5 nsew signal output
rlabel locali s 1263 51 1339 145 6 Y
port 5 nsew signal output
rlabel locali s 971 51 1047 145 6 Y
port 5 nsew signal output
rlabel locali s 783 51 859 145 6 Y
port 5 nsew signal output
rlabel locali s 653 181 687 283 6 Y
port 5 nsew signal output
rlabel locali s 595 51 671 145 6 Y
port 5 nsew signal output
rlabel locali s 407 145 1903 181 6 Y
port 5 nsew signal output
rlabel locali s 407 51 483 145 6 Y
port 5 nsew signal output
rlabel locali s 388 283 687 341 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -48 2024 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 2024 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2024 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2561144
string GDS_START 2546800
<< end >>
