magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 103 333 179 493
rect 291 333 367 493
rect 479 333 555 493
rect 667 333 743 493
rect 103 299 743 333
rect 22 215 376 265
rect 479 161 539 299
rect 573 215 823 265
rect 479 127 743 161
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 18 299 69 527
rect 223 367 257 527
rect 411 367 445 527
rect 599 367 633 527
rect 787 367 837 527
rect 18 143 445 181
rect 18 51 85 143
rect 129 17 163 109
rect 197 51 273 143
rect 317 17 351 109
rect 385 93 445 143
rect 787 93 837 177
rect 385 51 837 93
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
rlabel locali s 573 215 823 265 6 A
port 1 nsew signal input
rlabel locali s 22 215 376 265 6 B
port 2 nsew signal input
rlabel locali s 667 333 743 493 6 Y
port 3 nsew signal output
rlabel locali s 479 333 555 493 6 Y
port 3 nsew signal output
rlabel locali s 479 161 539 299 6 Y
port 3 nsew signal output
rlabel locali s 479 127 743 161 6 Y
port 3 nsew signal output
rlabel locali s 291 333 367 493 6 Y
port 3 nsew signal output
rlabel locali s 103 333 179 493 6 Y
port 3 nsew signal output
rlabel locali s 103 299 743 333 6 Y
port 3 nsew signal output
rlabel metal1 s 0 -48 920 48 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 496 920 592 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 920 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2204542
string GDS_START 2196624
<< end >>
