magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 2484 561
rect 113 452 186 527
rect 413 447 479 527
rect 190 215 288 255
rect 403 282 438 345
rect 398 255 438 282
rect 398 215 499 255
rect 119 17 153 109
rect 402 17 436 109
rect 1135 199 1185 265
rect 1968 455 2035 527
rect 1895 215 1973 265
rect 1938 187 1973 215
rect 1938 147 2002 187
rect 1981 17 2015 113
rect 2174 299 2278 493
rect 2312 357 2363 527
rect 2397 357 2467 493
rect 2174 165 2208 299
rect 2422 165 2467 357
rect 2174 54 2262 165
rect 2296 17 2362 165
rect 2396 51 2467 165
rect 0 -17 2484 17
<< obsli1 >>
rect 17 413 79 493
rect 527 459 990 493
rect 1025 459 1512 493
rect 527 413 561 459
rect 17 379 561 413
rect 606 391 864 425
rect 17 300 89 379
rect 197 323 263 343
rect 17 161 51 300
rect 123 291 263 323
rect 122 289 263 291
rect 298 300 368 345
rect 298 289 364 300
rect 122 276 163 289
rect 122 265 156 276
rect 85 199 156 265
rect 119 181 156 199
rect 323 181 364 289
rect 472 323 572 343
rect 472 289 490 323
rect 524 289 572 323
rect 17 51 85 161
rect 119 147 264 181
rect 198 51 264 147
rect 300 177 364 181
rect 300 143 504 177
rect 300 51 368 143
rect 470 85 504 143
rect 538 119 572 289
rect 606 93 640 391
rect 831 357 864 391
rect 674 291 763 357
rect 674 187 708 291
rect 814 289 873 323
rect 814 232 907 289
rect 814 215 880 232
rect 941 185 975 459
rect 1025 264 1059 459
rect 1095 391 1175 406
rect 1095 357 1114 391
rect 1148 357 1175 391
rect 1095 340 1175 357
rect 1258 391 1444 425
rect 1258 323 1292 391
rect 1221 289 1230 323
rect 1264 289 1292 323
rect 1025 230 1101 264
rect 1064 185 1101 230
rect 1342 255 1376 357
rect 1221 187 1287 255
rect 896 181 1029 185
rect 814 161 1029 181
rect 1064 173 1104 185
rect 1067 168 1104 173
rect 708 153 780 161
rect 674 127 780 153
rect 814 156 1031 161
rect 814 151 1034 156
rect 814 147 912 151
rect 985 148 1034 151
rect 985 147 1036 148
rect 814 129 880 147
rect 990 143 1036 147
rect 996 138 1036 143
rect 1000 131 1036 138
rect 930 93 968 117
rect 606 85 968 93
rect 470 51 968 85
rect 1002 85 1036 131
rect 1070 119 1104 168
rect 1221 153 1230 187
rect 1264 153 1287 187
rect 1221 148 1287 153
rect 1356 221 1376 255
rect 1322 185 1376 221
rect 1410 235 1444 391
rect 1478 285 1512 459
rect 1546 459 1931 493
rect 1546 302 1592 459
rect 1629 391 1850 425
rect 1478 280 1515 285
rect 1478 275 1519 280
rect 1478 255 1524 275
rect 1410 226 1449 235
rect 1410 212 1456 226
rect 1413 209 1456 212
rect 1418 202 1456 209
rect 1322 151 1388 185
rect 1354 119 1388 151
rect 1422 153 1456 202
rect 1490 199 1524 255
rect 1558 165 1592 302
rect 1645 323 1782 357
rect 1645 289 1692 323
rect 1726 289 1782 323
rect 1645 185 1681 289
rect 1816 255 1850 357
rect 1884 341 1931 459
rect 2069 391 2138 493
rect 2069 375 2104 391
rect 1884 299 2070 341
rect 1422 119 1489 153
rect 1150 85 1220 113
rect 1002 51 1220 85
rect 1254 85 1320 114
rect 1541 85 1592 165
rect 1631 119 1681 185
rect 1715 221 1850 255
rect 1715 119 1749 221
rect 2036 199 2070 299
rect 1818 153 1860 187
rect 1784 137 1860 153
rect 2104 165 2138 357
rect 1880 85 1947 103
rect 1254 51 1947 85
rect 2049 57 2138 165
rect 2326 289 2336 323
rect 2370 289 2388 323
rect 2242 255 2292 265
rect 2242 221 2244 255
rect 2278 221 2292 255
rect 2242 199 2292 221
rect 2326 199 2388 289
<< obsli1c >>
rect 490 289 524 323
rect 797 357 831 391
rect 873 289 907 323
rect 674 153 708 187
rect 1114 357 1148 391
rect 1230 289 1264 323
rect 1230 153 1264 187
rect 1322 221 1356 255
rect 1816 357 1850 391
rect 1692 289 1726 323
rect 2104 357 2138 391
rect 1784 153 1818 187
rect 2336 289 2370 323
rect 2244 221 2278 255
<< metal1 >>
rect 0 496 2484 592
rect 386 252 444 261
rect 1124 252 1182 261
rect 386 224 1182 252
rect 386 215 444 224
rect 1124 215 1182 224
rect 0 -48 2484 48
<< obsm1 >>
rect 785 391 843 397
rect 785 357 797 391
rect 831 388 843 391
rect 1102 391 1160 397
rect 1102 388 1114 391
rect 831 360 1114 388
rect 831 357 843 360
rect 785 351 843 357
rect 1102 357 1114 360
rect 1148 357 1160 391
rect 1102 351 1160 357
rect 1804 391 1862 397
rect 1804 357 1816 391
rect 1850 388 1862 391
rect 2092 391 2150 397
rect 2092 388 2104 391
rect 1850 360 2104 388
rect 1850 357 1862 360
rect 1804 351 1862 357
rect 2092 357 2104 360
rect 2138 357 2150 391
rect 2092 351 2150 357
rect 478 323 536 329
rect 478 289 490 323
rect 524 320 536 323
rect 861 323 919 329
rect 861 320 873 323
rect 524 292 873 320
rect 524 289 536 292
rect 478 283 536 289
rect 861 289 873 292
rect 907 320 919 323
rect 1218 323 1276 329
rect 1218 320 1230 323
rect 907 292 1230 320
rect 907 289 919 292
rect 861 283 919 289
rect 1218 289 1230 292
rect 1264 289 1276 323
rect 1218 283 1276 289
rect 1680 323 1738 329
rect 1680 289 1692 323
rect 1726 320 1738 323
rect 2324 323 2382 329
rect 2324 320 2336 323
rect 1726 292 2336 320
rect 1726 289 1738 292
rect 1680 283 1738 289
rect 2324 289 2336 292
rect 2370 289 2382 323
rect 2324 283 2382 289
rect 1310 255 1368 261
rect 1310 221 1322 255
rect 1356 252 1368 255
rect 2232 255 2290 261
rect 2232 252 2244 255
rect 1356 224 2244 252
rect 1356 221 1368 224
rect 1310 215 1368 221
rect 2232 221 2244 224
rect 2278 221 2290 255
rect 2232 215 2290 221
rect 662 187 720 193
rect 662 153 674 187
rect 708 184 720 187
rect 1218 187 1276 193
rect 1218 184 1230 187
rect 708 156 1230 184
rect 708 153 720 156
rect 662 147 720 153
rect 1218 153 1230 156
rect 1264 184 1276 187
rect 1772 187 1830 193
rect 1772 184 1784 187
rect 1264 156 1784 184
rect 1264 153 1276 156
rect 1218 147 1276 153
rect 1772 153 1784 156
rect 1818 153 1830 187
rect 1772 147 1830 153
<< labels >>
rlabel locali s 190 215 288 255 6 A
port 1 nsew signal input
rlabel locali s 403 282 438 345 6 B
port 2 nsew signal input
rlabel locali s 398 255 438 282 6 B
port 2 nsew signal input
rlabel locali s 398 215 499 255 6 B
port 2 nsew signal input
rlabel locali s 1135 199 1185 265 6 B
port 2 nsew signal input
rlabel metal1 s 1124 252 1182 261 6 B
port 2 nsew signal input
rlabel metal1 s 1124 215 1182 224 6 B
port 2 nsew signal input
rlabel metal1 s 386 252 444 261 6 B
port 2 nsew signal input
rlabel metal1 s 386 224 1182 252 6 B
port 2 nsew signal input
rlabel metal1 s 386 215 444 224 6 B
port 2 nsew signal input
rlabel locali s 1938 187 1973 215 6 CI
port 3 nsew signal input
rlabel locali s 1938 147 2002 187 6 CI
port 3 nsew signal input
rlabel locali s 1895 215 1973 265 6 CI
port 3 nsew signal input
rlabel locali s 2174 299 2278 493 6 COUT
port 4 nsew signal output
rlabel locali s 2174 165 2208 299 6 COUT
port 4 nsew signal output
rlabel locali s 2174 54 2262 165 6 COUT
port 4 nsew signal output
rlabel locali s 2422 165 2467 357 6 SUM
port 5 nsew signal output
rlabel locali s 2397 357 2467 493 6 SUM
port 5 nsew signal output
rlabel locali s 2396 51 2467 165 6 SUM
port 5 nsew signal output
rlabel locali s 2296 17 2362 165 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1981 17 2015 113 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 402 17 436 109 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 119 17 153 109 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 2484 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 2484 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 2312 357 2363 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1968 455 2035 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 413 447 479 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 113 452 186 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 2484 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 2484 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2484 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2067956
string GDS_START 2048516
<< end >>
