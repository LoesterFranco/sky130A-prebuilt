magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 19 359 69 459
rect 19 297 331 359
rect 17 200 119 263
rect 153 200 247 263
rect 281 163 331 297
rect 377 200 449 266
rect 483 200 547 266
rect 581 200 661 266
rect 695 200 799 266
rect 19 129 595 163
rect 19 51 85 129
rect 482 59 595 129
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 113 459 493 493
rect 113 411 179 459
rect 434 427 493 459
rect 537 366 587 450
rect 631 381 697 527
rect 365 347 587 366
rect 753 347 805 450
rect 365 300 805 347
rect 185 17 341 93
rect 711 17 793 163
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
rlabel locali s 581 200 661 266 6 A1
port 1 nsew signal input
rlabel locali s 695 200 799 266 6 A2
port 2 nsew signal input
rlabel locali s 483 200 547 266 6 B1
port 3 nsew signal input
rlabel locali s 377 200 449 266 6 B2
port 4 nsew signal input
rlabel locali s 17 200 119 263 6 C1
port 5 nsew signal input
rlabel locali s 153 200 247 263 6 C2
port 6 nsew signal input
rlabel locali s 482 59 595 129 6 Y
port 7 nsew signal output
rlabel locali s 281 163 331 297 6 Y
port 7 nsew signal output
rlabel locali s 19 359 69 459 6 Y
port 7 nsew signal output
rlabel locali s 19 297 331 359 6 Y
port 7 nsew signal output
rlabel locali s 19 129 595 163 6 Y
port 7 nsew signal output
rlabel locali s 19 51 85 129 6 Y
port 7 nsew signal output
rlabel metal1 s 0 -48 828 48 8 VGND
port 8 nsew ground bidirectional
rlabel metal1 s 0 496 828 592 6 VPWR
port 9 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1252514
string GDS_START 1245430
<< end >>
