magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 1602 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 89 47 119 131
rect 174 47 204 131
rect 269 47 299 119
rect 385 47 415 119
rect 516 47 546 131
rect 635 47 665 177
rect 833 47 863 131
rect 927 47 957 131
rect 1155 47 1185 131
rect 1227 47 1257 131
rect 1344 47 1374 177
rect 1438 47 1468 177
<< pmoshvt >>
rect 81 369 117 497
rect 163 369 199 497
rect 268 413 304 497
rect 374 413 410 497
rect 486 413 522 497
rect 627 297 663 497
rect 825 303 861 431
rect 945 303 981 431
rect 1147 369 1183 497
rect 1241 369 1277 497
rect 1346 297 1382 497
rect 1440 297 1476 497
<< ndiff >>
rect 27 103 89 131
rect 27 69 35 103
rect 69 69 89 103
rect 27 47 89 69
rect 119 89 174 131
rect 119 55 129 89
rect 163 55 174 89
rect 119 47 174 55
rect 204 119 254 131
rect 570 131 635 177
rect 463 119 516 131
rect 204 101 269 119
rect 204 67 223 101
rect 257 67 269 101
rect 204 47 269 67
rect 299 89 385 119
rect 299 55 329 89
rect 363 55 385 89
rect 299 47 385 55
rect 415 47 516 119
rect 546 119 635 131
rect 546 85 582 119
rect 616 85 635 119
rect 546 47 635 85
rect 665 101 717 177
rect 1272 131 1344 177
rect 665 67 675 101
rect 709 67 717 101
rect 665 47 717 67
rect 771 110 833 131
rect 771 76 779 110
rect 813 76 833 110
rect 771 47 833 76
rect 863 89 927 131
rect 863 55 873 89
rect 907 55 927 89
rect 863 47 927 55
rect 957 110 1009 131
rect 957 76 967 110
rect 1001 76 1009 110
rect 957 47 1009 76
rect 1093 109 1155 131
rect 1093 75 1101 109
rect 1135 75 1155 109
rect 1093 47 1155 75
rect 1185 47 1227 131
rect 1257 89 1344 131
rect 1257 55 1284 89
rect 1318 55 1344 89
rect 1257 47 1344 55
rect 1374 89 1438 177
rect 1374 55 1384 89
rect 1418 55 1438 89
rect 1374 47 1438 55
rect 1468 93 1520 177
rect 1468 59 1478 93
rect 1512 59 1520 93
rect 1468 47 1520 59
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 369 81 383
rect 117 369 163 497
rect 199 475 268 497
rect 199 441 222 475
rect 256 441 268 475
rect 199 413 268 441
rect 304 475 374 497
rect 304 441 322 475
rect 356 441 374 475
rect 304 413 374 441
rect 410 413 486 497
rect 522 489 627 497
rect 522 455 560 489
rect 594 455 627 489
rect 522 413 627 455
rect 199 369 251 413
rect 575 297 627 413
rect 663 458 717 497
rect 663 424 675 458
rect 709 424 717 458
rect 878 485 928 497
rect 878 451 886 485
rect 920 451 928 485
rect 1089 489 1147 497
rect 878 431 928 451
rect 1089 455 1101 489
rect 1135 455 1147 489
rect 663 297 717 424
rect 771 349 825 431
rect 771 315 779 349
rect 813 315 825 349
rect 771 303 825 315
rect 861 303 945 431
rect 981 349 1035 431
rect 1089 369 1147 455
rect 1183 442 1241 497
rect 1183 408 1195 442
rect 1229 408 1241 442
rect 1183 369 1241 408
rect 1277 489 1346 497
rect 1277 455 1295 489
rect 1329 455 1346 489
rect 1277 369 1346 455
rect 981 315 993 349
rect 1027 315 1035 349
rect 981 303 1035 315
rect 1294 297 1346 369
rect 1382 448 1440 497
rect 1382 414 1394 448
rect 1428 414 1440 448
rect 1382 380 1440 414
rect 1382 346 1394 380
rect 1428 346 1440 380
rect 1382 297 1440 346
rect 1476 485 1530 497
rect 1476 451 1488 485
rect 1522 451 1530 485
rect 1476 417 1530 451
rect 1476 383 1488 417
rect 1522 383 1530 417
rect 1476 297 1530 383
<< ndiffc >>
rect 35 69 69 103
rect 129 55 163 89
rect 223 67 257 101
rect 329 55 363 89
rect 582 85 616 119
rect 675 67 709 101
rect 779 76 813 110
rect 873 55 907 89
rect 967 76 1001 110
rect 1101 75 1135 109
rect 1284 55 1318 89
rect 1384 55 1418 89
rect 1478 59 1512 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 222 441 256 475
rect 322 441 356 475
rect 560 455 594 489
rect 675 424 709 458
rect 886 451 920 485
rect 1101 455 1135 489
rect 779 315 813 349
rect 1195 408 1229 442
rect 1295 455 1329 489
rect 993 315 1027 349
rect 1394 414 1428 448
rect 1394 346 1428 380
rect 1488 451 1522 485
rect 1488 383 1522 417
<< poly >>
rect 81 497 117 523
rect 163 497 199 523
rect 268 497 304 523
rect 374 497 410 523
rect 486 497 522 523
rect 627 497 663 523
rect 268 398 304 413
rect 374 398 410 413
rect 486 398 522 413
rect 81 354 117 369
rect 163 354 199 369
rect 79 265 119 354
rect 22 249 119 265
rect 22 215 32 249
rect 66 215 119 249
rect 22 199 119 215
rect 161 265 201 354
rect 266 273 306 398
rect 372 381 412 398
rect 348 365 412 381
rect 348 331 358 365
rect 392 331 412 365
rect 348 315 412 331
rect 484 381 524 398
rect 484 365 546 381
rect 484 331 494 365
rect 528 331 546 365
rect 484 315 546 331
rect 161 249 222 265
rect 161 215 178 249
rect 212 215 222 249
rect 266 243 424 273
rect 161 199 222 215
rect 385 207 424 243
rect 89 131 119 199
rect 174 131 204 199
rect 269 191 343 201
rect 269 157 293 191
rect 327 157 343 191
rect 269 147 343 157
rect 385 191 448 207
rect 385 157 395 191
rect 429 157 448 191
rect 269 119 299 147
rect 385 141 448 157
rect 385 119 415 141
rect 516 131 546 315
rect 823 457 863 523
rect 825 431 861 457
rect 943 457 983 523
rect 1147 497 1183 523
rect 1241 497 1277 523
rect 1346 497 1382 523
rect 1440 497 1476 523
rect 945 431 981 457
rect 1147 354 1183 369
rect 1241 354 1277 369
rect 627 282 663 297
rect 825 288 861 303
rect 945 288 981 303
rect 625 265 665 282
rect 823 265 863 288
rect 943 265 983 288
rect 1145 265 1185 354
rect 1239 265 1279 354
rect 1346 282 1382 297
rect 1440 282 1476 297
rect 597 249 665 265
rect 597 215 607 249
rect 641 215 665 249
rect 597 199 665 215
rect 815 255 891 265
rect 815 221 831 255
rect 865 221 891 255
rect 815 211 891 221
rect 943 249 1037 265
rect 943 215 993 249
rect 1027 215 1037 249
rect 635 177 665 199
rect 833 131 863 211
rect 943 176 1037 215
rect 1099 249 1185 265
rect 1099 215 1109 249
rect 1143 215 1185 249
rect 1099 199 1185 215
rect 927 146 1037 176
rect 927 131 957 146
rect 1155 131 1185 199
rect 1227 249 1291 265
rect 1227 215 1237 249
rect 1271 215 1291 249
rect 1227 199 1291 215
rect 1344 259 1384 282
rect 1438 259 1478 282
rect 1344 249 1478 259
rect 1344 215 1360 249
rect 1394 215 1478 249
rect 1344 205 1478 215
rect 1227 131 1257 199
rect 1344 177 1374 205
rect 1438 177 1468 205
rect 89 21 119 47
rect 174 21 204 47
rect 269 21 299 47
rect 385 21 415 47
rect 516 21 546 47
rect 635 21 665 47
rect 833 21 863 47
rect 927 21 957 47
rect 1155 21 1185 47
rect 1227 21 1257 47
rect 1344 21 1374 47
rect 1438 21 1468 47
<< polycont >>
rect 32 215 66 249
rect 358 331 392 365
rect 494 331 528 365
rect 178 215 212 249
rect 293 157 327 191
rect 395 157 429 191
rect 607 215 641 249
rect 831 221 865 255
rect 993 215 1027 249
rect 1109 215 1143 249
rect 1237 215 1271 249
rect 1360 215 1394 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 17 485 69 527
rect 17 451 35 485
rect 17 417 69 451
rect 17 383 35 417
rect 17 367 69 383
rect 103 475 256 493
rect 103 441 222 475
rect 103 425 256 441
rect 322 475 460 493
rect 356 441 460 475
rect 322 425 460 441
rect 17 249 66 333
rect 17 215 32 249
rect 17 191 66 215
rect 103 157 144 425
rect 178 249 259 391
rect 212 215 259 249
rect 178 191 259 215
rect 293 365 392 391
rect 293 331 358 365
rect 293 323 392 331
rect 293 289 325 323
rect 359 289 392 323
rect 293 241 392 289
rect 426 275 460 425
rect 504 489 621 527
rect 504 455 560 489
rect 594 455 621 489
rect 504 415 621 455
rect 665 458 709 493
rect 665 424 675 458
rect 777 489 1151 527
rect 777 485 1101 489
rect 777 451 886 485
rect 920 455 1101 485
rect 1135 455 1151 489
rect 920 451 1151 455
rect 665 417 709 424
rect 1195 442 1229 493
rect 1279 489 1345 527
rect 1279 455 1295 489
rect 1329 455 1345 489
rect 1279 451 1345 455
rect 665 383 1151 417
rect 665 381 709 383
rect 494 365 709 381
rect 528 331 709 365
rect 494 327 709 331
rect 494 315 533 327
rect 426 249 641 275
rect 426 241 607 249
rect 293 191 360 241
rect 495 215 607 241
rect 327 157 360 191
rect 17 123 259 157
rect 293 141 360 157
rect 394 191 461 207
rect 394 157 395 191
rect 429 187 461 191
rect 394 153 427 157
rect 394 141 461 153
rect 495 199 641 215
rect 17 103 69 123
rect 17 69 35 103
rect 223 101 259 123
rect 495 107 529 199
rect 17 51 69 69
rect 103 55 129 89
rect 163 55 179 89
rect 103 17 179 55
rect 257 67 259 101
rect 223 51 259 67
rect 293 89 529 107
rect 293 55 329 89
rect 363 55 529 89
rect 293 51 529 55
rect 582 119 616 165
rect 582 17 616 85
rect 675 101 709 327
rect 675 51 709 67
rect 747 315 779 349
rect 813 315 829 349
rect 873 323 993 349
rect 747 187 781 315
rect 873 289 900 323
rect 934 315 993 323
rect 1027 315 1043 349
rect 934 299 1043 315
rect 873 255 934 289
rect 815 221 831 255
rect 865 221 934 255
rect 747 153 798 187
rect 876 157 934 221
rect 993 255 1037 265
rect 993 249 1002 255
rect 1036 221 1037 255
rect 1027 215 1037 221
rect 993 199 1037 215
rect 1081 249 1151 383
rect 1394 448 1444 493
rect 1229 408 1350 417
rect 1195 299 1350 408
rect 1081 215 1109 249
rect 1143 215 1151 249
rect 1081 199 1151 215
rect 1195 255 1281 265
rect 1195 221 1200 255
rect 1234 249 1281 255
rect 1234 221 1237 249
rect 1195 215 1237 221
rect 1271 215 1281 249
rect 1195 199 1281 215
rect 1316 263 1350 299
rect 1428 414 1444 448
rect 1394 380 1444 414
rect 1428 346 1444 380
rect 1488 485 1538 527
rect 1522 451 1538 485
rect 1488 417 1538 451
rect 1522 383 1538 417
rect 1488 365 1538 383
rect 1394 331 1444 346
rect 1394 297 1535 331
rect 1316 249 1454 263
rect 1316 215 1360 249
rect 1394 215 1454 249
rect 1316 211 1454 215
rect 1316 157 1350 211
rect 1498 177 1535 297
rect 747 110 813 153
rect 876 123 1017 157
rect 747 76 779 110
rect 967 110 1017 123
rect 747 51 813 76
rect 857 55 873 89
rect 907 55 923 89
rect 857 17 923 55
rect 1001 76 1017 110
rect 967 51 1017 76
rect 1101 123 1350 157
rect 1394 143 1535 177
rect 1101 109 1135 123
rect 1394 89 1434 143
rect 1101 51 1135 75
rect 1267 55 1284 89
rect 1318 55 1334 89
rect 1267 17 1334 55
rect 1368 55 1384 89
rect 1418 55 1434 89
rect 1368 51 1434 55
rect 1478 93 1512 109
rect 1478 17 1512 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 325 289 359 323
rect 427 157 429 187
rect 429 157 461 187
rect 427 153 461 157
rect 900 289 934 323
rect 798 153 832 187
rect 1002 249 1036 255
rect 1002 221 1027 249
rect 1027 221 1036 249
rect 1200 221 1234 255
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
<< metal1 >>
rect 0 561 1564 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 0 496 1564 527
rect 313 323 371 329
rect 313 289 325 323
rect 359 320 371 323
rect 888 323 946 329
rect 888 320 900 323
rect 359 292 900 320
rect 359 289 371 292
rect 313 283 371 289
rect 888 289 900 292
rect 934 289 946 323
rect 888 283 946 289
rect 990 255 1048 261
rect 990 221 1002 255
rect 1036 252 1048 255
rect 1188 255 1246 261
rect 1188 252 1200 255
rect 1036 224 1200 252
rect 1036 221 1048 224
rect 990 215 1048 221
rect 1188 221 1200 224
rect 1234 221 1246 255
rect 1188 215 1246 221
rect 415 187 473 193
rect 415 153 427 187
rect 461 184 473 187
rect 786 187 844 193
rect 786 184 798 187
rect 461 156 798 184
rect 461 153 473 156
rect 415 147 473 153
rect 786 153 798 156
rect 832 153 844 187
rect 786 147 844 153
rect 0 17 1564 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
rect 0 -48 1564 -17
<< labels >>
rlabel comment s 0 0 0 0 4 sdlclkp_2
flabel metal1 s 994 221 1028 255 0 FreeSans 200 0 0 0 CLK
port 1 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel corelocali s 1501 221 1535 255 0 FreeSans 200 0 0 0 GCLK
port 8 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 200 0 0 0 SCE
port 3 nsew
flabel corelocali s 214 289 248 323 0 FreeSans 200 0 0 0 GATE
port 2 nsew
flabel corelocali s 214 357 248 391 0 FreeSans 200 0 0 0 GATE
port 2 nsew
flabel corelocali s 1409 357 1443 391 0 FreeSans 200 0 0 0 GCLK
port 8 nsew
flabel corelocali s 1409 425 1443 459 0 FreeSans 200 0 0 0 GCLK
port 8 nsew
flabel corelocali s 30 289 64 323 0 FreeSans 200 0 0 0 SCE
port 3 nsew
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 1564 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 393366
string GDS_START 381334
<< end >>
