magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 17 191 69 333
rect 181 289 268 391
rect 181 191 259 289
rect 1426 331 1476 493
rect 1426 297 1564 331
rect 1530 263 1564 297
rect 1641 263 1719 493
rect 1530 211 1811 263
rect 1530 177 1564 211
rect 1426 143 1564 177
rect 1426 89 1476 143
rect 1400 51 1476 89
rect 1641 51 1719 211
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 17 367 69 527
rect 103 425 272 493
rect 306 425 481 493
rect 103 157 147 425
rect 302 323 403 391
rect 302 289 336 323
rect 370 289 403 323
rect 302 265 403 289
rect 293 241 403 265
rect 447 275 481 425
rect 515 415 653 527
rect 697 417 741 493
rect 779 451 1183 527
rect 1227 417 1261 493
rect 1311 451 1377 527
rect 697 383 1183 417
rect 697 381 741 383
rect 515 327 741 381
rect 515 315 559 327
rect 447 241 653 275
rect 17 123 259 157
rect 293 141 371 241
rect 405 187 472 207
rect 405 153 438 187
rect 405 141 472 153
rect 506 199 653 241
rect 17 51 69 123
rect 103 17 179 89
rect 223 51 259 123
rect 506 107 540 199
rect 293 51 540 107
rect 584 17 653 165
rect 697 51 741 327
rect 779 315 861 349
rect 905 323 1075 349
rect 779 187 813 315
rect 905 289 932 323
rect 966 299 1075 323
rect 905 255 966 289
rect 847 221 966 255
rect 779 153 830 187
rect 908 157 966 221
rect 1011 255 1069 265
rect 1011 221 1023 255
rect 1057 221 1069 255
rect 1011 199 1069 221
rect 1113 199 1183 383
rect 1227 299 1382 417
rect 1227 255 1313 265
rect 1227 221 1232 255
rect 1266 221 1313 255
rect 1227 199 1313 221
rect 1348 263 1382 299
rect 1520 365 1570 527
rect 1753 297 1807 527
rect 1348 211 1486 263
rect 1348 157 1382 211
rect 779 51 845 153
rect 908 123 1049 157
rect 879 17 955 89
rect 999 51 1049 123
rect 1083 123 1382 157
rect 1083 51 1167 123
rect 1201 17 1366 89
rect 1520 17 1570 109
rect 1753 17 1807 177
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 336 289 370 323
rect 438 153 472 187
rect 932 289 966 323
rect 830 153 864 187
rect 1023 221 1057 255
rect 1232 221 1266 255
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
<< metal1 >>
rect 0 561 1840 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 0 496 1840 527
rect 1011 255 1069 261
rect 1011 221 1023 255
rect 1057 252 1069 255
rect 1220 255 1278 261
rect 1220 252 1232 255
rect 1057 224 1232 252
rect 1057 221 1069 224
rect 1011 215 1069 221
rect 1220 221 1232 224
rect 1266 221 1278 255
rect 1220 215 1278 221
rect 0 17 1840 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
rect 0 -48 1840 -17
<< obsm1 >>
rect 324 323 382 329
rect 324 289 336 323
rect 370 320 382 323
rect 920 323 978 329
rect 920 320 932 323
rect 370 292 932 320
rect 370 289 382 292
rect 324 283 382 289
rect 920 289 932 292
rect 966 289 978 323
rect 920 283 978 289
rect 426 187 484 193
rect 426 153 438 187
rect 472 184 484 187
rect 818 187 876 193
rect 818 184 830 187
rect 472 156 830 184
rect 472 153 484 156
rect 426 147 484 153
rect 818 153 830 156
rect 864 153 876 187
rect 818 147 876 153
<< labels >>
rlabel metal1 s 1220 252 1278 261 6 CLK
port 1 nsew signal input
rlabel metal1 s 1220 215 1278 224 6 CLK
port 1 nsew signal input
rlabel metal1 s 1011 252 1069 261 6 CLK
port 1 nsew signal input
rlabel metal1 s 1011 224 1278 252 6 CLK
port 1 nsew signal input
rlabel metal1 s 1011 215 1069 224 6 CLK
port 1 nsew signal input
rlabel locali s 181 289 268 391 6 GATE
port 2 nsew signal input
rlabel locali s 181 191 259 289 6 GATE
port 2 nsew signal input
rlabel locali s 1641 263 1719 493 6 GCLK
port 3 nsew signal output
rlabel locali s 1641 51 1719 211 6 GCLK
port 3 nsew signal output
rlabel locali s 1530 263 1564 297 6 GCLK
port 3 nsew signal output
rlabel locali s 1530 211 1811 263 6 GCLK
port 3 nsew signal output
rlabel locali s 1530 177 1564 211 6 GCLK
port 3 nsew signal output
rlabel locali s 1426 331 1476 493 6 GCLK
port 3 nsew signal output
rlabel locali s 1426 297 1564 331 6 GCLK
port 3 nsew signal output
rlabel locali s 1426 143 1564 177 6 GCLK
port 3 nsew signal output
rlabel locali s 1426 89 1476 143 6 GCLK
port 3 nsew signal output
rlabel locali s 1400 51 1476 89 6 GCLK
port 3 nsew signal output
rlabel locali s 17 191 69 333 6 SCE
port 4 nsew signal input
rlabel metal1 s 0 -48 1840 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 1840 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1840 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 407202
string GDS_START 393426
<< end >>
