magic
tech sky130A
magscale 1 2
timestamp 1604502693
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 79 47 109 177
rect 176 47 206 177
rect 366 47 396 177
rect 460 47 490 177
rect 659 47 689 177
rect 743 47 773 177
rect 827 47 857 177
rect 911 47 941 177
rect 995 47 1025 177
<< pmoshvt >>
rect 79 297 109 497
rect 174 297 204 497
rect 366 297 396 497
rect 460 297 490 497
rect 659 297 689 497
rect 743 297 773 497
rect 827 297 857 497
rect 911 297 941 497
rect 995 297 1025 497
<< ndiff >>
rect 27 109 79 177
rect 27 75 35 109
rect 69 75 79 109
rect 27 47 79 75
rect 109 93 176 177
rect 109 59 119 93
rect 153 59 176 93
rect 109 47 176 59
rect 206 47 366 177
rect 396 93 460 177
rect 396 59 411 93
rect 445 59 460 93
rect 396 47 460 59
rect 490 47 659 177
rect 689 93 743 177
rect 689 59 699 93
rect 733 59 743 93
rect 689 47 743 59
rect 773 101 827 177
rect 773 67 783 101
rect 817 67 827 101
rect 773 47 827 67
rect 857 93 911 177
rect 857 59 867 93
rect 901 59 911 93
rect 857 47 911 59
rect 941 101 995 177
rect 941 67 951 101
rect 985 67 995 101
rect 941 47 995 67
rect 1025 93 1077 177
rect 1025 59 1035 93
rect 1069 59 1077 93
rect 1025 47 1077 59
<< pdiff >>
rect 27 477 79 497
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 297 79 375
rect 109 485 174 497
rect 109 451 119 485
rect 153 451 174 485
rect 109 417 174 451
rect 109 383 119 417
rect 153 383 174 417
rect 109 297 174 383
rect 204 489 260 497
rect 204 455 214 489
rect 248 455 260 489
rect 204 421 260 455
rect 204 387 218 421
rect 252 387 260 421
rect 204 297 260 387
rect 314 421 366 497
rect 314 387 322 421
rect 356 387 366 421
rect 314 297 366 387
rect 396 353 460 497
rect 396 319 412 353
rect 446 319 460 353
rect 396 297 460 319
rect 490 489 550 497
rect 490 455 504 489
rect 538 455 550 489
rect 490 297 550 455
rect 607 477 659 497
rect 607 443 615 477
rect 649 443 659 477
rect 607 297 659 443
rect 689 485 743 497
rect 689 451 699 485
rect 733 451 743 485
rect 689 297 743 451
rect 773 477 827 497
rect 773 443 783 477
rect 817 443 827 477
rect 773 409 827 443
rect 773 375 783 409
rect 817 375 827 409
rect 773 297 827 375
rect 857 485 911 497
rect 857 451 867 485
rect 901 451 911 485
rect 857 417 911 451
rect 857 383 867 417
rect 901 383 911 417
rect 857 297 911 383
rect 941 477 995 497
rect 941 443 951 477
rect 985 443 995 477
rect 941 409 995 443
rect 941 375 951 409
rect 985 375 995 409
rect 941 297 995 375
rect 1025 485 1077 497
rect 1025 451 1035 485
rect 1069 451 1077 485
rect 1025 417 1077 451
rect 1025 383 1035 417
rect 1069 383 1077 417
rect 1025 297 1077 383
<< ndiffc >>
rect 35 75 69 109
rect 119 59 153 93
rect 411 59 445 93
rect 699 59 733 93
rect 783 67 817 101
rect 867 59 901 93
rect 951 67 985 101
rect 1035 59 1069 93
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 451 153 485
rect 119 383 153 417
rect 214 455 248 489
rect 218 387 252 421
rect 322 387 356 421
rect 412 319 446 353
rect 504 455 538 489
rect 615 443 649 477
rect 699 451 733 485
rect 783 443 817 477
rect 783 375 817 409
rect 867 451 901 485
rect 867 383 901 417
rect 951 443 985 477
rect 951 375 985 409
rect 1035 451 1069 485
rect 1035 383 1069 417
<< poly >>
rect 79 497 109 523
rect 174 497 204 523
rect 366 497 396 523
rect 460 497 490 523
rect 659 497 689 523
rect 743 497 773 523
rect 827 497 857 523
rect 911 497 941 523
rect 995 497 1025 523
rect 79 265 109 297
rect 174 265 204 297
rect 366 265 396 297
rect 460 265 490 297
rect 659 265 689 297
rect 76 249 130 265
rect 76 215 86 249
rect 120 215 130 249
rect 76 199 130 215
rect 172 249 226 265
rect 172 215 182 249
rect 216 215 226 249
rect 172 199 226 215
rect 306 249 396 265
rect 306 215 316 249
rect 350 215 396 249
rect 306 199 396 215
rect 443 249 497 265
rect 443 215 453 249
rect 487 215 497 249
rect 443 199 497 215
rect 567 249 689 265
rect 743 265 773 297
rect 827 265 857 297
rect 911 265 941 297
rect 995 265 1025 297
rect 743 259 1025 265
rect 567 215 577 249
rect 611 215 645 249
rect 679 215 689 249
rect 567 199 689 215
rect 736 249 1025 259
rect 736 215 752 249
rect 786 215 820 249
rect 854 215 888 249
rect 922 215 956 249
rect 990 215 1025 249
rect 736 205 1025 215
rect 79 177 109 199
rect 176 177 206 199
rect 366 177 396 199
rect 460 177 490 199
rect 659 177 689 199
rect 743 199 1025 205
rect 743 177 773 199
rect 827 177 857 199
rect 911 177 941 199
rect 995 177 1025 199
rect 79 21 109 47
rect 176 21 206 47
rect 366 21 396 47
rect 460 21 490 47
rect 659 21 689 47
rect 743 21 773 47
rect 827 21 857 47
rect 911 21 941 47
rect 995 21 1025 47
<< polycont >>
rect 86 215 120 249
rect 182 215 216 249
rect 316 215 350 249
rect 453 215 487 249
rect 577 215 611 249
rect 645 215 679 249
rect 752 215 786 249
rect 820 215 854 249
rect 888 215 922 249
rect 956 215 990 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 18 477 69 493
rect 18 443 35 477
rect 18 409 69 443
rect 18 375 35 409
rect 18 333 69 375
rect 103 485 164 527
rect 103 451 119 485
rect 153 451 164 485
rect 103 417 164 451
rect 103 383 119 417
rect 153 383 164 417
rect 198 455 214 489
rect 248 455 504 489
rect 538 455 554 489
rect 615 477 649 493
rect 198 421 268 455
rect 683 485 749 527
rect 683 451 699 485
rect 733 451 749 485
rect 783 477 817 493
rect 615 421 649 443
rect 198 387 218 421
rect 252 387 268 421
rect 306 387 322 421
rect 356 387 649 421
rect 783 409 817 443
rect 103 367 164 383
rect 851 485 917 527
rect 851 451 867 485
rect 901 451 917 485
rect 851 417 917 451
rect 851 383 867 417
rect 901 383 917 417
rect 951 477 985 493
rect 951 409 985 443
rect 713 353 747 357
rect 18 299 216 333
rect 18 125 52 299
rect 86 249 148 265
rect 120 215 148 249
rect 86 199 148 215
rect 182 249 216 299
rect 182 199 216 215
rect 296 249 350 323
rect 396 319 412 353
rect 446 319 747 353
rect 296 215 316 249
rect 296 199 350 215
rect 393 249 487 265
rect 393 215 453 249
rect 393 199 487 215
rect 536 249 679 265
rect 536 215 577 249
rect 611 215 645 249
rect 536 199 679 215
rect 713 249 747 319
rect 783 349 817 375
rect 1019 485 1085 527
rect 1019 451 1035 485
rect 1069 451 1085 485
rect 1019 417 1085 451
rect 1019 383 1035 417
rect 1069 383 1085 417
rect 951 349 985 375
rect 783 315 1086 349
rect 713 215 752 249
rect 786 215 820 249
rect 854 215 888 249
rect 922 215 956 249
rect 990 215 1006 249
rect 114 161 148 199
rect 536 161 570 199
rect 713 165 747 215
rect 114 127 570 161
rect 612 131 747 165
rect 1040 161 1086 315
rect 18 109 69 125
rect 18 75 35 109
rect 612 93 646 131
rect 783 127 1086 161
rect 783 101 817 127
rect 18 59 69 75
rect 103 59 119 93
rect 153 59 169 93
rect 395 59 411 93
rect 445 59 646 93
rect 683 59 699 93
rect 733 59 749 93
rect 103 17 169 59
rect 683 17 749 59
rect 951 101 985 127
rect 783 51 817 67
rect 851 59 867 93
rect 901 59 917 93
rect 851 17 917 59
rect 951 51 985 67
rect 1019 59 1035 93
rect 1069 59 1085 93
rect 1019 17 1085 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
flabel corelocali s 1040 153 1074 187 0 FreeSans 200 0 0 0 X
port 8 nsew
flabel corelocali s 1040 221 1074 255 0 FreeSans 200 0 0 0 X
port 8 nsew
flabel corelocali s 1040 289 1074 323 0 FreeSans 200 0 0 0 X
port 8 nsew
flabel corelocali s 580 221 614 255 0 FreeSans 200 0 0 0 S
port 3 nsew
flabel corelocali s 304 221 338 255 0 FreeSans 200 0 0 0 A0
port 1 nsew
flabel corelocali s 396 221 430 255 0 FreeSans 200 0 0 0 A1
port 2 nsew
flabel corelocali s 304 289 338 323 0 FreeSans 200 0 0 0 A0
port 1 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
rlabel comment s 0 0 0 0 4 mux2_4
<< properties >>
string FIXED_BBOX 0 0 1104 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1659120
string GDS_START 1650786
string path 0.000 0.000 27.600 0.000 
<< end >>
