magic
tech sky130A
magscale 1 2
timestamp 1604502697
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 360 -17 404 17
<< scnmos >>
rect 87 47 117 151
rect 171 47 201 151
rect 275 47 305 151
rect 359 47 389 151
rect 495 47 525 131
rect 593 47 623 131
rect 724 47 754 131
rect 925 47 955 131
rect 1049 47 1079 151
<< pmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 487 309 523 497
rect 602 309 638 497
rect 839 309 875 497
rect 927 309 963 497
rect 1041 309 1077 497
<< ndiff >>
rect 35 115 87 151
rect 35 81 43 115
rect 77 81 87 115
rect 35 47 87 81
rect 117 115 171 151
rect 117 81 127 115
rect 161 81 171 115
rect 117 47 171 81
rect 201 115 275 151
rect 201 81 219 115
rect 253 81 275 115
rect 201 47 275 81
rect 305 112 359 151
rect 305 78 315 112
rect 349 78 359 112
rect 305 47 359 78
rect 389 131 447 151
rect 999 131 1049 151
rect 389 93 495 131
rect 389 59 405 93
rect 439 59 495 93
rect 389 47 495 59
rect 525 47 593 131
rect 623 108 724 131
rect 623 74 666 108
rect 700 74 724 108
rect 623 47 724 74
rect 754 47 925 131
rect 955 89 1049 131
rect 955 55 985 89
rect 1019 55 1049 89
rect 955 47 1049 55
rect 1079 108 1131 151
rect 1079 74 1089 108
rect 1123 74 1131 108
rect 1079 47 1131 74
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 485 175 497
rect 117 451 129 485
rect 163 451 175 485
rect 117 417 175 451
rect 117 383 129 417
rect 163 383 175 417
rect 117 349 175 383
rect 117 315 129 349
rect 163 315 175 349
rect 117 297 175 315
rect 211 485 269 497
rect 211 451 223 485
rect 257 451 269 485
rect 211 417 269 451
rect 211 383 223 417
rect 257 383 269 417
rect 211 349 269 383
rect 211 315 223 349
rect 257 315 269 349
rect 211 297 269 315
rect 305 485 363 497
rect 305 451 317 485
rect 351 451 363 485
rect 305 417 363 451
rect 305 383 317 417
rect 351 383 363 417
rect 305 349 363 383
rect 305 315 317 349
rect 351 315 363 349
rect 305 297 363 315
rect 399 485 487 497
rect 399 451 411 485
rect 445 451 487 485
rect 399 417 487 451
rect 399 383 411 417
rect 445 383 487 417
rect 399 349 487 383
rect 399 315 411 349
rect 445 315 487 349
rect 399 309 487 315
rect 523 309 602 497
rect 638 425 839 497
rect 638 391 650 425
rect 684 391 725 425
rect 759 391 793 425
rect 827 391 839 425
rect 638 309 839 391
rect 875 309 927 497
rect 963 485 1041 497
rect 963 451 993 485
rect 1027 451 1041 485
rect 963 417 1041 451
rect 963 383 993 417
rect 1027 383 1041 417
rect 963 309 1041 383
rect 1077 485 1135 497
rect 1077 451 1089 485
rect 1123 451 1135 485
rect 1077 417 1135 451
rect 1077 383 1089 417
rect 1123 383 1135 417
rect 1077 309 1135 383
rect 399 297 461 309
<< ndiffc >>
rect 43 81 77 115
rect 127 81 161 115
rect 219 81 253 115
rect 315 78 349 112
rect 405 59 439 93
rect 666 74 700 108
rect 985 55 1019 89
rect 1089 74 1123 108
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 451 163 485
rect 129 383 163 417
rect 129 315 163 349
rect 223 451 257 485
rect 223 383 257 417
rect 223 315 257 349
rect 317 451 351 485
rect 317 383 351 417
rect 317 315 351 349
rect 411 451 445 485
rect 411 383 445 417
rect 411 315 445 349
rect 650 391 684 425
rect 725 391 759 425
rect 793 391 827 425
rect 993 451 1027 485
rect 993 383 1027 417
rect 1089 451 1123 485
rect 1089 383 1123 417
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 487 497 523 523
rect 602 497 638 523
rect 839 497 875 523
rect 927 497 963 523
rect 1041 497 1077 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 487 294 523 309
rect 602 294 638 309
rect 839 294 875 309
rect 927 294 963 309
rect 1041 294 1077 309
rect 79 265 119 282
rect 173 265 213 282
rect 267 265 307 282
rect 361 265 401 282
rect 485 265 525 294
rect 79 249 427 265
rect 79 215 383 249
rect 417 215 427 249
rect 79 199 427 215
rect 469 249 525 265
rect 600 264 764 294
rect 837 277 877 294
rect 469 215 479 249
rect 513 215 525 249
rect 724 229 764 264
rect 823 261 877 277
rect 469 199 525 215
rect 87 151 117 199
rect 171 151 201 199
rect 275 151 305 199
rect 359 151 389 199
rect 495 131 525 199
rect 593 212 682 222
rect 593 178 632 212
rect 666 178 682 212
rect 593 168 682 178
rect 724 213 778 229
rect 724 179 734 213
rect 768 179 778 213
rect 823 227 833 261
rect 867 227 877 261
rect 823 211 877 227
rect 925 237 965 294
rect 1039 277 1079 294
rect 1027 261 1081 277
rect 925 221 985 237
rect 593 131 623 168
rect 724 163 778 179
rect 925 187 941 221
rect 975 187 985 221
rect 1027 227 1037 261
rect 1071 227 1081 261
rect 1027 211 1081 227
rect 925 171 985 187
rect 724 131 754 163
rect 925 131 955 171
rect 1049 151 1079 211
rect 87 21 117 47
rect 171 21 201 47
rect 275 21 305 47
rect 359 21 389 47
rect 495 21 525 47
rect 593 21 623 47
rect 724 21 754 47
rect 925 21 955 47
rect 1049 21 1079 47
<< polycont >>
rect 383 215 417 249
rect 479 215 513 249
rect 632 178 666 212
rect 734 179 768 213
rect 833 227 867 261
rect 941 187 975 221
rect 1037 227 1071 261
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 27 485 79 527
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 299 79 315
rect 113 485 179 493
rect 113 451 129 485
rect 163 451 179 485
rect 113 417 179 451
rect 113 383 129 417
rect 163 383 179 417
rect 113 349 179 383
rect 113 315 129 349
rect 163 315 179 349
rect 113 299 179 315
rect 213 485 261 527
rect 213 451 223 485
rect 257 451 261 485
rect 213 417 261 451
rect 213 383 223 417
rect 257 383 261 417
rect 213 349 261 383
rect 213 315 223 349
rect 257 315 261 349
rect 213 299 261 315
rect 295 485 367 493
rect 295 451 317 485
rect 351 451 367 485
rect 295 417 367 451
rect 295 383 317 417
rect 351 383 367 417
rect 295 349 367 383
rect 295 315 317 349
rect 351 315 367 349
rect 295 299 367 315
rect 401 485 456 527
rect 401 451 411 485
rect 445 451 456 485
rect 401 417 456 451
rect 401 383 411 417
rect 445 383 456 417
rect 401 349 456 383
rect 401 315 411 349
rect 445 315 456 349
rect 401 299 456 315
rect 490 459 959 493
rect 118 265 170 299
rect 295 265 349 299
rect 490 265 530 459
rect 118 213 349 265
rect 35 115 84 131
rect 35 81 43 115
rect 77 81 84 115
rect 35 17 84 81
rect 118 115 170 213
rect 118 81 127 115
rect 161 81 170 115
rect 118 51 170 81
rect 211 115 261 131
rect 211 81 219 115
rect 253 81 261 115
rect 211 17 261 81
rect 295 112 349 213
rect 383 249 417 265
rect 383 165 417 215
rect 475 249 530 265
rect 475 215 479 249
rect 513 215 530 249
rect 475 199 530 215
rect 564 391 650 425
rect 684 391 725 425
rect 759 391 793 425
rect 827 391 853 425
rect 564 165 598 391
rect 383 131 598 165
rect 632 323 891 357
rect 632 212 666 323
rect 632 162 666 178
rect 734 213 799 283
rect 768 179 799 213
rect 295 78 315 112
rect 563 124 598 131
rect 563 108 700 124
rect 295 51 349 78
rect 383 93 455 97
rect 383 59 405 93
rect 439 59 455 93
rect 383 17 455 59
rect 563 74 666 108
rect 563 51 700 74
rect 734 51 799 179
rect 833 261 891 323
rect 925 326 959 459
rect 993 485 1039 527
rect 1027 451 1039 485
rect 993 417 1039 451
rect 1027 383 1039 417
rect 993 367 1039 383
rect 1073 485 1153 493
rect 1073 451 1089 485
rect 1123 451 1153 485
rect 1073 417 1153 451
rect 1073 383 1089 417
rect 1123 383 1153 417
rect 1073 367 1153 383
rect 925 288 1075 326
rect 867 227 891 261
rect 1037 261 1075 288
rect 833 51 891 227
rect 941 221 975 237
rect 1071 227 1075 261
rect 1037 211 1075 227
rect 941 173 975 187
rect 1119 173 1153 367
rect 941 139 1153 173
rect 1083 108 1132 139
rect 926 89 1029 105
rect 926 55 985 89
rect 1019 55 1029 89
rect 926 17 1029 55
rect 1083 74 1089 108
rect 1123 74 1132 108
rect 1083 51 1132 74
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
flabel metal1 s 306 -17 340 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 306 527 340 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
flabel corelocali s 948 289 982 323 0 FreeSans 250 0 0 0 S
port 3 nsew
flabel corelocali s 857 153 891 187 0 FreeSans 250 0 0 0 A1
port 2 nsew
flabel corelocali s 857 221 891 255 0 FreeSans 250 0 0 0 A1
port 2 nsew
flabel corelocali s 765 221 799 255 0 FreeSans 250 0 0 0 A0
port 1 nsew
flabel corelocali s 305 85 339 119 0 FreeSans 250 0 0 0 X
port 8 nsew
flabel corelocali s 305 357 339 391 0 FreeSans 250 0 0 0 X
port 8 nsew
flabel corelocali s 305 425 339 459 0 FreeSans 250 0 0 0 X
port 8 nsew
flabel corelocali s 1037 289 1071 323 0 FreeSans 250 0 0 0 S
port 3 nsew
flabel nbase s 350 527 384 561 0 FreeSans 250 0 0 0 VPB
port 6 nsew
flabel pwell s 360 -17 404 17 0 FreeSans 250 0 0 0 VNB
port 5 nsew
rlabel comment s 0 0 0 0 4 clkmux2_2
<< properties >>
string FIXED_BBOX 0 0 1196 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3293112
string GDS_START 3284120
<< end >>
