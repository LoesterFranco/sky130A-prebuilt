magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 1326 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 113 47 143 177
rect 197 47 227 177
rect 291 47 321 177
rect 385 47 415 177
rect 489 47 519 177
rect 687 47 717 177
rect 781 47 811 177
rect 875 47 905 177
rect 979 47 1009 177
rect 1063 47 1093 177
rect 1167 47 1197 177
<< pmoshvt >>
rect 105 297 141 497
rect 199 297 235 497
rect 293 297 329 497
rect 387 297 423 497
rect 481 297 517 497
rect 575 297 611 497
rect 669 297 705 497
rect 877 297 913 497
rect 971 297 1007 497
rect 1065 297 1101 497
rect 1159 297 1195 497
<< ndiff >>
rect 42 163 113 177
rect 42 129 59 163
rect 93 129 113 163
rect 42 95 113 129
rect 42 61 59 95
rect 93 61 113 95
rect 42 47 113 61
rect 143 163 197 177
rect 143 129 153 163
rect 187 129 197 163
rect 143 95 197 129
rect 143 61 153 95
rect 187 61 197 95
rect 143 47 197 61
rect 227 163 291 177
rect 227 129 247 163
rect 281 129 291 163
rect 227 95 291 129
rect 227 61 247 95
rect 281 61 291 95
rect 227 47 291 61
rect 321 95 385 177
rect 321 61 341 95
rect 375 61 385 95
rect 321 47 385 61
rect 415 163 489 177
rect 415 129 435 163
rect 469 129 489 163
rect 415 95 489 129
rect 415 61 425 95
rect 459 61 489 95
rect 415 47 489 61
rect 519 95 571 177
rect 519 61 529 95
rect 563 61 571 95
rect 519 47 571 61
rect 635 95 687 177
rect 635 61 643 95
rect 677 61 687 95
rect 635 47 687 61
rect 717 163 781 177
rect 717 129 737 163
rect 771 129 781 163
rect 717 47 781 129
rect 811 163 875 177
rect 811 129 831 163
rect 865 129 875 163
rect 811 95 875 129
rect 811 61 831 95
rect 865 61 875 95
rect 811 47 875 61
rect 905 95 979 177
rect 905 61 925 95
rect 959 61 979 95
rect 905 47 979 61
rect 1009 163 1063 177
rect 1009 129 1019 163
rect 1053 129 1063 163
rect 1009 95 1063 129
rect 1009 61 1019 95
rect 1053 61 1063 95
rect 1009 47 1063 61
rect 1093 95 1167 177
rect 1093 61 1113 95
rect 1147 61 1167 95
rect 1093 47 1167 61
rect 1197 163 1253 177
rect 1197 129 1207 163
rect 1241 129 1253 163
rect 1197 95 1253 129
rect 1197 61 1207 95
rect 1241 61 1253 95
rect 1197 47 1253 61
<< pdiff >>
rect 27 477 105 497
rect 27 443 53 477
rect 87 443 105 477
rect 27 409 105 443
rect 27 375 53 409
rect 87 375 105 409
rect 27 341 105 375
rect 27 307 53 341
rect 87 307 105 341
rect 27 297 105 307
rect 141 477 199 497
rect 141 443 153 477
rect 187 443 199 477
rect 141 297 199 443
rect 235 341 293 497
rect 235 307 247 341
rect 281 307 293 341
rect 235 297 293 307
rect 329 477 387 497
rect 329 443 341 477
rect 375 443 387 477
rect 329 297 387 443
rect 423 341 481 497
rect 423 307 435 341
rect 469 307 481 341
rect 423 297 481 307
rect 517 477 575 497
rect 517 443 529 477
rect 563 443 575 477
rect 517 297 575 443
rect 611 477 669 497
rect 611 443 623 477
rect 657 443 669 477
rect 611 409 669 443
rect 611 375 623 409
rect 657 375 669 409
rect 611 297 669 375
rect 705 477 759 497
rect 705 443 717 477
rect 751 443 759 477
rect 705 297 759 443
rect 823 477 877 497
rect 823 443 831 477
rect 865 443 877 477
rect 823 297 877 443
rect 913 409 971 497
rect 913 375 925 409
rect 959 375 971 409
rect 913 341 971 375
rect 913 307 925 341
rect 959 307 971 341
rect 913 297 971 307
rect 1007 477 1065 497
rect 1007 443 1019 477
rect 1053 443 1065 477
rect 1007 409 1065 443
rect 1007 375 1019 409
rect 1053 375 1065 409
rect 1007 341 1065 375
rect 1007 307 1019 341
rect 1053 307 1065 341
rect 1007 297 1065 307
rect 1101 485 1159 497
rect 1101 451 1113 485
rect 1147 451 1159 485
rect 1101 417 1159 451
rect 1101 383 1113 417
rect 1147 383 1159 417
rect 1101 297 1159 383
rect 1195 477 1253 497
rect 1195 443 1207 477
rect 1241 443 1253 477
rect 1195 409 1253 443
rect 1195 375 1207 409
rect 1241 375 1253 409
rect 1195 341 1253 375
rect 1195 307 1207 341
rect 1241 307 1253 341
rect 1195 297 1253 307
<< ndiffc >>
rect 59 129 93 163
rect 59 61 93 95
rect 153 129 187 163
rect 153 61 187 95
rect 247 129 281 163
rect 247 61 281 95
rect 341 61 375 95
rect 435 129 469 163
rect 425 61 459 95
rect 529 61 563 95
rect 643 61 677 95
rect 737 129 771 163
rect 831 129 865 163
rect 831 61 865 95
rect 925 61 959 95
rect 1019 129 1053 163
rect 1019 61 1053 95
rect 1113 61 1147 95
rect 1207 129 1241 163
rect 1207 61 1241 95
<< pdiffc >>
rect 53 443 87 477
rect 53 375 87 409
rect 53 307 87 341
rect 153 443 187 477
rect 247 307 281 341
rect 341 443 375 477
rect 435 307 469 341
rect 529 443 563 477
rect 623 443 657 477
rect 623 375 657 409
rect 717 443 751 477
rect 831 443 865 477
rect 925 375 959 409
rect 925 307 959 341
rect 1019 443 1053 477
rect 1019 375 1053 409
rect 1019 307 1053 341
rect 1113 451 1147 485
rect 1113 383 1147 417
rect 1207 443 1241 477
rect 1207 375 1241 409
rect 1207 307 1241 341
<< poly >>
rect 105 497 141 523
rect 199 497 235 523
rect 293 497 329 523
rect 387 497 423 523
rect 481 497 517 523
rect 575 497 611 523
rect 669 497 705 523
rect 877 497 913 523
rect 971 497 1007 523
rect 1065 497 1101 523
rect 1159 497 1195 523
rect 105 282 141 297
rect 199 282 235 297
rect 293 282 329 297
rect 387 282 423 297
rect 481 282 517 297
rect 575 282 611 297
rect 669 282 705 297
rect 877 282 913 297
rect 971 282 1007 297
rect 1065 282 1101 297
rect 1159 282 1195 297
rect 103 265 143 282
rect 197 265 237 282
rect 291 265 331 282
rect 385 265 425 282
rect 479 265 519 282
rect 91 249 155 265
rect 91 215 101 249
rect 135 215 155 249
rect 91 199 155 215
rect 197 250 519 265
rect 197 216 391 250
rect 425 216 469 250
rect 503 216 519 250
rect 197 199 519 216
rect 573 265 613 282
rect 667 265 707 282
rect 875 265 915 282
rect 969 265 1009 282
rect 573 249 811 265
rect 573 215 637 249
rect 671 215 811 249
rect 573 199 811 215
rect 113 177 143 199
rect 197 177 227 199
rect 291 177 321 199
rect 385 177 415 199
rect 489 177 519 199
rect 687 177 717 199
rect 781 177 811 199
rect 875 249 1009 265
rect 875 215 925 249
rect 959 215 1009 249
rect 875 199 1009 215
rect 875 177 905 199
rect 979 177 1009 199
rect 1063 265 1103 282
rect 1157 265 1197 282
rect 1063 249 1197 265
rect 1063 215 1124 249
rect 1158 215 1197 249
rect 1063 199 1197 215
rect 1063 177 1093 199
rect 1167 177 1197 199
rect 113 21 143 47
rect 197 21 227 47
rect 291 21 321 47
rect 385 21 415 47
rect 489 21 519 47
rect 687 21 717 47
rect 781 21 811 47
rect 875 21 905 47
rect 979 21 1009 47
rect 1063 21 1093 47
rect 1167 21 1197 47
<< polycont >>
rect 101 215 135 249
rect 391 216 425 250
rect 469 216 503 250
rect 637 215 671 249
rect 925 215 959 249
rect 1124 215 1158 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 17 477 87 493
rect 17 443 53 477
rect 127 477 203 527
rect 127 443 153 477
rect 187 443 203 477
rect 315 477 391 527
rect 315 443 341 477
rect 375 443 391 477
rect 503 477 579 527
rect 503 443 529 477
rect 563 443 579 477
rect 623 477 657 493
rect 17 409 87 443
rect 623 409 657 443
rect 710 477 760 527
rect 710 443 717 477
rect 751 443 760 477
rect 710 427 760 443
rect 807 477 1053 493
rect 807 443 831 477
rect 865 459 1019 477
rect 807 427 865 443
rect 17 375 53 409
rect 87 375 563 409
rect 17 341 87 375
rect 17 307 53 341
rect 17 291 87 307
rect 17 171 51 291
rect 121 257 187 341
rect 85 249 187 257
rect 85 215 101 249
rect 135 215 187 249
rect 231 307 247 341
rect 281 307 435 341
rect 469 307 485 341
rect 231 289 485 307
rect 529 323 563 375
rect 917 409 966 425
rect 917 393 925 409
rect 657 375 925 393
rect 959 375 966 409
rect 623 359 966 375
rect 529 289 641 323
rect 231 182 341 289
rect 375 216 391 250
rect 425 216 469 250
rect 503 216 563 250
rect 17 163 109 171
rect 17 129 59 163
rect 93 129 109 163
rect 17 95 109 129
rect 17 61 59 95
rect 93 61 109 95
rect 17 53 109 61
rect 153 163 187 181
rect 153 95 187 129
rect 153 17 187 61
rect 231 163 475 182
rect 231 129 247 163
rect 281 145 435 163
rect 281 129 297 145
rect 231 95 297 129
rect 409 129 435 145
rect 469 129 475 163
rect 529 179 563 216
rect 597 249 641 289
rect 597 215 637 249
rect 671 215 687 249
rect 749 179 787 359
rect 917 341 966 359
rect 917 307 925 341
rect 959 307 966 341
rect 917 289 966 307
rect 1019 409 1053 443
rect 1019 341 1053 375
rect 1087 485 1163 527
rect 1087 451 1113 485
rect 1147 451 1163 485
rect 1087 417 1163 451
rect 1087 383 1113 417
rect 1147 383 1163 417
rect 1087 367 1163 383
rect 1207 477 1262 493
rect 1241 443 1262 477
rect 1207 409 1262 443
rect 1241 375 1262 409
rect 1207 341 1262 375
rect 1053 307 1207 333
rect 1241 307 1262 341
rect 1019 291 1262 307
rect 836 249 1064 255
rect 836 215 925 249
rect 959 215 1064 249
rect 1108 249 1271 255
rect 1108 215 1124 249
rect 1158 215 1271 249
rect 529 163 787 179
rect 529 129 737 163
rect 771 129 787 163
rect 831 163 1262 181
rect 865 145 1019 163
rect 865 129 881 145
rect 231 61 247 95
rect 281 61 297 95
rect 231 51 297 61
rect 341 95 375 111
rect 341 17 375 61
rect 409 95 475 129
rect 831 95 881 129
rect 993 129 1019 145
rect 1053 145 1207 163
rect 1053 129 1069 145
rect 409 61 425 95
rect 459 61 475 95
rect 409 51 475 61
rect 513 61 529 95
rect 563 61 579 95
rect 513 17 579 61
rect 621 61 643 95
rect 677 61 831 95
rect 865 61 881 95
rect 621 51 881 61
rect 925 95 959 111
rect 925 17 959 61
rect 993 95 1069 129
rect 1181 129 1207 145
rect 1241 129 1262 163
rect 993 61 1019 95
rect 1053 61 1069 95
rect 993 51 1069 61
rect 1113 95 1147 111
rect 1113 17 1147 61
rect 1181 95 1262 129
rect 1181 61 1207 95
rect 1241 61 1262 95
rect 1181 53 1262 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
flabel corelocali s 121 221 155 255 0 FreeSans 400 180 0 0 B1_N
port 3 nsew
flabel corelocali s 1151 221 1185 255 0 FreeSans 400 180 0 0 A1
port 1 nsew
flabel corelocali s 874 238 874 238 0 FreeSans 400 180 0 0 A2
port 2 nsew
flabel corelocali s 420 85 454 119 0 FreeSans 400 180 0 0 X
port 8 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
rlabel comment s 0 0 0 0 4 o21ba_4
<< properties >>
string FIXED_BBOX 0 0 1288 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1070004
string GDS_START 1060508
<< end >>
