magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1196 561
rect 144 455 210 527
rect 316 455 382 527
rect 487 455 554 527
rect 847 455 913 527
rect 1015 455 1081 527
rect 100 202 166 325
rect 200 319 482 353
rect 200 157 247 319
rect 849 319 1078 353
rect 849 255 884 319
rect 805 202 884 255
rect 918 202 991 272
rect 1044 258 1078 319
rect 1044 211 1140 258
rect 200 123 468 157
rect 142 17 210 89
rect 316 17 382 89
rect 503 17 657 89
rect 771 17 837 89
rect 1109 17 1165 177
rect 0 -17 1196 17
<< obsli1 >>
rect 21 421 110 493
rect 611 442 813 476
rect 21 387 574 421
rect 21 359 113 387
rect 21 168 66 359
rect 21 51 108 168
rect 540 305 574 387
rect 611 339 645 442
rect 777 421 813 442
rect 777 387 1165 421
rect 540 271 661 305
rect 281 237 506 265
rect 281 199 562 237
rect 599 199 661 271
rect 528 160 562 199
rect 695 168 729 361
rect 777 289 813 387
rect 1114 292 1165 387
rect 528 157 602 160
rect 695 157 993 168
rect 528 134 993 157
rect 528 123 729 134
rect 695 51 729 123
rect 937 81 993 134
<< metal1 >>
rect 0 496 1196 592
rect 0 -48 1196 48
<< labels >>
rlabel locali s 918 202 991 272 6 A1
port 1 nsew signal input
rlabel locali s 1044 258 1078 319 6 A2
port 2 nsew signal input
rlabel locali s 1044 211 1140 258 6 A2
port 2 nsew signal input
rlabel locali s 849 319 1078 353 6 A2
port 2 nsew signal input
rlabel locali s 849 255 884 319 6 A2
port 2 nsew signal input
rlabel locali s 805 202 884 255 6 A2
port 2 nsew signal input
rlabel locali s 100 202 166 325 6 B1_N
port 3 nsew signal input
rlabel locali s 200 319 482 353 6 X
port 4 nsew signal output
rlabel locali s 200 157 247 319 6 X
port 4 nsew signal output
rlabel locali s 200 123 468 157 6 X
port 4 nsew signal output
rlabel locali s 1109 17 1165 177 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 771 17 837 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 503 17 657 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 316 17 382 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 142 17 210 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 1196 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1196 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 1015 455 1081 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 847 455 913 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 487 455 554 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 316 455 382 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 144 455 210 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 1196 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 1196 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3997818
string GDS_START 3989570
<< end >>
