magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 520 424 586 547
rect 700 424 750 596
rect 896 424 930 596
rect 1060 424 1126 596
rect 520 390 1126 424
rect 25 270 167 356
rect 217 270 455 356
rect 505 270 647 356
rect 697 270 839 356
rect 880 226 946 390
rect 985 260 1127 356
rect 880 192 1129 226
rect 880 119 941 192
rect 1079 70 1129 192
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 24 424 90 596
rect 130 458 180 649
rect 214 424 280 596
rect 318 581 660 615
rect 318 458 384 581
rect 424 424 474 547
rect 24 390 474 424
rect 626 458 660 581
rect 790 458 856 649
rect 970 458 1020 649
rect 23 202 845 236
rect 23 70 73 202
rect 109 17 175 168
rect 223 70 273 202
rect 307 17 373 168
rect 409 70 459 202
rect 493 17 559 168
rect 595 70 645 202
rect 679 85 745 168
rect 779 119 845 202
rect 977 85 1043 158
rect 679 51 1043 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
rlabel locali s 25 270 167 356 6 A1
port 1 nsew signal input
rlabel locali s 217 270 455 356 6 A2
port 2 nsew signal input
rlabel locali s 505 270 647 356 6 A3
port 3 nsew signal input
rlabel locali s 697 270 839 356 6 B1
port 4 nsew signal input
rlabel locali s 985 260 1127 356 6 C1
port 5 nsew signal input
rlabel locali s 1079 70 1129 192 6 Y
port 6 nsew signal output
rlabel locali s 1060 424 1126 596 6 Y
port 6 nsew signal output
rlabel locali s 896 424 930 596 6 Y
port 6 nsew signal output
rlabel locali s 880 226 946 390 6 Y
port 6 nsew signal output
rlabel locali s 880 192 1129 226 6 Y
port 6 nsew signal output
rlabel locali s 880 119 941 192 6 Y
port 6 nsew signal output
rlabel locali s 700 424 750 596 6 Y
port 6 nsew signal output
rlabel locali s 520 424 586 547 6 Y
port 6 nsew signal output
rlabel locali s 520 390 1126 424 6 Y
port 6 nsew signal output
rlabel metal1 s 0 -49 1152 49 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1152 715 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 782804
string GDS_START 772050
<< end >>
