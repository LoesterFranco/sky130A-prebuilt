magic
tech sky130A
magscale 1 2
timestamp 1599588238
<< locali >>
rect 121 310 172 596
rect 138 70 172 310
rect 313 270 455 356
rect 489 270 555 578
rect 597 270 663 356
rect 697 270 839 356
rect 873 270 939 356
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 31 364 81 649
rect 211 458 277 649
rect 351 424 417 596
rect 238 390 417 424
rect 238 310 272 390
rect 36 17 102 226
rect 206 244 272 310
rect 627 424 701 596
rect 735 458 809 649
rect 843 424 909 596
rect 627 390 909 424
rect 238 236 272 244
rect 238 202 904 236
rect 208 17 274 168
rect 356 70 406 202
rect 442 17 516 168
rect 552 70 602 202
rect 636 17 746 168
rect 838 70 904 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
rlabel locali s 873 270 939 356 6 A1
port 1 nsew signal input
rlabel locali s 697 270 839 356 6 A2
port 2 nsew signal input
rlabel locali s 597 270 663 356 6 B1
port 3 nsew signal input
rlabel locali s 489 270 555 578 6 C1
port 4 nsew signal input
rlabel locali s 313 270 455 356 6 D1
port 5 nsew signal input
rlabel locali s 138 70 172 310 6 X
port 6 nsew signal output
rlabel locali s 121 310 172 596 6 X
port 6 nsew signal output
rlabel metal1 s 0 -49 960 49 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 617 960 715 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3893854
string GDS_START 3884908
<< end >>
