magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 422 704
<< pwell >>
rect 0 0 384 49
<< ndiff >>
rect 27 116 357 222
rect 27 82 43 116
rect 77 82 111 116
rect 145 82 239 116
rect 273 82 307 116
rect 341 82 357 116
rect 27 74 357 82
<< pdiff >>
rect 27 584 357 592
rect 27 550 43 584
rect 77 550 111 584
rect 145 550 239 584
rect 273 550 307 584
rect 341 550 357 584
rect 27 368 357 550
<< ndiffc >>
rect 43 82 77 116
rect 111 82 145 116
rect 239 82 273 116
rect 307 82 341 116
<< pdiffc >>
rect 43 550 77 584
rect 111 550 145 584
rect 239 550 273 584
rect 307 550 341 584
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 384 683
rect 27 584 357 649
rect 27 550 43 584
rect 77 550 111 584
rect 145 550 239 584
rect 273 550 307 584
rect 341 550 357 584
rect 27 82 43 116
rect 77 82 111 116
rect 145 82 239 116
rect 273 82 307 116
rect 341 82 357 116
rect 27 17 357 82
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 384 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
<< metal1 >>
rect 0 683 384 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 384 683
rect 0 617 384 649
rect 0 17 384 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 384 17
rect 0 -49 384 -17
<< labels >>
flabel pwell s 0 0 384 49 0 FreeSans 200 0 0 0 VNB
port 2 nsew
flabel nbase s 0 617 384 666 0 FreeSans 200 0 0 0 VPB
port 3 nsew
rlabel comment s 0 0 0 0 4 fill_4
flabel metal1 s 0 617 384 666 0 FreeSans 200 0 0 0 VPWR
port 4 nsew
flabel metal1 s 0 0 384 49 0 FreeSans 200 0 0 0 VGND
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 384 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2390060
string GDS_START 2387616
<< end >>
