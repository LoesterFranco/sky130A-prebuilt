magic
tech sky130A
magscale 1 2
timestamp 1599588209
<< nwell >>
rect -38 332 614 704
<< pwell >>
rect 0 0 576 49
<< scpmos >>
rect 148 368 178 592
rect 238 368 268 592
rect 360 368 390 592
rect 460 368 490 592
<< nmoslvt >>
rect 151 74 181 222
rect 229 74 259 222
rect 343 74 373 222
rect 457 74 487 222
<< ndiff >>
rect 101 132 151 222
rect 27 120 151 132
rect 27 86 38 120
rect 72 86 106 120
rect 140 86 151 120
rect 27 74 151 86
rect 181 74 229 222
rect 259 74 343 222
rect 373 74 457 222
rect 487 202 540 222
rect 487 168 498 202
rect 532 198 540 202
rect 532 168 544 198
rect 487 120 544 168
rect 487 86 498 120
rect 532 86 544 120
rect 487 74 544 86
<< pdiff >>
rect 79 582 148 592
rect 79 548 91 582
rect 125 548 148 582
rect 79 514 148 548
rect 79 480 91 514
rect 125 480 148 514
rect 79 446 148 480
rect 79 412 91 446
rect 125 412 148 446
rect 79 368 148 412
rect 178 580 238 592
rect 178 546 191 580
rect 225 546 238 580
rect 178 497 238 546
rect 178 463 191 497
rect 225 463 238 497
rect 178 414 238 463
rect 178 380 191 414
rect 225 380 238 414
rect 178 368 238 380
rect 268 584 360 592
rect 268 550 296 584
rect 330 550 360 584
rect 268 498 360 550
rect 268 464 296 498
rect 330 464 360 498
rect 268 368 360 464
rect 390 580 460 592
rect 390 546 403 580
rect 437 546 460 580
rect 390 497 460 546
rect 390 463 403 497
rect 437 463 460 497
rect 390 414 460 463
rect 390 380 403 414
rect 437 380 460 414
rect 390 368 460 380
rect 490 580 549 592
rect 490 546 503 580
rect 537 546 549 580
rect 490 497 549 546
rect 490 463 503 497
rect 537 463 549 497
rect 490 414 549 463
rect 490 380 503 414
rect 537 380 549 414
rect 490 368 549 380
<< ndiffc >>
rect 38 86 72 120
rect 106 86 140 120
rect 498 168 532 202
rect 498 86 532 120
<< pdiffc >>
rect 91 548 125 582
rect 91 480 125 514
rect 91 412 125 446
rect 191 546 225 580
rect 191 463 225 497
rect 191 380 225 414
rect 296 550 330 584
rect 296 464 330 498
rect 403 546 437 580
rect 403 463 437 497
rect 403 380 437 414
rect 503 546 537 580
rect 503 463 537 497
rect 503 380 537 414
<< poly >>
rect 148 592 178 618
rect 238 592 268 618
rect 360 592 390 618
rect 460 592 490 618
rect 148 353 178 368
rect 238 353 268 368
rect 360 353 390 368
rect 460 353 490 368
rect 145 310 181 353
rect 235 310 271 353
rect 357 310 393 353
rect 457 310 493 353
rect 115 294 181 310
rect 115 260 131 294
rect 165 260 181 294
rect 115 244 181 260
rect 151 222 181 244
rect 229 294 295 310
rect 229 260 245 294
rect 279 260 295 294
rect 229 244 295 260
rect 343 294 409 310
rect 343 260 359 294
rect 393 260 409 294
rect 343 244 409 260
rect 457 294 555 310
rect 457 260 505 294
rect 539 260 555 294
rect 457 244 555 260
rect 229 222 259 244
rect 343 222 373 244
rect 457 222 487 244
rect 151 48 181 74
rect 229 48 259 74
rect 343 48 373 74
rect 457 48 487 74
<< polycont >>
rect 131 260 165 294
rect 245 260 279 294
rect 359 260 393 294
rect 505 260 539 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 75 582 141 649
rect 75 548 91 582
rect 125 548 141 582
rect 75 514 141 548
rect 75 480 91 514
rect 125 480 141 514
rect 75 446 141 480
rect 75 412 91 446
rect 125 412 141 446
rect 175 580 241 596
rect 175 546 191 580
rect 225 546 241 580
rect 175 497 241 546
rect 175 463 191 497
rect 225 463 241 497
rect 280 584 346 649
rect 280 550 296 584
rect 330 550 346 584
rect 280 498 346 550
rect 280 464 296 498
rect 330 464 346 498
rect 387 580 453 596
rect 387 546 403 580
rect 437 546 453 580
rect 387 497 453 546
rect 175 430 241 463
rect 387 463 403 497
rect 437 463 453 497
rect 387 430 453 463
rect 175 414 453 430
rect 175 380 191 414
rect 225 380 403 414
rect 437 380 453 414
rect 175 378 453 380
rect 47 364 453 378
rect 487 580 553 649
rect 487 546 503 580
rect 537 546 553 580
rect 487 497 553 546
rect 487 463 503 497
rect 537 463 553 497
rect 487 414 553 463
rect 487 380 503 414
rect 537 380 553 414
rect 487 364 553 380
rect 47 344 241 364
rect 47 202 81 344
rect 115 294 181 310
rect 115 260 131 294
rect 165 260 181 294
rect 115 236 181 260
rect 217 294 295 310
rect 217 260 245 294
rect 279 260 295 294
rect 217 236 295 260
rect 343 294 455 310
rect 343 260 359 294
rect 393 260 455 294
rect 343 236 455 260
rect 489 294 555 310
rect 489 260 505 294
rect 539 260 555 294
rect 489 236 555 260
rect 47 168 498 202
rect 532 168 548 202
rect 482 120 548 168
rect 22 86 38 120
rect 72 86 106 120
rect 140 86 157 120
rect 22 17 157 86
rect 482 86 498 120
rect 532 86 548 120
rect 482 70 548 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
rlabel comment s 0 0 0 0 4 nand4_1
flabel pwell s 0 0 576 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nwell s 0 617 576 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 576 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 576 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 223 242 257 276 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 319 390 353 424 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 127 242 161 276 0 FreeSans 340 0 0 0 D
port 4 nsew
flabel corelocali s 415 242 449 276 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 511 242 545 276 0 FreeSans 340 0 0 0 A
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 576 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 2127420
string GDS_START 2122040
<< end >>
