magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 231 333 297 493
rect 438 401 516 493
rect 438 333 536 401
rect 86 215 165 331
rect 231 299 536 333
rect 199 215 265 265
rect 299 147 352 265
rect 482 165 536 299
rect 482 51 600 165
rect 660 145 742 323
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 17 413 85 493
rect 17 181 52 413
rect 129 367 195 527
rect 339 367 403 527
rect 550 435 704 527
rect 748 401 811 493
rect 17 143 244 181
rect 17 97 85 143
rect 210 111 244 143
rect 398 111 448 265
rect 129 17 176 109
rect 210 73 448 111
rect 570 367 811 401
rect 570 199 625 367
rect 777 109 811 367
rect 638 17 708 109
rect 742 51 811 109
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
rlabel locali s 660 145 742 323 6 A_N
port 1 nsew signal input
rlabel locali s 86 215 165 331 6 B_N
port 2 nsew signal input
rlabel locali s 299 147 352 265 6 C
port 3 nsew signal input
rlabel locali s 199 215 265 265 6 D
port 4 nsew signal input
rlabel locali s 482 165 536 299 6 Y
port 5 nsew signal output
rlabel locali s 482 51 600 165 6 Y
port 5 nsew signal output
rlabel locali s 438 401 516 493 6 Y
port 5 nsew signal output
rlabel locali s 438 333 536 401 6 Y
port 5 nsew signal output
rlabel locali s 231 333 297 493 6 Y
port 5 nsew signal output
rlabel locali s 231 299 536 333 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -48 828 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 828 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2354726
string GDS_START 2347394
<< end >>
