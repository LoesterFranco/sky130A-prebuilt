magic
tech sky130A
magscale 1 2
timestamp 1599588238
<< locali >>
rect 113 394 179 596
rect 293 394 359 596
rect 25 360 359 394
rect 504 390 779 424
rect 25 226 71 360
rect 442 270 551 390
rect 585 290 651 356
rect 718 290 779 390
rect 25 192 340 226
rect 109 70 159 192
rect 281 70 340 192
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 23 428 73 649
rect 219 428 253 649
rect 399 424 449 649
rect 490 581 746 615
rect 490 458 556 581
rect 596 492 646 547
rect 680 526 746 581
rect 786 526 841 649
rect 596 458 847 492
rect 119 260 408 326
rect 374 236 408 260
rect 813 236 847 458
rect 374 202 847 236
rect 23 17 73 158
rect 195 17 245 158
rect 384 17 450 168
rect 484 70 550 202
rect 584 17 841 168
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel locali s 718 290 779 390 6 A
port 1 nsew signal input
rlabel locali s 504 390 779 424 6 A
port 1 nsew signal input
rlabel locali s 442 270 551 390 6 A
port 1 nsew signal input
rlabel locali s 585 290 651 356 6 B
port 2 nsew signal input
rlabel locali s 293 394 359 596 6 X
port 3 nsew signal output
rlabel locali s 281 70 340 192 6 X
port 3 nsew signal output
rlabel locali s 113 394 179 596 6 X
port 3 nsew signal output
rlabel locali s 109 70 159 192 6 X
port 3 nsew signal output
rlabel locali s 25 360 359 394 6 X
port 3 nsew signal output
rlabel locali s 25 226 71 360 6 X
port 3 nsew signal output
rlabel locali s 25 192 340 226 6 X
port 3 nsew signal output
rlabel metal1 s 0 -49 864 49 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 617 864 715 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1016712
string GDS_START 1009396
<< end >>
