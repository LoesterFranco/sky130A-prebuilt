magic
tech sky130A
magscale 1 2
timestamp 1599588209
<< nwell >>
rect -38 332 2150 704
<< pwell >>
rect 0 0 2112 49
<< scpmos >>
rect 87 368 117 592
rect 177 368 207 592
rect 267 368 297 592
rect 367 368 397 592
rect 457 368 487 592
rect 547 368 577 592
rect 647 368 677 592
rect 744 368 774 592
rect 837 368 867 592
rect 947 368 977 592
rect 1037 368 1067 592
rect 1147 368 1177 592
rect 1237 368 1267 592
rect 1347 368 1377 592
rect 1437 368 1467 592
rect 1561 368 1591 592
rect 1806 368 1836 592
rect 1906 368 1936 592
rect 1996 368 2026 592
<< nmoslvt >>
rect 84 74 114 222
rect 170 74 200 222
rect 261 74 291 222
rect 347 74 377 222
rect 447 74 477 222
rect 547 74 577 222
rect 650 74 680 222
rect 747 74 777 222
rect 833 74 863 222
rect 919 74 949 222
rect 1005 74 1035 222
rect 1091 74 1121 222
rect 1177 74 1207 222
rect 1263 74 1293 222
rect 1349 74 1379 222
rect 1435 74 1465 222
rect 1825 74 1855 222
rect 1911 74 1941 222
rect 1997 74 2027 222
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 169 170 222
rect 114 135 125 169
rect 159 135 170 169
rect 114 74 170 135
rect 200 143 261 222
rect 200 109 211 143
rect 245 109 261 143
rect 200 74 261 109
rect 291 169 347 222
rect 291 135 302 169
rect 336 135 347 169
rect 291 74 347 135
rect 377 146 447 222
rect 377 112 402 146
rect 436 112 447 146
rect 377 74 447 112
rect 477 169 547 222
rect 477 135 502 169
rect 536 135 547 169
rect 477 74 547 135
rect 577 146 650 222
rect 577 112 602 146
rect 636 112 650 146
rect 577 74 650 112
rect 680 169 747 222
rect 680 135 702 169
rect 736 135 747 169
rect 680 74 747 135
rect 777 210 833 222
rect 777 176 788 210
rect 822 176 833 210
rect 777 120 833 176
rect 777 86 788 120
rect 822 86 833 120
rect 777 74 833 86
rect 863 184 919 222
rect 863 150 874 184
rect 908 150 919 184
rect 863 116 919 150
rect 863 82 874 116
rect 908 82 919 116
rect 863 74 919 82
rect 949 210 1005 222
rect 949 176 960 210
rect 994 176 1005 210
rect 949 120 1005 176
rect 949 86 960 120
rect 994 86 1005 120
rect 949 74 1005 86
rect 1035 210 1091 222
rect 1035 176 1046 210
rect 1080 176 1091 210
rect 1035 120 1091 176
rect 1035 86 1046 120
rect 1080 86 1091 120
rect 1035 74 1091 86
rect 1121 210 1177 222
rect 1121 176 1132 210
rect 1166 176 1177 210
rect 1121 120 1177 176
rect 1121 86 1132 120
rect 1166 86 1177 120
rect 1121 74 1177 86
rect 1207 210 1263 222
rect 1207 176 1218 210
rect 1252 176 1263 210
rect 1207 120 1263 176
rect 1207 86 1218 120
rect 1252 86 1263 120
rect 1207 74 1263 86
rect 1293 210 1349 222
rect 1293 176 1304 210
rect 1338 176 1349 210
rect 1293 120 1349 176
rect 1293 86 1304 120
rect 1338 86 1349 120
rect 1293 74 1349 86
rect 1379 210 1435 222
rect 1379 176 1390 210
rect 1424 176 1435 210
rect 1379 120 1435 176
rect 1379 86 1390 120
rect 1424 86 1435 120
rect 1379 74 1435 86
rect 1465 210 1522 222
rect 1465 176 1476 210
rect 1510 176 1522 210
rect 1465 120 1522 176
rect 1465 86 1476 120
rect 1510 86 1522 120
rect 1465 74 1522 86
rect 1768 197 1825 222
rect 1768 163 1780 197
rect 1814 163 1825 197
rect 1768 120 1825 163
rect 1768 86 1780 120
rect 1814 86 1825 120
rect 1768 74 1825 86
rect 1855 186 1911 222
rect 1855 152 1866 186
rect 1900 152 1911 186
rect 1855 118 1911 152
rect 1855 84 1866 118
rect 1900 84 1911 118
rect 1855 74 1911 84
rect 1941 202 1997 222
rect 1941 168 1952 202
rect 1986 168 1997 202
rect 1941 118 1997 168
rect 1941 84 1952 118
rect 1986 84 1997 118
rect 1941 74 1997 84
rect 2027 120 2085 222
rect 2027 86 2038 120
rect 2072 86 2085 120
rect 2027 74 2085 86
<< pdiff >>
rect 1485 614 1543 626
rect 1485 592 1497 614
rect 28 580 87 592
rect 28 546 40 580
rect 74 546 87 580
rect 28 497 87 546
rect 28 463 40 497
rect 74 463 87 497
rect 28 414 87 463
rect 28 380 40 414
rect 74 380 87 414
rect 28 368 87 380
rect 117 547 177 592
rect 117 513 130 547
rect 164 513 177 547
rect 117 479 177 513
rect 117 445 130 479
rect 164 445 177 479
rect 117 411 177 445
rect 117 377 130 411
rect 164 377 177 411
rect 117 368 177 377
rect 207 580 267 592
rect 207 546 220 580
rect 254 546 267 580
rect 207 482 267 546
rect 207 448 220 482
rect 254 448 267 482
rect 207 368 267 448
rect 297 547 367 592
rect 297 513 320 547
rect 354 513 367 547
rect 297 479 367 513
rect 297 445 320 479
rect 354 445 367 479
rect 297 411 367 445
rect 297 377 320 411
rect 354 377 367 411
rect 297 368 367 377
rect 397 580 457 592
rect 397 546 410 580
rect 444 546 457 580
rect 397 482 457 546
rect 397 448 410 482
rect 444 448 457 482
rect 397 368 457 448
rect 487 547 547 592
rect 487 513 500 547
rect 534 513 547 547
rect 487 479 547 513
rect 487 445 500 479
rect 534 445 547 479
rect 487 411 547 445
rect 487 377 500 411
rect 534 377 547 411
rect 487 368 547 377
rect 577 580 647 592
rect 577 546 600 580
rect 634 546 647 580
rect 577 482 647 546
rect 577 448 600 482
rect 634 448 647 482
rect 577 368 647 448
rect 677 547 744 592
rect 677 513 690 547
rect 724 513 744 547
rect 677 479 744 513
rect 677 445 690 479
rect 724 445 744 479
rect 677 411 744 445
rect 677 377 690 411
rect 724 377 744 411
rect 677 368 744 377
rect 774 580 837 592
rect 774 546 790 580
rect 824 546 837 580
rect 774 512 837 546
rect 774 478 790 512
rect 824 478 837 512
rect 774 368 837 478
rect 867 580 947 592
rect 867 546 890 580
rect 924 546 947 580
rect 867 368 947 546
rect 977 580 1037 592
rect 977 546 990 580
rect 1024 546 1037 580
rect 977 512 1037 546
rect 977 478 990 512
rect 1024 478 1037 512
rect 977 368 1037 478
rect 1067 580 1147 592
rect 1067 546 1090 580
rect 1124 546 1147 580
rect 1067 368 1147 546
rect 1177 580 1237 592
rect 1177 546 1190 580
rect 1224 546 1237 580
rect 1177 512 1237 546
rect 1177 478 1190 512
rect 1224 478 1237 512
rect 1177 368 1237 478
rect 1267 580 1347 592
rect 1267 546 1290 580
rect 1324 546 1347 580
rect 1267 368 1347 546
rect 1377 580 1437 592
rect 1377 546 1390 580
rect 1424 546 1437 580
rect 1377 512 1437 546
rect 1377 478 1390 512
rect 1424 478 1437 512
rect 1377 368 1437 478
rect 1467 580 1497 592
rect 1531 592 1543 614
rect 1531 580 1561 592
rect 1467 368 1561 580
rect 1591 571 1650 592
rect 1591 537 1604 571
rect 1638 537 1650 571
rect 1591 368 1650 537
rect 1704 410 1806 592
rect 1704 376 1737 410
rect 1771 376 1806 410
rect 1704 368 1806 376
rect 1836 561 1906 592
rect 1836 527 1849 561
rect 1883 527 1906 561
rect 1836 368 1906 527
rect 1936 580 1996 592
rect 1936 546 1949 580
rect 1983 546 1996 580
rect 1936 497 1996 546
rect 1936 463 1949 497
rect 1983 463 1996 497
rect 1936 414 1996 463
rect 1936 380 1949 414
rect 1983 380 1996 414
rect 1936 368 1996 380
rect 2026 582 2085 592
rect 2026 548 2039 582
rect 2073 548 2085 582
rect 2026 514 2085 548
rect 2026 480 2039 514
rect 2073 480 2085 514
rect 2026 446 2085 480
rect 2026 412 2039 446
rect 2073 412 2085 446
rect 2026 368 2085 412
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 125 135 159 169
rect 211 109 245 143
rect 302 135 336 169
rect 402 112 436 146
rect 502 135 536 169
rect 602 112 636 146
rect 702 135 736 169
rect 788 176 822 210
rect 788 86 822 120
rect 874 150 908 184
rect 874 82 908 116
rect 960 176 994 210
rect 960 86 994 120
rect 1046 176 1080 210
rect 1046 86 1080 120
rect 1132 176 1166 210
rect 1132 86 1166 120
rect 1218 176 1252 210
rect 1218 86 1252 120
rect 1304 176 1338 210
rect 1304 86 1338 120
rect 1390 176 1424 210
rect 1390 86 1424 120
rect 1476 176 1510 210
rect 1476 86 1510 120
rect 1780 163 1814 197
rect 1780 86 1814 120
rect 1866 152 1900 186
rect 1866 84 1900 118
rect 1952 168 1986 202
rect 1952 84 1986 118
rect 2038 86 2072 120
<< pdiffc >>
rect 40 546 74 580
rect 40 463 74 497
rect 40 380 74 414
rect 130 513 164 547
rect 130 445 164 479
rect 130 377 164 411
rect 220 546 254 580
rect 220 448 254 482
rect 320 513 354 547
rect 320 445 354 479
rect 320 377 354 411
rect 410 546 444 580
rect 410 448 444 482
rect 500 513 534 547
rect 500 445 534 479
rect 500 377 534 411
rect 600 546 634 580
rect 600 448 634 482
rect 690 513 724 547
rect 690 445 724 479
rect 690 377 724 411
rect 790 546 824 580
rect 790 478 824 512
rect 890 546 924 580
rect 990 546 1024 580
rect 990 478 1024 512
rect 1090 546 1124 580
rect 1190 546 1224 580
rect 1190 478 1224 512
rect 1290 546 1324 580
rect 1390 546 1424 580
rect 1390 478 1424 512
rect 1497 580 1531 614
rect 1604 537 1638 571
rect 1737 376 1771 410
rect 1849 527 1883 561
rect 1949 546 1983 580
rect 1949 463 1983 497
rect 1949 380 1983 414
rect 2039 548 2073 582
rect 2039 480 2073 514
rect 2039 412 2073 446
<< poly >>
rect 87 592 117 618
rect 177 592 207 618
rect 267 592 297 618
rect 367 592 397 618
rect 457 592 487 618
rect 547 592 577 618
rect 647 592 677 618
rect 744 592 774 618
rect 837 592 867 618
rect 947 592 977 618
rect 1037 592 1067 618
rect 1147 592 1177 618
rect 1237 592 1267 618
rect 1347 592 1377 618
rect 1437 592 1467 618
rect 1561 592 1591 618
rect 1806 592 1836 618
rect 1906 592 1936 618
rect 1996 592 2026 618
rect 87 353 117 368
rect 177 353 207 368
rect 267 353 297 368
rect 367 353 397 368
rect 457 353 487 368
rect 547 353 577 368
rect 647 353 677 368
rect 744 353 774 368
rect 837 353 867 368
rect 947 353 977 368
rect 1037 353 1067 368
rect 1147 353 1177 368
rect 1237 353 1267 368
rect 1347 353 1377 368
rect 1437 353 1467 368
rect 1561 353 1591 368
rect 1806 353 1836 368
rect 1906 353 1936 368
rect 1996 353 2026 368
rect 84 330 120 353
rect 174 330 210 353
rect 264 330 300 353
rect 364 330 400 353
rect 454 330 490 353
rect 544 330 580 353
rect 644 330 680 353
rect 741 330 777 353
rect 84 314 777 330
rect 834 323 1839 353
rect 84 280 211 314
rect 245 280 279 314
rect 313 280 347 314
rect 381 280 415 314
rect 449 280 483 314
rect 517 280 551 314
rect 585 280 619 314
rect 653 280 687 314
rect 721 280 777 314
rect 84 264 777 280
rect 1653 310 1839 323
rect 1903 310 1939 353
rect 1993 310 2029 353
rect 1653 294 1855 310
rect 84 222 114 264
rect 170 222 200 264
rect 261 222 291 264
rect 347 222 377 264
rect 447 222 477 264
rect 547 222 577 264
rect 650 222 680 264
rect 747 222 777 264
rect 833 237 1574 267
rect 1653 260 1669 294
rect 1703 260 1737 294
rect 1771 260 1805 294
rect 1839 260 1855 294
rect 1653 244 1855 260
rect 1903 294 2029 310
rect 1903 260 1945 294
rect 1979 260 2029 294
rect 1903 244 2029 260
rect 833 222 863 237
rect 919 222 949 237
rect 1005 222 1035 237
rect 1091 222 1121 237
rect 1177 222 1207 237
rect 1263 222 1293 237
rect 1349 222 1379 237
rect 1435 222 1465 237
rect 1544 134 1574 237
rect 1825 222 1855 244
rect 1911 222 1941 244
rect 1997 222 2027 244
rect 1544 118 1746 134
rect 1544 84 1560 118
rect 1594 84 1628 118
rect 1662 84 1696 118
rect 1730 84 1746 118
rect 84 48 114 74
rect 170 48 200 74
rect 261 48 291 74
rect 347 48 377 74
rect 447 48 477 74
rect 547 48 577 74
rect 650 48 680 74
rect 747 48 777 74
rect 833 48 863 74
rect 919 48 949 74
rect 1005 48 1035 74
rect 1091 48 1121 74
rect 1177 48 1207 74
rect 1263 48 1293 74
rect 1349 48 1379 74
rect 1435 48 1465 74
rect 1544 68 1746 84
rect 1825 48 1855 74
rect 1911 48 1941 74
rect 1997 48 2027 74
<< polycont >>
rect 211 280 245 314
rect 279 280 313 314
rect 347 280 381 314
rect 415 280 449 314
rect 483 280 517 314
rect 551 280 585 314
rect 619 280 653 314
rect 687 280 721 314
rect 1669 260 1703 294
rect 1737 260 1771 294
rect 1805 260 1839 294
rect 1945 260 1979 294
rect 1560 84 1594 118
rect 1628 84 1662 118
rect 1696 84 1730 118
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 24 581 840 615
rect 24 580 74 581
rect 24 546 40 580
rect 217 580 270 581
rect 24 497 74 546
rect 24 463 40 497
rect 24 414 74 463
rect 24 380 40 414
rect 24 364 74 380
rect 109 513 130 547
rect 164 513 180 547
rect 109 479 180 513
rect 109 445 130 479
rect 164 445 180 479
rect 109 411 180 445
rect 217 546 220 580
rect 254 546 270 580
rect 410 580 444 581
rect 217 482 270 546
rect 217 448 220 482
rect 254 448 270 482
rect 217 432 270 448
rect 304 513 320 547
rect 354 513 370 547
rect 304 479 370 513
rect 304 445 320 479
rect 354 445 370 479
rect 109 377 130 411
rect 164 398 180 411
rect 304 411 370 445
rect 584 580 638 581
rect 410 482 444 546
rect 410 432 444 448
rect 484 513 500 547
rect 534 513 550 547
rect 484 479 550 513
rect 484 445 500 479
rect 534 445 550 479
rect 304 398 320 411
rect 164 377 320 398
rect 354 398 370 411
rect 484 411 550 445
rect 584 546 600 580
rect 634 546 638 580
rect 774 580 840 581
rect 584 482 638 546
rect 584 448 600 482
rect 634 448 638 482
rect 584 432 638 448
rect 674 513 690 547
rect 724 513 740 547
rect 674 479 740 513
rect 674 445 690 479
rect 724 445 740 479
rect 774 546 790 580
rect 824 546 840 580
rect 874 580 940 649
rect 874 546 890 580
rect 924 546 940 580
rect 974 580 1040 596
rect 974 546 990 580
rect 1024 546 1040 580
rect 1074 580 1140 649
rect 1074 546 1090 580
rect 1124 546 1140 580
rect 1174 580 1240 596
rect 1174 546 1190 580
rect 1224 546 1240 580
rect 1274 580 1340 649
rect 1481 614 1547 649
rect 1274 546 1290 580
rect 1324 546 1340 580
rect 1374 580 1440 596
rect 1481 580 1497 614
rect 1531 580 1547 614
rect 1374 546 1390 580
rect 1424 546 1440 580
rect 1588 571 1654 596
rect 1588 546 1604 571
rect 774 512 840 546
rect 974 512 1040 546
rect 1174 512 1240 546
rect 1374 537 1604 546
rect 1638 537 1654 571
rect 1374 512 1654 537
rect 1833 561 1899 649
rect 1833 527 1849 561
rect 1883 527 1899 561
rect 1833 512 1899 527
rect 1933 580 1989 596
rect 1933 546 1949 580
rect 1983 546 1989 580
rect 774 478 790 512
rect 824 478 990 512
rect 1024 478 1190 512
rect 1224 478 1390 512
rect 1424 478 1440 512
rect 1933 497 1989 546
rect 1933 478 1949 497
rect 484 398 500 411
rect 354 377 500 398
rect 534 398 550 411
rect 674 411 740 445
rect 1517 463 1949 478
rect 1983 463 1989 497
rect 1517 444 1989 463
rect 674 398 690 411
rect 534 377 690 398
rect 724 377 740 411
rect 109 364 740 377
rect 774 410 1551 444
rect 1933 414 1989 444
rect 109 230 167 364
rect 774 330 808 410
rect 207 314 808 330
rect 207 280 211 314
rect 245 280 279 314
rect 313 280 347 314
rect 381 280 415 314
rect 449 280 483 314
rect 517 280 551 314
rect 585 280 619 314
rect 653 280 687 314
rect 721 296 808 314
rect 1585 376 1737 410
rect 1771 376 1809 410
rect 1585 360 1809 376
rect 1933 380 1949 414
rect 1983 380 1989 414
rect 2023 582 2089 649
rect 2023 548 2039 582
rect 2073 548 2089 582
rect 2023 514 2089 548
rect 2023 480 2039 514
rect 2073 480 2089 514
rect 2023 446 2089 480
rect 2023 412 2039 446
rect 2073 412 2089 446
rect 1933 378 1989 380
rect 721 280 731 296
rect 207 264 731 280
rect 944 262 1510 294
rect 788 260 1510 262
rect 23 210 73 226
rect 23 176 39 210
rect 23 120 73 176
rect 23 86 39 120
rect 109 196 752 230
rect 109 169 175 196
rect 109 135 125 169
rect 159 135 175 169
rect 286 169 352 196
rect 109 119 175 135
rect 211 143 245 162
rect 23 85 73 86
rect 286 135 302 169
rect 336 135 352 169
rect 486 169 552 196
rect 286 119 352 135
rect 386 146 452 162
rect 211 85 245 109
rect 386 112 402 146
rect 436 112 452 146
rect 486 135 502 169
rect 536 135 552 169
rect 686 169 752 196
rect 486 119 552 135
rect 586 146 652 162
rect 386 85 452 112
rect 586 112 602 146
rect 636 112 652 146
rect 686 135 702 169
rect 736 135 752 169
rect 686 119 752 135
rect 788 228 1010 260
rect 788 210 822 228
rect 960 210 1010 228
rect 788 120 822 176
rect 586 85 652 112
rect 788 85 822 86
rect 23 51 822 85
rect 858 184 924 194
rect 858 150 874 184
rect 908 150 924 184
rect 858 116 924 150
rect 858 82 874 116
rect 908 82 924 116
rect 858 17 924 82
rect 994 176 1010 210
rect 960 120 1010 176
rect 994 86 1010 120
rect 960 70 1010 86
rect 1046 210 1080 226
rect 1046 120 1080 176
rect 1046 17 1080 86
rect 1116 210 1166 260
rect 1116 176 1132 210
rect 1116 120 1166 176
rect 1116 86 1132 120
rect 1116 70 1166 86
rect 1202 210 1252 226
rect 1202 176 1218 210
rect 1202 120 1252 176
rect 1202 86 1218 120
rect 1202 17 1252 86
rect 1288 210 1338 260
rect 1288 176 1304 210
rect 1288 120 1338 176
rect 1288 86 1304 120
rect 1288 70 1338 86
rect 1374 210 1424 226
rect 1374 176 1390 210
rect 1374 120 1424 176
rect 1374 86 1390 120
rect 1374 17 1424 86
rect 1460 210 1510 260
rect 1460 176 1476 210
rect 1460 120 1510 176
rect 1585 202 1619 360
rect 1933 344 2063 378
rect 1653 294 1895 310
rect 1653 260 1669 294
rect 1703 260 1737 294
rect 1771 260 1805 294
rect 1839 260 1895 294
rect 1653 236 1895 260
rect 1929 294 1995 310
rect 1929 260 1945 294
rect 1979 260 1995 294
rect 1929 236 1995 260
rect 2029 202 2063 344
rect 1585 197 1830 202
rect 1585 163 1780 197
rect 1814 163 1830 197
rect 1585 134 1830 163
rect 1460 86 1476 120
rect 1460 70 1510 86
rect 1544 120 1830 134
rect 1544 118 1780 120
rect 1544 84 1560 118
rect 1594 84 1628 118
rect 1662 84 1696 118
rect 1730 86 1780 118
rect 1814 86 1830 120
rect 1730 84 1830 86
rect 1544 68 1830 84
rect 1866 186 1900 202
rect 1866 118 1900 152
rect 1866 17 1900 84
rect 1936 168 1952 202
rect 1986 168 2063 202
rect 1936 118 1986 168
rect 1936 84 1952 118
rect 1936 68 1986 84
rect 2022 86 2038 120
rect 2072 86 2089 120
rect 2022 17 2089 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
<< metal1 >>
rect 0 683 2112 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 0 617 2112 649
rect 0 17 2112 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
rect 0 -49 2112 -17
<< labels >>
rlabel comment s 0 0 0 0 4 ebufn_8
flabel pwell s 0 0 2112 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nwell s 0 617 2112 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 0 617 2112 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 2112 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 1663 242 1697 276 0 FreeSans 340 0 0 0 TE_B
port 2 nsew
flabel corelocali s 1759 242 1793 276 0 FreeSans 340 0 0 0 TE_B
port 2 nsew
flabel corelocali s 1855 242 1889 276 0 FreeSans 340 0 0 0 TE_B
port 2 nsew
flabel corelocali s 1951 242 1985 276 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 127 168 161 202 0 FreeSans 340 0 0 0 Z
port 7 nsew
flabel corelocali s 127 242 161 276 0 FreeSans 340 0 0 0 Z
port 7 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 Z
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 2112 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 2408520
string GDS_START 2393746
<< end >>
