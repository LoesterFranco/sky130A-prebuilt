magic
tech sky130A
magscale 1 2
timestamp 1604502693
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 79 47 109 177
rect 171 47 201 177
rect 359 47 389 131
rect 443 47 473 131
rect 527 47 557 131
rect 736 47 766 131
rect 808 47 838 131
rect 903 47 933 177
rect 995 47 1025 177
<< pmoshvt >>
rect 79 297 109 497
rect 171 297 201 497
rect 354 369 384 497
rect 438 369 468 497
rect 548 369 578 497
rect 720 369 750 497
rect 808 369 838 497
rect 903 297 933 497
rect 995 297 1025 497
<< ndiff >>
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 165 171 177
rect 109 131 127 165
rect 161 131 171 165
rect 109 97 171 131
rect 109 63 127 97
rect 161 63 171 97
rect 109 47 171 63
rect 201 161 253 177
rect 201 127 211 161
rect 245 127 253 161
rect 853 131 903 177
rect 201 93 253 127
rect 201 59 211 93
rect 245 59 253 93
rect 201 47 253 59
rect 307 119 359 131
rect 307 85 315 119
rect 349 85 359 119
rect 307 47 359 85
rect 389 119 443 131
rect 389 85 399 119
rect 433 85 443 119
rect 389 47 443 85
rect 473 93 527 131
rect 473 59 483 93
rect 517 59 527 93
rect 473 47 527 59
rect 557 119 609 131
rect 557 85 567 119
rect 601 85 609 119
rect 557 47 609 85
rect 684 119 736 131
rect 684 85 692 119
rect 726 85 736 119
rect 684 47 736 85
rect 766 47 808 131
rect 838 93 903 131
rect 838 59 859 93
rect 893 59 903 93
rect 838 47 903 59
rect 933 165 995 177
rect 933 131 943 165
rect 977 131 995 165
rect 933 97 995 131
rect 933 63 943 97
rect 977 63 995 97
rect 933 47 995 63
rect 1025 161 1077 177
rect 1025 127 1035 161
rect 1069 127 1077 161
rect 1025 93 1077 127
rect 1025 59 1035 93
rect 1069 59 1077 93
rect 1025 47 1077 59
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 483 171 497
rect 109 449 127 483
rect 161 449 171 483
rect 109 415 171 449
rect 109 381 127 415
rect 161 381 171 415
rect 109 347 171 381
rect 109 313 127 347
rect 161 313 171 347
rect 109 297 171 313
rect 201 489 354 497
rect 201 455 211 489
rect 245 455 354 489
rect 201 421 354 455
rect 201 387 211 421
rect 245 387 354 421
rect 201 369 354 387
rect 384 475 438 497
rect 384 441 394 475
rect 428 441 438 475
rect 384 369 438 441
rect 468 369 548 497
rect 578 475 720 497
rect 578 441 598 475
rect 632 441 666 475
rect 700 441 720 475
rect 578 369 720 441
rect 750 455 808 497
rect 750 421 762 455
rect 796 421 808 455
rect 750 369 808 421
rect 838 475 903 497
rect 838 441 859 475
rect 893 441 903 475
rect 838 369 903 441
rect 201 353 253 369
rect 201 319 211 353
rect 245 319 253 353
rect 201 297 253 319
rect 853 297 903 369
rect 933 467 995 497
rect 933 433 943 467
rect 977 433 995 467
rect 933 359 995 433
rect 933 325 943 359
rect 977 325 995 359
rect 933 297 995 325
rect 1025 485 1077 497
rect 1025 451 1035 485
rect 1069 451 1077 485
rect 1025 417 1077 451
rect 1025 383 1035 417
rect 1069 383 1077 417
rect 1025 349 1077 383
rect 1025 315 1035 349
rect 1069 315 1077 349
rect 1025 297 1077 315
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 127 131 161 165
rect 127 63 161 97
rect 211 127 245 161
rect 211 59 245 93
rect 315 85 349 119
rect 399 85 433 119
rect 483 59 517 93
rect 567 85 601 119
rect 692 85 726 119
rect 859 59 893 93
rect 943 131 977 165
rect 943 63 977 97
rect 1035 127 1069 161
rect 1035 59 1069 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 127 449 161 483
rect 127 381 161 415
rect 127 313 161 347
rect 211 455 245 489
rect 211 387 245 421
rect 394 441 428 475
rect 598 441 632 475
rect 666 441 700 475
rect 762 421 796 455
rect 859 441 893 475
rect 211 319 245 353
rect 943 433 977 467
rect 943 325 977 359
rect 1035 451 1069 485
rect 1035 383 1069 417
rect 1035 315 1069 349
<< poly >>
rect 79 497 109 523
rect 171 497 201 523
rect 354 497 384 523
rect 438 497 468 523
rect 548 497 578 523
rect 720 497 750 523
rect 808 497 838 523
rect 903 497 933 523
rect 995 497 1025 523
rect 79 265 109 297
rect 171 265 201 297
rect 354 265 384 369
rect 438 285 468 369
rect 438 269 506 285
rect 79 249 250 265
rect 79 215 206 249
rect 240 215 250 249
rect 79 199 250 215
rect 342 249 396 265
rect 342 215 352 249
rect 386 215 396 249
rect 438 235 462 269
rect 496 235 506 269
rect 438 219 506 235
rect 548 261 578 369
rect 720 349 750 369
rect 683 337 750 349
rect 659 321 750 337
rect 659 287 669 321
rect 703 319 750 321
rect 703 287 713 319
rect 659 271 713 287
rect 808 273 838 369
rect 548 245 618 261
rect 342 199 396 215
rect 79 177 109 199
rect 171 177 201 199
rect 359 131 389 199
rect 443 131 473 219
rect 548 211 574 245
rect 608 211 618 245
rect 548 195 618 211
rect 548 177 583 195
rect 527 147 583 177
rect 683 177 713 271
rect 755 263 838 273
rect 903 265 933 297
rect 995 265 1025 297
rect 755 229 771 263
rect 805 229 838 263
rect 755 219 838 229
rect 683 147 766 177
rect 527 131 557 147
rect 736 131 766 147
rect 808 131 838 219
rect 880 249 1025 265
rect 880 215 890 249
rect 924 215 1025 249
rect 880 199 1025 215
rect 903 177 933 199
rect 995 177 1025 199
rect 79 21 109 47
rect 171 21 201 47
rect 359 21 389 47
rect 443 21 473 47
rect 527 21 557 47
rect 736 21 766 47
rect 808 21 838 47
rect 903 21 933 47
rect 995 21 1025 47
<< polycont >>
rect 206 215 240 249
rect 352 215 386 249
rect 462 235 496 269
rect 669 287 703 321
rect 574 211 608 245
rect 771 229 805 263
rect 890 215 924 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 27 485 75 527
rect 27 451 35 485
rect 69 451 75 485
rect 211 489 250 527
rect 27 417 75 451
rect 27 383 35 417
rect 69 383 75 417
rect 27 349 75 383
rect 27 315 35 349
rect 69 315 75 349
rect 27 299 75 315
rect 111 449 127 483
rect 161 449 177 483
rect 111 415 177 449
rect 111 381 127 415
rect 161 381 177 415
rect 111 347 177 381
rect 111 313 127 347
rect 161 313 177 347
rect 245 455 250 489
rect 570 475 728 527
rect 211 421 250 455
rect 245 387 250 421
rect 211 353 250 387
rect 245 319 250 353
rect 27 161 75 177
rect 27 127 35 161
rect 69 127 75 161
rect 27 93 75 127
rect 27 59 35 93
rect 69 59 75 93
rect 111 165 156 313
rect 211 303 250 319
rect 284 441 394 475
rect 428 441 444 475
rect 570 441 598 475
rect 632 441 666 475
rect 700 441 728 475
rect 843 475 909 527
rect 1029 485 1077 527
rect 762 455 796 471
rect 284 249 318 441
rect 843 441 859 475
rect 893 441 909 475
rect 943 467 993 483
rect 762 405 796 421
rect 977 433 993 467
rect 190 215 206 249
rect 240 215 318 249
rect 111 131 127 165
rect 161 131 177 165
rect 111 97 177 131
rect 111 63 127 97
rect 161 63 177 97
rect 211 161 250 177
rect 245 127 250 161
rect 211 93 250 127
rect 27 17 75 59
rect 245 59 250 93
rect 284 135 318 215
rect 352 371 893 405
rect 352 249 386 371
rect 352 199 386 215
rect 462 321 719 335
rect 462 287 669 321
rect 703 287 719 321
rect 462 279 719 287
rect 462 269 523 279
rect 496 235 523 269
rect 764 263 809 335
rect 764 245 771 263
rect 462 201 523 235
rect 558 211 574 245
rect 608 229 771 245
rect 805 229 809 263
rect 608 211 809 229
rect 859 265 893 371
rect 943 359 993 433
rect 977 325 993 359
rect 943 309 993 325
rect 859 249 924 265
rect 859 215 890 249
rect 859 199 924 215
rect 859 177 893 199
rect 284 119 349 135
rect 284 85 315 119
rect 284 69 349 85
rect 399 127 601 161
rect 399 119 433 127
rect 567 119 601 127
rect 399 69 433 85
rect 211 17 250 59
rect 467 59 483 93
rect 517 59 533 93
rect 567 69 601 85
rect 692 143 893 177
rect 958 165 993 309
rect 1029 451 1035 485
rect 1069 451 1077 485
rect 1029 417 1077 451
rect 1029 383 1035 417
rect 1069 383 1077 417
rect 1029 349 1077 383
rect 1029 315 1035 349
rect 1069 315 1077 349
rect 1029 299 1077 315
rect 692 119 726 143
rect 927 131 943 165
rect 977 131 993 165
rect 692 69 726 85
rect 843 93 893 109
rect 467 17 533 59
rect 843 59 859 93
rect 927 97 993 131
rect 927 63 943 97
rect 977 63 993 97
rect 1029 161 1077 177
rect 1029 127 1035 161
rect 1069 127 1077 161
rect 1029 93 1077 127
rect 843 17 893 59
rect 1029 59 1035 93
rect 1069 59 1077 93
rect 1029 17 1077 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew
flabel corelocali s 764 221 798 255 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 948 357 982 391 0 FreeSans 340 0 0 0 COUT
port 7 nsew
flabel corelocali s 948 85 982 119 0 FreeSans 340 0 0 0 COUT
port 7 nsew
flabel corelocali s 122 85 156 119 0 FreeSans 340 0 0 0 SUM
port 8 nsew
flabel corelocali s 122 153 156 187 0 FreeSans 340 0 0 0 SUM
port 8 nsew
flabel corelocali s 122 221 156 255 0 FreeSans 340 0 0 0 SUM
port 8 nsew
flabel corelocali s 122 289 156 323 0 FreeSans 340 0 0 0 SUM
port 8 nsew
flabel corelocali s 122 357 156 391 0 FreeSans 340 0 0 0 SUM
port 8 nsew
flabel corelocali s 122 425 156 459 0 FreeSans 340 0 0 0 SUM
port 8 nsew
flabel corelocali s 948 425 982 459 0 FreeSans 340 0 0 0 COUT
port 7 nsew
flabel corelocali s 764 289 798 323 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 489 289 523 323 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 489 221 523 255 0 FreeSans 340 0 0 0 B
port 2 nsew
rlabel comment s 0 0 0 0 4 ha_2
<< properties >>
string FIXED_BBOX 0 0 1104 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2131262
string GDS_START 2121692
string path 14.600 1.725 14.600 3.600 10.400 3.600 10.400 1.725 
<< end >>
