magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1288 561
rect 103 427 169 527
rect 290 439 363 527
rect 17 197 66 325
rect 103 17 169 89
rect 305 287 437 337
rect 296 17 362 181
rect 397 77 437 287
rect 679 427 739 527
rect 862 402 919 527
rect 1114 426 1184 527
rect 1038 221 1102 287
rect 1218 299 1271 491
rect 779 17 829 122
rect 1234 119 1271 299
rect 1134 17 1168 109
rect 1211 51 1271 119
rect 0 -17 1288 17
<< obsli1 >>
rect 35 393 69 493
rect 203 405 248 493
rect 495 451 645 485
rect 35 359 156 393
rect 122 278 156 359
rect 203 371 518 405
rect 122 212 168 278
rect 122 157 156 212
rect 35 123 156 157
rect 35 52 69 123
rect 203 52 256 371
rect 478 197 518 371
rect 611 265 645 451
rect 782 373 826 487
rect 686 368 826 373
rect 1001 379 1067 493
rect 686 307 942 368
rect 1001 345 1184 379
rect 869 265 942 307
rect 611 231 835 265
rect 711 199 835 231
rect 869 199 948 265
rect 1150 265 1184 345
rect 478 163 644 197
rect 711 112 745 199
rect 869 123 916 199
rect 1150 187 1200 265
rect 987 153 1200 187
rect 987 124 1031 153
rect 558 78 745 112
rect 864 51 916 123
rect 968 58 1031 124
<< metal1 >>
rect 0 496 1288 592
rect 17 252 76 261
rect 1030 252 1088 261
rect 17 224 1088 252
rect 17 215 76 224
rect 1030 215 1088 224
rect 0 -48 1288 48
<< labels >>
rlabel locali s 397 77 437 287 6 GATE
port 1 nsew signal input
rlabel locali s 305 287 437 337 6 GATE
port 1 nsew signal input
rlabel locali s 1234 119 1271 299 6 GCLK
port 2 nsew signal output
rlabel locali s 1218 299 1271 491 6 GCLK
port 2 nsew signal output
rlabel locali s 1211 51 1271 119 6 GCLK
port 2 nsew signal output
rlabel locali s 17 197 66 325 6 CLK
port 3 nsew clock input
rlabel locali s 1038 221 1102 287 6 CLK
port 3 nsew clock input
rlabel metal1 s 1030 252 1088 261 6 CLK
port 3 nsew clock input
rlabel metal1 s 1030 215 1088 224 6 CLK
port 3 nsew clock input
rlabel metal1 s 17 252 76 261 6 CLK
port 3 nsew clock input
rlabel metal1 s 17 224 1088 252 6 CLK
port 3 nsew clock input
rlabel metal1 s 17 215 76 224 6 CLK
port 3 nsew clock input
rlabel locali s 1134 17 1168 109 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 779 17 829 122 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 296 17 362 181 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 103 17 169 89 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 1288 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1288 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 1114 426 1184 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 862 402 919 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 679 427 739 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 290 439 363 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 103 427 169 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 1288 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 1288 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1288 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2575634
string GDS_START 2565668
<< end >>
