magic
tech sky130A
magscale 1 2
timestamp 1604502710
<< nwell >>
rect -38 332 1670 704
<< pwell >>
rect 0 0 1632 49
<< scpmos >>
rect 149 368 185 592
rect 239 368 275 592
rect 329 368 365 592
rect 419 368 455 592
rect 526 386 562 554
rect 616 386 652 554
rect 818 368 854 592
rect 908 368 944 592
rect 1000 368 1036 592
rect 1090 368 1126 592
rect 1180 368 1216 592
rect 1270 368 1306 592
rect 1368 368 1404 592
rect 1468 368 1504 592
<< nmoslvt >>
rect 110 74 140 222
rect 196 74 226 222
rect 296 74 326 222
rect 382 74 412 222
rect 580 124 610 252
rect 666 124 696 252
rect 770 124 800 252
rect 920 120 950 248
rect 1006 120 1036 248
rect 1092 120 1122 248
rect 1180 120 1210 248
rect 1266 120 1296 248
rect 1352 120 1382 248
rect 1452 123 1482 251
<< ndiff >>
rect 39 128 110 222
rect 39 94 51 128
rect 85 94 110 128
rect 39 74 110 94
rect 140 204 196 222
rect 140 170 151 204
rect 185 170 196 204
rect 140 120 196 170
rect 140 86 151 120
rect 185 86 196 120
rect 140 74 196 86
rect 226 128 296 222
rect 226 94 237 128
rect 271 94 296 128
rect 226 74 296 94
rect 326 204 382 222
rect 326 170 337 204
rect 371 170 382 204
rect 326 120 382 170
rect 326 86 337 120
rect 371 86 382 120
rect 326 74 382 86
rect 412 204 469 222
rect 412 170 423 204
rect 457 170 469 204
rect 412 120 469 170
rect 523 170 580 252
rect 523 136 535 170
rect 569 136 580 170
rect 523 124 580 136
rect 610 238 666 252
rect 610 204 621 238
rect 655 204 666 238
rect 610 170 666 204
rect 610 136 621 170
rect 655 136 666 170
rect 610 124 666 136
rect 696 238 770 252
rect 696 204 707 238
rect 741 204 770 238
rect 696 170 770 204
rect 696 136 707 170
rect 741 136 770 170
rect 696 124 770 136
rect 800 248 850 252
rect 1402 248 1452 251
rect 800 167 920 248
rect 800 133 875 167
rect 909 133 920 167
rect 800 124 920 133
rect 412 86 423 120
rect 457 86 469 120
rect 863 120 920 124
rect 950 235 1006 248
rect 950 201 961 235
rect 995 201 1006 235
rect 950 166 1006 201
rect 950 132 961 166
rect 995 132 1006 166
rect 950 120 1006 132
rect 1036 166 1092 248
rect 1036 132 1047 166
rect 1081 132 1092 166
rect 1036 120 1092 132
rect 1122 235 1180 248
rect 1122 201 1134 235
rect 1168 201 1180 235
rect 1122 166 1180 201
rect 1122 132 1134 166
rect 1168 132 1180 166
rect 1122 120 1180 132
rect 1210 166 1266 248
rect 1210 132 1221 166
rect 1255 132 1266 166
rect 1210 120 1266 132
rect 1296 234 1352 248
rect 1296 200 1307 234
rect 1341 200 1352 234
rect 1296 166 1352 200
rect 1296 132 1307 166
rect 1341 132 1352 166
rect 1296 120 1352 132
rect 1382 166 1452 248
rect 1382 132 1393 166
rect 1427 132 1452 166
rect 1382 123 1452 132
rect 1482 212 1539 251
rect 1482 178 1493 212
rect 1527 178 1539 212
rect 1482 123 1539 178
rect 1382 120 1432 123
rect 412 74 469 86
<< pdiff >>
rect 93 580 149 592
rect 93 546 105 580
rect 139 546 149 580
rect 93 472 149 546
rect 93 438 105 472
rect 139 438 149 472
rect 93 368 149 438
rect 185 580 239 592
rect 185 546 195 580
rect 229 546 239 580
rect 185 497 239 546
rect 185 463 195 497
rect 229 463 239 497
rect 185 414 239 463
rect 185 380 195 414
rect 229 380 239 414
rect 185 368 239 380
rect 275 580 329 592
rect 275 546 285 580
rect 319 546 329 580
rect 275 472 329 546
rect 275 438 285 472
rect 319 438 329 472
rect 275 368 329 438
rect 365 580 419 592
rect 365 546 375 580
rect 409 546 419 580
rect 365 497 419 546
rect 365 463 375 497
rect 409 463 419 497
rect 365 414 419 463
rect 365 380 375 414
rect 409 380 419 414
rect 365 368 419 380
rect 455 554 505 592
rect 762 580 818 592
rect 455 542 526 554
rect 455 508 465 542
rect 499 508 526 542
rect 455 432 526 508
rect 455 398 465 432
rect 499 398 526 432
rect 455 386 526 398
rect 562 542 616 554
rect 562 508 572 542
rect 606 508 616 542
rect 562 432 616 508
rect 562 398 572 432
rect 606 398 616 432
rect 562 386 616 398
rect 652 525 708 554
rect 652 491 662 525
rect 696 491 708 525
rect 652 386 708 491
rect 762 546 774 580
rect 808 546 818 580
rect 762 508 818 546
rect 762 474 774 508
rect 808 474 818 508
rect 455 368 511 386
rect 762 368 818 474
rect 854 578 908 592
rect 854 544 864 578
rect 898 544 908 578
rect 854 368 908 544
rect 944 424 1000 592
rect 944 390 955 424
rect 989 390 1000 424
rect 944 368 1000 390
rect 1036 578 1090 592
rect 1036 544 1046 578
rect 1080 544 1090 578
rect 1036 368 1090 544
rect 1126 580 1180 592
rect 1126 546 1136 580
rect 1170 546 1180 580
rect 1126 497 1180 546
rect 1126 463 1136 497
rect 1170 463 1180 497
rect 1126 414 1180 463
rect 1126 380 1136 414
rect 1170 380 1180 414
rect 1126 368 1180 380
rect 1216 580 1270 592
rect 1216 546 1226 580
rect 1260 546 1270 580
rect 1216 508 1270 546
rect 1216 474 1226 508
rect 1260 474 1270 508
rect 1216 368 1270 474
rect 1306 580 1368 592
rect 1306 546 1320 580
rect 1354 546 1368 580
rect 1306 368 1368 546
rect 1404 580 1468 592
rect 1404 546 1424 580
rect 1458 546 1468 580
rect 1404 508 1468 546
rect 1404 474 1424 508
rect 1458 474 1468 508
rect 1404 368 1468 474
rect 1504 580 1570 592
rect 1504 546 1524 580
rect 1558 546 1570 580
rect 1504 497 1570 546
rect 1504 463 1524 497
rect 1558 463 1570 497
rect 1504 414 1570 463
rect 1504 380 1524 414
rect 1558 380 1570 414
rect 1504 368 1570 380
<< ndiffc >>
rect 51 94 85 128
rect 151 170 185 204
rect 151 86 185 120
rect 237 94 271 128
rect 337 170 371 204
rect 337 86 371 120
rect 423 170 457 204
rect 535 136 569 170
rect 621 204 655 238
rect 621 136 655 170
rect 707 204 741 238
rect 707 136 741 170
rect 875 133 909 167
rect 423 86 457 120
rect 961 201 995 235
rect 961 132 995 166
rect 1047 132 1081 166
rect 1134 201 1168 235
rect 1134 132 1168 166
rect 1221 132 1255 166
rect 1307 200 1341 234
rect 1307 132 1341 166
rect 1393 132 1427 166
rect 1493 178 1527 212
<< pdiffc >>
rect 105 546 139 580
rect 105 438 139 472
rect 195 546 229 580
rect 195 463 229 497
rect 195 380 229 414
rect 285 546 319 580
rect 285 438 319 472
rect 375 546 409 580
rect 375 463 409 497
rect 375 380 409 414
rect 465 508 499 542
rect 465 398 499 432
rect 572 508 606 542
rect 572 398 606 432
rect 662 491 696 525
rect 774 546 808 580
rect 774 474 808 508
rect 864 544 898 578
rect 955 390 989 424
rect 1046 544 1080 578
rect 1136 546 1170 580
rect 1136 463 1170 497
rect 1136 380 1170 414
rect 1226 546 1260 580
rect 1226 474 1260 508
rect 1320 546 1354 580
rect 1424 546 1458 580
rect 1424 474 1458 508
rect 1524 546 1558 580
rect 1524 463 1558 497
rect 1524 380 1558 414
<< poly >>
rect 149 592 185 618
rect 239 592 275 618
rect 329 592 365 618
rect 419 592 455 618
rect 818 592 854 618
rect 908 592 944 618
rect 1000 592 1036 618
rect 1090 592 1126 618
rect 1180 592 1216 618
rect 1270 592 1306 618
rect 1368 592 1404 618
rect 1468 592 1504 618
rect 526 554 562 580
rect 616 554 652 580
rect 149 320 185 368
rect 239 320 275 368
rect 329 320 365 368
rect 419 320 455 368
rect 110 304 455 320
rect 110 270 133 304
rect 167 270 201 304
rect 235 270 269 304
rect 303 270 337 304
rect 371 270 405 304
rect 439 270 455 304
rect 526 318 562 386
rect 616 354 652 386
rect 616 338 722 354
rect 616 318 672 338
rect 526 304 672 318
rect 706 304 722 338
rect 526 288 722 304
rect 818 297 854 368
rect 908 336 944 368
rect 1000 336 1036 368
rect 110 254 455 270
rect 110 222 140 254
rect 196 222 226 254
rect 296 222 326 254
rect 382 222 412 254
rect 580 252 610 288
rect 666 252 696 288
rect 770 267 854 297
rect 902 320 1036 336
rect 902 286 918 320
rect 952 286 986 320
rect 1020 286 1036 320
rect 902 270 1036 286
rect 770 252 800 267
rect 920 248 950 270
rect 1006 248 1036 270
rect 1090 263 1126 368
rect 1180 263 1216 368
rect 1270 336 1306 368
rect 1368 336 1404 368
rect 1266 320 1404 336
rect 1266 286 1282 320
rect 1316 306 1404 320
rect 1316 286 1382 306
rect 1468 296 1504 368
rect 1266 270 1382 286
rect 1092 248 1122 263
rect 1180 248 1210 263
rect 1266 248 1296 270
rect 1352 248 1382 270
rect 1452 266 1504 296
rect 1452 251 1482 266
rect 580 98 610 124
rect 666 98 696 124
rect 770 102 800 124
rect 770 86 841 102
rect 920 94 950 120
rect 1006 94 1036 120
rect 110 48 140 74
rect 196 48 226 74
rect 296 48 326 74
rect 382 48 412 74
rect 770 52 791 86
rect 825 52 841 86
rect 1092 52 1122 120
rect 770 22 1122 52
rect 1180 52 1210 120
rect 1266 94 1296 120
rect 1352 94 1382 120
rect 1452 101 1482 123
rect 1452 85 1527 101
rect 1452 52 1477 85
rect 1180 51 1477 52
rect 1511 51 1527 85
rect 1180 22 1527 51
<< polycont >>
rect 133 270 167 304
rect 201 270 235 304
rect 269 270 303 304
rect 337 270 371 304
rect 405 270 439 304
rect 672 304 706 338
rect 918 286 952 320
rect 986 286 1020 320
rect 1282 286 1316 320
rect 791 52 825 86
rect 1477 51 1511 85
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 105 580 139 649
rect 25 388 71 578
rect 105 472 139 546
rect 105 422 139 438
rect 179 580 245 596
rect 179 546 195 580
rect 229 546 245 580
rect 179 497 245 546
rect 179 463 195 497
rect 229 463 245 497
rect 179 414 245 463
rect 285 580 319 649
rect 285 472 319 546
rect 285 422 319 438
rect 359 580 425 596
rect 359 546 375 580
rect 409 546 425 580
rect 359 497 425 546
rect 359 463 375 497
rect 409 463 425 497
rect 179 388 195 414
rect 25 380 195 388
rect 229 388 245 414
rect 359 414 425 463
rect 359 388 375 414
rect 229 380 375 388
rect 409 380 425 414
rect 465 542 515 649
rect 499 508 515 542
rect 465 432 515 508
rect 499 398 515 432
rect 465 382 515 398
rect 556 542 622 558
rect 556 508 572 542
rect 606 508 622 542
rect 556 432 622 508
rect 662 525 712 649
rect 696 491 712 525
rect 662 458 712 491
rect 758 580 808 596
rect 758 546 774 580
rect 758 508 808 546
rect 848 578 1096 596
rect 848 544 864 578
rect 898 544 1046 578
rect 1080 544 1096 578
rect 848 526 1096 544
rect 1136 580 1170 596
rect 758 474 774 508
rect 1136 497 1170 546
rect 808 474 1136 492
rect 758 463 1136 474
rect 758 458 1170 463
rect 1210 580 1276 596
rect 1210 546 1226 580
rect 1260 546 1276 580
rect 1210 508 1276 546
rect 1316 580 1374 649
rect 1316 546 1320 580
rect 1354 546 1374 580
rect 1316 530 1374 546
rect 1408 580 1474 596
rect 1408 546 1424 580
rect 1458 546 1474 580
rect 1210 474 1226 508
rect 1260 492 1276 508
rect 1408 508 1474 546
rect 1408 492 1424 508
rect 1260 474 1424 492
rect 1458 474 1474 508
rect 1210 458 1474 474
rect 1508 580 1574 596
rect 1508 546 1524 580
rect 1558 546 1574 580
rect 1508 497 1574 546
rect 1508 463 1524 497
rect 1558 463 1574 497
rect 556 398 572 432
rect 606 424 622 432
rect 1136 424 1170 458
rect 1508 424 1574 463
rect 606 398 955 424
rect 556 390 955 398
rect 989 390 1006 424
rect 1136 414 1574 424
rect 25 354 425 380
rect 25 220 59 354
rect 556 320 622 390
rect 1170 390 1524 414
rect 1136 364 1170 380
rect 1508 380 1524 390
rect 1558 380 1574 414
rect 1508 364 1574 380
rect 117 304 622 320
rect 117 270 133 304
rect 167 270 201 304
rect 235 270 269 304
rect 303 270 337 304
rect 371 270 405 304
rect 439 270 622 304
rect 656 338 839 356
rect 656 304 672 338
rect 706 304 839 338
rect 656 288 839 304
rect 889 320 1036 356
rect 889 286 918 320
rect 952 286 986 320
rect 1020 286 1036 320
rect 889 285 1036 286
rect 1266 320 1415 356
rect 1266 286 1282 320
rect 1316 286 1415 320
rect 1266 284 1415 286
rect 117 254 622 270
rect 588 238 655 254
rect 588 220 621 238
rect 25 204 371 220
rect 25 186 151 204
rect 135 170 151 186
rect 185 186 337 204
rect 35 128 101 152
rect 35 94 51 128
rect 85 94 101 128
rect 35 17 101 94
rect 135 120 185 170
rect 321 170 337 186
rect 135 86 151 120
rect 135 70 185 86
rect 221 128 287 152
rect 221 94 237 128
rect 271 94 287 128
rect 221 17 287 94
rect 321 120 371 170
rect 321 86 337 120
rect 321 70 371 86
rect 407 204 473 220
rect 407 170 423 204
rect 457 170 473 204
rect 407 120 473 170
rect 407 86 423 120
rect 457 86 473 120
rect 407 17 473 86
rect 519 170 585 186
rect 519 136 535 170
rect 569 136 585 170
rect 519 86 585 136
rect 621 170 655 204
rect 621 120 655 136
rect 691 251 741 254
rect 691 250 1169 251
rect 1477 250 1527 255
rect 691 238 1527 250
rect 691 204 707 238
rect 741 235 1527 238
rect 741 217 961 235
rect 691 170 741 204
rect 945 201 961 217
rect 995 217 1134 235
rect 691 136 707 170
rect 691 86 741 136
rect 875 167 909 183
rect 519 52 741 86
rect 775 86 841 134
rect 775 52 791 86
rect 825 52 841 86
rect 775 51 841 52
rect 875 17 909 133
rect 945 166 995 201
rect 1133 201 1134 217
rect 1168 234 1527 235
rect 1168 216 1307 234
rect 1168 201 1169 216
rect 945 132 961 166
rect 945 116 995 132
rect 1031 166 1097 183
rect 1031 132 1047 166
rect 1081 132 1097 166
rect 1031 17 1097 132
rect 1133 166 1169 201
rect 1291 200 1307 216
rect 1341 216 1527 234
rect 1133 132 1134 166
rect 1168 132 1169 166
rect 1133 116 1169 132
rect 1205 166 1255 182
rect 1205 132 1221 166
rect 1205 17 1255 132
rect 1291 166 1341 200
rect 1477 212 1527 216
rect 1291 132 1307 166
rect 1291 116 1341 132
rect 1377 166 1427 182
rect 1377 132 1393 166
rect 1477 178 1493 212
rect 1477 135 1527 178
rect 1377 17 1427 132
rect 1561 101 1607 134
rect 1461 85 1607 101
rect 1461 51 1477 85
rect 1511 67 1607 85
rect 1511 51 1527 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
rlabel comment s 0 0 0 0 4 o41a_4
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 B1
port 5 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 B1
port 5 nsew
flabel corelocali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 10 nsew
flabel corelocali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 10 nsew
flabel corelocali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 10 nsew
flabel corelocali s 1279 316 1313 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 1375 316 1409 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 1567 94 1601 128 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 799 94 833 128 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 A4
port 4 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 A4
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 1632 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 721824
string GDS_START 709130
<< end >>
