magic
tech sky130A
magscale 1 2
timestamp 1601050056
<< nwell >>
rect -38 332 1766 704
<< pwell >>
rect 0 0 1728 49
<< scpmos >>
rect 92 392 128 592
rect 192 392 228 592
rect 282 392 318 592
rect 372 392 408 592
rect 567 368 603 592
rect 657 368 693 592
rect 747 368 783 592
rect 837 368 873 592
rect 927 368 963 592
rect 1045 368 1081 592
rect 1135 368 1171 592
rect 1251 368 1287 592
rect 1341 368 1377 592
rect 1431 368 1467 592
rect 1521 368 1557 592
rect 1611 368 1647 592
<< nmoslvt >>
rect 130 98 160 246
rect 216 98 246 246
rect 334 98 364 246
rect 442 98 472 246
rect 560 98 590 246
rect 703 98 733 246
rect 934 74 964 222
rect 1052 74 1082 222
rect 1138 74 1168 222
rect 1256 74 1286 222
rect 1342 74 1372 222
rect 1428 74 1458 222
rect 1528 74 1558 222
rect 1614 74 1644 222
<< ndiff >>
rect 27 234 130 246
rect 27 200 35 234
rect 69 200 130 234
rect 27 144 130 200
rect 27 110 35 144
rect 69 110 130 144
rect 27 98 130 110
rect 160 234 216 246
rect 160 200 171 234
rect 205 200 216 234
rect 160 98 216 200
rect 246 98 334 246
rect 364 222 442 246
rect 364 188 386 222
rect 420 188 442 222
rect 364 98 442 188
rect 472 98 560 246
rect 590 149 703 246
rect 590 115 658 149
rect 692 115 703 149
rect 590 98 703 115
rect 733 98 823 246
rect 261 82 319 98
rect 261 48 273 82
rect 307 48 319 82
rect 487 84 545 98
rect 261 36 319 48
rect 487 50 499 84
rect 533 50 545 84
rect 748 86 823 98
rect 487 36 545 50
rect 748 52 768 86
rect 802 52 823 86
rect 877 152 934 222
rect 877 118 889 152
rect 923 118 934 152
rect 877 74 934 118
rect 964 84 1052 222
rect 964 74 991 84
rect 748 40 823 52
rect 979 50 991 74
rect 1025 74 1052 84
rect 1082 152 1138 222
rect 1082 118 1093 152
rect 1127 118 1138 152
rect 1082 74 1138 118
rect 1168 84 1256 222
rect 1168 74 1195 84
rect 1025 50 1037 74
rect 979 38 1037 50
rect 1183 50 1195 74
rect 1229 74 1256 84
rect 1286 152 1342 222
rect 1286 118 1297 152
rect 1331 118 1342 152
rect 1286 74 1342 118
rect 1372 169 1428 222
rect 1372 135 1383 169
rect 1417 135 1428 169
rect 1372 74 1428 135
rect 1458 152 1528 222
rect 1458 118 1483 152
rect 1517 118 1528 152
rect 1458 74 1528 118
rect 1558 178 1614 222
rect 1558 144 1569 178
rect 1603 144 1614 178
rect 1558 74 1614 144
rect 1644 152 1701 222
rect 1644 118 1655 152
rect 1689 118 1701 152
rect 1644 74 1701 118
rect 1229 50 1241 74
rect 1183 38 1241 50
<< pdiff >>
rect 978 627 1030 639
rect 978 593 987 627
rect 1021 593 1030 627
rect 1186 627 1236 639
rect 978 592 1030 593
rect 1186 593 1194 627
rect 1228 593 1236 627
rect 1186 592 1236 593
rect 36 580 92 592
rect 36 546 48 580
rect 82 546 92 580
rect 36 509 92 546
rect 36 475 48 509
rect 82 475 92 509
rect 36 438 92 475
rect 36 404 48 438
rect 82 404 92 438
rect 36 392 92 404
rect 128 580 192 592
rect 128 546 138 580
rect 172 546 192 580
rect 128 502 192 546
rect 128 468 138 502
rect 172 468 192 502
rect 128 392 192 468
rect 228 580 282 592
rect 228 546 238 580
rect 272 546 282 580
rect 228 509 282 546
rect 228 475 238 509
rect 272 475 282 509
rect 228 438 282 475
rect 228 404 238 438
rect 272 404 282 438
rect 228 392 282 404
rect 318 531 372 592
rect 318 497 328 531
rect 362 497 372 531
rect 318 438 372 497
rect 318 404 328 438
rect 362 404 372 438
rect 318 392 372 404
rect 408 580 460 592
rect 408 546 418 580
rect 452 546 460 580
rect 408 488 460 546
rect 408 454 418 488
rect 452 454 460 488
rect 408 392 460 454
rect 514 580 567 592
rect 514 546 523 580
rect 557 546 567 580
rect 514 488 567 546
rect 514 454 523 488
rect 557 454 567 488
rect 514 368 567 454
rect 603 547 657 592
rect 603 513 613 547
rect 647 513 657 547
rect 603 472 657 513
rect 603 438 613 472
rect 647 438 657 472
rect 603 368 657 438
rect 693 577 747 592
rect 693 543 703 577
rect 737 543 747 577
rect 693 368 747 543
rect 783 519 837 592
rect 783 485 793 519
rect 827 485 837 519
rect 783 368 837 485
rect 873 577 927 592
rect 873 543 883 577
rect 917 543 927 577
rect 873 368 927 543
rect 963 368 1045 592
rect 1081 577 1135 592
rect 1081 543 1091 577
rect 1125 543 1135 577
rect 1081 368 1135 543
rect 1171 368 1251 592
rect 1287 580 1341 592
rect 1287 546 1297 580
rect 1331 546 1341 580
rect 1287 508 1341 546
rect 1287 474 1297 508
rect 1331 474 1341 508
rect 1287 368 1341 474
rect 1377 578 1431 592
rect 1377 544 1387 578
rect 1421 544 1431 578
rect 1377 368 1431 544
rect 1467 580 1521 592
rect 1467 546 1477 580
rect 1511 546 1521 580
rect 1467 508 1521 546
rect 1467 474 1477 508
rect 1511 474 1521 508
rect 1467 368 1521 474
rect 1557 578 1611 592
rect 1557 544 1567 578
rect 1601 544 1611 578
rect 1557 368 1611 544
rect 1647 580 1701 592
rect 1647 546 1657 580
rect 1691 546 1701 580
rect 1647 508 1701 546
rect 1647 474 1657 508
rect 1691 474 1701 508
rect 1647 368 1701 474
<< ndiffc >>
rect 35 200 69 234
rect 35 110 69 144
rect 171 200 205 234
rect 386 188 420 222
rect 658 115 692 149
rect 273 48 307 82
rect 499 50 533 84
rect 768 52 802 86
rect 889 118 923 152
rect 991 50 1025 84
rect 1093 118 1127 152
rect 1195 50 1229 84
rect 1297 118 1331 152
rect 1383 135 1417 169
rect 1483 118 1517 152
rect 1569 144 1603 178
rect 1655 118 1689 152
<< pdiffc >>
rect 987 593 1021 627
rect 1194 593 1228 627
rect 48 546 82 580
rect 48 475 82 509
rect 48 404 82 438
rect 138 546 172 580
rect 138 468 172 502
rect 238 546 272 580
rect 238 475 272 509
rect 238 404 272 438
rect 328 497 362 531
rect 328 404 362 438
rect 418 546 452 580
rect 418 454 452 488
rect 523 546 557 580
rect 523 454 557 488
rect 613 513 647 547
rect 613 438 647 472
rect 703 543 737 577
rect 793 485 827 519
rect 883 543 917 577
rect 1091 543 1125 577
rect 1297 546 1331 580
rect 1297 474 1331 508
rect 1387 544 1421 578
rect 1477 546 1511 580
rect 1477 474 1511 508
rect 1567 544 1601 578
rect 1657 546 1691 580
rect 1657 474 1691 508
<< poly >>
rect 92 592 128 618
rect 192 592 228 618
rect 282 592 318 618
rect 372 592 408 618
rect 567 592 603 618
rect 657 592 693 618
rect 747 592 783 618
rect 837 592 873 618
rect 927 592 963 618
rect 1045 592 1081 618
rect 1135 592 1171 618
rect 1251 592 1287 618
rect 1341 592 1377 618
rect 1431 592 1467 618
rect 1521 592 1557 618
rect 1611 592 1647 618
rect 92 350 128 392
rect 192 350 228 392
rect 282 362 318 392
rect 88 334 228 350
rect 88 300 104 334
rect 138 300 172 334
rect 206 314 228 334
rect 288 358 318 362
rect 372 369 408 392
rect 372 358 472 369
rect 288 344 472 358
rect 206 300 246 314
rect 88 284 246 300
rect 288 310 422 344
rect 456 310 472 344
rect 567 336 603 368
rect 657 336 693 368
rect 747 336 783 368
rect 837 336 873 368
rect 927 336 963 368
rect 1045 336 1081 368
rect 1135 336 1171 368
rect 288 294 472 310
rect 130 246 160 284
rect 216 246 246 284
rect 334 246 364 294
rect 442 246 472 294
rect 517 320 873 336
rect 517 286 533 320
rect 567 286 601 320
rect 635 286 669 320
rect 703 306 873 320
rect 921 324 1171 336
rect 1251 324 1287 368
rect 921 320 1287 324
rect 703 286 733 306
rect 517 270 733 286
rect 921 286 937 320
rect 971 286 1005 320
rect 1039 286 1073 320
rect 1107 286 1287 320
rect 921 270 1287 286
rect 560 246 590 270
rect 703 246 733 270
rect 934 222 964 270
rect 1052 222 1082 270
rect 1138 222 1168 270
rect 1256 222 1286 270
rect 1341 237 1377 368
rect 1431 336 1467 368
rect 1521 336 1557 368
rect 1611 336 1647 368
rect 1431 320 1647 336
rect 1431 286 1447 320
rect 1481 286 1515 320
rect 1549 286 1583 320
rect 1617 286 1647 320
rect 1431 270 1647 286
rect 1431 267 1461 270
rect 1428 237 1461 267
rect 1342 222 1372 237
rect 1428 222 1458 237
rect 1528 222 1558 270
rect 1614 222 1644 270
rect 130 72 160 98
rect 216 72 246 98
rect 334 72 364 98
rect 442 72 472 98
rect 560 72 590 98
rect 703 72 733 98
rect 934 48 964 74
rect 1052 48 1082 74
rect 1138 48 1168 74
rect 1256 48 1286 74
rect 1342 59 1372 74
rect 1428 59 1458 74
rect 1342 29 1458 59
rect 1528 48 1558 74
rect 1614 48 1644 74
<< polycont >>
rect 104 300 138 334
rect 172 300 206 334
rect 422 310 456 344
rect 533 286 567 320
rect 601 286 635 320
rect 669 286 703 320
rect 937 286 971 320
rect 1005 286 1039 320
rect 1073 286 1107 320
rect 1447 286 1481 320
rect 1515 286 1549 320
rect 1583 286 1617 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 32 580 98 596
rect 32 546 48 580
rect 82 546 98 580
rect 32 509 98 546
rect 32 475 48 509
rect 82 475 98 509
rect 32 438 98 475
rect 138 580 188 649
rect 971 627 1037 649
rect 172 546 188 580
rect 138 502 188 546
rect 172 468 188 502
rect 138 452 188 468
rect 222 581 468 615
rect 222 580 272 581
rect 222 546 238 580
rect 402 580 468 581
rect 222 509 272 546
rect 222 475 238 509
rect 32 404 48 438
rect 82 418 98 438
rect 222 438 272 475
rect 222 418 238 438
rect 82 404 238 418
rect 32 384 272 404
rect 312 531 362 547
rect 312 497 328 531
rect 312 438 362 497
rect 402 546 418 580
rect 452 546 468 580
rect 402 488 468 546
rect 402 454 418 488
rect 452 454 468 488
rect 402 438 468 454
rect 507 581 933 615
rect 971 593 987 627
rect 1021 593 1037 627
rect 1178 627 1244 649
rect 507 580 557 581
rect 507 546 523 580
rect 703 577 737 581
rect 507 488 557 546
rect 507 454 523 488
rect 507 438 557 454
rect 597 513 613 547
rect 647 513 663 547
rect 883 577 933 581
rect 703 525 737 543
rect 597 491 663 513
rect 777 519 843 547
rect 917 559 933 577
rect 1075 577 1141 596
rect 1178 593 1194 627
rect 1228 593 1244 627
rect 1075 559 1091 577
rect 917 543 1091 559
rect 1125 559 1141 577
rect 1297 580 1331 596
rect 1125 546 1297 559
rect 1125 543 1331 546
rect 883 525 1331 543
rect 1371 578 1421 649
rect 1371 544 1387 578
rect 1371 526 1421 544
rect 1461 580 1527 596
rect 1461 546 1477 580
rect 1511 546 1527 580
rect 777 491 793 519
rect 597 485 793 491
rect 827 491 843 519
rect 1297 508 1331 525
rect 827 485 1263 491
rect 597 472 1263 485
rect 597 438 613 472
rect 647 457 1263 472
rect 1461 508 1527 546
rect 1567 578 1601 649
rect 1567 526 1601 544
rect 1641 580 1707 596
rect 1641 546 1657 580
rect 1691 546 1707 580
rect 1461 492 1477 508
rect 1331 474 1477 492
rect 1511 492 1527 508
rect 1641 508 1707 546
rect 1641 492 1657 508
rect 1511 474 1657 492
rect 1691 474 1707 508
rect 1297 458 1707 474
rect 647 438 663 457
rect 312 404 328 438
rect 1229 424 1263 457
rect 697 404 1195 423
rect 88 334 222 350
rect 88 300 104 334
rect 138 300 172 334
rect 206 300 222 334
rect 88 284 222 300
rect 19 234 69 250
rect 19 200 35 234
rect 19 144 69 200
rect 19 110 35 144
rect 103 150 137 284
rect 171 238 221 250
rect 312 238 362 404
rect 406 389 1195 404
rect 1229 390 1701 424
rect 406 370 731 389
rect 406 344 472 370
rect 1161 356 1195 389
rect 406 310 422 344
rect 456 310 472 344
rect 406 294 472 310
rect 506 320 719 336
rect 506 286 533 320
rect 567 286 601 320
rect 635 286 669 320
rect 703 286 719 320
rect 793 320 1127 355
rect 793 304 937 320
rect 506 272 719 286
rect 753 286 937 304
rect 971 286 1005 320
rect 1039 286 1073 320
rect 1107 286 1127 320
rect 1161 320 1633 356
rect 1161 310 1447 320
rect 506 238 540 272
rect 753 270 1127 286
rect 1177 286 1447 310
rect 1481 286 1515 320
rect 1549 286 1583 320
rect 1617 286 1633 320
rect 1177 270 1633 286
rect 753 238 787 270
rect 171 234 540 238
rect 205 222 540 234
rect 205 200 386 222
rect 171 188 386 200
rect 420 188 540 222
rect 574 204 787 238
rect 1667 236 1701 390
rect 171 184 221 188
rect 574 154 608 204
rect 821 202 1701 236
rect 821 170 855 202
rect 255 150 608 154
rect 103 120 608 150
rect 642 149 855 170
rect 1367 169 1433 202
rect 103 116 289 120
rect 19 17 69 110
rect 642 115 658 149
rect 692 136 855 149
rect 889 152 1331 168
rect 692 115 708 136
rect 642 94 708 115
rect 923 134 1093 152
rect 923 118 939 134
rect 744 86 827 102
rect 483 84 549 86
rect 257 48 273 82
rect 307 48 323 82
rect 257 17 323 48
rect 483 50 499 84
rect 533 50 549 84
rect 483 17 549 50
rect 744 52 768 86
rect 802 52 827 86
rect 889 70 939 118
rect 1077 118 1093 134
rect 1127 134 1297 152
rect 1127 118 1143 134
rect 975 84 1041 100
rect 744 17 827 52
rect 975 50 991 84
rect 1025 50 1041 84
rect 1077 70 1143 118
rect 1281 118 1297 134
rect 1367 135 1383 169
rect 1417 135 1433 169
rect 1569 178 1603 202
rect 1367 119 1433 135
rect 1467 152 1533 168
rect 1179 84 1245 100
rect 975 17 1041 50
rect 1179 50 1195 84
rect 1229 50 1245 84
rect 1281 85 1331 118
rect 1467 118 1483 152
rect 1517 118 1533 152
rect 1569 119 1603 144
rect 1639 152 1705 168
rect 1467 85 1533 118
rect 1639 118 1655 152
rect 1689 118 1705 152
rect 1639 85 1705 118
rect 1281 51 1705 85
rect 1179 17 1245 50
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
<< metal1 >>
rect 0 683 1728 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 0 617 1728 649
rect 0 17 1728 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
rect 0 -49 1728 -17
<< labels >>
flabel pwell s 0 0 1728 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 0 617 1728 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
rlabel comment s 0 0 0 0 4 xor2_4
flabel metal1 s 0 617 1728 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 1728 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 1183 316 1217 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 1279 316 1313 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 1375 316 1409 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 1471 316 1505 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 1567 316 1601 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 799 464 833 498 0 FreeSans 340 0 0 0 X
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 1728 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 558948
string GDS_START 546588
<< end >>
