magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 113 364 187 430
rect 145 230 187 364
rect 123 66 187 230
rect 289 270 355 356
rect 403 270 469 356
rect 505 270 583 356
rect 631 270 743 356
rect 777 260 843 356
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 23 532 89 649
rect 220 532 302 649
rect 45 464 255 498
rect 45 330 79 464
rect 45 264 111 330
rect 23 17 89 226
rect 221 424 255 464
rect 343 492 409 572
rect 453 526 529 649
rect 575 581 841 615
rect 575 492 641 581
rect 343 458 641 492
rect 675 424 741 547
rect 221 390 741 424
rect 775 390 841 581
rect 221 236 255 390
rect 221 202 621 236
rect 237 17 303 168
rect 555 70 621 202
rect 770 17 836 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel locali s 505 270 583 356 6 A1
port 1 nsew signal input
rlabel locali s 403 270 469 356 6 A2
port 2 nsew signal input
rlabel locali s 289 270 355 356 6 A3
port 3 nsew signal input
rlabel locali s 631 270 743 356 6 B1
port 4 nsew signal input
rlabel locali s 777 260 843 356 6 B2
port 5 nsew signal input
rlabel locali s 145 230 187 364 6 X
port 6 nsew signal output
rlabel locali s 123 66 187 230 6 X
port 6 nsew signal output
rlabel locali s 113 364 187 430 6 X
port 6 nsew signal output
rlabel metal1 s 0 -49 864 49 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 617 864 715 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3719660
string GDS_START 3712684
<< end >>
