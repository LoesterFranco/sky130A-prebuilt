magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 736 561
rect 115 359 165 527
rect 567 325 609 425
rect 475 257 528 325
rect 567 291 719 325
rect 27 215 193 257
rect 227 215 437 257
rect 475 215 593 257
rect 627 181 719 291
rect 18 17 73 181
rect 107 145 719 181
rect 107 51 173 145
rect 207 17 241 111
rect 275 51 341 145
rect 375 17 517 111
rect 551 51 617 145
rect 651 17 709 111
rect 0 -17 736 17
<< obsli1 >>
rect 30 325 81 493
rect 199 325 249 493
rect 283 459 693 493
rect 283 359 333 459
rect 367 325 417 425
rect 483 359 525 459
rect 643 359 693 459
rect 30 291 417 325
<< metal1 >>
rect 0 496 736 592
rect 0 -48 736 48
<< labels >>
rlabel locali s 27 215 193 257 6 A
port 1 nsew signal input
rlabel locali s 227 215 437 257 6 B
port 2 nsew signal input
rlabel locali s 475 257 528 325 6 C
port 3 nsew signal input
rlabel locali s 475 215 593 257 6 C
port 3 nsew signal input
rlabel locali s 627 181 719 291 6 Y
port 4 nsew signal output
rlabel locali s 567 325 609 425 6 Y
port 4 nsew signal output
rlabel locali s 567 291 719 325 6 Y
port 4 nsew signal output
rlabel locali s 551 51 617 145 6 Y
port 4 nsew signal output
rlabel locali s 275 51 341 145 6 Y
port 4 nsew signal output
rlabel locali s 107 145 719 181 6 Y
port 4 nsew signal output
rlabel locali s 107 51 173 145 6 Y
port 4 nsew signal output
rlabel locali s 651 17 709 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 375 17 517 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 207 17 241 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 18 17 73 181 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 736 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 736 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 115 359 165 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 736 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 736 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1979216
string GDS_START 1972668
<< end >>
