magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 2054 704
<< pwell >>
rect 0 0 2016 49
<< scnmos >>
rect 184 74 214 222
rect 273 74 303 222
rect 375 74 405 222
rect 475 74 505 222
rect 561 74 591 222
rect 675 74 705 222
rect 761 74 791 222
rect 956 74 986 222
rect 1042 74 1072 222
rect 1225 74 1255 222
rect 1325 74 1355 222
rect 1425 74 1455 222
rect 1511 74 1541 222
rect 1630 74 1660 222
rect 1716 74 1746 222
rect 1802 74 1832 222
rect 1888 74 1918 222
<< pmoshvt >>
rect 86 424 116 592
rect 176 424 206 592
rect 378 368 408 592
rect 468 368 498 592
rect 568 368 598 592
rect 658 368 688 592
rect 748 368 778 592
rect 848 368 878 592
rect 953 368 983 592
rect 1048 368 1078 592
rect 1250 368 1280 592
rect 1350 368 1380 592
rect 1450 368 1480 592
rect 1540 368 1570 592
rect 1630 368 1660 592
rect 1720 368 1750 592
rect 1810 368 1840 592
rect 1900 368 1930 592
<< ndiff >>
rect 134 146 184 222
rect 47 134 184 146
rect 47 100 71 134
rect 105 100 139 134
rect 173 100 184 134
rect 47 88 184 100
rect 134 74 184 88
rect 214 210 273 222
rect 214 176 228 210
rect 262 176 273 210
rect 214 120 273 176
rect 214 86 228 120
rect 262 86 273 120
rect 214 74 273 86
rect 303 210 375 222
rect 303 176 330 210
rect 364 176 375 210
rect 303 120 375 176
rect 303 86 330 120
rect 364 86 375 120
rect 303 74 375 86
rect 405 142 475 222
rect 405 108 416 142
rect 450 108 475 142
rect 405 74 475 108
rect 505 210 561 222
rect 505 176 516 210
rect 550 176 561 210
rect 505 120 561 176
rect 505 86 516 120
rect 550 86 561 120
rect 505 74 561 86
rect 591 210 675 222
rect 591 176 616 210
rect 650 176 675 210
rect 591 120 675 176
rect 591 86 616 120
rect 650 86 675 120
rect 591 74 675 86
rect 705 210 761 222
rect 705 176 716 210
rect 750 176 761 210
rect 705 120 761 176
rect 705 86 716 120
rect 750 86 761 120
rect 705 74 761 86
rect 791 152 956 222
rect 791 118 802 152
rect 836 118 911 152
rect 945 118 956 152
rect 791 74 956 118
rect 986 210 1042 222
rect 986 176 997 210
rect 1031 176 1042 210
rect 986 120 1042 176
rect 986 86 997 120
rect 1031 86 1042 120
rect 986 74 1042 86
rect 1072 152 1225 222
rect 1072 118 1083 152
rect 1117 118 1180 152
rect 1214 118 1225 152
rect 1072 74 1225 118
rect 1255 210 1325 222
rect 1255 176 1266 210
rect 1300 176 1325 210
rect 1255 120 1325 176
rect 1255 86 1266 120
rect 1300 86 1325 120
rect 1255 74 1325 86
rect 1355 145 1425 222
rect 1355 111 1366 145
rect 1400 111 1425 145
rect 1355 74 1425 111
rect 1455 210 1511 222
rect 1455 176 1466 210
rect 1500 176 1511 210
rect 1455 120 1511 176
rect 1455 86 1466 120
rect 1500 86 1511 120
rect 1455 74 1511 86
rect 1541 145 1630 222
rect 1541 111 1568 145
rect 1602 111 1630 145
rect 1541 74 1630 111
rect 1660 210 1716 222
rect 1660 176 1671 210
rect 1705 176 1716 210
rect 1660 120 1716 176
rect 1660 86 1671 120
rect 1705 86 1716 120
rect 1660 74 1716 86
rect 1746 145 1802 222
rect 1746 111 1757 145
rect 1791 111 1802 145
rect 1746 74 1802 111
rect 1832 210 1888 222
rect 1832 176 1843 210
rect 1877 176 1888 210
rect 1832 120 1888 176
rect 1832 86 1843 120
rect 1877 86 1888 120
rect 1832 74 1888 86
rect 1918 210 1989 222
rect 1918 176 1943 210
rect 1977 176 1989 210
rect 1918 120 1989 176
rect 1918 86 1943 120
rect 1977 86 1989 120
rect 1918 74 1989 86
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 470 86 546
rect 27 436 39 470
rect 73 436 86 470
rect 27 424 86 436
rect 116 580 176 592
rect 116 546 129 580
rect 163 546 176 580
rect 116 470 176 546
rect 116 436 129 470
rect 163 436 176 470
rect 116 424 176 436
rect 206 575 265 592
rect 206 541 219 575
rect 253 541 265 575
rect 206 470 265 541
rect 206 436 219 470
rect 253 436 265 470
rect 206 424 265 436
rect 319 580 378 592
rect 319 546 331 580
rect 365 546 378 580
rect 319 497 378 546
rect 319 463 331 497
rect 365 463 378 497
rect 319 414 378 463
rect 319 380 331 414
rect 365 380 378 414
rect 319 368 378 380
rect 408 547 468 592
rect 408 513 421 547
rect 455 513 468 547
rect 408 479 468 513
rect 408 445 421 479
rect 455 445 468 479
rect 408 411 468 445
rect 408 377 421 411
rect 455 377 468 411
rect 408 368 468 377
rect 498 584 568 592
rect 498 550 515 584
rect 549 550 568 584
rect 498 482 568 550
rect 498 448 515 482
rect 549 448 568 482
rect 498 368 568 448
rect 598 547 658 592
rect 598 513 611 547
rect 645 513 658 547
rect 598 479 658 513
rect 598 445 611 479
rect 645 445 658 479
rect 598 411 658 445
rect 598 377 611 411
rect 645 377 658 411
rect 598 368 658 377
rect 688 584 748 592
rect 688 550 701 584
rect 735 550 748 584
rect 688 514 748 550
rect 688 480 701 514
rect 735 480 748 514
rect 688 368 748 480
rect 778 573 848 592
rect 778 539 801 573
rect 835 539 848 573
rect 778 368 848 539
rect 878 519 953 592
rect 878 485 901 519
rect 935 485 953 519
rect 878 368 953 485
rect 983 570 1048 592
rect 983 536 1001 570
rect 1035 536 1048 570
rect 983 368 1048 536
rect 1078 492 1137 592
rect 1078 458 1091 492
rect 1125 458 1137 492
rect 1078 368 1137 458
rect 1191 531 1250 592
rect 1191 497 1203 531
rect 1237 497 1250 531
rect 1191 424 1250 497
rect 1191 390 1203 424
rect 1237 390 1250 424
rect 1191 368 1250 390
rect 1280 580 1350 592
rect 1280 546 1303 580
rect 1337 546 1350 580
rect 1280 508 1350 546
rect 1280 474 1303 508
rect 1337 474 1350 508
rect 1280 368 1350 474
rect 1380 531 1450 592
rect 1380 497 1403 531
rect 1437 497 1450 531
rect 1380 424 1450 497
rect 1380 390 1403 424
rect 1437 390 1450 424
rect 1380 368 1450 390
rect 1480 576 1540 592
rect 1480 542 1493 576
rect 1527 542 1540 576
rect 1480 508 1540 542
rect 1480 474 1493 508
rect 1527 474 1540 508
rect 1480 368 1540 474
rect 1570 580 1630 592
rect 1570 546 1583 580
rect 1617 546 1630 580
rect 1570 505 1630 546
rect 1570 471 1583 505
rect 1617 471 1630 505
rect 1570 424 1630 471
rect 1570 390 1583 424
rect 1617 390 1630 424
rect 1570 368 1630 390
rect 1660 580 1720 592
rect 1660 546 1673 580
rect 1707 546 1720 580
rect 1660 508 1720 546
rect 1660 474 1673 508
rect 1707 474 1720 508
rect 1660 368 1720 474
rect 1750 580 1810 592
rect 1750 546 1763 580
rect 1797 546 1810 580
rect 1750 505 1810 546
rect 1750 471 1763 505
rect 1797 471 1810 505
rect 1750 424 1810 471
rect 1750 390 1763 424
rect 1797 390 1810 424
rect 1750 368 1810 390
rect 1840 580 1900 592
rect 1840 546 1853 580
rect 1887 546 1900 580
rect 1840 508 1900 546
rect 1840 474 1853 508
rect 1887 474 1900 508
rect 1840 368 1900 474
rect 1930 580 1989 592
rect 1930 546 1943 580
rect 1977 546 1989 580
rect 1930 497 1989 546
rect 1930 463 1943 497
rect 1977 463 1989 497
rect 1930 414 1989 463
rect 1930 380 1943 414
rect 1977 380 1989 414
rect 1930 368 1989 380
<< ndiffc >>
rect 71 100 105 134
rect 139 100 173 134
rect 228 176 262 210
rect 228 86 262 120
rect 330 176 364 210
rect 330 86 364 120
rect 416 108 450 142
rect 516 176 550 210
rect 516 86 550 120
rect 616 176 650 210
rect 616 86 650 120
rect 716 176 750 210
rect 716 86 750 120
rect 802 118 836 152
rect 911 118 945 152
rect 997 176 1031 210
rect 997 86 1031 120
rect 1083 118 1117 152
rect 1180 118 1214 152
rect 1266 176 1300 210
rect 1266 86 1300 120
rect 1366 111 1400 145
rect 1466 176 1500 210
rect 1466 86 1500 120
rect 1568 111 1602 145
rect 1671 176 1705 210
rect 1671 86 1705 120
rect 1757 111 1791 145
rect 1843 176 1877 210
rect 1843 86 1877 120
rect 1943 176 1977 210
rect 1943 86 1977 120
<< pdiffc >>
rect 39 546 73 580
rect 39 436 73 470
rect 129 546 163 580
rect 129 436 163 470
rect 219 541 253 575
rect 219 436 253 470
rect 331 546 365 580
rect 331 463 365 497
rect 331 380 365 414
rect 421 513 455 547
rect 421 445 455 479
rect 421 377 455 411
rect 515 550 549 584
rect 515 448 549 482
rect 611 513 645 547
rect 611 445 645 479
rect 611 377 645 411
rect 701 550 735 584
rect 701 480 735 514
rect 801 539 835 573
rect 901 485 935 519
rect 1001 536 1035 570
rect 1091 458 1125 492
rect 1203 497 1237 531
rect 1203 390 1237 424
rect 1303 546 1337 580
rect 1303 474 1337 508
rect 1403 497 1437 531
rect 1403 390 1437 424
rect 1493 542 1527 576
rect 1493 474 1527 508
rect 1583 546 1617 580
rect 1583 471 1617 505
rect 1583 390 1617 424
rect 1673 546 1707 580
rect 1673 474 1707 508
rect 1763 546 1797 580
rect 1763 471 1797 505
rect 1763 390 1797 424
rect 1853 546 1887 580
rect 1853 474 1887 508
rect 1943 546 1977 580
rect 1943 463 1977 497
rect 1943 380 1977 414
<< poly >>
rect 86 592 116 618
rect 176 592 206 618
rect 378 592 408 618
rect 468 592 498 618
rect 568 592 598 618
rect 658 592 688 618
rect 748 592 778 618
rect 848 592 878 618
rect 953 592 983 618
rect 1048 592 1078 618
rect 1250 592 1280 618
rect 1350 592 1380 618
rect 1450 592 1480 618
rect 1540 592 1570 618
rect 1630 592 1660 618
rect 1720 592 1750 618
rect 1810 592 1840 618
rect 1900 592 1930 618
rect 86 409 116 424
rect 176 409 206 424
rect 83 386 119 409
rect 44 377 119 386
rect 173 377 209 409
rect 44 370 209 377
rect 44 336 60 370
rect 94 336 209 370
rect 378 353 408 368
rect 468 353 498 368
rect 568 353 598 368
rect 658 353 688 368
rect 748 353 778 368
rect 848 353 878 368
rect 953 353 983 368
rect 1048 353 1078 368
rect 1250 353 1280 368
rect 1350 353 1380 368
rect 1450 353 1480 368
rect 1540 353 1570 368
rect 1630 353 1660 368
rect 1720 353 1750 368
rect 1810 353 1840 368
rect 1900 353 1930 368
rect 375 345 411 353
rect 465 345 501 353
rect 565 345 601 353
rect 655 345 691 353
rect 44 302 209 336
rect 44 268 60 302
rect 94 268 209 302
rect 44 267 209 268
rect 264 315 691 345
rect 745 336 781 353
rect 845 336 881 353
rect 950 336 986 353
rect 745 320 986 336
rect 264 314 591 315
rect 264 280 280 314
rect 314 280 348 314
rect 382 280 416 314
rect 450 280 591 314
rect 44 237 214 267
rect 264 264 591 280
rect 745 286 800 320
rect 834 286 868 320
rect 902 286 936 320
rect 970 286 986 320
rect 745 267 986 286
rect 1045 267 1081 353
rect 1247 336 1283 353
rect 1347 336 1383 353
rect 1447 336 1483 353
rect 1537 336 1573 353
rect 44 234 119 237
rect 44 200 60 234
rect 94 200 119 234
rect 184 222 214 237
rect 273 222 303 264
rect 375 222 405 264
rect 475 222 505 264
rect 561 222 591 264
rect 675 237 1081 267
rect 1225 320 1573 336
rect 1225 286 1241 320
rect 1275 286 1309 320
rect 1343 286 1377 320
rect 1411 286 1445 320
rect 1479 286 1573 320
rect 1627 336 1663 353
rect 1717 336 1753 353
rect 1807 336 1843 353
rect 1897 336 1933 353
rect 1627 320 1933 336
rect 1627 300 1646 320
rect 1225 270 1573 286
rect 1630 286 1646 300
rect 1680 286 1714 320
rect 1748 286 1782 320
rect 1816 286 1850 320
rect 1884 286 1933 320
rect 1630 270 1933 286
rect 675 222 705 237
rect 761 222 791 237
rect 956 222 986 237
rect 1042 222 1072 237
rect 1225 222 1255 270
rect 1325 222 1355 270
rect 1425 222 1455 270
rect 1511 222 1541 270
rect 1630 222 1660 270
rect 1716 222 1746 270
rect 1802 222 1832 270
rect 1888 222 1918 270
rect 44 184 119 200
rect 184 48 214 74
rect 273 48 303 74
rect 375 48 405 74
rect 475 48 505 74
rect 561 48 591 74
rect 675 48 705 74
rect 761 48 791 74
rect 956 48 986 74
rect 1042 48 1072 74
rect 1225 48 1255 74
rect 1325 48 1355 74
rect 1425 48 1455 74
rect 1511 48 1541 74
rect 1630 48 1660 74
rect 1716 48 1746 74
rect 1802 48 1832 74
rect 1888 48 1918 74
<< polycont >>
rect 60 336 94 370
rect 60 268 94 302
rect 280 280 314 314
rect 348 280 382 314
rect 416 280 450 314
rect 800 286 834 320
rect 868 286 902 320
rect 936 286 970 320
rect 60 200 94 234
rect 1241 286 1275 320
rect 1309 286 1343 320
rect 1377 286 1411 320
rect 1445 286 1479 320
rect 1646 286 1680 320
rect 1714 286 1748 320
rect 1782 286 1816 320
rect 1850 286 1884 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 23 580 73 649
rect 23 546 39 580
rect 23 470 73 546
rect 23 436 39 470
rect 23 420 73 436
rect 113 580 179 596
rect 113 546 129 580
rect 163 546 179 580
rect 113 470 179 546
rect 113 436 129 470
rect 163 436 179 470
rect 113 420 179 436
rect 215 575 269 649
rect 215 541 219 575
rect 253 541 269 575
rect 215 470 269 541
rect 215 436 219 470
rect 253 436 269 470
rect 215 420 269 436
rect 315 584 751 615
rect 315 581 515 584
rect 315 580 365 581
rect 315 546 331 580
rect 505 550 515 581
rect 549 581 701 584
rect 549 550 561 581
rect 315 497 365 546
rect 315 463 331 497
rect 25 370 110 386
rect 25 336 60 370
rect 94 336 110 370
rect 25 302 110 336
rect 25 268 60 302
rect 94 268 110 302
rect 25 234 110 268
rect 25 200 60 234
rect 94 200 110 234
rect 25 184 110 200
rect 144 330 178 420
rect 315 414 365 463
rect 315 380 331 414
rect 315 364 365 380
rect 405 513 421 547
rect 455 513 471 547
rect 405 479 471 513
rect 405 445 421 479
rect 455 445 471 479
rect 405 411 471 445
rect 505 482 561 550
rect 695 550 701 581
rect 735 550 751 584
rect 505 448 515 482
rect 549 448 561 482
rect 505 432 561 448
rect 595 513 611 547
rect 645 513 661 547
rect 595 479 661 513
rect 595 445 611 479
rect 645 445 661 479
rect 695 514 751 550
rect 785 581 1543 615
rect 785 573 851 581
rect 785 539 801 573
rect 835 539 851 573
rect 985 570 1051 581
rect 785 532 851 539
rect 695 480 701 514
rect 735 498 751 514
rect 885 519 951 544
rect 985 536 1001 570
rect 1035 536 1051 570
rect 1287 580 1353 581
rect 985 526 1051 536
rect 1187 531 1253 547
rect 885 498 901 519
rect 735 485 901 498
rect 935 492 951 519
rect 1088 492 1141 508
rect 935 485 1091 492
rect 735 480 1091 485
rect 695 464 1091 480
rect 885 458 1091 464
rect 1125 458 1141 492
rect 1187 497 1203 531
rect 1237 497 1253 531
rect 405 377 421 411
rect 455 398 471 411
rect 595 424 661 445
rect 1187 424 1253 497
rect 1287 546 1303 580
rect 1337 546 1353 580
rect 1493 576 1543 581
rect 1287 508 1353 546
rect 1287 474 1303 508
rect 1337 474 1353 508
rect 1287 458 1353 474
rect 1387 531 1453 547
rect 1387 497 1403 531
rect 1437 497 1453 531
rect 1387 424 1453 497
rect 1527 542 1543 576
rect 1493 508 1543 542
rect 1527 474 1543 508
rect 1493 458 1543 474
rect 1577 580 1623 596
rect 1577 546 1583 580
rect 1617 546 1623 580
rect 1577 505 1623 546
rect 1577 471 1583 505
rect 1617 471 1623 505
rect 1577 424 1623 471
rect 1657 580 1707 649
rect 1657 546 1673 580
rect 1657 508 1707 546
rect 1657 474 1673 508
rect 1657 458 1707 474
rect 1747 580 1813 596
rect 1747 546 1763 580
rect 1797 546 1813 580
rect 1747 505 1813 546
rect 1747 471 1763 505
rect 1797 471 1813 505
rect 1747 424 1813 471
rect 1853 580 1903 649
rect 1887 546 1903 580
rect 1853 508 1903 546
rect 1887 474 1903 508
rect 1853 458 1903 474
rect 1943 580 1993 596
rect 1977 546 1993 580
rect 1943 497 1993 546
rect 1977 463 1993 497
rect 1943 424 1993 463
rect 595 411 1127 424
rect 595 398 611 411
rect 455 377 611 398
rect 645 390 1127 411
rect 1187 390 1203 424
rect 1237 390 1403 424
rect 1437 390 1583 424
rect 1617 390 1763 424
rect 1797 414 1993 424
rect 1797 390 1943 414
rect 645 377 661 390
rect 405 364 661 377
rect 144 314 466 330
rect 144 280 280 314
rect 314 280 348 314
rect 382 280 416 314
rect 450 280 466 314
rect 784 320 1031 356
rect 144 264 466 280
rect 144 150 178 264
rect 500 260 750 294
rect 784 286 800 320
rect 834 286 868 320
rect 902 286 936 320
rect 970 286 1031 320
rect 784 270 1031 286
rect 500 230 566 260
rect 55 134 178 150
rect 55 100 71 134
rect 105 100 139 134
rect 173 100 178 134
rect 55 84 178 100
rect 212 210 278 226
rect 212 176 228 210
rect 262 176 278 210
rect 212 120 278 176
rect 212 86 228 120
rect 262 86 278 120
rect 212 17 278 86
rect 314 210 566 230
rect 700 236 750 260
rect 1081 236 1127 390
rect 1977 380 1993 414
rect 1943 364 1993 380
rect 1177 320 1511 356
rect 1177 286 1241 320
rect 1275 286 1309 320
rect 1343 286 1377 320
rect 1411 286 1445 320
rect 1479 286 1511 320
rect 1177 270 1511 286
rect 1561 320 1895 356
rect 1561 286 1646 320
rect 1680 286 1714 320
rect 1748 286 1782 320
rect 1816 286 1850 320
rect 1884 286 1895 320
rect 1561 270 1895 286
rect 314 176 330 210
rect 364 196 516 210
rect 314 120 364 176
rect 500 176 516 196
rect 550 176 566 210
rect 314 86 330 120
rect 314 70 364 86
rect 400 142 466 158
rect 400 108 416 142
rect 450 108 466 142
rect 400 17 466 108
rect 500 120 566 176
rect 500 86 516 120
rect 550 86 566 120
rect 500 70 566 86
rect 600 210 666 226
rect 600 176 616 210
rect 650 176 666 210
rect 600 120 666 176
rect 600 86 616 120
rect 650 86 666 120
rect 600 17 666 86
rect 700 210 1893 236
rect 700 176 716 210
rect 750 202 997 210
rect 700 120 750 176
rect 981 176 997 202
rect 1031 202 1266 210
rect 1031 176 1047 202
rect 700 86 716 120
rect 700 70 750 86
rect 786 152 947 168
rect 786 118 802 152
rect 836 118 911 152
rect 945 118 947 152
rect 786 17 947 118
rect 981 120 1047 176
rect 1250 176 1266 202
rect 1300 202 1466 210
rect 1300 176 1316 202
rect 981 86 997 120
rect 1031 86 1047 120
rect 981 70 1047 86
rect 1081 152 1216 168
rect 1081 118 1083 152
rect 1117 118 1180 152
rect 1214 118 1216 152
rect 1081 17 1216 118
rect 1250 120 1316 176
rect 1450 176 1466 202
rect 1500 202 1671 210
rect 1500 176 1516 202
rect 1250 86 1266 120
rect 1300 86 1316 120
rect 1250 70 1316 86
rect 1350 145 1416 161
rect 1350 111 1366 145
rect 1400 111 1416 145
rect 1350 17 1416 111
rect 1450 120 1516 176
rect 1655 176 1671 202
rect 1705 202 1843 210
rect 1450 86 1466 120
rect 1500 86 1516 120
rect 1450 70 1516 86
rect 1550 145 1621 161
rect 1550 111 1568 145
rect 1602 111 1621 145
rect 1550 17 1621 111
rect 1655 120 1705 176
rect 1877 176 1893 210
rect 1655 86 1671 120
rect 1655 70 1705 86
rect 1741 145 1807 161
rect 1741 111 1757 145
rect 1791 111 1807 145
rect 1741 17 1807 111
rect 1843 120 1893 176
rect 1877 86 1893 120
rect 1843 70 1893 86
rect 1927 210 1993 226
rect 1927 176 1943 210
rect 1977 176 1993 210
rect 1927 120 1993 176
rect 1927 86 1943 120
rect 1977 86 1993 120
rect 1927 17 1993 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
rlabel comment s 0 0 0 0 4 nor4b_4
flabel pwell s 0 0 2016 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 2016 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 2016 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 2016 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 D_N
port 4 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 D_N
port 4 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 1183 316 1217 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 1279 316 1313 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 1375 316 1409 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 1471 316 1505 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 1567 316 1601 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 1663 316 1697 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 1759 316 1793 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 1855 316 1889 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 1087 242 1121 276 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 1087 316 1121 350 0 FreeSans 340 0 0 0 Y
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 2016 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1175886
string GDS_START 1159914
<< end >>
