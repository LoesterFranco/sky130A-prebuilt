magic
tech sky130A
magscale 1 2
timestamp 1599588244
<< locali >>
rect 217 384 305 596
rect 24 51 90 321
rect 255 378 305 384
rect 255 344 375 378
rect 341 236 375 344
rect 409 270 459 356
rect 501 236 647 310
rect 341 202 412 236
rect 362 70 412 202
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 21 389 87 596
rect 127 423 177 649
rect 21 355 183 389
rect 345 446 404 596
rect 438 480 504 649
rect 538 446 597 596
rect 345 412 597 446
rect 149 310 183 355
rect 531 364 597 412
rect 149 244 307 310
rect 149 210 190 244
rect 124 108 190 210
rect 224 152 290 210
rect 224 17 326 152
rect 526 17 592 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel locali s 409 270 459 356 6 A1
port 1 nsew signal input
rlabel locali s 501 236 647 310 6 A2
port 2 nsew signal input
rlabel locali s 24 51 90 321 6 B1_N
port 3 nsew signal input
rlabel locali s 362 70 412 202 6 Y
port 4 nsew signal output
rlabel locali s 341 236 375 344 6 Y
port 4 nsew signal output
rlabel locali s 341 202 412 236 6 Y
port 4 nsew signal output
rlabel locali s 255 378 305 384 6 Y
port 4 nsew signal output
rlabel locali s 255 344 375 378 6 Y
port 4 nsew signal output
rlabel locali s 217 384 305 596 6 Y
port 4 nsew signal output
rlabel metal1 s 0 -49 672 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 6 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 617 672 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3915634
string GDS_START 3908960
<< end >>
