magic
tech sky130A
magscale 1 2
timestamp 1604502710
<< nwell >>
rect -38 332 710 704
<< pwell >>
rect 0 0 672 49
<< scpmos >>
rect 123 368 159 592
rect 201 368 237 592
rect 309 368 345 592
rect 417 368 453 592
rect 525 368 561 592
<< nmoslvt >>
rect 129 74 159 222
rect 215 74 245 222
rect 345 74 375 222
rect 431 74 461 222
rect 525 74 555 222
<< ndiff >>
rect 76 152 129 222
rect 76 118 84 152
rect 118 118 129 152
rect 76 74 129 118
rect 159 210 215 222
rect 159 176 170 210
rect 204 176 215 210
rect 159 120 215 176
rect 159 86 170 120
rect 204 86 215 120
rect 159 74 215 86
rect 245 152 345 222
rect 245 118 278 152
rect 312 118 345 152
rect 245 74 345 118
rect 375 210 431 222
rect 375 176 386 210
rect 420 176 431 210
rect 375 120 431 176
rect 375 86 386 120
rect 420 86 431 120
rect 375 74 431 86
rect 461 74 525 222
rect 555 197 612 222
rect 555 163 566 197
rect 600 163 612 197
rect 555 120 612 163
rect 555 86 566 120
rect 600 86 612 120
rect 555 74 612 86
<< pdiff >>
rect 71 580 123 592
rect 71 546 79 580
rect 113 546 123 580
rect 71 503 123 546
rect 71 469 79 503
rect 113 469 123 503
rect 71 424 123 469
rect 71 390 79 424
rect 113 390 123 424
rect 71 368 123 390
rect 159 368 201 592
rect 237 368 309 592
rect 345 580 417 592
rect 345 546 359 580
rect 393 546 417 580
rect 345 504 417 546
rect 345 470 359 504
rect 393 470 417 504
rect 345 424 417 470
rect 345 390 359 424
rect 393 390 417 424
rect 345 368 417 390
rect 453 580 525 592
rect 453 546 467 580
rect 501 546 525 580
rect 453 499 525 546
rect 453 465 467 499
rect 501 465 525 499
rect 453 368 525 465
rect 561 580 613 592
rect 561 546 571 580
rect 605 546 613 580
rect 561 497 613 546
rect 561 463 571 497
rect 605 463 613 497
rect 561 414 613 463
rect 561 380 571 414
rect 605 380 613 414
rect 561 368 613 380
<< ndiffc >>
rect 84 118 118 152
rect 170 176 204 210
rect 170 86 204 120
rect 278 118 312 152
rect 386 176 420 210
rect 386 86 420 120
rect 566 163 600 197
rect 566 86 600 120
<< pdiffc >>
rect 79 546 113 580
rect 79 469 113 503
rect 79 390 113 424
rect 359 546 393 580
rect 359 470 393 504
rect 359 390 393 424
rect 467 546 501 580
rect 467 465 501 499
rect 571 546 605 580
rect 571 463 605 497
rect 571 380 605 414
<< poly >>
rect 123 592 159 618
rect 201 592 237 618
rect 309 592 345 618
rect 417 592 453 618
rect 525 592 561 618
rect 123 336 159 368
rect 93 320 159 336
rect 93 286 109 320
rect 143 286 159 320
rect 93 270 159 286
rect 201 336 237 368
rect 309 336 345 368
rect 417 336 453 368
rect 201 320 267 336
rect 201 286 217 320
rect 251 286 267 320
rect 201 270 267 286
rect 309 320 375 336
rect 309 286 325 320
rect 359 286 375 320
rect 309 270 375 286
rect 417 320 483 336
rect 417 286 433 320
rect 467 286 483 320
rect 417 270 483 286
rect 525 310 561 368
rect 525 294 591 310
rect 129 222 159 270
rect 215 222 245 270
rect 345 222 375 270
rect 431 222 461 270
rect 525 260 541 294
rect 575 260 591 294
rect 525 244 591 260
rect 525 222 555 244
rect 129 48 159 74
rect 215 48 245 74
rect 345 48 375 74
rect 431 48 461 74
rect 525 48 555 74
<< polycont >>
rect 109 286 143 320
rect 217 286 251 320
rect 325 286 359 320
rect 433 286 467 320
rect 541 260 575 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 25 580 263 596
rect 25 546 79 580
rect 113 546 263 580
rect 25 503 263 546
rect 25 469 79 503
rect 113 469 263 503
rect 25 424 263 469
rect 25 390 79 424
rect 113 390 263 424
rect 339 580 413 596
rect 339 546 359 580
rect 393 546 413 580
rect 339 504 413 546
rect 339 470 359 504
rect 393 470 413 504
rect 339 424 413 470
rect 447 580 521 649
rect 447 546 467 580
rect 501 546 521 580
rect 447 499 521 546
rect 447 465 467 499
rect 501 465 521 499
rect 447 458 521 465
rect 555 580 621 596
rect 555 546 571 580
rect 605 546 621 580
rect 555 497 621 546
rect 555 463 571 497
rect 605 463 621 497
rect 555 424 621 463
rect 339 390 359 424
rect 393 414 621 424
rect 393 390 571 414
rect 25 236 59 390
rect 555 380 571 390
rect 605 380 621 414
rect 555 364 621 380
rect 93 320 167 356
rect 93 286 109 320
rect 143 286 167 320
rect 93 270 167 286
rect 201 320 267 356
rect 201 286 217 320
rect 251 286 267 320
rect 201 270 267 286
rect 309 320 375 356
rect 309 286 325 320
rect 359 286 375 320
rect 309 270 375 286
rect 409 320 483 356
rect 409 286 433 320
rect 467 286 483 320
rect 409 270 483 286
rect 525 294 647 310
rect 525 260 541 294
rect 575 260 647 294
rect 525 236 647 260
rect 25 210 436 236
rect 25 202 170 210
rect 204 202 386 210
rect 204 176 220 202
rect 68 152 134 168
rect 68 118 84 152
rect 118 118 134 152
rect 68 17 134 118
rect 170 120 220 176
rect 370 176 386 202
rect 420 176 436 210
rect 204 86 220 120
rect 170 70 220 86
rect 254 152 336 168
rect 254 118 278 152
rect 312 118 336 152
rect 254 17 336 118
rect 370 120 436 176
rect 370 86 386 120
rect 420 86 436 120
rect 370 70 436 86
rect 550 197 616 202
rect 550 163 566 197
rect 600 163 616 197
rect 550 120 616 163
rect 550 86 566 120
rect 600 86 616 120
rect 550 17 616 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
rlabel comment s 0 0 0 0 4 a2111oi_1
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 D1
port 5 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 607 242 641 276 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 31 464 65 498 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 31 538 65 572 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 127 464 161 498 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 127 538 161 572 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 223 464 257 498 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 223 538 257 572 0 FreeSans 340 0 0 0 Y
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 672 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3852498
string GDS_START 3845976
<< end >>
