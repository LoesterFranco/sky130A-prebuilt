magic
tech sky130A
magscale 1 2
timestamp 1601050047
<< nwell >>
rect -38 332 902 704
<< pwell >>
rect 0 0 864 49
<< scpmos >>
rect 90 387 120 587
rect 200 387 230 587
rect 290 387 320 587
rect 506 387 536 587
rect 620 387 650 587
rect 744 368 774 592
<< nmoslvt >>
rect 101 74 131 202
rect 179 74 209 202
rect 287 74 317 202
rect 431 74 461 202
rect 647 74 677 202
rect 749 74 779 222
<< ndiff >>
rect 699 202 749 222
rect 44 188 101 202
rect 44 154 56 188
rect 90 154 101 188
rect 44 120 101 154
rect 44 86 56 120
rect 90 86 101 120
rect 44 74 101 86
rect 131 74 179 202
rect 209 188 287 202
rect 209 154 228 188
rect 262 154 287 188
rect 209 120 287 154
rect 209 86 228 120
rect 262 86 287 120
rect 209 74 287 86
rect 317 190 431 202
rect 317 156 357 190
rect 391 156 431 190
rect 317 74 431 156
rect 461 122 647 202
rect 461 88 472 122
rect 506 88 586 122
rect 620 88 647 122
rect 461 74 647 88
rect 677 190 749 202
rect 677 156 688 190
rect 722 156 749 190
rect 677 120 749 156
rect 677 86 688 120
rect 722 86 749 120
rect 677 74 749 86
rect 779 210 836 222
rect 779 176 790 210
rect 824 176 836 210
rect 779 120 836 176
rect 779 86 790 120
rect 824 86 836 120
rect 779 74 836 86
<< pdiff >>
rect 675 587 744 592
rect 31 575 90 587
rect 31 541 43 575
rect 77 541 90 575
rect 31 504 90 541
rect 31 470 43 504
rect 77 470 90 504
rect 31 433 90 470
rect 31 399 43 433
rect 77 399 90 433
rect 31 387 90 399
rect 120 575 200 587
rect 120 541 143 575
rect 177 541 200 575
rect 120 507 200 541
rect 120 473 143 507
rect 177 473 200 507
rect 120 439 200 473
rect 120 405 143 439
rect 177 405 200 439
rect 120 387 200 405
rect 230 575 290 587
rect 230 541 243 575
rect 277 541 290 575
rect 230 504 290 541
rect 230 470 243 504
rect 277 470 290 504
rect 230 433 290 470
rect 230 399 243 433
rect 277 399 290 433
rect 230 387 290 399
rect 320 387 506 587
rect 536 387 620 587
rect 650 580 744 587
rect 650 546 687 580
rect 721 546 744 580
rect 650 511 744 546
rect 650 477 687 511
rect 721 477 744 511
rect 650 442 744 477
rect 650 408 687 442
rect 721 408 744 442
rect 650 387 744 408
rect 691 368 744 387
rect 774 580 833 592
rect 774 546 787 580
rect 821 546 833 580
rect 774 511 833 546
rect 774 477 787 511
rect 821 477 833 511
rect 774 442 833 477
rect 774 408 787 442
rect 821 408 833 442
rect 774 368 833 408
<< ndiffc >>
rect 56 154 90 188
rect 56 86 90 120
rect 228 154 262 188
rect 228 86 262 120
rect 357 156 391 190
rect 472 88 506 122
rect 586 88 620 122
rect 688 156 722 190
rect 688 86 722 120
rect 790 176 824 210
rect 790 86 824 120
<< pdiffc >>
rect 43 541 77 575
rect 43 470 77 504
rect 43 399 77 433
rect 143 541 177 575
rect 143 473 177 507
rect 143 405 177 439
rect 243 541 277 575
rect 243 470 277 504
rect 243 399 277 433
rect 687 546 721 580
rect 687 477 721 511
rect 687 408 721 442
rect 787 546 821 580
rect 787 477 821 511
rect 787 408 821 442
<< poly >>
rect 90 587 120 613
rect 200 587 230 613
rect 290 587 320 613
rect 506 587 536 613
rect 620 587 650 613
rect 744 592 774 618
rect 90 372 120 387
rect 200 372 230 387
rect 290 372 320 387
rect 506 372 536 387
rect 620 372 650 387
rect 87 294 123 372
rect 197 294 233 372
rect 287 342 425 372
rect 21 278 131 294
rect 21 244 37 278
rect 71 244 131 278
rect 21 228 131 244
rect 101 202 131 228
rect 179 278 245 294
rect 179 244 195 278
rect 229 244 245 278
rect 179 228 245 244
rect 287 278 353 294
rect 287 244 303 278
rect 337 244 353 278
rect 287 228 353 244
rect 395 290 425 342
rect 503 355 539 372
rect 503 339 569 355
rect 503 305 519 339
rect 553 305 569 339
rect 395 274 461 290
rect 503 289 569 305
rect 617 290 653 372
rect 744 353 774 368
rect 741 336 777 353
rect 719 320 785 336
rect 395 240 411 274
rect 445 240 461 274
rect 179 202 209 228
rect 287 202 317 228
rect 395 217 461 240
rect 611 274 677 290
rect 611 240 627 274
rect 661 240 677 274
rect 719 286 735 320
rect 769 286 785 320
rect 719 270 785 286
rect 611 224 677 240
rect 431 202 461 217
rect 647 202 677 224
rect 749 222 779 270
rect 101 48 131 74
rect 179 48 209 74
rect 287 48 317 74
rect 431 48 461 74
rect 647 48 677 74
rect 749 48 779 74
<< polycont >>
rect 37 244 71 278
rect 195 244 229 278
rect 303 244 337 278
rect 519 305 553 339
rect 411 240 445 274
rect 627 240 661 274
rect 735 286 769 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 27 575 93 591
rect 27 541 43 575
rect 77 541 93 575
rect 27 504 93 541
rect 27 470 43 504
rect 77 470 93 504
rect 27 433 93 470
rect 27 399 43 433
rect 77 399 93 433
rect 27 362 93 399
rect 127 575 193 649
rect 127 541 143 575
rect 177 541 193 575
rect 127 507 193 541
rect 127 473 143 507
rect 177 473 193 507
rect 127 439 193 473
rect 127 405 143 439
rect 177 405 193 439
rect 127 396 193 405
rect 227 575 637 591
rect 227 541 243 575
rect 277 557 637 575
rect 277 541 293 557
rect 227 504 293 541
rect 227 470 243 504
rect 277 470 293 504
rect 227 433 293 470
rect 227 399 243 433
rect 277 399 293 433
rect 227 362 293 399
rect 27 328 293 362
rect 327 464 569 498
rect 21 278 82 294
rect 21 244 37 278
rect 71 244 82 278
rect 21 228 82 244
rect 116 194 150 328
rect 327 294 361 464
rect 184 278 257 294
rect 184 244 195 278
rect 229 244 257 278
rect 184 228 257 244
rect 291 278 361 294
rect 291 244 303 278
rect 337 244 361 278
rect 291 228 361 244
rect 395 274 461 430
rect 503 339 569 464
rect 503 305 519 339
rect 553 305 569 339
rect 603 358 637 557
rect 671 580 737 649
rect 671 546 687 580
rect 721 546 737 580
rect 671 511 737 546
rect 671 477 687 511
rect 721 477 737 511
rect 671 442 737 477
rect 671 408 687 442
rect 721 408 737 442
rect 671 392 737 408
rect 771 580 847 596
rect 771 546 787 580
rect 821 546 847 580
rect 771 511 847 546
rect 771 477 787 511
rect 821 477 847 511
rect 771 442 847 477
rect 771 408 787 442
rect 821 408 847 442
rect 771 392 847 408
rect 603 324 779 358
rect 503 289 569 305
rect 719 320 779 324
rect 395 240 411 274
rect 445 240 461 274
rect 395 224 461 240
rect 603 274 677 290
rect 603 240 627 274
rect 661 240 677 274
rect 719 286 735 320
rect 769 286 779 320
rect 719 270 779 286
rect 603 224 677 240
rect 813 226 847 392
rect 774 210 847 226
rect 40 188 150 194
rect 40 154 56 188
rect 90 160 150 188
rect 212 188 278 194
rect 90 154 106 160
rect 40 120 106 154
rect 40 86 56 120
rect 90 86 106 120
rect 40 70 106 86
rect 212 154 228 188
rect 262 154 278 188
rect 312 156 357 190
rect 391 156 688 190
rect 722 156 738 190
rect 212 122 278 154
rect 212 120 472 122
rect 212 86 228 120
rect 262 88 472 120
rect 506 88 586 122
rect 620 88 636 122
rect 262 86 636 88
rect 212 56 636 86
rect 672 120 738 156
rect 672 86 688 120
rect 722 86 738 120
rect 672 17 738 86
rect 774 176 790 210
rect 824 176 847 210
rect 774 120 847 176
rect 774 86 790 120
rect 824 86 847 120
rect 774 70 847 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o311a_1
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 C1
port 5 nsew
flabel corelocali s 223 242 257 276 0 FreeSans 340 0 0 0 B1
port 4 nsew
flabel corelocali s 415 242 449 276 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 415 390 449 424 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 319 242 353 276 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 607 242 641 276 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 799 94 833 128 0 FreeSans 340 0 0 0 X
port 10 nsew
flabel corelocali s 799 168 833 202 0 FreeSans 340 0 0 0 X
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 864 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1324100
string GDS_START 1316248
<< end >>
