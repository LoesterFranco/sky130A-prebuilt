magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 3442 827
<< pwell >>
rect 29 1071 63 1105
rect 857 1071 891 1105
rect 1685 1071 1719 1105
rect 2513 1071 2547 1105
rect 3341 1071 3375 1105
rect 29 -17 63 17
rect 857 -17 891 17
rect 1685 -17 1719 17
rect 2513 -17 2547 17
rect 3341 -17 3375 17
<< scnmos >>
rect 79 911 109 1041
rect 174 937 204 1041
rect 387 937 417 1041
rect 503 937 533 1041
rect 716 937 746 1041
rect 811 911 841 1041
rect 907 911 937 1041
rect 1002 937 1032 1041
rect 1215 937 1245 1041
rect 1331 937 1361 1041
rect 1544 937 1574 1041
rect 1639 911 1669 1041
rect 1735 911 1765 1041
rect 1830 937 1860 1041
rect 2043 937 2073 1041
rect 2159 937 2189 1041
rect 2372 937 2402 1041
rect 2467 911 2497 1041
rect 2563 911 2593 1041
rect 2658 937 2688 1041
rect 2871 937 2901 1041
rect 2987 937 3017 1041
rect 3200 937 3230 1041
rect 3295 911 3325 1041
rect 79 47 109 177
rect 174 47 204 151
rect 387 47 417 151
rect 503 47 533 151
rect 716 47 746 151
rect 811 47 841 177
rect 907 47 937 177
rect 1002 47 1032 151
rect 1215 47 1245 151
rect 1331 47 1361 151
rect 1544 47 1574 151
rect 1639 47 1669 177
rect 1735 47 1765 177
rect 1830 47 1860 151
rect 2043 47 2073 151
rect 2159 47 2189 151
rect 2372 47 2402 151
rect 2467 47 2497 177
rect 2563 47 2593 177
rect 2658 47 2688 151
rect 2871 47 2901 151
rect 2987 47 3017 151
rect 3200 47 3230 151
rect 3295 47 3325 177
<< pmoshvt >>
rect 81 591 117 791
rect 186 591 222 755
rect 384 591 420 791
rect 500 591 536 791
rect 698 591 734 755
rect 803 591 839 791
rect 909 591 945 791
rect 1014 591 1050 755
rect 1212 591 1248 791
rect 1328 591 1364 791
rect 1526 591 1562 755
rect 1631 591 1667 791
rect 1737 591 1773 791
rect 1842 591 1878 755
rect 2040 591 2076 791
rect 2156 591 2192 791
rect 2354 591 2390 755
rect 2459 591 2495 791
rect 2565 591 2601 791
rect 2670 591 2706 755
rect 2868 591 2904 791
rect 2984 591 3020 791
rect 3182 591 3218 755
rect 3287 591 3323 791
rect 81 297 117 497
rect 186 333 222 497
rect 384 297 420 497
rect 500 297 536 497
rect 698 333 734 497
rect 803 297 839 497
rect 909 297 945 497
rect 1014 333 1050 497
rect 1212 297 1248 497
rect 1328 297 1364 497
rect 1526 333 1562 497
rect 1631 297 1667 497
rect 1737 297 1773 497
rect 1842 333 1878 497
rect 2040 297 2076 497
rect 2156 297 2192 497
rect 2354 333 2390 497
rect 2459 297 2495 497
rect 2565 297 2601 497
rect 2670 333 2706 497
rect 2868 297 2904 497
rect 2984 297 3020 497
rect 3182 333 3218 497
rect 3287 297 3323 497
<< ndiff >>
rect 27 1029 79 1041
rect 27 995 35 1029
rect 69 995 79 1029
rect 27 961 79 995
rect 27 927 35 961
rect 69 927 79 961
rect 27 911 79 927
rect 109 937 174 1041
rect 204 1006 256 1041
rect 204 972 214 1006
rect 248 972 256 1006
rect 204 937 256 972
rect 330 1006 387 1041
rect 330 972 338 1006
rect 372 972 387 1006
rect 330 937 387 972
rect 417 1006 503 1041
rect 417 972 443 1006
rect 477 972 503 1006
rect 417 937 503 972
rect 533 1006 590 1041
rect 533 972 548 1006
rect 582 972 590 1006
rect 533 937 590 972
rect 664 1006 716 1041
rect 664 972 672 1006
rect 706 972 716 1006
rect 664 937 716 972
rect 746 937 811 1041
rect 109 911 159 937
rect 761 911 811 937
rect 841 1029 907 1041
rect 841 995 857 1029
rect 891 995 907 1029
rect 841 961 907 995
rect 841 927 857 961
rect 891 927 907 961
rect 841 911 907 927
rect 937 937 1002 1041
rect 1032 1006 1084 1041
rect 1032 972 1042 1006
rect 1076 972 1084 1006
rect 1032 937 1084 972
rect 1158 1006 1215 1041
rect 1158 972 1166 1006
rect 1200 972 1215 1006
rect 1158 937 1215 972
rect 1245 1006 1331 1041
rect 1245 972 1271 1006
rect 1305 972 1331 1006
rect 1245 937 1331 972
rect 1361 1006 1418 1041
rect 1361 972 1376 1006
rect 1410 972 1418 1006
rect 1361 937 1418 972
rect 1492 1006 1544 1041
rect 1492 972 1500 1006
rect 1534 972 1544 1006
rect 1492 937 1544 972
rect 1574 937 1639 1041
rect 937 911 987 937
rect 1589 911 1639 937
rect 1669 1029 1735 1041
rect 1669 995 1685 1029
rect 1719 995 1735 1029
rect 1669 961 1735 995
rect 1669 927 1685 961
rect 1719 927 1735 961
rect 1669 911 1735 927
rect 1765 937 1830 1041
rect 1860 1006 1912 1041
rect 1860 972 1870 1006
rect 1904 972 1912 1006
rect 1860 937 1912 972
rect 1986 1006 2043 1041
rect 1986 972 1994 1006
rect 2028 972 2043 1006
rect 1986 937 2043 972
rect 2073 1006 2159 1041
rect 2073 972 2099 1006
rect 2133 972 2159 1006
rect 2073 937 2159 972
rect 2189 1006 2246 1041
rect 2189 972 2204 1006
rect 2238 972 2246 1006
rect 2189 937 2246 972
rect 2320 1006 2372 1041
rect 2320 972 2328 1006
rect 2362 972 2372 1006
rect 2320 937 2372 972
rect 2402 937 2467 1041
rect 1765 911 1815 937
rect 2417 911 2467 937
rect 2497 1029 2563 1041
rect 2497 995 2513 1029
rect 2547 995 2563 1029
rect 2497 961 2563 995
rect 2497 927 2513 961
rect 2547 927 2563 961
rect 2497 911 2563 927
rect 2593 937 2658 1041
rect 2688 1006 2740 1041
rect 2688 972 2698 1006
rect 2732 972 2740 1006
rect 2688 937 2740 972
rect 2814 1006 2871 1041
rect 2814 972 2822 1006
rect 2856 972 2871 1006
rect 2814 937 2871 972
rect 2901 1006 2987 1041
rect 2901 972 2927 1006
rect 2961 972 2987 1006
rect 2901 937 2987 972
rect 3017 1006 3074 1041
rect 3017 972 3032 1006
rect 3066 972 3074 1006
rect 3017 937 3074 972
rect 3148 1006 3200 1041
rect 3148 972 3156 1006
rect 3190 972 3200 1006
rect 3148 937 3200 972
rect 3230 937 3295 1041
rect 2593 911 2643 937
rect 3245 911 3295 937
rect 3325 1029 3377 1041
rect 3325 995 3335 1029
rect 3369 995 3377 1029
rect 3325 961 3377 995
rect 3325 927 3335 961
rect 3369 927 3377 961
rect 3325 911 3377 927
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 151 159 177
rect 761 151 811 177
rect 109 47 174 151
rect 204 116 256 151
rect 204 82 214 116
rect 248 82 256 116
rect 204 47 256 82
rect 330 116 387 151
rect 330 82 338 116
rect 372 82 387 116
rect 330 47 387 82
rect 417 116 503 151
rect 417 82 443 116
rect 477 82 503 116
rect 417 47 503 82
rect 533 116 590 151
rect 533 82 548 116
rect 582 82 590 116
rect 533 47 590 82
rect 664 116 716 151
rect 664 82 672 116
rect 706 82 716 116
rect 664 47 716 82
rect 746 47 811 151
rect 841 161 907 177
rect 841 127 857 161
rect 891 127 907 161
rect 841 93 907 127
rect 841 59 857 93
rect 891 59 907 93
rect 841 47 907 59
rect 937 151 987 177
rect 1589 151 1639 177
rect 937 47 1002 151
rect 1032 116 1084 151
rect 1032 82 1042 116
rect 1076 82 1084 116
rect 1032 47 1084 82
rect 1158 116 1215 151
rect 1158 82 1166 116
rect 1200 82 1215 116
rect 1158 47 1215 82
rect 1245 116 1331 151
rect 1245 82 1271 116
rect 1305 82 1331 116
rect 1245 47 1331 82
rect 1361 116 1418 151
rect 1361 82 1376 116
rect 1410 82 1418 116
rect 1361 47 1418 82
rect 1492 116 1544 151
rect 1492 82 1500 116
rect 1534 82 1544 116
rect 1492 47 1544 82
rect 1574 47 1639 151
rect 1669 161 1735 177
rect 1669 127 1685 161
rect 1719 127 1735 161
rect 1669 93 1735 127
rect 1669 59 1685 93
rect 1719 59 1735 93
rect 1669 47 1735 59
rect 1765 151 1815 177
rect 2417 151 2467 177
rect 1765 47 1830 151
rect 1860 116 1912 151
rect 1860 82 1870 116
rect 1904 82 1912 116
rect 1860 47 1912 82
rect 1986 116 2043 151
rect 1986 82 1994 116
rect 2028 82 2043 116
rect 1986 47 2043 82
rect 2073 116 2159 151
rect 2073 82 2099 116
rect 2133 82 2159 116
rect 2073 47 2159 82
rect 2189 116 2246 151
rect 2189 82 2204 116
rect 2238 82 2246 116
rect 2189 47 2246 82
rect 2320 116 2372 151
rect 2320 82 2328 116
rect 2362 82 2372 116
rect 2320 47 2372 82
rect 2402 47 2467 151
rect 2497 161 2563 177
rect 2497 127 2513 161
rect 2547 127 2563 161
rect 2497 93 2563 127
rect 2497 59 2513 93
rect 2547 59 2563 93
rect 2497 47 2563 59
rect 2593 151 2643 177
rect 3245 151 3295 177
rect 2593 47 2658 151
rect 2688 116 2740 151
rect 2688 82 2698 116
rect 2732 82 2740 116
rect 2688 47 2740 82
rect 2814 116 2871 151
rect 2814 82 2822 116
rect 2856 82 2871 116
rect 2814 47 2871 82
rect 2901 116 2987 151
rect 2901 82 2927 116
rect 2961 82 2987 116
rect 2901 47 2987 82
rect 3017 116 3074 151
rect 3017 82 3032 116
rect 3066 82 3074 116
rect 3017 47 3074 82
rect 3148 116 3200 151
rect 3148 82 3156 116
rect 3190 82 3200 116
rect 3148 47 3200 82
rect 3230 47 3295 151
rect 3325 161 3377 177
rect 3325 127 3335 161
rect 3369 127 3377 161
rect 3325 93 3377 127
rect 3325 59 3335 93
rect 3369 59 3377 93
rect 3325 47 3377 59
<< pdiff >>
rect 27 773 81 791
rect 27 739 35 773
rect 69 739 81 773
rect 27 705 81 739
rect 27 671 35 705
rect 69 671 81 705
rect 27 637 81 671
rect 27 603 35 637
rect 69 603 81 637
rect 27 591 81 603
rect 117 755 169 791
rect 330 779 384 791
rect 117 591 186 755
rect 222 705 276 755
rect 222 671 234 705
rect 268 671 276 705
rect 222 637 276 671
rect 222 603 234 637
rect 268 603 276 637
rect 222 591 276 603
rect 330 745 338 779
rect 372 745 384 779
rect 330 711 384 745
rect 330 677 338 711
rect 372 677 384 711
rect 330 643 384 677
rect 330 609 338 643
rect 372 609 384 643
rect 330 591 384 609
rect 420 779 500 791
rect 420 745 443 779
rect 477 745 500 779
rect 420 711 500 745
rect 420 677 443 711
rect 477 677 500 711
rect 420 643 500 677
rect 420 609 443 643
rect 477 609 500 643
rect 420 591 500 609
rect 536 779 590 791
rect 536 745 548 779
rect 582 745 590 779
rect 751 755 803 791
rect 536 711 590 745
rect 536 677 548 711
rect 582 677 590 711
rect 536 643 590 677
rect 536 609 548 643
rect 582 609 590 643
rect 536 591 590 609
rect 644 705 698 755
rect 644 671 652 705
rect 686 671 698 705
rect 644 637 698 671
rect 644 603 652 637
rect 686 603 698 637
rect 644 591 698 603
rect 734 591 803 755
rect 839 773 909 791
rect 839 739 857 773
rect 891 739 909 773
rect 839 705 909 739
rect 839 671 857 705
rect 891 671 909 705
rect 839 637 909 671
rect 839 603 857 637
rect 891 603 909 637
rect 839 591 909 603
rect 945 755 997 791
rect 1158 779 1212 791
rect 945 591 1014 755
rect 1050 705 1104 755
rect 1050 671 1062 705
rect 1096 671 1104 705
rect 1050 637 1104 671
rect 1050 603 1062 637
rect 1096 603 1104 637
rect 1050 591 1104 603
rect 1158 745 1166 779
rect 1200 745 1212 779
rect 1158 711 1212 745
rect 1158 677 1166 711
rect 1200 677 1212 711
rect 1158 643 1212 677
rect 1158 609 1166 643
rect 1200 609 1212 643
rect 1158 591 1212 609
rect 1248 779 1328 791
rect 1248 745 1271 779
rect 1305 745 1328 779
rect 1248 711 1328 745
rect 1248 677 1271 711
rect 1305 677 1328 711
rect 1248 643 1328 677
rect 1248 609 1271 643
rect 1305 609 1328 643
rect 1248 591 1328 609
rect 1364 779 1418 791
rect 1364 745 1376 779
rect 1410 745 1418 779
rect 1579 755 1631 791
rect 1364 711 1418 745
rect 1364 677 1376 711
rect 1410 677 1418 711
rect 1364 643 1418 677
rect 1364 609 1376 643
rect 1410 609 1418 643
rect 1364 591 1418 609
rect 1472 705 1526 755
rect 1472 671 1480 705
rect 1514 671 1526 705
rect 1472 637 1526 671
rect 1472 603 1480 637
rect 1514 603 1526 637
rect 1472 591 1526 603
rect 1562 591 1631 755
rect 1667 773 1737 791
rect 1667 739 1685 773
rect 1719 739 1737 773
rect 1667 705 1737 739
rect 1667 671 1685 705
rect 1719 671 1737 705
rect 1667 637 1737 671
rect 1667 603 1685 637
rect 1719 603 1737 637
rect 1667 591 1737 603
rect 1773 755 1825 791
rect 1986 779 2040 791
rect 1773 591 1842 755
rect 1878 705 1932 755
rect 1878 671 1890 705
rect 1924 671 1932 705
rect 1878 637 1932 671
rect 1878 603 1890 637
rect 1924 603 1932 637
rect 1878 591 1932 603
rect 1986 745 1994 779
rect 2028 745 2040 779
rect 1986 711 2040 745
rect 1986 677 1994 711
rect 2028 677 2040 711
rect 1986 643 2040 677
rect 1986 609 1994 643
rect 2028 609 2040 643
rect 1986 591 2040 609
rect 2076 779 2156 791
rect 2076 745 2099 779
rect 2133 745 2156 779
rect 2076 711 2156 745
rect 2076 677 2099 711
rect 2133 677 2156 711
rect 2076 643 2156 677
rect 2076 609 2099 643
rect 2133 609 2156 643
rect 2076 591 2156 609
rect 2192 779 2246 791
rect 2192 745 2204 779
rect 2238 745 2246 779
rect 2407 755 2459 791
rect 2192 711 2246 745
rect 2192 677 2204 711
rect 2238 677 2246 711
rect 2192 643 2246 677
rect 2192 609 2204 643
rect 2238 609 2246 643
rect 2192 591 2246 609
rect 2300 705 2354 755
rect 2300 671 2308 705
rect 2342 671 2354 705
rect 2300 637 2354 671
rect 2300 603 2308 637
rect 2342 603 2354 637
rect 2300 591 2354 603
rect 2390 591 2459 755
rect 2495 773 2565 791
rect 2495 739 2513 773
rect 2547 739 2565 773
rect 2495 705 2565 739
rect 2495 671 2513 705
rect 2547 671 2565 705
rect 2495 637 2565 671
rect 2495 603 2513 637
rect 2547 603 2565 637
rect 2495 591 2565 603
rect 2601 755 2653 791
rect 2814 779 2868 791
rect 2601 591 2670 755
rect 2706 705 2760 755
rect 2706 671 2718 705
rect 2752 671 2760 705
rect 2706 637 2760 671
rect 2706 603 2718 637
rect 2752 603 2760 637
rect 2706 591 2760 603
rect 2814 745 2822 779
rect 2856 745 2868 779
rect 2814 711 2868 745
rect 2814 677 2822 711
rect 2856 677 2868 711
rect 2814 643 2868 677
rect 2814 609 2822 643
rect 2856 609 2868 643
rect 2814 591 2868 609
rect 2904 779 2984 791
rect 2904 745 2927 779
rect 2961 745 2984 779
rect 2904 711 2984 745
rect 2904 677 2927 711
rect 2961 677 2984 711
rect 2904 643 2984 677
rect 2904 609 2927 643
rect 2961 609 2984 643
rect 2904 591 2984 609
rect 3020 779 3074 791
rect 3020 745 3032 779
rect 3066 745 3074 779
rect 3235 755 3287 791
rect 3020 711 3074 745
rect 3020 677 3032 711
rect 3066 677 3074 711
rect 3020 643 3074 677
rect 3020 609 3032 643
rect 3066 609 3074 643
rect 3020 591 3074 609
rect 3128 705 3182 755
rect 3128 671 3136 705
rect 3170 671 3182 705
rect 3128 637 3182 671
rect 3128 603 3136 637
rect 3170 603 3182 637
rect 3128 591 3182 603
rect 3218 591 3287 755
rect 3323 773 3377 791
rect 3323 739 3335 773
rect 3369 739 3377 773
rect 3323 705 3377 739
rect 3323 671 3335 705
rect 3369 671 3377 705
rect 3323 637 3377 671
rect 3323 603 3335 637
rect 3369 603 3377 637
rect 3323 591 3377 603
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 333 186 497
rect 222 485 276 497
rect 222 451 234 485
rect 268 451 276 485
rect 222 417 276 451
rect 222 383 234 417
rect 268 383 276 417
rect 222 333 276 383
rect 330 479 384 497
rect 330 445 338 479
rect 372 445 384 479
rect 330 411 384 445
rect 330 377 338 411
rect 372 377 384 411
rect 330 343 384 377
rect 117 297 169 333
rect 330 309 338 343
rect 372 309 384 343
rect 330 297 384 309
rect 420 479 500 497
rect 420 445 443 479
rect 477 445 500 479
rect 420 411 500 445
rect 420 377 443 411
rect 477 377 500 411
rect 420 343 500 377
rect 420 309 443 343
rect 477 309 500 343
rect 420 297 500 309
rect 536 479 590 497
rect 536 445 548 479
rect 582 445 590 479
rect 536 411 590 445
rect 536 377 548 411
rect 582 377 590 411
rect 536 343 590 377
rect 536 309 548 343
rect 582 309 590 343
rect 644 485 698 497
rect 644 451 652 485
rect 686 451 698 485
rect 644 417 698 451
rect 644 383 652 417
rect 686 383 698 417
rect 644 333 698 383
rect 734 333 803 497
rect 536 297 590 309
rect 751 297 803 333
rect 839 485 909 497
rect 839 451 857 485
rect 891 451 909 485
rect 839 417 909 451
rect 839 383 857 417
rect 891 383 909 417
rect 839 349 909 383
rect 839 315 857 349
rect 891 315 909 349
rect 839 297 909 315
rect 945 333 1014 497
rect 1050 485 1104 497
rect 1050 451 1062 485
rect 1096 451 1104 485
rect 1050 417 1104 451
rect 1050 383 1062 417
rect 1096 383 1104 417
rect 1050 333 1104 383
rect 1158 479 1212 497
rect 1158 445 1166 479
rect 1200 445 1212 479
rect 1158 411 1212 445
rect 1158 377 1166 411
rect 1200 377 1212 411
rect 1158 343 1212 377
rect 945 297 997 333
rect 1158 309 1166 343
rect 1200 309 1212 343
rect 1158 297 1212 309
rect 1248 479 1328 497
rect 1248 445 1271 479
rect 1305 445 1328 479
rect 1248 411 1328 445
rect 1248 377 1271 411
rect 1305 377 1328 411
rect 1248 343 1328 377
rect 1248 309 1271 343
rect 1305 309 1328 343
rect 1248 297 1328 309
rect 1364 479 1418 497
rect 1364 445 1376 479
rect 1410 445 1418 479
rect 1364 411 1418 445
rect 1364 377 1376 411
rect 1410 377 1418 411
rect 1364 343 1418 377
rect 1364 309 1376 343
rect 1410 309 1418 343
rect 1472 485 1526 497
rect 1472 451 1480 485
rect 1514 451 1526 485
rect 1472 417 1526 451
rect 1472 383 1480 417
rect 1514 383 1526 417
rect 1472 333 1526 383
rect 1562 333 1631 497
rect 1364 297 1418 309
rect 1579 297 1631 333
rect 1667 485 1737 497
rect 1667 451 1685 485
rect 1719 451 1737 485
rect 1667 417 1737 451
rect 1667 383 1685 417
rect 1719 383 1737 417
rect 1667 349 1737 383
rect 1667 315 1685 349
rect 1719 315 1737 349
rect 1667 297 1737 315
rect 1773 333 1842 497
rect 1878 485 1932 497
rect 1878 451 1890 485
rect 1924 451 1932 485
rect 1878 417 1932 451
rect 1878 383 1890 417
rect 1924 383 1932 417
rect 1878 333 1932 383
rect 1986 479 2040 497
rect 1986 445 1994 479
rect 2028 445 2040 479
rect 1986 411 2040 445
rect 1986 377 1994 411
rect 2028 377 2040 411
rect 1986 343 2040 377
rect 1773 297 1825 333
rect 1986 309 1994 343
rect 2028 309 2040 343
rect 1986 297 2040 309
rect 2076 479 2156 497
rect 2076 445 2099 479
rect 2133 445 2156 479
rect 2076 411 2156 445
rect 2076 377 2099 411
rect 2133 377 2156 411
rect 2076 343 2156 377
rect 2076 309 2099 343
rect 2133 309 2156 343
rect 2076 297 2156 309
rect 2192 479 2246 497
rect 2192 445 2204 479
rect 2238 445 2246 479
rect 2192 411 2246 445
rect 2192 377 2204 411
rect 2238 377 2246 411
rect 2192 343 2246 377
rect 2192 309 2204 343
rect 2238 309 2246 343
rect 2300 485 2354 497
rect 2300 451 2308 485
rect 2342 451 2354 485
rect 2300 417 2354 451
rect 2300 383 2308 417
rect 2342 383 2354 417
rect 2300 333 2354 383
rect 2390 333 2459 497
rect 2192 297 2246 309
rect 2407 297 2459 333
rect 2495 485 2565 497
rect 2495 451 2513 485
rect 2547 451 2565 485
rect 2495 417 2565 451
rect 2495 383 2513 417
rect 2547 383 2565 417
rect 2495 349 2565 383
rect 2495 315 2513 349
rect 2547 315 2565 349
rect 2495 297 2565 315
rect 2601 333 2670 497
rect 2706 485 2760 497
rect 2706 451 2718 485
rect 2752 451 2760 485
rect 2706 417 2760 451
rect 2706 383 2718 417
rect 2752 383 2760 417
rect 2706 333 2760 383
rect 2814 479 2868 497
rect 2814 445 2822 479
rect 2856 445 2868 479
rect 2814 411 2868 445
rect 2814 377 2822 411
rect 2856 377 2868 411
rect 2814 343 2868 377
rect 2601 297 2653 333
rect 2814 309 2822 343
rect 2856 309 2868 343
rect 2814 297 2868 309
rect 2904 479 2984 497
rect 2904 445 2927 479
rect 2961 445 2984 479
rect 2904 411 2984 445
rect 2904 377 2927 411
rect 2961 377 2984 411
rect 2904 343 2984 377
rect 2904 309 2927 343
rect 2961 309 2984 343
rect 2904 297 2984 309
rect 3020 479 3074 497
rect 3020 445 3032 479
rect 3066 445 3074 479
rect 3020 411 3074 445
rect 3020 377 3032 411
rect 3066 377 3074 411
rect 3020 343 3074 377
rect 3020 309 3032 343
rect 3066 309 3074 343
rect 3128 485 3182 497
rect 3128 451 3136 485
rect 3170 451 3182 485
rect 3128 417 3182 451
rect 3128 383 3136 417
rect 3170 383 3182 417
rect 3128 333 3182 383
rect 3218 333 3287 497
rect 3020 297 3074 309
rect 3235 297 3287 333
rect 3323 485 3377 497
rect 3323 451 3335 485
rect 3369 451 3377 485
rect 3323 417 3377 451
rect 3323 383 3335 417
rect 3369 383 3377 417
rect 3323 349 3377 383
rect 3323 315 3335 349
rect 3369 315 3377 349
rect 3323 297 3377 315
<< ndiffc >>
rect 35 995 69 1029
rect 35 927 69 961
rect 214 972 248 1006
rect 338 972 372 1006
rect 443 972 477 1006
rect 548 972 582 1006
rect 672 972 706 1006
rect 857 995 891 1029
rect 857 927 891 961
rect 1042 972 1076 1006
rect 1166 972 1200 1006
rect 1271 972 1305 1006
rect 1376 972 1410 1006
rect 1500 972 1534 1006
rect 1685 995 1719 1029
rect 1685 927 1719 961
rect 1870 972 1904 1006
rect 1994 972 2028 1006
rect 2099 972 2133 1006
rect 2204 972 2238 1006
rect 2328 972 2362 1006
rect 2513 995 2547 1029
rect 2513 927 2547 961
rect 2698 972 2732 1006
rect 2822 972 2856 1006
rect 2927 972 2961 1006
rect 3032 972 3066 1006
rect 3156 972 3190 1006
rect 3335 995 3369 1029
rect 3335 927 3369 961
rect 35 127 69 161
rect 35 59 69 93
rect 214 82 248 116
rect 338 82 372 116
rect 443 82 477 116
rect 548 82 582 116
rect 672 82 706 116
rect 857 127 891 161
rect 857 59 891 93
rect 1042 82 1076 116
rect 1166 82 1200 116
rect 1271 82 1305 116
rect 1376 82 1410 116
rect 1500 82 1534 116
rect 1685 127 1719 161
rect 1685 59 1719 93
rect 1870 82 1904 116
rect 1994 82 2028 116
rect 2099 82 2133 116
rect 2204 82 2238 116
rect 2328 82 2362 116
rect 2513 127 2547 161
rect 2513 59 2547 93
rect 2698 82 2732 116
rect 2822 82 2856 116
rect 2927 82 2961 116
rect 3032 82 3066 116
rect 3156 82 3190 116
rect 3335 127 3369 161
rect 3335 59 3369 93
<< pdiffc >>
rect 35 739 69 773
rect 35 671 69 705
rect 35 603 69 637
rect 234 671 268 705
rect 234 603 268 637
rect 338 745 372 779
rect 338 677 372 711
rect 338 609 372 643
rect 443 745 477 779
rect 443 677 477 711
rect 443 609 477 643
rect 548 745 582 779
rect 548 677 582 711
rect 548 609 582 643
rect 652 671 686 705
rect 652 603 686 637
rect 857 739 891 773
rect 857 671 891 705
rect 857 603 891 637
rect 1062 671 1096 705
rect 1062 603 1096 637
rect 1166 745 1200 779
rect 1166 677 1200 711
rect 1166 609 1200 643
rect 1271 745 1305 779
rect 1271 677 1305 711
rect 1271 609 1305 643
rect 1376 745 1410 779
rect 1376 677 1410 711
rect 1376 609 1410 643
rect 1480 671 1514 705
rect 1480 603 1514 637
rect 1685 739 1719 773
rect 1685 671 1719 705
rect 1685 603 1719 637
rect 1890 671 1924 705
rect 1890 603 1924 637
rect 1994 745 2028 779
rect 1994 677 2028 711
rect 1994 609 2028 643
rect 2099 745 2133 779
rect 2099 677 2133 711
rect 2099 609 2133 643
rect 2204 745 2238 779
rect 2204 677 2238 711
rect 2204 609 2238 643
rect 2308 671 2342 705
rect 2308 603 2342 637
rect 2513 739 2547 773
rect 2513 671 2547 705
rect 2513 603 2547 637
rect 2718 671 2752 705
rect 2718 603 2752 637
rect 2822 745 2856 779
rect 2822 677 2856 711
rect 2822 609 2856 643
rect 2927 745 2961 779
rect 2927 677 2961 711
rect 2927 609 2961 643
rect 3032 745 3066 779
rect 3032 677 3066 711
rect 3032 609 3066 643
rect 3136 671 3170 705
rect 3136 603 3170 637
rect 3335 739 3369 773
rect 3335 671 3369 705
rect 3335 603 3369 637
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 234 451 268 485
rect 234 383 268 417
rect 338 445 372 479
rect 338 377 372 411
rect 338 309 372 343
rect 443 445 477 479
rect 443 377 477 411
rect 443 309 477 343
rect 548 445 582 479
rect 548 377 582 411
rect 548 309 582 343
rect 652 451 686 485
rect 652 383 686 417
rect 857 451 891 485
rect 857 383 891 417
rect 857 315 891 349
rect 1062 451 1096 485
rect 1062 383 1096 417
rect 1166 445 1200 479
rect 1166 377 1200 411
rect 1166 309 1200 343
rect 1271 445 1305 479
rect 1271 377 1305 411
rect 1271 309 1305 343
rect 1376 445 1410 479
rect 1376 377 1410 411
rect 1376 309 1410 343
rect 1480 451 1514 485
rect 1480 383 1514 417
rect 1685 451 1719 485
rect 1685 383 1719 417
rect 1685 315 1719 349
rect 1890 451 1924 485
rect 1890 383 1924 417
rect 1994 445 2028 479
rect 1994 377 2028 411
rect 1994 309 2028 343
rect 2099 445 2133 479
rect 2099 377 2133 411
rect 2099 309 2133 343
rect 2204 445 2238 479
rect 2204 377 2238 411
rect 2204 309 2238 343
rect 2308 451 2342 485
rect 2308 383 2342 417
rect 2513 451 2547 485
rect 2513 383 2547 417
rect 2513 315 2547 349
rect 2718 451 2752 485
rect 2718 383 2752 417
rect 2822 445 2856 479
rect 2822 377 2856 411
rect 2822 309 2856 343
rect 2927 445 2961 479
rect 2927 377 2961 411
rect 2927 309 2961 343
rect 3032 445 3066 479
rect 3032 377 3066 411
rect 3032 309 3066 343
rect 3136 451 3170 485
rect 3136 383 3170 417
rect 3335 451 3369 485
rect 3335 383 3369 417
rect 3335 315 3369 349
<< poly >>
rect 79 1041 109 1067
rect 174 1041 204 1067
rect 387 1041 417 1067
rect 503 1041 533 1067
rect 716 1041 746 1067
rect 811 1041 841 1067
rect 907 1041 937 1067
rect 1002 1041 1032 1067
rect 1215 1041 1245 1067
rect 1331 1041 1361 1067
rect 1544 1041 1574 1067
rect 1639 1041 1669 1067
rect 1735 1041 1765 1067
rect 1830 1041 1860 1067
rect 2043 1041 2073 1067
rect 2159 1041 2189 1067
rect 2372 1041 2402 1067
rect 2467 1041 2497 1067
rect 2563 1041 2593 1067
rect 2658 1041 2688 1067
rect 2871 1041 2901 1067
rect 2987 1041 3017 1067
rect 3200 1041 3230 1067
rect 3295 1041 3325 1067
rect 174 922 204 937
rect 387 922 417 937
rect 174 915 417 922
rect 503 922 533 937
rect 716 922 746 937
rect 503 915 746 922
rect 79 889 109 911
rect 174 899 422 915
rect 174 892 378 899
rect 73 873 127 889
rect 73 839 83 873
rect 117 839 127 873
rect 368 865 378 892
rect 412 865 422 899
rect 368 849 422 865
rect 73 823 127 839
rect 232 837 298 847
rect 232 823 248 837
rect 79 806 119 823
rect 81 791 117 806
rect 184 803 248 823
rect 282 803 298 837
rect 382 806 422 849
rect 498 899 746 915
rect 1002 922 1032 937
rect 1215 922 1245 937
rect 1002 915 1245 922
rect 1331 922 1361 937
rect 1544 922 1574 937
rect 1331 915 1574 922
rect 498 865 508 899
rect 542 892 746 899
rect 542 865 552 892
rect 811 889 841 911
rect 907 889 937 911
rect 1002 899 1250 915
rect 1002 892 1206 899
rect 498 849 552 865
rect 793 873 847 889
rect 498 806 538 849
rect 622 837 688 847
rect 184 793 298 803
rect 186 755 222 793
rect 384 791 420 806
rect 500 791 536 806
rect 622 803 638 837
rect 672 823 688 837
rect 793 839 803 873
rect 837 839 847 873
rect 793 823 847 839
rect 901 873 955 889
rect 901 839 911 873
rect 945 839 955 873
rect 1196 865 1206 892
rect 1240 865 1250 899
rect 1196 849 1250 865
rect 901 823 955 839
rect 1060 837 1126 847
rect 1060 823 1076 837
rect 672 803 736 823
rect 801 806 841 823
rect 907 806 947 823
rect 622 793 736 803
rect 698 755 734 793
rect 803 791 839 806
rect 909 791 945 806
rect 1012 803 1076 823
rect 1110 803 1126 837
rect 1210 806 1250 849
rect 1326 899 1574 915
rect 1830 922 1860 937
rect 2043 922 2073 937
rect 1830 915 2073 922
rect 2159 922 2189 937
rect 2372 922 2402 937
rect 2159 915 2402 922
rect 1326 865 1336 899
rect 1370 892 1574 899
rect 1370 865 1380 892
rect 1639 889 1669 911
rect 1735 889 1765 911
rect 1830 899 2078 915
rect 1830 892 2034 899
rect 1326 849 1380 865
rect 1621 873 1675 889
rect 1326 806 1366 849
rect 1450 837 1516 847
rect 1012 793 1126 803
rect 1014 755 1050 793
rect 1212 791 1248 806
rect 1328 791 1364 806
rect 1450 803 1466 837
rect 1500 823 1516 837
rect 1621 839 1631 873
rect 1665 839 1675 873
rect 1621 823 1675 839
rect 1729 873 1783 889
rect 1729 839 1739 873
rect 1773 839 1783 873
rect 2024 865 2034 892
rect 2068 865 2078 899
rect 2024 849 2078 865
rect 1729 823 1783 839
rect 1888 837 1954 847
rect 1888 823 1904 837
rect 1500 803 1564 823
rect 1629 806 1669 823
rect 1735 806 1775 823
rect 1450 793 1564 803
rect 1526 755 1562 793
rect 1631 791 1667 806
rect 1737 791 1773 806
rect 1840 803 1904 823
rect 1938 803 1954 837
rect 2038 806 2078 849
rect 2154 899 2402 915
rect 2658 922 2688 937
rect 2871 922 2901 937
rect 2658 915 2901 922
rect 2987 922 3017 937
rect 3200 922 3230 937
rect 2987 915 3230 922
rect 2154 865 2164 899
rect 2198 892 2402 899
rect 2198 865 2208 892
rect 2467 889 2497 911
rect 2563 889 2593 911
rect 2658 899 2906 915
rect 2658 892 2862 899
rect 2154 849 2208 865
rect 2449 873 2503 889
rect 2154 806 2194 849
rect 2278 837 2344 847
rect 1840 793 1954 803
rect 1842 755 1878 793
rect 2040 791 2076 806
rect 2156 791 2192 806
rect 2278 803 2294 837
rect 2328 823 2344 837
rect 2449 839 2459 873
rect 2493 839 2503 873
rect 2449 823 2503 839
rect 2557 873 2611 889
rect 2557 839 2567 873
rect 2601 839 2611 873
rect 2852 865 2862 892
rect 2896 865 2906 899
rect 2852 849 2906 865
rect 2557 823 2611 839
rect 2716 837 2782 847
rect 2716 823 2732 837
rect 2328 803 2392 823
rect 2457 806 2497 823
rect 2563 806 2603 823
rect 2278 793 2392 803
rect 2354 755 2390 793
rect 2459 791 2495 806
rect 2565 791 2601 806
rect 2668 803 2732 823
rect 2766 803 2782 837
rect 2866 806 2906 849
rect 2982 899 3230 915
rect 2982 865 2992 899
rect 3026 892 3230 899
rect 3026 865 3036 892
rect 3295 889 3325 911
rect 2982 849 3036 865
rect 3277 873 3331 889
rect 2982 806 3022 849
rect 3106 837 3172 847
rect 2668 793 2782 803
rect 2670 755 2706 793
rect 2868 791 2904 806
rect 2984 791 3020 806
rect 3106 803 3122 837
rect 3156 823 3172 837
rect 3277 839 3287 873
rect 3321 839 3331 873
rect 3277 823 3331 839
rect 3156 803 3220 823
rect 3285 806 3325 823
rect 3106 793 3220 803
rect 3182 755 3218 793
rect 3287 791 3323 806
rect 81 565 117 591
rect 186 565 222 591
rect 384 565 420 591
rect 500 565 536 591
rect 698 565 734 591
rect 803 565 839 591
rect 909 565 945 591
rect 1014 565 1050 591
rect 1212 565 1248 591
rect 1328 565 1364 591
rect 1526 565 1562 591
rect 1631 565 1667 591
rect 1737 565 1773 591
rect 1842 565 1878 591
rect 2040 565 2076 591
rect 2156 565 2192 591
rect 2354 565 2390 591
rect 2459 565 2495 591
rect 2565 565 2601 591
rect 2670 565 2706 591
rect 2868 565 2904 591
rect 2984 565 3020 591
rect 3182 565 3218 591
rect 3287 565 3323 591
rect 81 497 117 523
rect 186 497 222 523
rect 384 497 420 523
rect 500 497 536 523
rect 698 497 734 523
rect 803 497 839 523
rect 909 497 945 523
rect 1014 497 1050 523
rect 1212 497 1248 523
rect 1328 497 1364 523
rect 1526 497 1562 523
rect 1631 497 1667 523
rect 1737 497 1773 523
rect 1842 497 1878 523
rect 2040 497 2076 523
rect 2156 497 2192 523
rect 2354 497 2390 523
rect 2459 497 2495 523
rect 2565 497 2601 523
rect 2670 497 2706 523
rect 2868 497 2904 523
rect 2984 497 3020 523
rect 3182 497 3218 523
rect 3287 497 3323 523
rect 81 282 117 297
rect 186 295 222 333
rect 184 285 298 295
rect 79 265 119 282
rect 184 265 248 285
rect 73 249 127 265
rect 73 215 83 249
rect 117 215 127 249
rect 232 251 248 265
rect 282 251 298 285
rect 384 282 420 297
rect 500 282 536 297
rect 698 295 734 333
rect 622 285 736 295
rect 232 241 298 251
rect 382 239 422 282
rect 73 199 127 215
rect 368 223 422 239
rect 79 177 109 199
rect 368 196 378 223
rect 174 189 378 196
rect 412 189 422 223
rect 174 173 422 189
rect 498 239 538 282
rect 622 251 638 285
rect 672 265 736 285
rect 803 282 839 297
rect 909 282 945 297
rect 1014 295 1050 333
rect 1012 285 1126 295
rect 801 265 841 282
rect 907 265 947 282
rect 1012 265 1076 285
rect 672 251 688 265
rect 622 241 688 251
rect 793 249 847 265
rect 498 223 552 239
rect 498 189 508 223
rect 542 196 552 223
rect 793 215 803 249
rect 837 215 847 249
rect 793 199 847 215
rect 901 249 955 265
rect 901 215 911 249
rect 945 215 955 249
rect 1060 251 1076 265
rect 1110 251 1126 285
rect 1212 282 1248 297
rect 1328 282 1364 297
rect 1526 295 1562 333
rect 1450 285 1564 295
rect 1060 241 1126 251
rect 1210 239 1250 282
rect 901 199 955 215
rect 1196 223 1250 239
rect 542 189 746 196
rect 498 173 746 189
rect 811 177 841 199
rect 907 177 937 199
rect 1196 196 1206 223
rect 1002 189 1206 196
rect 1240 189 1250 223
rect 174 166 417 173
rect 174 151 204 166
rect 387 151 417 166
rect 503 166 746 173
rect 503 151 533 166
rect 716 151 746 166
rect 1002 173 1250 189
rect 1326 239 1366 282
rect 1450 251 1466 285
rect 1500 265 1564 285
rect 1631 282 1667 297
rect 1737 282 1773 297
rect 1842 295 1878 333
rect 1840 285 1954 295
rect 1629 265 1669 282
rect 1735 265 1775 282
rect 1840 265 1904 285
rect 1500 251 1516 265
rect 1450 241 1516 251
rect 1621 249 1675 265
rect 1326 223 1380 239
rect 1326 189 1336 223
rect 1370 196 1380 223
rect 1621 215 1631 249
rect 1665 215 1675 249
rect 1621 199 1675 215
rect 1729 249 1783 265
rect 1729 215 1739 249
rect 1773 215 1783 249
rect 1888 251 1904 265
rect 1938 251 1954 285
rect 2040 282 2076 297
rect 2156 282 2192 297
rect 2354 295 2390 333
rect 2278 285 2392 295
rect 1888 241 1954 251
rect 2038 239 2078 282
rect 1729 199 1783 215
rect 2024 223 2078 239
rect 1370 189 1574 196
rect 1326 173 1574 189
rect 1639 177 1669 199
rect 1735 177 1765 199
rect 2024 196 2034 223
rect 1830 189 2034 196
rect 2068 189 2078 223
rect 1002 166 1245 173
rect 1002 151 1032 166
rect 1215 151 1245 166
rect 1331 166 1574 173
rect 1331 151 1361 166
rect 1544 151 1574 166
rect 1830 173 2078 189
rect 2154 239 2194 282
rect 2278 251 2294 285
rect 2328 265 2392 285
rect 2459 282 2495 297
rect 2565 282 2601 297
rect 2670 295 2706 333
rect 2668 285 2782 295
rect 2457 265 2497 282
rect 2563 265 2603 282
rect 2668 265 2732 285
rect 2328 251 2344 265
rect 2278 241 2344 251
rect 2449 249 2503 265
rect 2154 223 2208 239
rect 2154 189 2164 223
rect 2198 196 2208 223
rect 2449 215 2459 249
rect 2493 215 2503 249
rect 2449 199 2503 215
rect 2557 249 2611 265
rect 2557 215 2567 249
rect 2601 215 2611 249
rect 2716 251 2732 265
rect 2766 251 2782 285
rect 2868 282 2904 297
rect 2984 282 3020 297
rect 3182 295 3218 333
rect 3106 285 3220 295
rect 2716 241 2782 251
rect 2866 239 2906 282
rect 2557 199 2611 215
rect 2852 223 2906 239
rect 2198 189 2402 196
rect 2154 173 2402 189
rect 2467 177 2497 199
rect 2563 177 2593 199
rect 2852 196 2862 223
rect 2658 189 2862 196
rect 2896 189 2906 223
rect 1830 166 2073 173
rect 1830 151 1860 166
rect 2043 151 2073 166
rect 2159 166 2402 173
rect 2159 151 2189 166
rect 2372 151 2402 166
rect 2658 173 2906 189
rect 2982 239 3022 282
rect 3106 251 3122 285
rect 3156 265 3220 285
rect 3287 282 3323 297
rect 3285 265 3325 282
rect 3156 251 3172 265
rect 3106 241 3172 251
rect 3277 249 3331 265
rect 2982 223 3036 239
rect 2982 189 2992 223
rect 3026 196 3036 223
rect 3277 215 3287 249
rect 3321 215 3331 249
rect 3277 199 3331 215
rect 3026 189 3230 196
rect 2982 173 3230 189
rect 3295 177 3325 199
rect 2658 166 2901 173
rect 2658 151 2688 166
rect 2871 151 2901 166
rect 2987 166 3230 173
rect 2987 151 3017 166
rect 3200 151 3230 166
rect 79 21 109 47
rect 174 21 204 47
rect 387 21 417 47
rect 503 21 533 47
rect 716 21 746 47
rect 811 21 841 47
rect 907 21 937 47
rect 1002 21 1032 47
rect 1215 21 1245 47
rect 1331 21 1361 47
rect 1544 21 1574 47
rect 1639 21 1669 47
rect 1735 21 1765 47
rect 1830 21 1860 47
rect 2043 21 2073 47
rect 2159 21 2189 47
rect 2372 21 2402 47
rect 2467 21 2497 47
rect 2563 21 2593 47
rect 2658 21 2688 47
rect 2871 21 2901 47
rect 2987 21 3017 47
rect 3200 21 3230 47
rect 3295 21 3325 47
<< polycont >>
rect 83 839 117 873
rect 378 865 412 899
rect 248 803 282 837
rect 508 865 542 899
rect 638 803 672 837
rect 803 839 837 873
rect 911 839 945 873
rect 1206 865 1240 899
rect 1076 803 1110 837
rect 1336 865 1370 899
rect 1466 803 1500 837
rect 1631 839 1665 873
rect 1739 839 1773 873
rect 2034 865 2068 899
rect 1904 803 1938 837
rect 2164 865 2198 899
rect 2294 803 2328 837
rect 2459 839 2493 873
rect 2567 839 2601 873
rect 2862 865 2896 899
rect 2732 803 2766 837
rect 2992 865 3026 899
rect 3122 803 3156 837
rect 3287 839 3321 873
rect 83 215 117 249
rect 248 251 282 285
rect 378 189 412 223
rect 638 251 672 285
rect 508 189 542 223
rect 803 215 837 249
rect 911 215 945 249
rect 1076 251 1110 285
rect 1206 189 1240 223
rect 1466 251 1500 285
rect 1336 189 1370 223
rect 1631 215 1665 249
rect 1739 215 1773 249
rect 1904 251 1938 285
rect 2034 189 2068 223
rect 2294 251 2328 285
rect 2164 189 2198 223
rect 2459 215 2493 249
rect 2567 215 2601 249
rect 2732 251 2766 285
rect 2862 189 2896 223
rect 3122 251 3156 285
rect 2992 189 3026 223
rect 3287 215 3321 249
<< locali >>
rect 0 1071 29 1105
rect 63 1071 121 1105
rect 155 1071 213 1105
rect 247 1071 305 1105
rect 339 1071 397 1105
rect 431 1071 489 1105
rect 523 1071 581 1105
rect 615 1071 673 1105
rect 707 1071 765 1105
rect 799 1071 857 1105
rect 891 1071 949 1105
rect 983 1071 1041 1105
rect 1075 1071 1133 1105
rect 1167 1071 1225 1105
rect 1259 1071 1317 1105
rect 1351 1071 1409 1105
rect 1443 1071 1501 1105
rect 1535 1071 1593 1105
rect 1627 1071 1685 1105
rect 1719 1071 1777 1105
rect 1811 1071 1869 1105
rect 1903 1071 1961 1105
rect 1995 1071 2053 1105
rect 2087 1071 2145 1105
rect 2179 1071 2237 1105
rect 2271 1071 2329 1105
rect 2363 1071 2421 1105
rect 2455 1071 2513 1105
rect 2547 1071 2605 1105
rect 2639 1071 2697 1105
rect 2731 1071 2789 1105
rect 2823 1071 2881 1105
rect 2915 1071 2973 1105
rect 3007 1071 3065 1105
rect 3099 1071 3157 1105
rect 3191 1071 3249 1105
rect 3283 1071 3341 1105
rect 3375 1071 3404 1105
rect 26 1029 78 1071
rect 26 995 35 1029
rect 69 995 78 1029
rect 26 961 78 995
rect 26 927 35 961
rect 69 927 78 961
rect 26 911 78 927
rect 112 963 167 1009
rect 209 1006 258 1022
rect 209 972 214 1006
rect 248 972 258 1006
rect 112 877 146 963
rect 209 921 258 972
rect 330 1006 380 1022
rect 330 972 338 1006
rect 372 972 380 1006
rect 330 971 380 972
rect 67 873 146 877
rect 67 839 83 873
rect 117 839 146 873
rect 67 823 146 839
rect 180 887 258 921
rect 292 937 380 971
rect 427 1006 493 1071
rect 842 1029 906 1071
rect 427 972 443 1006
rect 477 972 493 1006
rect 427 956 493 972
rect 540 1006 590 1022
rect 540 972 548 1006
rect 582 972 590 1006
rect 540 971 590 972
rect 662 1006 711 1022
rect 662 972 672 1006
rect 706 972 711 1006
rect 540 937 628 971
rect 19 773 85 789
rect 19 739 35 773
rect 69 739 85 773
rect 19 705 85 739
rect 19 671 35 705
rect 69 671 85 705
rect 180 737 214 887
rect 292 853 326 937
rect 248 837 326 853
rect 282 803 326 837
rect 361 865 378 899
rect 412 865 441 899
rect 361 829 441 865
rect 479 865 508 899
rect 542 865 559 899
rect 479 829 559 865
rect 594 853 628 937
rect 662 921 711 972
rect 753 963 808 1009
rect 662 887 740 921
rect 594 837 672 853
rect 248 795 326 803
rect 594 803 638 837
rect 594 795 672 803
rect 248 787 388 795
rect 292 779 388 787
rect 292 761 338 779
rect 322 745 338 761
rect 372 745 388 779
rect 180 731 259 737
rect 180 697 213 731
rect 247 727 259 731
rect 247 705 284 727
rect 180 691 234 697
rect 19 637 85 671
rect 19 603 35 637
rect 69 603 85 637
rect 19 561 85 603
rect 218 671 234 691
rect 268 671 284 705
rect 218 637 284 671
rect 218 603 234 637
rect 268 603 284 637
rect 218 595 284 603
rect 322 711 388 745
rect 322 677 338 711
rect 372 677 388 711
rect 322 643 388 677
rect 322 609 338 643
rect 372 609 388 643
rect 322 595 388 609
rect 427 779 493 795
rect 427 745 443 779
rect 477 745 493 779
rect 427 711 493 745
rect 427 677 443 711
rect 477 677 493 711
rect 427 643 493 677
rect 427 609 443 643
rect 477 609 493 643
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 184 561
rect 19 485 85 527
rect 19 451 35 485
rect 69 451 85 485
rect 19 417 85 451
rect 19 383 35 417
rect 69 383 85 417
rect 218 493 259 595
rect 427 561 493 609
rect 532 787 672 795
rect 532 779 628 787
rect 532 745 548 779
rect 582 761 628 779
rect 582 745 598 761
rect 532 711 598 745
rect 706 737 740 887
rect 774 877 808 963
rect 842 995 857 1029
rect 891 995 906 1029
rect 842 961 906 995
rect 842 927 857 961
rect 891 927 906 961
rect 842 911 906 927
rect 940 963 995 1009
rect 1037 1006 1086 1022
rect 1037 972 1042 1006
rect 1076 972 1086 1006
rect 940 877 974 963
rect 1037 921 1086 972
rect 1158 1006 1208 1022
rect 1158 972 1166 1006
rect 1200 972 1208 1006
rect 1158 971 1208 972
rect 774 873 853 877
rect 774 839 803 873
rect 837 839 853 873
rect 774 823 853 839
rect 895 873 974 877
rect 895 839 911 873
rect 945 839 974 873
rect 895 823 974 839
rect 1008 887 1086 921
rect 1120 937 1208 971
rect 1255 1006 1321 1071
rect 1670 1029 1734 1071
rect 1255 972 1271 1006
rect 1305 972 1321 1006
rect 1255 956 1321 972
rect 1368 1006 1418 1022
rect 1368 972 1376 1006
rect 1410 972 1418 1006
rect 1368 971 1418 972
rect 1490 1006 1539 1022
rect 1490 972 1500 1006
rect 1534 972 1539 1006
rect 1368 937 1456 971
rect 661 731 740 737
rect 661 727 673 731
rect 532 677 548 711
rect 582 677 598 711
rect 532 643 598 677
rect 532 609 548 643
rect 582 609 598 643
rect 532 595 598 609
rect 636 705 673 727
rect 636 671 652 705
rect 707 697 740 731
rect 686 691 740 697
rect 835 773 913 789
rect 835 739 857 773
rect 891 739 913 773
rect 835 705 913 739
rect 686 671 702 691
rect 636 637 702 671
rect 636 603 652 637
rect 686 603 702 637
rect 636 595 702 603
rect 293 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 627 561
rect 218 485 284 493
rect 218 451 234 485
rect 268 451 284 485
rect 218 417 284 451
rect 218 397 234 417
rect 19 349 85 383
rect 19 315 35 349
rect 69 315 85 349
rect 19 299 85 315
rect 180 391 234 397
rect 180 357 213 391
rect 268 383 284 417
rect 247 361 284 383
rect 322 479 388 493
rect 322 445 338 479
rect 372 445 388 479
rect 322 411 388 445
rect 322 377 338 411
rect 372 377 388 411
rect 247 357 259 361
rect 180 351 259 357
rect 67 249 146 265
rect 67 215 83 249
rect 117 215 146 249
rect 67 211 146 215
rect 26 161 78 177
rect 26 127 35 161
rect 69 127 78 161
rect 26 93 78 127
rect 26 59 35 93
rect 69 59 78 93
rect 112 125 146 211
rect 180 201 214 351
rect 322 343 388 377
rect 322 327 338 343
rect 292 309 338 327
rect 372 309 388 343
rect 292 301 388 309
rect 248 293 388 301
rect 427 479 493 527
rect 661 493 702 595
rect 835 671 857 705
rect 891 671 913 705
rect 1008 737 1042 887
rect 1120 853 1154 937
rect 1076 837 1154 853
rect 1110 803 1154 837
rect 1189 865 1206 899
rect 1240 865 1269 899
rect 1189 829 1269 865
rect 1307 865 1336 899
rect 1370 865 1387 899
rect 1307 829 1387 865
rect 1422 853 1456 937
rect 1490 921 1539 972
rect 1581 963 1636 1009
rect 1490 887 1568 921
rect 1422 837 1500 853
rect 1076 795 1154 803
rect 1422 803 1466 837
rect 1422 795 1500 803
rect 1076 787 1216 795
rect 1120 779 1216 787
rect 1120 761 1166 779
rect 1150 745 1166 761
rect 1200 745 1216 779
rect 1008 731 1087 737
rect 1008 697 1041 731
rect 1075 727 1087 731
rect 1075 705 1112 727
rect 1008 691 1062 697
rect 835 637 913 671
rect 835 603 857 637
rect 891 603 913 637
rect 835 561 913 603
rect 1046 671 1062 691
rect 1096 671 1112 705
rect 1046 637 1112 671
rect 1046 603 1062 637
rect 1096 603 1112 637
rect 1046 595 1112 603
rect 1150 711 1216 745
rect 1150 677 1166 711
rect 1200 677 1216 711
rect 1150 643 1216 677
rect 1150 609 1166 643
rect 1200 609 1216 643
rect 1150 595 1216 609
rect 1255 779 1321 795
rect 1255 745 1271 779
rect 1305 745 1321 779
rect 1255 711 1321 745
rect 1255 677 1271 711
rect 1305 677 1321 711
rect 1255 643 1321 677
rect 1255 609 1271 643
rect 1305 609 1321 643
rect 736 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 427 445 443 479
rect 477 445 493 479
rect 427 411 493 445
rect 427 377 443 411
rect 477 377 493 411
rect 427 343 493 377
rect 427 309 443 343
rect 477 309 493 343
rect 427 293 493 309
rect 532 479 598 493
rect 532 445 548 479
rect 582 445 598 479
rect 532 411 598 445
rect 532 377 548 411
rect 582 377 598 411
rect 532 343 598 377
rect 636 485 702 493
rect 636 451 652 485
rect 686 451 702 485
rect 636 417 702 451
rect 636 383 652 417
rect 686 397 702 417
rect 835 485 913 527
rect 835 451 857 485
rect 891 451 913 485
rect 835 417 913 451
rect 686 391 740 397
rect 636 361 673 383
rect 661 357 673 361
rect 707 357 740 391
rect 661 351 740 357
rect 532 309 548 343
rect 582 327 598 343
rect 582 309 628 327
rect 532 301 628 309
rect 532 293 672 301
rect 248 285 326 293
rect 282 251 326 285
rect 594 285 672 293
rect 248 235 326 251
rect 180 167 258 201
rect 112 79 167 125
rect 209 116 258 167
rect 292 151 326 235
rect 361 223 441 259
rect 361 189 378 223
rect 412 189 441 223
rect 479 223 559 259
rect 479 189 508 223
rect 542 189 559 223
rect 594 251 638 285
rect 594 235 672 251
rect 594 151 628 235
rect 706 201 740 351
rect 835 383 857 417
rect 891 383 913 417
rect 1046 493 1087 595
rect 1255 561 1321 609
rect 1360 787 1500 795
rect 1360 779 1456 787
rect 1360 745 1376 779
rect 1410 761 1456 779
rect 1410 745 1426 761
rect 1360 711 1426 745
rect 1534 737 1568 887
rect 1602 877 1636 963
rect 1670 995 1685 1029
rect 1719 995 1734 1029
rect 1670 961 1734 995
rect 1670 927 1685 961
rect 1719 927 1734 961
rect 1670 911 1734 927
rect 1768 963 1823 1009
rect 1865 1006 1914 1022
rect 1865 972 1870 1006
rect 1904 972 1914 1006
rect 1768 877 1802 963
rect 1865 921 1914 972
rect 1986 1006 2036 1022
rect 1986 972 1994 1006
rect 2028 972 2036 1006
rect 1986 971 2036 972
rect 1602 873 1681 877
rect 1602 839 1631 873
rect 1665 839 1681 873
rect 1602 823 1681 839
rect 1723 873 1802 877
rect 1723 839 1739 873
rect 1773 839 1802 873
rect 1723 823 1802 839
rect 1836 887 1914 921
rect 1948 937 2036 971
rect 2083 1006 2149 1071
rect 2498 1029 2562 1071
rect 2083 972 2099 1006
rect 2133 972 2149 1006
rect 2083 956 2149 972
rect 2196 1006 2246 1022
rect 2196 972 2204 1006
rect 2238 972 2246 1006
rect 2196 971 2246 972
rect 2318 1006 2367 1022
rect 2318 972 2328 1006
rect 2362 972 2367 1006
rect 2196 937 2284 971
rect 1489 731 1568 737
rect 1489 727 1501 731
rect 1360 677 1376 711
rect 1410 677 1426 711
rect 1360 643 1426 677
rect 1360 609 1376 643
rect 1410 609 1426 643
rect 1360 595 1426 609
rect 1464 705 1501 727
rect 1464 671 1480 705
rect 1535 697 1568 731
rect 1514 691 1568 697
rect 1663 773 1741 789
rect 1663 739 1685 773
rect 1719 739 1741 773
rect 1663 705 1741 739
rect 1514 671 1530 691
rect 1464 637 1530 671
rect 1464 603 1480 637
rect 1514 603 1530 637
rect 1464 595 1530 603
rect 1121 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1455 561
rect 1046 485 1112 493
rect 1046 451 1062 485
rect 1096 451 1112 485
rect 1046 417 1112 451
rect 1046 397 1062 417
rect 835 349 913 383
rect 835 315 857 349
rect 891 315 913 349
rect 835 299 913 315
rect 1008 391 1062 397
rect 1008 357 1041 391
rect 1096 383 1112 417
rect 1075 361 1112 383
rect 1150 479 1216 493
rect 1150 445 1166 479
rect 1200 445 1216 479
rect 1150 411 1216 445
rect 1150 377 1166 411
rect 1200 377 1216 411
rect 1075 357 1087 361
rect 1008 351 1087 357
rect 292 117 380 151
rect 209 82 214 116
rect 248 82 258 116
rect 209 66 258 82
rect 330 116 380 117
rect 330 82 338 116
rect 372 82 380 116
rect 330 66 380 82
rect 427 116 493 132
rect 427 82 443 116
rect 477 82 493 116
rect 26 17 78 59
rect 427 17 493 82
rect 540 117 628 151
rect 662 167 740 201
rect 774 249 853 265
rect 774 215 803 249
rect 837 215 853 249
rect 774 211 853 215
rect 895 249 974 265
rect 895 215 911 249
rect 945 215 974 249
rect 895 211 974 215
rect 540 116 590 117
rect 540 82 548 116
rect 582 82 590 116
rect 540 66 590 82
rect 662 116 711 167
rect 774 125 808 211
rect 662 82 672 116
rect 706 82 711 116
rect 662 66 711 82
rect 753 79 808 125
rect 842 161 906 177
rect 842 127 857 161
rect 891 127 906 161
rect 842 93 906 127
rect 842 59 857 93
rect 891 59 906 93
rect 940 125 974 211
rect 1008 201 1042 351
rect 1150 343 1216 377
rect 1150 327 1166 343
rect 1120 309 1166 327
rect 1200 309 1216 343
rect 1120 301 1216 309
rect 1076 293 1216 301
rect 1255 479 1321 527
rect 1489 493 1530 595
rect 1663 671 1685 705
rect 1719 671 1741 705
rect 1836 737 1870 887
rect 1948 853 1982 937
rect 1904 837 1982 853
rect 1938 803 1982 837
rect 2017 865 2034 899
rect 2068 865 2097 899
rect 2017 829 2097 865
rect 2135 865 2164 899
rect 2198 865 2215 899
rect 2135 829 2215 865
rect 2250 853 2284 937
rect 2318 921 2367 972
rect 2409 963 2464 1009
rect 2318 887 2396 921
rect 2250 837 2328 853
rect 1904 795 1982 803
rect 2250 803 2294 837
rect 2250 795 2328 803
rect 1904 787 2044 795
rect 1948 779 2044 787
rect 1948 761 1994 779
rect 1978 745 1994 761
rect 2028 745 2044 779
rect 1836 731 1915 737
rect 1836 697 1869 731
rect 1903 727 1915 731
rect 1903 705 1940 727
rect 1836 691 1890 697
rect 1663 637 1741 671
rect 1663 603 1685 637
rect 1719 603 1741 637
rect 1663 561 1741 603
rect 1874 671 1890 691
rect 1924 671 1940 705
rect 1874 637 1940 671
rect 1874 603 1890 637
rect 1924 603 1940 637
rect 1874 595 1940 603
rect 1978 711 2044 745
rect 1978 677 1994 711
rect 2028 677 2044 711
rect 1978 643 2044 677
rect 1978 609 1994 643
rect 2028 609 2044 643
rect 1978 595 2044 609
rect 2083 779 2149 795
rect 2083 745 2099 779
rect 2133 745 2149 779
rect 2083 711 2149 745
rect 2083 677 2099 711
rect 2133 677 2149 711
rect 2083 643 2149 677
rect 2083 609 2099 643
rect 2133 609 2149 643
rect 1564 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 1255 445 1271 479
rect 1305 445 1321 479
rect 1255 411 1321 445
rect 1255 377 1271 411
rect 1305 377 1321 411
rect 1255 343 1321 377
rect 1255 309 1271 343
rect 1305 309 1321 343
rect 1255 293 1321 309
rect 1360 479 1426 493
rect 1360 445 1376 479
rect 1410 445 1426 479
rect 1360 411 1426 445
rect 1360 377 1376 411
rect 1410 377 1426 411
rect 1360 343 1426 377
rect 1464 485 1530 493
rect 1464 451 1480 485
rect 1514 451 1530 485
rect 1464 417 1530 451
rect 1464 383 1480 417
rect 1514 397 1530 417
rect 1663 485 1741 527
rect 1663 451 1685 485
rect 1719 451 1741 485
rect 1663 417 1741 451
rect 1514 391 1568 397
rect 1464 361 1501 383
rect 1489 357 1501 361
rect 1535 357 1568 391
rect 1489 351 1568 357
rect 1360 309 1376 343
rect 1410 327 1426 343
rect 1410 309 1456 327
rect 1360 301 1456 309
rect 1360 293 1500 301
rect 1076 285 1154 293
rect 1110 251 1154 285
rect 1422 285 1500 293
rect 1076 235 1154 251
rect 1008 167 1086 201
rect 940 79 995 125
rect 1037 116 1086 167
rect 1120 151 1154 235
rect 1189 223 1269 259
rect 1189 189 1206 223
rect 1240 189 1269 223
rect 1307 223 1387 259
rect 1307 189 1336 223
rect 1370 189 1387 223
rect 1422 251 1466 285
rect 1422 235 1500 251
rect 1422 151 1456 235
rect 1534 201 1568 351
rect 1663 383 1685 417
rect 1719 383 1741 417
rect 1874 493 1915 595
rect 2083 561 2149 609
rect 2188 787 2328 795
rect 2188 779 2284 787
rect 2188 745 2204 779
rect 2238 761 2284 779
rect 2238 745 2254 761
rect 2188 711 2254 745
rect 2362 737 2396 887
rect 2430 877 2464 963
rect 2498 995 2513 1029
rect 2547 995 2562 1029
rect 2498 961 2562 995
rect 2498 927 2513 961
rect 2547 927 2562 961
rect 2498 911 2562 927
rect 2596 963 2651 1009
rect 2693 1006 2742 1022
rect 2693 972 2698 1006
rect 2732 972 2742 1006
rect 2596 877 2630 963
rect 2693 921 2742 972
rect 2814 1006 2864 1022
rect 2814 972 2822 1006
rect 2856 972 2864 1006
rect 2814 971 2864 972
rect 2430 873 2509 877
rect 2430 839 2459 873
rect 2493 839 2509 873
rect 2430 823 2509 839
rect 2551 873 2630 877
rect 2551 839 2567 873
rect 2601 839 2630 873
rect 2551 823 2630 839
rect 2664 887 2742 921
rect 2776 937 2864 971
rect 2911 1006 2977 1071
rect 3326 1029 3378 1071
rect 2911 972 2927 1006
rect 2961 972 2977 1006
rect 2911 956 2977 972
rect 3024 1006 3074 1022
rect 3024 972 3032 1006
rect 3066 972 3074 1006
rect 3024 971 3074 972
rect 3146 1006 3195 1022
rect 3146 972 3156 1006
rect 3190 972 3195 1006
rect 3024 937 3112 971
rect 2317 731 2396 737
rect 2317 727 2329 731
rect 2188 677 2204 711
rect 2238 677 2254 711
rect 2188 643 2254 677
rect 2188 609 2204 643
rect 2238 609 2254 643
rect 2188 595 2254 609
rect 2292 705 2329 727
rect 2292 671 2308 705
rect 2363 697 2396 731
rect 2342 691 2396 697
rect 2491 773 2569 789
rect 2491 739 2513 773
rect 2547 739 2569 773
rect 2491 705 2569 739
rect 2342 671 2358 691
rect 2292 637 2358 671
rect 2292 603 2308 637
rect 2342 603 2358 637
rect 2292 595 2358 603
rect 1949 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2283 561
rect 1874 485 1940 493
rect 1874 451 1890 485
rect 1924 451 1940 485
rect 1874 417 1940 451
rect 1874 397 1890 417
rect 1663 349 1741 383
rect 1663 315 1685 349
rect 1719 315 1741 349
rect 1663 299 1741 315
rect 1836 391 1890 397
rect 1836 357 1869 391
rect 1924 383 1940 417
rect 1903 361 1940 383
rect 1978 479 2044 493
rect 1978 445 1994 479
rect 2028 445 2044 479
rect 1978 411 2044 445
rect 1978 377 1994 411
rect 2028 377 2044 411
rect 1903 357 1915 361
rect 1836 351 1915 357
rect 1120 117 1208 151
rect 1037 82 1042 116
rect 1076 82 1086 116
rect 1037 66 1086 82
rect 1158 116 1208 117
rect 1158 82 1166 116
rect 1200 82 1208 116
rect 1158 66 1208 82
rect 1255 116 1321 132
rect 1255 82 1271 116
rect 1305 82 1321 116
rect 842 17 906 59
rect 1255 17 1321 82
rect 1368 117 1456 151
rect 1490 167 1568 201
rect 1602 249 1681 265
rect 1602 215 1631 249
rect 1665 215 1681 249
rect 1602 211 1681 215
rect 1723 249 1802 265
rect 1723 215 1739 249
rect 1773 215 1802 249
rect 1723 211 1802 215
rect 1368 116 1418 117
rect 1368 82 1376 116
rect 1410 82 1418 116
rect 1368 66 1418 82
rect 1490 116 1539 167
rect 1602 125 1636 211
rect 1490 82 1500 116
rect 1534 82 1539 116
rect 1490 66 1539 82
rect 1581 79 1636 125
rect 1670 161 1734 177
rect 1670 127 1685 161
rect 1719 127 1734 161
rect 1670 93 1734 127
rect 1670 59 1685 93
rect 1719 59 1734 93
rect 1768 125 1802 211
rect 1836 201 1870 351
rect 1978 343 2044 377
rect 1978 327 1994 343
rect 1948 309 1994 327
rect 2028 309 2044 343
rect 1948 301 2044 309
rect 1904 293 2044 301
rect 2083 479 2149 527
rect 2317 493 2358 595
rect 2491 671 2513 705
rect 2547 671 2569 705
rect 2664 737 2698 887
rect 2776 853 2810 937
rect 2732 837 2810 853
rect 2766 803 2810 837
rect 2845 865 2862 899
rect 2896 865 2925 899
rect 2845 829 2925 865
rect 2963 865 2992 899
rect 3026 865 3043 899
rect 2963 829 3043 865
rect 3078 853 3112 937
rect 3146 921 3195 972
rect 3237 963 3292 1009
rect 3146 887 3224 921
rect 3078 837 3156 853
rect 2732 795 2810 803
rect 3078 803 3122 837
rect 3078 795 3156 803
rect 2732 787 2872 795
rect 2776 779 2872 787
rect 2776 761 2822 779
rect 2806 745 2822 761
rect 2856 745 2872 779
rect 2664 731 2743 737
rect 2664 697 2697 731
rect 2731 727 2743 731
rect 2731 705 2768 727
rect 2664 691 2718 697
rect 2491 637 2569 671
rect 2491 603 2513 637
rect 2547 603 2569 637
rect 2491 561 2569 603
rect 2702 671 2718 691
rect 2752 671 2768 705
rect 2702 637 2768 671
rect 2702 603 2718 637
rect 2752 603 2768 637
rect 2702 595 2768 603
rect 2806 711 2872 745
rect 2806 677 2822 711
rect 2856 677 2872 711
rect 2806 643 2872 677
rect 2806 609 2822 643
rect 2856 609 2872 643
rect 2806 595 2872 609
rect 2911 779 2977 795
rect 2911 745 2927 779
rect 2961 745 2977 779
rect 2911 711 2977 745
rect 2911 677 2927 711
rect 2961 677 2977 711
rect 2911 643 2977 677
rect 2911 609 2927 643
rect 2961 609 2977 643
rect 2392 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2668 561
rect 2083 445 2099 479
rect 2133 445 2149 479
rect 2083 411 2149 445
rect 2083 377 2099 411
rect 2133 377 2149 411
rect 2083 343 2149 377
rect 2083 309 2099 343
rect 2133 309 2149 343
rect 2083 293 2149 309
rect 2188 479 2254 493
rect 2188 445 2204 479
rect 2238 445 2254 479
rect 2188 411 2254 445
rect 2188 377 2204 411
rect 2238 377 2254 411
rect 2188 343 2254 377
rect 2292 485 2358 493
rect 2292 451 2308 485
rect 2342 451 2358 485
rect 2292 417 2358 451
rect 2292 383 2308 417
rect 2342 397 2358 417
rect 2491 485 2569 527
rect 2491 451 2513 485
rect 2547 451 2569 485
rect 2491 417 2569 451
rect 2342 391 2396 397
rect 2292 361 2329 383
rect 2317 357 2329 361
rect 2363 357 2396 391
rect 2317 351 2396 357
rect 2188 309 2204 343
rect 2238 327 2254 343
rect 2238 309 2284 327
rect 2188 301 2284 309
rect 2188 293 2328 301
rect 1904 285 1982 293
rect 1938 251 1982 285
rect 2250 285 2328 293
rect 1904 235 1982 251
rect 1836 167 1914 201
rect 1768 79 1823 125
rect 1865 116 1914 167
rect 1948 151 1982 235
rect 2017 223 2097 259
rect 2017 189 2034 223
rect 2068 189 2097 223
rect 2135 223 2215 259
rect 2135 189 2164 223
rect 2198 189 2215 223
rect 2250 251 2294 285
rect 2250 235 2328 251
rect 2250 151 2284 235
rect 2362 201 2396 351
rect 2491 383 2513 417
rect 2547 383 2569 417
rect 2702 493 2743 595
rect 2911 561 2977 609
rect 3016 787 3156 795
rect 3016 779 3112 787
rect 3016 745 3032 779
rect 3066 761 3112 779
rect 3066 745 3082 761
rect 3016 711 3082 745
rect 3190 737 3224 887
rect 3258 877 3292 963
rect 3326 995 3335 1029
rect 3369 995 3378 1029
rect 3326 961 3378 995
rect 3326 927 3335 961
rect 3369 927 3378 961
rect 3326 911 3378 927
rect 3258 873 3337 877
rect 3258 839 3287 873
rect 3321 839 3337 873
rect 3258 823 3337 839
rect 3145 731 3224 737
rect 3145 727 3157 731
rect 3016 677 3032 711
rect 3066 677 3082 711
rect 3016 643 3082 677
rect 3016 609 3032 643
rect 3066 609 3082 643
rect 3016 595 3082 609
rect 3120 705 3157 727
rect 3120 671 3136 705
rect 3191 697 3224 731
rect 3170 691 3224 697
rect 3319 773 3385 789
rect 3319 739 3335 773
rect 3369 739 3385 773
rect 3319 705 3385 739
rect 3170 671 3186 691
rect 3120 637 3186 671
rect 3120 603 3136 637
rect 3170 603 3186 637
rect 3120 595 3186 603
rect 2777 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3111 561
rect 2702 485 2768 493
rect 2702 451 2718 485
rect 2752 451 2768 485
rect 2702 417 2768 451
rect 2702 397 2718 417
rect 2491 349 2569 383
rect 2491 315 2513 349
rect 2547 315 2569 349
rect 2491 299 2569 315
rect 2664 391 2718 397
rect 2664 357 2697 391
rect 2752 383 2768 417
rect 2731 361 2768 383
rect 2806 479 2872 493
rect 2806 445 2822 479
rect 2856 445 2872 479
rect 2806 411 2872 445
rect 2806 377 2822 411
rect 2856 377 2872 411
rect 2731 357 2743 361
rect 2664 351 2743 357
rect 1948 117 2036 151
rect 1865 82 1870 116
rect 1904 82 1914 116
rect 1865 66 1914 82
rect 1986 116 2036 117
rect 1986 82 1994 116
rect 2028 82 2036 116
rect 1986 66 2036 82
rect 2083 116 2149 132
rect 2083 82 2099 116
rect 2133 82 2149 116
rect 1670 17 1734 59
rect 2083 17 2149 82
rect 2196 117 2284 151
rect 2318 167 2396 201
rect 2430 249 2509 265
rect 2430 215 2459 249
rect 2493 215 2509 249
rect 2430 211 2509 215
rect 2551 249 2630 265
rect 2551 215 2567 249
rect 2601 215 2630 249
rect 2551 211 2630 215
rect 2196 116 2246 117
rect 2196 82 2204 116
rect 2238 82 2246 116
rect 2196 66 2246 82
rect 2318 116 2367 167
rect 2430 125 2464 211
rect 2318 82 2328 116
rect 2362 82 2367 116
rect 2318 66 2367 82
rect 2409 79 2464 125
rect 2498 161 2562 177
rect 2498 127 2513 161
rect 2547 127 2562 161
rect 2498 93 2562 127
rect 2498 59 2513 93
rect 2547 59 2562 93
rect 2596 125 2630 211
rect 2664 201 2698 351
rect 2806 343 2872 377
rect 2806 327 2822 343
rect 2776 309 2822 327
rect 2856 309 2872 343
rect 2776 301 2872 309
rect 2732 293 2872 301
rect 2911 479 2977 527
rect 3145 493 3186 595
rect 3319 671 3335 705
rect 3369 671 3385 705
rect 3319 637 3385 671
rect 3319 603 3335 637
rect 3369 603 3385 637
rect 3319 561 3385 603
rect 3220 527 3249 561
rect 3283 527 3341 561
rect 3375 527 3404 561
rect 2911 445 2927 479
rect 2961 445 2977 479
rect 2911 411 2977 445
rect 2911 377 2927 411
rect 2961 377 2977 411
rect 2911 343 2977 377
rect 2911 309 2927 343
rect 2961 309 2977 343
rect 2911 293 2977 309
rect 3016 479 3082 493
rect 3016 445 3032 479
rect 3066 445 3082 479
rect 3016 411 3082 445
rect 3016 377 3032 411
rect 3066 377 3082 411
rect 3016 343 3082 377
rect 3120 485 3186 493
rect 3120 451 3136 485
rect 3170 451 3186 485
rect 3120 417 3186 451
rect 3120 383 3136 417
rect 3170 397 3186 417
rect 3319 485 3385 527
rect 3319 451 3335 485
rect 3369 451 3385 485
rect 3319 417 3385 451
rect 3170 391 3224 397
rect 3120 361 3157 383
rect 3145 357 3157 361
rect 3191 357 3224 391
rect 3145 351 3224 357
rect 3016 309 3032 343
rect 3066 327 3082 343
rect 3066 309 3112 327
rect 3016 301 3112 309
rect 3016 293 3156 301
rect 2732 285 2810 293
rect 2766 251 2810 285
rect 3078 285 3156 293
rect 2732 235 2810 251
rect 2664 167 2742 201
rect 2596 79 2651 125
rect 2693 116 2742 167
rect 2776 151 2810 235
rect 2845 223 2925 259
rect 2845 189 2862 223
rect 2896 189 2925 223
rect 2963 223 3043 259
rect 2963 189 2992 223
rect 3026 189 3043 223
rect 3078 251 3122 285
rect 3078 235 3156 251
rect 3078 151 3112 235
rect 3190 201 3224 351
rect 3319 383 3335 417
rect 3369 383 3385 417
rect 3319 349 3385 383
rect 3319 315 3335 349
rect 3369 315 3385 349
rect 3319 299 3385 315
rect 2776 117 2864 151
rect 2693 82 2698 116
rect 2732 82 2742 116
rect 2693 66 2742 82
rect 2814 116 2864 117
rect 2814 82 2822 116
rect 2856 82 2864 116
rect 2814 66 2864 82
rect 2911 116 2977 132
rect 2911 82 2927 116
rect 2961 82 2977 116
rect 2498 17 2562 59
rect 2911 17 2977 82
rect 3024 117 3112 151
rect 3146 167 3224 201
rect 3258 249 3337 265
rect 3258 215 3287 249
rect 3321 215 3337 249
rect 3258 211 3337 215
rect 3024 116 3074 117
rect 3024 82 3032 116
rect 3066 82 3074 116
rect 3024 66 3074 82
rect 3146 116 3195 167
rect 3258 125 3292 211
rect 3146 82 3156 116
rect 3190 82 3195 116
rect 3146 66 3195 82
rect 3237 79 3292 125
rect 3326 161 3378 177
rect 3326 127 3335 161
rect 3369 127 3378 161
rect 3326 93 3378 127
rect 3326 59 3335 93
rect 3369 59 3378 93
rect 3326 17 3378 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3341 17
rect 3375 -17 3404 17
<< viali >>
rect 29 1071 63 1105
rect 121 1071 155 1105
rect 213 1071 247 1105
rect 305 1071 339 1105
rect 397 1071 431 1105
rect 489 1071 523 1105
rect 581 1071 615 1105
rect 673 1071 707 1105
rect 765 1071 799 1105
rect 857 1071 891 1105
rect 949 1071 983 1105
rect 1041 1071 1075 1105
rect 1133 1071 1167 1105
rect 1225 1071 1259 1105
rect 1317 1071 1351 1105
rect 1409 1071 1443 1105
rect 1501 1071 1535 1105
rect 1593 1071 1627 1105
rect 1685 1071 1719 1105
rect 1777 1071 1811 1105
rect 1869 1071 1903 1105
rect 1961 1071 1995 1105
rect 2053 1071 2087 1105
rect 2145 1071 2179 1105
rect 2237 1071 2271 1105
rect 2329 1071 2363 1105
rect 2421 1071 2455 1105
rect 2513 1071 2547 1105
rect 2605 1071 2639 1105
rect 2697 1071 2731 1105
rect 2789 1071 2823 1105
rect 2881 1071 2915 1105
rect 2973 1071 3007 1105
rect 3065 1071 3099 1105
rect 3157 1071 3191 1105
rect 3249 1071 3283 1105
rect 3341 1071 3375 1105
rect 213 705 247 731
rect 213 697 234 705
rect 234 697 247 705
rect 29 527 63 561
rect 121 527 155 561
rect 673 705 707 731
rect 673 697 686 705
rect 686 697 707 705
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 213 383 234 391
rect 234 383 247 391
rect 213 357 247 383
rect 1041 705 1075 731
rect 1041 697 1062 705
rect 1062 697 1075 705
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 673 383 686 391
rect 686 383 707 391
rect 673 357 707 383
rect 1501 705 1535 731
rect 1501 697 1514 705
rect 1514 697 1535 705
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1041 383 1062 391
rect 1062 383 1075 391
rect 1041 357 1075 383
rect 1869 705 1903 731
rect 1869 697 1890 705
rect 1890 697 1903 705
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1501 383 1514 391
rect 1514 383 1535 391
rect 1501 357 1535 383
rect 2329 705 2363 731
rect 2329 697 2342 705
rect 2342 697 2363 705
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 1869 383 1890 391
rect 1890 383 1903 391
rect 1869 357 1903 383
rect 2697 705 2731 731
rect 2697 697 2718 705
rect 2718 697 2731 705
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2329 383 2342 391
rect 2342 383 2363 391
rect 2329 357 2363 383
rect 3157 705 3191 731
rect 3157 697 3170 705
rect 3170 697 3191 705
rect 2789 527 2823 561
rect 2881 527 2915 561
rect 2973 527 3007 561
rect 3065 527 3099 561
rect 2697 383 2718 391
rect 2718 383 2731 391
rect 2697 357 2731 383
rect 3249 527 3283 561
rect 3341 527 3375 561
rect 3157 383 3170 391
rect 3170 383 3191 391
rect 3157 357 3191 383
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
rect 2881 -17 2915 17
rect 2973 -17 3007 17
rect 3065 -17 3099 17
rect 3157 -17 3191 17
rect 3249 -17 3283 17
rect 3341 -17 3375 17
<< metal1 >>
rect 0 1105 3404 1136
rect 0 1071 29 1105
rect 63 1071 121 1105
rect 155 1071 213 1105
rect 247 1071 305 1105
rect 339 1071 397 1105
rect 431 1071 489 1105
rect 523 1071 581 1105
rect 615 1071 673 1105
rect 707 1071 765 1105
rect 799 1071 857 1105
rect 891 1071 949 1105
rect 983 1071 1041 1105
rect 1075 1071 1133 1105
rect 1167 1071 1225 1105
rect 1259 1071 1317 1105
rect 1351 1071 1409 1105
rect 1443 1071 1501 1105
rect 1535 1071 1593 1105
rect 1627 1071 1685 1105
rect 1719 1071 1777 1105
rect 1811 1071 1869 1105
rect 1903 1071 1961 1105
rect 1995 1071 2053 1105
rect 2087 1071 2145 1105
rect 2179 1071 2237 1105
rect 2271 1071 2329 1105
rect 2363 1071 2421 1105
rect 2455 1071 2513 1105
rect 2547 1071 2605 1105
rect 2639 1071 2697 1105
rect 2731 1071 2789 1105
rect 2823 1071 2881 1105
rect 2915 1071 2973 1105
rect 3007 1071 3065 1105
rect 3099 1071 3157 1105
rect 3191 1071 3249 1105
rect 3283 1071 3341 1105
rect 3375 1071 3404 1105
rect 0 1040 3404 1071
rect 201 731 259 737
rect 201 697 213 731
rect 247 728 259 731
rect 661 731 719 737
rect 661 728 673 731
rect 247 700 673 728
rect 247 697 259 700
rect 201 691 259 697
rect 661 697 673 700
rect 707 728 719 731
rect 1029 731 1087 737
rect 1029 728 1041 731
rect 707 700 1041 728
rect 707 697 719 700
rect 661 691 719 697
rect 1029 697 1041 700
rect 1075 728 1087 731
rect 1489 731 1547 737
rect 1489 728 1501 731
rect 1075 700 1501 728
rect 1075 697 1087 700
rect 1029 691 1087 697
rect 1489 697 1501 700
rect 1535 728 1547 731
rect 1857 731 1915 737
rect 1857 728 1869 731
rect 1535 700 1869 728
rect 1535 697 1547 700
rect 1489 691 1547 697
rect 1857 697 1869 700
rect 1903 728 1915 731
rect 2317 731 2375 737
rect 2317 728 2329 731
rect 1903 700 2329 728
rect 1903 697 1915 700
rect 1857 691 1915 697
rect 2317 697 2329 700
rect 2363 728 2375 731
rect 2685 731 2743 737
rect 2685 728 2697 731
rect 2363 700 2697 728
rect 2363 697 2375 700
rect 2317 691 2375 697
rect 2685 697 2697 700
rect 2731 728 2743 731
rect 3145 731 3203 737
rect 3145 728 3157 731
rect 2731 700 3157 728
rect 2731 697 2743 700
rect 2685 691 2743 697
rect 3145 697 3157 700
rect 3191 697 3203 731
rect 3145 691 3203 697
rect 0 561 3404 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3249 561
rect 3283 527 3341 561
rect 3375 527 3404 561
rect 0 496 3404 527
rect 201 391 259 397
rect 201 357 213 391
rect 247 388 259 391
rect 661 391 719 397
rect 661 388 673 391
rect 247 360 673 388
rect 247 357 259 360
rect 201 351 259 357
rect 661 357 673 360
rect 707 388 719 391
rect 1029 391 1087 397
rect 1029 388 1041 391
rect 707 360 1041 388
rect 707 357 719 360
rect 661 351 719 357
rect 1029 357 1041 360
rect 1075 388 1087 391
rect 1489 391 1547 397
rect 1489 388 1501 391
rect 1075 360 1501 388
rect 1075 357 1087 360
rect 1029 351 1087 357
rect 1489 357 1501 360
rect 1535 388 1547 391
rect 1857 391 1915 397
rect 1857 388 1869 391
rect 1535 360 1869 388
rect 1535 357 1547 360
rect 1489 351 1547 357
rect 1857 357 1869 360
rect 1903 388 1915 391
rect 2317 391 2375 397
rect 2317 388 2329 391
rect 1903 360 2329 388
rect 1903 357 1915 360
rect 1857 351 1915 357
rect 2317 357 2329 360
rect 2363 388 2375 391
rect 2685 391 2743 397
rect 2685 388 2697 391
rect 2363 360 2697 388
rect 2363 357 2375 360
rect 2317 351 2375 357
rect 2685 357 2697 360
rect 2731 388 2743 391
rect 3145 391 3203 397
rect 3145 388 3157 391
rect 2731 360 3157 388
rect 2731 357 2743 360
rect 2685 351 2743 357
rect 3145 357 3157 360
rect 3191 357 3203 391
rect 3145 351 3203 357
rect 0 17 3404 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3341 17
rect 3375 -17 3404 17
rect 0 -48 3404 -17
<< labels >>
rlabel comment s 0 0 0 0 4 muxb16to1_1
flabel metal1 s 213 697 247 731 0 FreeSans 200 0 0 0 Z
port 37 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 33 nsew
flabel metal1 s 213 357 247 391 0 FreeSans 200 0 0 0 Z
port 37 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 36 nsew
flabel metal1 s 29 1071 63 1105 0 FreeSans 200 0 0 0 VGND
port 33 nsew
flabel metal1 s 1501 357 1535 391 0 FreeSans 200 180 0 0 Z
port 37 nsew
flabel metal1 s 1685 527 1719 561 0 FreeSans 200 180 0 0 VPWR
port 36 nsew
flabel metal1 s 1685 -17 1719 17 0 FreeSans 200 180 0 0 VGND
port 33 nsew
flabel metal1 s 1041 357 1075 391 0 FreeSans 200 0 0 0 Z
port 37 nsew
flabel metal1 s 857 527 891 561 0 FreeSans 200 0 0 0 VPWR
port 36 nsew
flabel metal1 s 857 -17 891 17 0 FreeSans 200 0 0 0 VGND
port 33 nsew
flabel metal1 s 1041 697 1075 731 0 FreeSans 200 0 0 0 Z
port 37 nsew
flabel metal1 s 874 544 874 544 0 FreeSans 200 0 0 0 VPWR
port 36 nsew
flabel metal1 s 857 1071 891 1105 0 FreeSans 200 0 0 0 VGND
port 33 nsew
flabel metal1 s 673 357 707 391 0 FreeSans 200 180 0 0 Z
port 37 nsew
flabel metal1 s 874 544 874 544 0 FreeSans 200 180 0 0 VPWR
port 36 nsew
flabel metal1 s 874 0 874 0 0 FreeSans 200 180 0 0 VGND
port 33 nsew
flabel metal1 s 673 697 707 731 0 FreeSans 200 180 0 0 Z
port 37 nsew
flabel metal1 s 874 544 874 544 0 FreeSans 200 180 0 0 VPWR
port 36 nsew
flabel metal1 s 874 1088 874 1088 0 FreeSans 200 180 0 0 VGND
port 33 nsew
flabel metal1 s 230 714 230 714 0 FreeSans 200 0 0 0 Z
port 37 nsew
flabel metal1 s 46 544 46 544 0 FreeSans 200 0 0 0 VPWR
port 36 nsew
flabel metal1 s 46 1088 46 1088 0 FreeSans 200 0 0 0 VGND
port 33 nsew
flabel metal1 s 230 374 230 374 0 FreeSans 200 0 0 0 Z
port 37 nsew
flabel metal1 s 46 544 46 544 0 FreeSans 200 0 0 0 VPWR
port 36 nsew
flabel metal1 s 46 0 46 0 0 FreeSans 200 0 0 0 VGND
port 33 nsew
flabel metal1 s 1501 697 1535 731 0 FreeSans 200 180 0 0 Z
port 37 nsew
flabel metal1 s 1702 544 1702 544 0 FreeSans 200 180 0 0 VPWR
port 36 nsew
flabel metal1 s 1685 1071 1719 1105 0 FreeSans 200 180 0 0 VGND
port 33 nsew
flabel metal1 s 1869 697 1903 731 0 FreeSans 200 0 0 0 Z
port 37 nsew
flabel metal1 s 1702 544 1702 544 0 FreeSans 200 0 0 0 VPWR
port 36 nsew
flabel metal1 s 1702 1088 1702 1088 0 FreeSans 200 0 0 0 VGND
port 33 nsew
flabel metal1 s 1869 357 1903 391 0 FreeSans 200 0 0 0 Z
port 37 nsew
flabel metal1 s 1702 544 1702 544 0 FreeSans 200 0 0 0 VPWR
port 36 nsew
flabel metal1 s 1702 0 1702 0 0 FreeSans 200 0 0 0 VGND
port 33 nsew
flabel metal1 s 2329 357 2363 391 0 FreeSans 200 180 0 0 Z
port 37 nsew
flabel metal1 s 2513 527 2547 561 0 FreeSans 200 180 0 0 VPWR
port 36 nsew
flabel metal1 s 2513 -17 2547 17 0 FreeSans 200 180 0 0 VGND
port 33 nsew
flabel metal1 s 2329 697 2363 731 0 FreeSans 200 180 0 0 Z
port 37 nsew
flabel metal1 s 2530 544 2530 544 0 FreeSans 200 180 0 0 VPWR
port 36 nsew
flabel metal1 s 2513 1071 2547 1105 0 FreeSans 200 180 0 0 VGND
port 33 nsew
flabel metal1 s 2697 697 2731 731 0 FreeSans 200 0 0 0 Z
port 37 nsew
flabel metal1 s 2530 544 2530 544 0 FreeSans 200 0 0 0 VPWR
port 36 nsew
flabel metal1 s 2530 1088 2530 1088 0 FreeSans 200 0 0 0 VGND
port 33 nsew
flabel metal1 s 2697 357 2731 391 0 FreeSans 200 0 0 0 Z
port 37 nsew
flabel metal1 s 2530 544 2530 544 0 FreeSans 200 0 0 0 VPWR
port 36 nsew
flabel metal1 s 2530 0 2530 0 0 FreeSans 200 0 0 0 VGND
port 33 nsew
flabel metal1 s 3157 357 3191 391 0 FreeSans 200 180 0 0 Z
port 37 nsew
flabel metal1 s 3341 527 3375 561 0 FreeSans 200 180 0 0 VPWR
port 36 nsew
flabel metal1 s 3341 -17 3375 17 0 FreeSans 200 180 0 0 VGND
port 33 nsew
flabel metal1 s 3157 697 3191 731 0 FreeSans 200 180 0 0 Z
port 37 nsew
flabel metal1 s 3358 544 3358 544 0 FreeSans 200 180 0 0 VPWR
port 36 nsew
flabel metal1 s 3341 1071 3375 1105 0 FreeSans 200 180 0 0 VGND
port 33 nsew
flabel pwell s 29 1071 63 1105 0 FreeSans 200 0 0 0 VNB
port 34 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 34 nsew
flabel pwell s 1685 -17 1719 17 0 FreeSans 200 180 0 0 VNB
port 34 nsew
flabel pwell s 857 -17 891 17 0 FreeSans 200 0 0 0 VNB
port 34 nsew
flabel pwell s 857 1071 891 1105 0 FreeSans 200 0 0 0 VNB
port 34 nsew
flabel pwell s 874 0 874 0 0 FreeSans 200 180 0 0 VNB
port 34 nsew
flabel pwell s 874 1088 874 1088 0 FreeSans 200 180 0 0 VNB
port 34 nsew
flabel pwell s 46 1088 46 1088 0 FreeSans 200 0 0 0 VNB
port 34 nsew
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
port 34 nsew
flabel pwell s 1685 1071 1719 1105 0 FreeSans 200 180 0 0 VNB
port 34 nsew
flabel pwell s 1702 1088 1702 1088 0 FreeSans 200 0 0 0 VNB
port 34 nsew
flabel pwell s 1702 0 1702 0 0 FreeSans 200 0 0 0 VNB
port 34 nsew
flabel pwell s 2513 -17 2547 17 0 FreeSans 200 180 0 0 VNB
port 34 nsew
flabel pwell s 2513 1071 2547 1105 0 FreeSans 200 180 0 0 VNB
port 34 nsew
flabel pwell s 2530 1088 2530 1088 0 FreeSans 200 0 0 0 VNB
port 34 nsew
flabel pwell s 2530 0 2530 0 0 FreeSans 200 0 0 0 VNB
port 34 nsew
flabel pwell s 3341 -17 3375 17 0 FreeSans 200 180 0 0 VNB
port 34 nsew
flabel pwell s 3341 1071 3375 1105 0 FreeSans 200 180 0 0 VNB
port 34 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 35 nsew
flabel nbase s 1685 527 1719 561 0 FreeSans 200 180 0 0 VPB
port 35 nsew
flabel nbase s 857 527 891 561 0 FreeSans 200 0 0 0 VPB
port 35 nsew
flabel nbase s 874 544 874 544 0 FreeSans 200 0 0 0 VPB
port 35 nsew
flabel nbase s 874 544 874 544 0 FreeSans 200 180 0 0 VPB
port 35 nsew
flabel nbase s 874 544 874 544 0 FreeSans 200 180 0 0 VPB
port 35 nsew
flabel nbase s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
port 35 nsew
flabel nbase s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
port 35 nsew
flabel nbase s 1702 544 1702 544 0 FreeSans 200 180 0 0 VPB
port 35 nsew
flabel nbase s 1702 544 1702 544 0 FreeSans 200 0 0 0 VPB
port 35 nsew
flabel nbase s 1702 544 1702 544 0 FreeSans 200 0 0 0 VPB
port 35 nsew
flabel nbase s 2513 527 2547 561 0 FreeSans 200 180 0 0 VPB
port 35 nsew
flabel nbase s 2530 544 2530 544 0 FreeSans 200 180 0 0 VPB
port 35 nsew
flabel nbase s 2530 544 2530 544 0 FreeSans 200 0 0 0 VPB
port 35 nsew
flabel nbase s 2530 544 2530 544 0 FreeSans 200 0 0 0 VPB
port 35 nsew
flabel nbase s 3341 527 3375 561 0 FreeSans 200 180 0 0 VPB
port 35 nsew
flabel nbase s 3358 544 3358 544 0 FreeSans 200 180 0 0 VPB
port 35 nsew
flabel corelocali s 121 85 155 119 0 FreeSans 200 0 0 0 D[0]
port 16 nsew
flabel corelocali s 2053 833 2087 867 0 FreeSans 200 0 0 0 S[12]
port 20 nsew
flabel corelocali s 2145 833 2179 867 0 FreeSans 200 0 0 0 S[13]
port 19 nsew
flabel corelocali s 397 833 431 867 0 FreeSans 200 0 0 0 S[8]
port 24 nsew
flabel corelocali s 489 833 523 867 0 FreeSans 200 0 0 0 S[9]
port 23 nsew
flabel corelocali s 1225 833 1259 867 0 FreeSans 200 0 0 0 S[10]
port 22 nsew
flabel corelocali s 1317 833 1351 867 0 FreeSans 200 0 0 0 S[11]
port 21 nsew
flabel corelocali s 2881 833 2915 867 0 FreeSans 200 0 0 0 S[14]
port 18 nsew
flabel corelocali s 2973 833 3007 867 0 FreeSans 200 0 0 0 S[15]
port 17 nsew
flabel corelocali s 1777 969 1811 1003 0 FreeSans 200 0 0 0 D[12]
port 4 nsew
flabel corelocali s 765 969 799 1003 0 FreeSans 200 0 0 0 D[9]
port 7 nsew
flabel corelocali s 949 969 983 1003 0 FreeSans 200 0 0 0 D[10]
port 6 nsew
flabel corelocali s 2421 969 2455 1003 0 FreeSans 200 0 0 0 D[13]
port 3 nsew
flabel corelocali s 2605 969 2639 1003 0 FreeSans 200 0 0 0 D[14]
port 2 nsew
flabel corelocali s 3249 969 3283 1003 0 FreeSans 200 0 0 0 D[15]
port 1 nsew
flabel corelocali s 121 969 155 1003 0 FreeSans 200 0 0 0 D[8]
port 8 nsew
flabel corelocali s 1593 969 1627 1003 0 FreeSans 200 0 0 0 D[11]
port 5 nsew
flabel corelocali s 397 221 431 255 0 FreeSans 200 0 0 0 S[0]
port 32 nsew
flabel corelocali s 489 221 523 255 0 FreeSans 200 0 0 0 S[1]
port 31 nsew
flabel corelocali s 765 85 799 119 0 FreeSans 200 0 0 0 D[1]
port 15 nsew
flabel corelocali s 949 85 983 119 0 FreeSans 200 0 0 0 D[2]
port 14 nsew
flabel corelocali s 1225 221 1259 255 0 FreeSans 200 0 0 0 S[2]
port 30 nsew
flabel corelocali s 1317 221 1351 255 0 FreeSans 200 0 0 0 S[3]
port 29 nsew
flabel corelocali s 1777 85 1811 119 0 FreeSans 200 0 0 0 D[4]
port 12 nsew
flabel corelocali s 2053 221 2087 255 0 FreeSans 200 0 0 0 S[4]
port 28 nsew
flabel corelocali s 2145 221 2179 255 0 FreeSans 200 0 0 0 S[5]
port 27 nsew
flabel corelocali s 2421 85 2455 119 0 FreeSans 200 0 0 0 D[5]
port 11 nsew
flabel corelocali s 2605 85 2639 119 0 FreeSans 200 0 0 0 D[6]
port 10 nsew
flabel corelocali s 2881 221 2915 255 0 FreeSans 200 0 0 0 S[6]
port 26 nsew
flabel corelocali s 2973 221 3007 255 0 FreeSans 200 0 0 0 S[7]
port 25 nsew
flabel corelocali s 3249 85 3283 119 0 FreeSans 200 0 0 0 D[7]
port 9 nsew
flabel corelocali s 1593 85 1627 119 0 FreeSans 200 0 0 0 D[3]
port 13 nsew
<< properties >>
string FIXED_BBOX 0 0 3404 1088
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3026090
string GDS_START 2964356
<< end >>
