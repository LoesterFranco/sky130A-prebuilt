magic
tech sky130A
magscale 1 2
timestamp 1599588209
<< nwell >>
rect -38 332 902 704
<< pwell >>
rect 0 0 864 49
<< scpmos >>
rect 87 368 117 592
rect 339 368 369 592
rect 439 368 469 592
rect 738 368 768 592
<< nmoslvt >>
rect 84 74 114 222
rect 170 74 200 222
rect 256 74 286 222
rect 342 74 372 222
rect 436 74 466 222
rect 528 74 558 222
rect 628 74 658 222
rect 741 74 771 222
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 142 170 222
rect 114 108 125 142
rect 159 108 170 142
rect 114 74 170 108
rect 200 210 256 222
rect 200 176 211 210
rect 245 176 256 210
rect 200 120 256 176
rect 200 86 211 120
rect 245 86 256 120
rect 200 74 256 86
rect 286 142 342 222
rect 286 108 297 142
rect 331 108 342 142
rect 286 74 342 108
rect 372 210 436 222
rect 372 176 383 210
rect 417 176 436 210
rect 372 120 436 176
rect 372 86 383 120
rect 417 86 436 120
rect 372 74 436 86
rect 466 174 528 222
rect 466 140 483 174
rect 517 140 528 174
rect 466 74 528 140
rect 558 142 628 222
rect 558 108 583 142
rect 617 108 628 142
rect 558 74 628 108
rect 658 174 741 222
rect 658 140 687 174
rect 721 140 741 174
rect 658 74 741 140
rect 771 142 837 222
rect 771 108 791 142
rect 825 108 837 142
rect 771 74 837 108
<< pdiff >>
rect 27 580 87 592
rect 27 546 39 580
rect 73 546 87 580
rect 27 500 87 546
rect 27 466 39 500
rect 73 466 87 500
rect 27 420 87 466
rect 27 386 39 420
rect 73 386 87 420
rect 27 368 87 386
rect 117 580 339 592
rect 117 546 130 580
rect 164 546 210 580
rect 244 546 292 580
rect 326 546 339 580
rect 117 511 339 546
rect 117 477 130 511
rect 164 477 210 511
rect 244 477 292 511
rect 326 477 339 511
rect 117 440 339 477
rect 117 406 130 440
rect 164 406 210 440
rect 244 406 292 440
rect 326 406 339 440
rect 117 368 339 406
rect 369 580 439 592
rect 369 546 382 580
rect 416 546 439 580
rect 369 501 439 546
rect 369 467 382 501
rect 416 467 439 501
rect 369 368 439 467
rect 469 580 738 592
rect 469 546 482 580
rect 516 546 551 580
rect 585 546 622 580
rect 656 546 691 580
rect 725 546 738 580
rect 469 511 738 546
rect 469 477 482 511
rect 516 477 551 511
rect 585 477 622 511
rect 656 477 691 511
rect 725 477 738 511
rect 469 440 738 477
rect 469 406 482 440
rect 516 406 551 440
rect 585 406 622 440
rect 656 406 691 440
rect 725 406 738 440
rect 469 368 738 406
rect 768 580 837 592
rect 768 546 791 580
rect 825 546 837 580
rect 768 501 837 546
rect 768 467 791 501
rect 825 467 837 501
rect 768 368 837 467
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 125 108 159 142
rect 211 176 245 210
rect 211 86 245 120
rect 297 108 331 142
rect 383 176 417 210
rect 383 86 417 120
rect 483 140 517 174
rect 583 108 617 142
rect 687 140 721 174
rect 791 108 825 142
<< pdiffc >>
rect 39 546 73 580
rect 39 466 73 500
rect 39 386 73 420
rect 130 546 164 580
rect 210 546 244 580
rect 292 546 326 580
rect 130 477 164 511
rect 210 477 244 511
rect 292 477 326 511
rect 130 406 164 440
rect 210 406 244 440
rect 292 406 326 440
rect 382 546 416 580
rect 382 467 416 501
rect 482 546 516 580
rect 551 546 585 580
rect 622 546 656 580
rect 691 546 725 580
rect 482 477 516 511
rect 551 477 585 511
rect 622 477 656 511
rect 691 477 725 511
rect 482 406 516 440
rect 551 406 585 440
rect 622 406 656 440
rect 691 406 725 440
rect 791 546 825 580
rect 791 467 825 501
<< poly >>
rect 87 592 117 618
rect 339 592 369 618
rect 439 592 469 618
rect 738 592 768 618
rect 87 353 117 368
rect 339 353 369 368
rect 439 353 469 368
rect 738 353 768 368
rect 84 336 120 353
rect 336 336 372 353
rect 84 320 372 336
rect 84 286 118 320
rect 152 286 186 320
rect 220 286 254 320
rect 288 286 322 320
rect 356 286 372 320
rect 84 270 372 286
rect 84 222 114 270
rect 170 222 200 270
rect 256 222 286 270
rect 342 222 372 270
rect 436 336 472 353
rect 735 336 771 353
rect 436 320 771 336
rect 436 286 505 320
rect 539 286 573 320
rect 607 286 641 320
rect 675 286 709 320
rect 743 286 771 320
rect 436 270 771 286
rect 436 222 466 270
rect 528 222 558 270
rect 628 222 658 270
rect 741 222 771 270
rect 84 48 114 74
rect 170 48 200 74
rect 256 48 286 74
rect 342 48 372 74
rect 436 48 466 74
rect 528 48 558 74
rect 628 48 658 74
rect 741 48 771 74
<< polycont >>
rect 118 286 152 320
rect 186 286 220 320
rect 254 286 288 320
rect 322 286 356 320
rect 505 286 539 320
rect 573 286 607 320
rect 641 286 675 320
rect 709 286 743 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 23 580 89 649
rect 23 546 39 580
rect 73 546 89 580
rect 23 500 89 546
rect 23 466 39 500
rect 73 466 89 500
rect 23 420 89 466
rect 23 386 39 420
rect 73 386 89 420
rect 123 580 332 596
rect 123 546 130 580
rect 164 546 210 580
rect 244 546 292 580
rect 326 546 332 580
rect 123 511 332 546
rect 123 477 130 511
rect 164 477 210 511
rect 244 477 292 511
rect 326 477 332 511
rect 123 440 332 477
rect 366 580 432 649
rect 366 546 382 580
rect 416 546 432 580
rect 366 501 432 546
rect 366 467 382 501
rect 416 467 432 501
rect 366 458 432 467
rect 466 580 741 596
rect 466 546 482 580
rect 516 546 551 580
rect 585 546 622 580
rect 656 546 691 580
rect 725 546 741 580
rect 466 511 741 546
rect 466 477 482 511
rect 516 477 551 511
rect 585 477 622 511
rect 656 477 691 511
rect 725 477 741 511
rect 123 406 130 440
rect 164 406 210 440
rect 244 406 292 440
rect 326 424 332 440
rect 466 440 741 477
rect 775 580 841 649
rect 775 546 791 580
rect 825 546 841 580
rect 775 501 841 546
rect 775 467 791 501
rect 825 467 841 501
rect 775 458 841 467
rect 466 424 482 440
rect 326 406 482 424
rect 516 406 551 440
rect 585 406 622 440
rect 656 406 691 440
rect 725 424 741 440
rect 725 406 839 424
rect 123 390 839 406
rect 23 370 89 386
rect 217 336 455 356
rect 102 320 455 336
rect 102 286 118 320
rect 152 286 186 320
rect 220 286 254 320
rect 288 286 322 320
rect 356 286 455 320
rect 102 270 455 286
rect 489 320 759 356
rect 489 286 505 320
rect 539 286 573 320
rect 607 286 641 320
rect 675 286 709 320
rect 743 286 759 320
rect 489 270 759 286
rect 793 236 839 390
rect 23 210 433 236
rect 23 176 39 210
rect 73 202 211 210
rect 23 120 73 176
rect 245 202 383 210
rect 23 86 39 120
rect 23 70 73 86
rect 109 142 175 161
rect 109 108 125 142
rect 159 108 175 142
rect 109 17 175 108
rect 211 120 245 176
rect 417 176 433 210
rect 211 70 245 86
rect 281 142 347 161
rect 281 108 297 142
rect 331 108 347 142
rect 281 17 347 108
rect 383 120 433 176
rect 467 202 839 236
rect 467 174 533 202
rect 467 140 483 174
rect 517 140 533 174
rect 667 174 741 202
rect 467 122 533 140
rect 567 142 633 161
rect 417 86 433 120
rect 383 85 433 86
rect 567 108 583 142
rect 617 108 633 142
rect 667 140 687 174
rect 721 140 741 174
rect 667 122 741 140
rect 775 142 841 161
rect 567 85 633 108
rect 775 108 791 142
rect 825 108 841 142
rect 775 85 841 108
rect 383 51 841 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel comment s 0 0 0 0 4 nand2_4
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 799 242 833 276 0 FreeSans 340 0 0 0 Y
port 7 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 Y
port 7 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 A
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 864 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1926168
string GDS_START 1918250
<< end >>
