magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 127 424 177 547
rect 323 424 357 547
rect 503 424 537 547
rect 683 424 723 547
rect 127 390 723 424
rect 121 270 391 356
rect 453 270 655 356
rect 689 304 723 390
rect 689 236 839 304
rect 889 270 1127 356
rect 1177 270 1493 356
rect 470 226 839 236
rect 470 202 1156 226
rect 470 119 536 202
rect 642 170 1156 202
rect 642 154 798 170
rect 1090 154 1156 170
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 37 581 807 615
rect 37 364 87 581
rect 217 458 283 581
rect 397 458 463 581
rect 577 458 643 581
rect 757 424 807 581
rect 847 458 913 649
rect 953 424 1003 596
rect 1037 458 1129 649
rect 1163 424 1213 596
rect 1253 458 1319 649
rect 1359 424 1393 596
rect 1433 458 1499 649
rect 1539 424 1589 596
rect 757 390 1589 424
rect 757 364 807 390
rect 1539 364 1589 390
rect 40 202 434 236
rect 40 70 90 202
rect 126 17 176 168
rect 212 70 262 202
rect 298 17 364 168
rect 400 85 434 202
rect 572 120 606 168
rect 1192 202 1586 236
rect 832 120 898 136
rect 1192 120 1226 202
rect 572 85 794 120
rect 400 51 794 85
rect 832 70 1226 120
rect 1262 17 1312 168
rect 1348 70 1398 202
rect 1434 17 1484 168
rect 1520 70 1586 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
rlabel locali s 889 270 1127 356 6 A1
port 1 nsew signal input
rlabel locali s 1177 270 1493 356 6 A2
port 2 nsew signal input
rlabel locali s 453 270 655 356 6 B1
port 3 nsew signal input
rlabel locali s 121 270 391 356 6 B2
port 4 nsew signal input
rlabel locali s 1090 154 1156 170 6 Y
port 5 nsew signal output
rlabel locali s 689 304 723 390 6 Y
port 5 nsew signal output
rlabel locali s 689 236 839 304 6 Y
port 5 nsew signal output
rlabel locali s 683 424 723 547 6 Y
port 5 nsew signal output
rlabel locali s 642 170 1156 202 6 Y
port 5 nsew signal output
rlabel locali s 642 154 798 170 6 Y
port 5 nsew signal output
rlabel locali s 503 424 537 547 6 Y
port 5 nsew signal output
rlabel locali s 470 226 839 236 6 Y
port 5 nsew signal output
rlabel locali s 470 202 1156 226 6 Y
port 5 nsew signal output
rlabel locali s 470 119 536 202 6 Y
port 5 nsew signal output
rlabel locali s 323 424 357 547 6 Y
port 5 nsew signal output
rlabel locali s 127 424 177 547 6 Y
port 5 nsew signal output
rlabel locali s 127 390 723 424 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -49 1632 49 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1632 715 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3514782
string GDS_START 3501242
<< end >>
