magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1104 561
rect 83 374 149 527
rect 183 340 221 493
rect 255 374 321 527
rect 355 340 391 493
rect 427 451 497 527
rect 603 455 737 527
rect 18 306 391 340
rect 1015 387 1087 527
rect 18 161 64 306
rect 497 215 631 323
rect 696 299 1080 341
rect 696 198 757 299
rect 828 199 938 265
rect 1006 199 1080 299
rect 18 127 343 161
rect 119 123 343 127
rect 19 17 85 93
rect 191 17 257 89
rect 363 17 429 93
rect 755 17 823 89
rect 929 17 995 89
rect 0 -17 1104 17
<< obsli1 >>
rect 531 421 569 493
rect 843 421 909 489
rect 531 417 909 421
rect 425 375 909 417
rect 425 366 569 375
rect 425 267 463 366
rect 98 199 463 267
rect 423 174 463 199
rect 423 131 619 174
rect 655 123 1081 157
rect 655 97 721 123
rect 467 51 721 97
<< metal1 >>
rect 0 496 1104 592
rect 0 -48 1104 48
<< labels >>
rlabel locali s 1006 199 1080 299 6 A1
port 1 nsew signal input
rlabel locali s 696 299 1080 341 6 A1
port 1 nsew signal input
rlabel locali s 696 198 757 299 6 A1
port 1 nsew signal input
rlabel locali s 828 199 938 265 6 A2
port 2 nsew signal input
rlabel locali s 497 215 631 323 6 B1
port 3 nsew signal input
rlabel locali s 355 340 391 493 6 X
port 4 nsew signal output
rlabel locali s 183 340 221 493 6 X
port 4 nsew signal output
rlabel locali s 119 123 343 127 6 X
port 4 nsew signal output
rlabel locali s 18 306 391 340 6 X
port 4 nsew signal output
rlabel locali s 18 161 64 306 6 X
port 4 nsew signal output
rlabel locali s 18 127 343 161 6 X
port 4 nsew signal output
rlabel locali s 929 17 995 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 755 17 823 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 363 17 429 93 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 191 17 257 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 19 17 85 93 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 1104 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1104 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 1015 387 1087 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 603 455 737 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 427 451 497 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 255 374 321 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 83 374 149 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 1104 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 1104 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1104 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1347106
string GDS_START 1339182
<< end >>
