magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 1510 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 89 47 119 131
rect 196 47 226 177
rect 390 47 420 177
rect 484 47 514 177
rect 588 47 618 177
rect 672 47 702 177
rect 766 47 796 177
rect 860 47 890 177
rect 954 47 984 177
rect 1048 47 1078 177
rect 1142 47 1172 177
rect 1236 47 1266 177
rect 1340 47 1370 177
<< pmoshvt >>
rect 81 297 117 425
rect 188 297 224 497
rect 392 297 428 497
rect 486 297 522 497
rect 580 297 616 497
rect 674 297 710 497
rect 768 297 804 497
rect 862 297 898 497
rect 956 297 992 497
rect 1050 297 1086 497
rect 1144 297 1180 497
rect 1238 297 1274 497
rect 1332 297 1368 497
<< ndiff >>
rect 134 131 196 177
rect 27 111 89 131
rect 27 77 35 111
rect 69 77 89 111
rect 27 47 89 77
rect 119 97 196 131
rect 119 63 129 97
rect 163 63 196 97
rect 119 47 196 63
rect 226 165 278 177
rect 226 131 236 165
rect 270 131 278 165
rect 226 97 278 131
rect 226 63 236 97
rect 270 63 278 97
rect 226 47 278 63
rect 338 165 390 177
rect 338 131 346 165
rect 380 131 390 165
rect 338 97 390 131
rect 338 63 346 97
rect 380 63 390 97
rect 338 47 390 63
rect 420 97 484 177
rect 420 63 440 97
rect 474 63 484 97
rect 420 47 484 63
rect 514 165 588 177
rect 514 131 534 165
rect 568 131 588 165
rect 514 97 588 131
rect 514 63 534 97
rect 568 63 588 97
rect 514 47 588 63
rect 618 97 672 177
rect 618 63 628 97
rect 662 63 672 97
rect 618 47 672 63
rect 702 165 766 177
rect 702 131 722 165
rect 756 131 766 165
rect 702 97 766 131
rect 702 63 722 97
rect 756 63 766 97
rect 702 47 766 63
rect 796 97 860 177
rect 796 63 816 97
rect 850 63 860 97
rect 796 47 860 63
rect 890 165 954 177
rect 890 131 910 165
rect 944 131 954 165
rect 890 97 954 131
rect 890 63 910 97
rect 944 63 954 97
rect 890 47 954 63
rect 984 97 1048 177
rect 984 63 1004 97
rect 1038 63 1048 97
rect 984 47 1048 63
rect 1078 165 1142 177
rect 1078 131 1098 165
rect 1132 131 1142 165
rect 1078 97 1142 131
rect 1078 63 1098 97
rect 1132 63 1142 97
rect 1078 47 1142 63
rect 1172 97 1236 177
rect 1172 63 1192 97
rect 1226 63 1236 97
rect 1172 47 1236 63
rect 1266 165 1340 177
rect 1266 131 1286 165
rect 1320 131 1340 165
rect 1266 97 1340 131
rect 1266 63 1286 97
rect 1320 63 1340 97
rect 1266 47 1340 63
rect 1370 97 1422 177
rect 1370 63 1380 97
rect 1414 63 1422 97
rect 1370 47 1422 63
<< pdiff >>
rect 134 425 188 497
rect 27 411 81 425
rect 27 377 35 411
rect 69 377 81 411
rect 27 343 81 377
rect 27 309 35 343
rect 69 309 81 343
rect 27 297 81 309
rect 117 407 188 425
rect 117 373 129 407
rect 163 373 188 407
rect 117 297 188 373
rect 224 479 278 497
rect 224 445 236 479
rect 270 445 278 479
rect 224 411 278 445
rect 224 377 236 411
rect 270 377 278 411
rect 224 343 278 377
rect 224 309 236 343
rect 270 309 278 343
rect 224 297 278 309
rect 338 479 392 497
rect 338 445 346 479
rect 380 445 392 479
rect 338 411 392 445
rect 338 377 346 411
rect 380 377 392 411
rect 338 343 392 377
rect 338 309 346 343
rect 380 309 392 343
rect 338 297 392 309
rect 428 485 486 497
rect 428 451 440 485
rect 474 451 486 485
rect 428 417 486 451
rect 428 383 440 417
rect 474 383 486 417
rect 428 297 486 383
rect 522 479 580 497
rect 522 445 534 479
rect 568 445 580 479
rect 522 411 580 445
rect 522 377 534 411
rect 568 377 580 411
rect 522 343 580 377
rect 522 309 534 343
rect 568 309 580 343
rect 522 297 580 309
rect 616 485 674 497
rect 616 451 628 485
rect 662 451 674 485
rect 616 417 674 451
rect 616 383 628 417
rect 662 383 674 417
rect 616 297 674 383
rect 710 479 768 497
rect 710 445 722 479
rect 756 445 768 479
rect 710 411 768 445
rect 710 377 722 411
rect 756 377 768 411
rect 710 343 768 377
rect 710 309 722 343
rect 756 309 768 343
rect 710 297 768 309
rect 804 485 862 497
rect 804 451 816 485
rect 850 451 862 485
rect 804 417 862 451
rect 804 383 816 417
rect 850 383 862 417
rect 804 297 862 383
rect 898 479 956 497
rect 898 445 910 479
rect 944 445 956 479
rect 898 411 956 445
rect 898 377 910 411
rect 944 377 956 411
rect 898 343 956 377
rect 898 309 910 343
rect 944 309 956 343
rect 898 297 956 309
rect 992 485 1050 497
rect 992 451 1004 485
rect 1038 451 1050 485
rect 992 417 1050 451
rect 992 383 1004 417
rect 1038 383 1050 417
rect 992 297 1050 383
rect 1086 479 1144 497
rect 1086 445 1098 479
rect 1132 445 1144 479
rect 1086 411 1144 445
rect 1086 377 1098 411
rect 1132 377 1144 411
rect 1086 343 1144 377
rect 1086 309 1098 343
rect 1132 309 1144 343
rect 1086 297 1144 309
rect 1180 485 1238 497
rect 1180 451 1192 485
rect 1226 451 1238 485
rect 1180 417 1238 451
rect 1180 383 1192 417
rect 1226 383 1238 417
rect 1180 297 1238 383
rect 1274 479 1332 497
rect 1274 445 1286 479
rect 1320 445 1332 479
rect 1274 411 1332 445
rect 1274 377 1286 411
rect 1320 377 1332 411
rect 1274 343 1332 377
rect 1274 309 1286 343
rect 1320 309 1332 343
rect 1274 297 1332 309
rect 1368 485 1422 497
rect 1368 451 1380 485
rect 1414 451 1422 485
rect 1368 417 1422 451
rect 1368 383 1380 417
rect 1414 383 1422 417
rect 1368 297 1422 383
<< ndiffc >>
rect 35 77 69 111
rect 129 63 163 97
rect 236 131 270 165
rect 236 63 270 97
rect 346 131 380 165
rect 346 63 380 97
rect 440 63 474 97
rect 534 131 568 165
rect 534 63 568 97
rect 628 63 662 97
rect 722 131 756 165
rect 722 63 756 97
rect 816 63 850 97
rect 910 131 944 165
rect 910 63 944 97
rect 1004 63 1038 97
rect 1098 131 1132 165
rect 1098 63 1132 97
rect 1192 63 1226 97
rect 1286 131 1320 165
rect 1286 63 1320 97
rect 1380 63 1414 97
<< pdiffc >>
rect 35 377 69 411
rect 35 309 69 343
rect 129 373 163 407
rect 236 445 270 479
rect 236 377 270 411
rect 236 309 270 343
rect 346 445 380 479
rect 346 377 380 411
rect 346 309 380 343
rect 440 451 474 485
rect 440 383 474 417
rect 534 445 568 479
rect 534 377 568 411
rect 534 309 568 343
rect 628 451 662 485
rect 628 383 662 417
rect 722 445 756 479
rect 722 377 756 411
rect 722 309 756 343
rect 816 451 850 485
rect 816 383 850 417
rect 910 445 944 479
rect 910 377 944 411
rect 910 309 944 343
rect 1004 451 1038 485
rect 1004 383 1038 417
rect 1098 445 1132 479
rect 1098 377 1132 411
rect 1098 309 1132 343
rect 1192 451 1226 485
rect 1192 383 1226 417
rect 1286 445 1320 479
rect 1286 377 1320 411
rect 1286 309 1320 343
rect 1380 451 1414 485
rect 1380 383 1414 417
<< poly >>
rect 188 497 224 523
rect 392 497 428 523
rect 486 497 522 523
rect 580 497 616 523
rect 674 497 710 523
rect 768 497 804 523
rect 862 497 898 523
rect 956 497 992 523
rect 1050 497 1086 523
rect 1144 497 1180 523
rect 1238 497 1274 523
rect 1332 497 1368 523
rect 81 425 117 451
rect 81 282 117 297
rect 188 282 224 297
rect 392 282 428 297
rect 486 282 522 297
rect 580 282 616 297
rect 674 282 710 297
rect 768 282 804 297
rect 862 282 898 297
rect 956 282 992 297
rect 1050 282 1086 297
rect 1144 282 1180 297
rect 1238 282 1274 297
rect 1332 282 1368 297
rect 79 265 119 282
rect 186 265 226 282
rect 22 249 119 265
rect 22 215 38 249
rect 72 215 119 249
rect 22 199 119 215
rect 171 249 238 265
rect 171 215 184 249
rect 218 215 238 249
rect 171 199 238 215
rect 390 259 430 282
rect 484 259 524 282
rect 578 259 618 282
rect 390 249 618 259
rect 390 215 440 249
rect 474 215 508 249
rect 542 215 618 249
rect 390 205 618 215
rect 89 131 119 199
rect 196 177 226 199
rect 390 177 420 205
rect 484 177 514 205
rect 588 177 618 205
rect 672 259 712 282
rect 766 259 806 282
rect 860 259 900 282
rect 954 259 994 282
rect 1048 259 1088 282
rect 1142 259 1182 282
rect 1236 259 1276 282
rect 1330 259 1370 282
rect 672 249 1370 259
rect 672 215 696 249
rect 730 215 774 249
rect 808 215 852 249
rect 886 215 930 249
rect 964 215 1008 249
rect 1042 215 1076 249
rect 1110 215 1370 249
rect 672 205 1370 215
rect 672 177 702 205
rect 766 177 796 205
rect 860 177 890 205
rect 954 177 984 205
rect 1048 177 1078 205
rect 1142 177 1172 205
rect 1236 177 1266 205
rect 1340 177 1370 205
rect 89 21 119 47
rect 196 21 226 47
rect 390 21 420 47
rect 484 21 514 47
rect 588 21 618 47
rect 672 21 702 47
rect 766 21 796 47
rect 860 21 890 47
rect 954 21 984 47
rect 1048 21 1078 47
rect 1142 21 1172 47
rect 1236 21 1266 47
rect 1340 21 1370 47
<< polycont >>
rect 38 215 72 249
rect 184 215 218 249
rect 440 215 474 249
rect 508 215 542 249
rect 696 215 730 249
rect 774 215 808 249
rect 852 215 886 249
rect 930 215 964 249
rect 1008 215 1042 249
rect 1076 215 1110 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 19 411 85 432
rect 19 377 35 411
rect 69 377 85 411
rect 19 343 85 377
rect 129 407 163 527
rect 129 357 163 373
rect 210 479 296 493
rect 210 445 236 479
rect 270 445 296 479
rect 210 411 296 445
rect 210 377 236 411
rect 270 377 296 411
rect 19 309 35 343
rect 69 323 85 343
rect 210 343 296 377
rect 69 309 166 323
rect 210 309 236 343
rect 270 309 296 343
rect 19 289 166 309
rect 132 265 166 289
rect 22 249 88 255
rect 22 215 38 249
rect 72 215 88 249
rect 132 249 228 265
rect 132 215 184 249
rect 218 215 228 249
rect 132 199 228 215
rect 262 255 296 309
rect 330 479 396 493
rect 330 445 346 479
rect 380 445 396 479
rect 330 411 396 445
rect 330 377 346 411
rect 380 377 396 411
rect 330 343 396 377
rect 440 485 474 527
rect 440 417 474 451
rect 440 357 474 383
rect 508 479 584 493
rect 508 445 534 479
rect 568 445 584 479
rect 508 411 584 445
rect 508 377 534 411
rect 568 377 584 411
rect 330 309 346 343
rect 380 323 396 343
rect 508 343 584 377
rect 628 485 662 527
rect 628 417 662 451
rect 628 357 662 383
rect 696 479 772 493
rect 696 445 722 479
rect 756 445 772 479
rect 696 411 772 445
rect 696 377 722 411
rect 756 377 772 411
rect 508 323 534 343
rect 380 309 534 323
rect 568 323 584 343
rect 696 343 772 377
rect 816 485 850 527
rect 816 417 850 451
rect 816 367 850 383
rect 884 479 960 493
rect 884 445 910 479
rect 944 445 960 479
rect 884 411 960 445
rect 884 377 910 411
rect 944 377 960 411
rect 568 309 662 323
rect 330 289 662 309
rect 696 309 722 343
rect 756 323 772 343
rect 884 343 960 377
rect 1004 485 1038 527
rect 1004 417 1038 451
rect 1004 367 1038 383
rect 1072 479 1148 493
rect 1072 445 1098 479
rect 1132 445 1148 479
rect 1072 411 1148 445
rect 1072 377 1098 411
rect 1132 377 1148 411
rect 884 323 910 343
rect 756 309 910 323
rect 944 323 960 343
rect 1072 343 1148 377
rect 1192 485 1226 527
rect 1192 417 1226 451
rect 1192 367 1226 383
rect 1260 479 1336 493
rect 1260 445 1286 479
rect 1320 445 1336 479
rect 1260 411 1336 445
rect 1260 377 1286 411
rect 1320 377 1336 411
rect 1072 323 1098 343
rect 944 309 1098 323
rect 1132 323 1148 343
rect 1260 343 1336 377
rect 1380 485 1414 527
rect 1380 417 1414 451
rect 1380 367 1414 383
rect 1260 323 1286 343
rect 1132 309 1286 323
rect 1320 323 1336 343
rect 1320 309 1448 323
rect 696 289 1448 309
rect 628 255 662 289
rect 262 249 584 255
rect 262 215 440 249
rect 474 215 508 249
rect 542 215 584 249
rect 628 249 1182 255
rect 628 215 696 249
rect 730 215 774 249
rect 808 215 852 249
rect 886 215 930 249
rect 964 215 1008 249
rect 1042 215 1076 249
rect 1110 215 1182 249
rect 132 181 166 199
rect 19 147 166 181
rect 262 165 296 215
rect 628 181 662 215
rect 1372 181 1448 289
rect 19 111 85 147
rect 210 131 236 165
rect 270 131 296 165
rect 19 77 35 111
rect 69 77 85 111
rect 19 52 85 77
rect 129 97 163 113
rect 129 17 163 63
rect 210 97 296 131
rect 210 63 236 97
rect 270 63 296 97
rect 210 52 296 63
rect 330 165 662 181
rect 330 131 346 165
rect 380 147 534 165
rect 380 131 396 147
rect 330 97 396 131
rect 508 131 534 147
rect 568 147 662 165
rect 696 165 1448 181
rect 568 131 584 147
rect 330 63 346 97
rect 380 63 396 97
rect 330 52 396 63
rect 440 97 474 113
rect 440 17 474 63
rect 508 97 584 131
rect 696 131 722 165
rect 756 147 910 165
rect 756 131 772 147
rect 508 63 534 97
rect 568 63 584 97
rect 508 52 584 63
rect 628 97 662 113
rect 628 17 662 63
rect 696 97 772 131
rect 884 131 910 147
rect 944 147 1098 165
rect 944 131 960 147
rect 696 63 722 97
rect 756 63 772 97
rect 696 52 772 63
rect 816 97 850 113
rect 816 17 850 63
rect 884 97 960 131
rect 1072 131 1098 147
rect 1132 147 1286 165
rect 1132 131 1148 147
rect 884 63 910 97
rect 944 63 960 97
rect 884 52 960 63
rect 1004 97 1038 113
rect 1004 17 1038 63
rect 1072 97 1148 131
rect 1260 131 1286 147
rect 1320 147 1448 165
rect 1320 131 1336 147
rect 1072 63 1098 97
rect 1132 63 1148 97
rect 1072 52 1148 63
rect 1192 97 1226 113
rect 1192 17 1226 63
rect 1260 97 1336 131
rect 1260 63 1286 97
rect 1320 63 1336 97
rect 1260 52 1336 63
rect 1380 97 1414 113
rect 1380 17 1414 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< labels >>
flabel corelocali s 30 221 64 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 1390 238 1390 238 0 FreeSans 200 0 0 0 X
port 6 nsew
flabel corelocali s 1390 306 1390 306 0 FreeSans 200 0 0 0 X
port 6 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 1472 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1714314
string GDS_START 1703340
<< end >>
