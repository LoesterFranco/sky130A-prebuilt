magic
tech sky130A
magscale 1 2
timestamp 1604502711
<< locali >>
rect 18 195 88 325
rect 354 201 436 325
rect 722 187 804 213
rect 722 153 770 187
rect 722 147 804 153
rect 1336 201 1402 213
rect 1336 187 1468 201
rect 1336 153 1422 187
rect 1456 153 1468 187
rect 1336 147 1468 153
rect 1789 331 1840 465
rect 1804 159 1840 331
rect 1789 53 1840 159
<< viali >>
rect 770 153 804 187
rect 1422 153 1456 187
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 35 393 69 493
rect 103 427 169 527
rect 35 359 168 393
rect 122 161 168 359
rect 35 127 168 161
rect 35 69 69 127
rect 103 17 169 93
rect 203 69 248 493
rect 291 427 357 527
rect 391 393 425 493
rect 472 450 638 484
rect 686 451 762 527
rect 286 359 425 393
rect 286 165 320 359
rect 470 315 570 391
rect 286 127 425 165
rect 470 141 514 315
rect 604 281 638 450
rect 798 417 832 475
rect 866 451 932 527
rect 1026 433 1152 483
rect 1188 451 1272 527
rect 1118 417 1152 433
rect 1312 417 1360 475
rect 672 367 946 417
rect 672 315 722 367
rect 824 281 874 313
rect 604 247 874 281
rect 604 239 688 247
rect 550 129 620 203
rect 291 17 357 93
rect 391 61 425 127
rect 654 93 688 239
rect 908 213 946 367
rect 862 145 946 213
rect 980 331 1084 393
rect 1118 383 1360 417
rect 1406 389 1472 527
rect 980 179 1014 331
rect 1048 213 1084 295
rect 1118 281 1152 383
rect 1506 353 1540 475
rect 1594 383 1660 485
rect 1506 349 1570 353
rect 1186 315 1570 349
rect 1118 247 1498 281
rect 1164 179 1230 203
rect 980 145 1230 179
rect 485 53 688 93
rect 722 17 804 105
rect 862 59 912 145
rect 952 17 1016 109
rect 1264 95 1298 247
rect 1432 235 1498 247
rect 1532 136 1570 315
rect 1128 61 1298 95
rect 1338 17 1470 113
rect 1506 70 1570 136
rect 1610 265 1660 383
rect 1696 367 1753 527
rect 1610 199 1770 265
rect 1610 69 1660 199
rect 1696 17 1753 109
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
rect 758 187 816 193
rect 758 153 770 187
rect 804 184 816 187
rect 1410 187 1468 193
rect 1410 184 1422 187
rect 804 156 1422 184
rect 804 153 816 156
rect 758 147 816 153
rect 1410 153 1422 156
rect 1456 153 1468 187
rect 1410 147 1468 153
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< obsm1 >>
rect 110 388 168 397
rect 482 388 540 397
rect 1038 388 1096 397
rect 110 360 1096 388
rect 110 351 168 360
rect 482 351 540 360
rect 1038 351 1096 360
rect 1038 252 1096 261
rect 589 224 1096 252
rect 589 193 632 224
rect 1038 215 1096 224
rect 202 184 260 193
rect 574 184 632 193
rect 202 156 632 184
rect 202 147 260 156
rect 574 147 632 156
<< labels >>
rlabel locali s 354 201 436 325 6 D
port 1 nsew signal input
rlabel locali s 1804 159 1840 331 6 Q
port 2 nsew signal output
rlabel locali s 1789 331 1840 465 6 Q
port 2 nsew signal output
rlabel locali s 1789 53 1840 159 6 Q
port 2 nsew signal output
rlabel viali s 770 153 804 187 6 SET_B
port 3 nsew signal input
rlabel locali s 722 147 804 213 6 SET_B
port 3 nsew signal input
rlabel viali s 1422 153 1456 187 6 SET_B
port 3 nsew signal input
rlabel locali s 1336 201 1402 213 6 SET_B
port 3 nsew signal input
rlabel locali s 1336 147 1468 201 6 SET_B
port 3 nsew signal input
rlabel metal1 s 1410 184 1468 193 6 SET_B
port 3 nsew signal input
rlabel metal1 s 1410 147 1468 156 6 SET_B
port 3 nsew signal input
rlabel metal1 s 758 184 816 193 6 SET_B
port 3 nsew signal input
rlabel metal1 s 758 156 1468 184 6 SET_B
port 3 nsew signal input
rlabel metal1 s 758 147 816 156 6 SET_B
port 3 nsew signal input
rlabel locali s 18 195 88 325 6 CLK
port 4 nsew clock input
rlabel metal1 s 0 -48 1932 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1932 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1932 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2460222
string GDS_START 2444680
<< end >>
