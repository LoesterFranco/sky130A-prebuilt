magic
tech sky130A
magscale 1 2
timestamp 1601050056
<< nwell >>
rect -38 332 710 704
<< pwell >>
rect 0 0 672 49
<< scpmos >>
rect 83 424 119 592
rect 320 368 356 568
rect 404 368 440 568
rect 521 368 557 592
<< nmoslvt >>
rect 161 112 191 222
rect 318 112 348 222
rect 404 112 434 222
rect 550 74 580 222
<< ndiff >>
rect 27 186 161 222
rect 27 152 39 186
rect 73 152 116 186
rect 150 152 161 186
rect 27 112 161 152
rect 191 184 318 222
rect 191 150 202 184
rect 236 150 270 184
rect 304 150 318 184
rect 191 112 318 150
rect 348 184 404 222
rect 348 150 359 184
rect 393 150 404 184
rect 348 112 404 150
rect 434 154 550 222
rect 434 120 476 154
rect 510 120 550 154
rect 434 112 550 120
rect 479 74 550 112
rect 580 210 637 222
rect 580 176 591 210
rect 625 176 637 210
rect 580 120 637 176
rect 580 86 591 120
rect 625 86 637 120
rect 580 74 637 86
<< pdiff >>
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 470 83 546
rect 27 436 39 470
rect 73 436 83 470
rect 27 424 83 436
rect 119 580 185 592
rect 119 546 139 580
rect 173 546 185 580
rect 455 580 521 592
rect 455 568 467 580
rect 119 470 185 546
rect 119 436 139 470
rect 173 436 185 470
rect 119 424 185 436
rect 264 556 320 568
rect 264 522 276 556
rect 310 522 320 556
rect 264 485 320 522
rect 264 451 276 485
rect 310 451 320 485
rect 264 414 320 451
rect 264 380 276 414
rect 310 380 320 414
rect 264 368 320 380
rect 356 368 404 568
rect 440 546 467 568
rect 501 546 521 580
rect 440 510 521 546
rect 440 476 467 510
rect 501 476 521 510
rect 440 440 521 476
rect 440 406 467 440
rect 501 406 521 440
rect 440 368 521 406
rect 557 580 613 592
rect 557 546 567 580
rect 601 546 613 580
rect 557 497 613 546
rect 557 463 567 497
rect 601 463 613 497
rect 557 414 613 463
rect 557 380 567 414
rect 601 380 613 414
rect 557 368 613 380
<< ndiffc >>
rect 39 152 73 186
rect 116 152 150 186
rect 202 150 236 184
rect 270 150 304 184
rect 359 150 393 184
rect 476 120 510 154
rect 591 176 625 210
rect 591 86 625 120
<< pdiffc >>
rect 39 546 73 580
rect 39 436 73 470
rect 139 546 173 580
rect 139 436 173 470
rect 276 522 310 556
rect 276 451 310 485
rect 276 380 310 414
rect 467 546 501 580
rect 467 476 501 510
rect 467 406 501 440
rect 567 546 601 580
rect 567 463 601 497
rect 567 380 601 414
<< poly >>
rect 83 592 119 618
rect 320 568 356 594
rect 404 568 440 594
rect 521 592 557 618
rect 83 322 119 424
rect 320 326 356 368
rect 83 310 113 322
rect 25 294 113 310
rect 25 260 41 294
rect 75 274 113 294
rect 239 310 356 326
rect 239 276 255 310
rect 289 296 356 310
rect 404 336 440 368
rect 404 320 473 336
rect 289 276 348 296
rect 75 260 191 274
rect 239 260 348 276
rect 25 244 191 260
rect 161 222 191 244
rect 318 222 348 260
rect 404 286 423 320
rect 457 286 473 320
rect 404 270 473 286
rect 521 326 557 368
rect 521 310 587 326
rect 521 276 537 310
rect 571 276 587 310
rect 404 222 434 270
rect 521 260 587 276
rect 550 222 580 260
rect 161 86 191 112
rect 318 86 348 112
rect 404 86 434 112
rect 550 48 580 74
<< polycont >>
rect 41 260 75 294
rect 255 276 289 310
rect 423 286 457 320
rect 537 276 571 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 23 580 89 596
rect 23 546 39 580
rect 73 546 89 580
rect 23 470 89 546
rect 23 436 39 470
rect 73 436 89 470
rect 23 386 89 436
rect 123 580 189 649
rect 123 546 139 580
rect 173 546 189 580
rect 451 580 517 649
rect 123 470 189 546
rect 123 436 139 470
rect 173 436 189 470
rect 123 420 189 436
rect 260 556 326 572
rect 260 522 276 556
rect 310 522 326 556
rect 260 485 326 522
rect 260 451 276 485
rect 310 451 326 485
rect 260 414 326 451
rect 23 352 166 386
rect 260 380 276 414
rect 310 398 326 414
rect 451 546 467 580
rect 501 546 517 580
rect 451 510 517 546
rect 451 476 467 510
rect 501 476 517 510
rect 451 440 517 476
rect 451 406 467 440
rect 501 406 517 440
rect 310 380 373 398
rect 451 390 517 406
rect 551 580 655 596
rect 551 546 567 580
rect 601 546 655 580
rect 551 497 655 546
rect 551 463 567 497
rect 601 463 655 497
rect 551 414 655 463
rect 260 364 373 380
rect 551 380 567 414
rect 601 380 655 414
rect 551 364 655 380
rect 132 326 166 352
rect 132 310 305 326
rect 25 294 91 310
rect 25 260 41 294
rect 75 260 91 294
rect 25 236 91 260
rect 132 276 255 310
rect 289 276 305 310
rect 132 260 305 276
rect 132 202 166 260
rect 339 236 373 364
rect 407 320 473 356
rect 407 286 423 320
rect 457 286 473 320
rect 407 270 473 286
rect 507 310 587 326
rect 507 276 537 310
rect 571 276 587 310
rect 507 260 587 276
rect 507 236 541 260
rect 23 186 166 202
rect 23 152 39 186
rect 73 152 116 186
rect 150 152 166 186
rect 23 136 166 152
rect 200 184 305 226
rect 200 150 202 184
rect 236 150 270 184
rect 304 150 305 184
rect 200 17 305 150
rect 339 202 541 236
rect 621 226 655 364
rect 575 210 655 226
rect 339 184 409 202
rect 339 150 359 184
rect 393 150 409 184
rect 575 176 591 210
rect 625 176 655 210
rect 339 108 409 150
rect 453 154 536 168
rect 453 120 476 154
rect 510 120 536 154
rect 453 17 536 120
rect 575 120 655 176
rect 575 86 591 120
rect 625 86 655 120
rect 575 70 655 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
rlabel comment s 0 0 0 0 4 or2b_1
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 607 390 641 424 0 FreeSans 340 0 0 0 X
port 7 nsew
flabel corelocali s 607 464 641 498 0 FreeSans 340 0 0 0 X
port 7 nsew
flabel corelocali s 607 538 641 572 0 FreeSans 340 0 0 0 X
port 7 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 B_N
port 2 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 672 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 761892
string GDS_START 756080
<< end >>
