magic
tech sky130A
magscale 1 2
timestamp 1601050056
<< nwell >>
rect -38 332 902 704
<< pwell >>
rect 0 0 864 49
<< scpmos >>
rect 83 368 119 592
rect 173 368 209 592
rect 273 368 309 592
rect 363 368 399 592
rect 453 368 489 592
rect 543 368 579 592
rect 643 368 679 592
rect 733 368 769 592
<< nmoslvt >>
rect 87 74 117 222
rect 173 74 203 222
rect 259 74 289 222
rect 345 74 375 222
rect 445 74 475 222
rect 531 74 561 222
rect 645 74 675 222
rect 731 74 761 222
<< ndiff >>
rect 30 210 87 222
rect 30 176 42 210
rect 76 176 87 210
rect 30 120 87 176
rect 30 86 42 120
rect 76 86 87 120
rect 30 74 87 86
rect 117 210 173 222
rect 117 176 128 210
rect 162 176 173 210
rect 117 120 173 176
rect 117 86 128 120
rect 162 86 173 120
rect 117 74 173 86
rect 203 152 259 222
rect 203 118 214 152
rect 248 118 259 152
rect 203 74 259 118
rect 289 210 345 222
rect 289 176 300 210
rect 334 176 345 210
rect 289 120 345 176
rect 289 86 300 120
rect 334 86 345 120
rect 289 74 345 86
rect 375 152 445 222
rect 375 118 386 152
rect 420 118 445 152
rect 375 74 445 118
rect 475 210 531 222
rect 475 176 486 210
rect 520 176 531 210
rect 475 120 531 176
rect 475 86 486 120
rect 520 86 531 120
rect 475 74 531 86
rect 561 192 645 222
rect 561 158 586 192
rect 620 158 645 192
rect 561 116 645 158
rect 561 82 586 116
rect 620 82 645 116
rect 561 74 645 82
rect 675 210 731 222
rect 675 176 686 210
rect 720 176 731 210
rect 675 120 731 176
rect 675 86 686 120
rect 720 86 731 120
rect 675 74 731 86
rect 761 194 819 222
rect 761 160 772 194
rect 806 160 819 194
rect 761 120 819 160
rect 761 86 772 120
rect 806 86 819 120
rect 761 74 819 86
<< pdiff >>
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 497 83 546
rect 27 463 39 497
rect 73 463 83 497
rect 27 414 83 463
rect 27 380 39 414
rect 73 380 83 414
rect 27 368 83 380
rect 119 580 173 592
rect 119 546 129 580
rect 163 546 173 580
rect 119 510 173 546
rect 119 476 129 510
rect 163 476 173 510
rect 119 440 173 476
rect 119 406 129 440
rect 163 406 173 440
rect 119 368 173 406
rect 209 580 273 592
rect 209 546 219 580
rect 253 546 273 580
rect 209 508 273 546
rect 209 474 219 508
rect 253 474 273 508
rect 209 368 273 474
rect 309 580 363 592
rect 309 546 319 580
rect 353 546 363 580
rect 309 510 363 546
rect 309 476 319 510
rect 353 476 363 510
rect 309 440 363 476
rect 309 406 319 440
rect 353 406 363 440
rect 309 368 363 406
rect 399 580 453 592
rect 399 546 409 580
rect 443 546 453 580
rect 399 508 453 546
rect 399 474 409 508
rect 443 474 453 508
rect 399 368 453 474
rect 489 580 543 592
rect 489 546 499 580
rect 533 546 543 580
rect 489 497 543 546
rect 489 463 499 497
rect 533 463 543 497
rect 489 414 543 463
rect 489 380 499 414
rect 533 380 543 414
rect 489 368 543 380
rect 579 580 643 592
rect 579 546 589 580
rect 623 546 643 580
rect 579 497 643 546
rect 579 463 589 497
rect 623 463 643 497
rect 579 414 643 463
rect 579 380 589 414
rect 623 380 643 414
rect 579 368 643 380
rect 679 580 733 592
rect 679 546 689 580
rect 723 546 733 580
rect 679 497 733 546
rect 679 463 689 497
rect 723 463 733 497
rect 679 414 733 463
rect 679 380 689 414
rect 723 380 733 414
rect 679 368 733 380
rect 769 580 835 592
rect 769 546 789 580
rect 823 546 835 580
rect 769 497 835 546
rect 769 463 789 497
rect 823 463 835 497
rect 769 414 835 463
rect 769 380 789 414
rect 823 380 835 414
rect 769 368 835 380
<< ndiffc >>
rect 42 176 76 210
rect 42 86 76 120
rect 128 176 162 210
rect 128 86 162 120
rect 214 118 248 152
rect 300 176 334 210
rect 300 86 334 120
rect 386 118 420 152
rect 486 176 520 210
rect 486 86 520 120
rect 586 158 620 192
rect 586 82 620 116
rect 686 176 720 210
rect 686 86 720 120
rect 772 160 806 194
rect 772 86 806 120
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 129 546 163 580
rect 129 476 163 510
rect 129 406 163 440
rect 219 546 253 580
rect 219 474 253 508
rect 319 546 353 580
rect 319 476 353 510
rect 319 406 353 440
rect 409 546 443 580
rect 409 474 443 508
rect 499 546 533 580
rect 499 463 533 497
rect 499 380 533 414
rect 589 546 623 580
rect 589 463 623 497
rect 589 380 623 414
rect 689 546 723 580
rect 689 463 723 497
rect 689 380 723 414
rect 789 546 823 580
rect 789 463 823 497
rect 789 380 823 414
<< poly >>
rect 83 592 119 618
rect 173 592 209 618
rect 273 592 309 618
rect 363 592 399 618
rect 453 592 489 618
rect 543 592 579 618
rect 643 592 679 618
rect 733 592 769 618
rect 83 336 119 368
rect 173 336 209 368
rect 273 336 309 368
rect 363 336 399 368
rect 453 336 489 368
rect 543 336 579 368
rect 643 336 679 368
rect 733 336 769 368
rect 83 320 769 336
rect 83 286 128 320
rect 162 286 196 320
rect 230 286 264 320
rect 298 286 332 320
rect 366 286 400 320
rect 434 286 769 320
rect 83 270 769 286
rect 83 240 203 270
rect 87 222 117 240
rect 173 222 203 240
rect 259 222 289 270
rect 345 222 375 270
rect 445 222 475 270
rect 531 222 561 270
rect 645 222 675 270
rect 731 222 761 270
rect 87 48 117 74
rect 173 48 203 74
rect 259 48 289 74
rect 345 48 375 74
rect 445 48 475 74
rect 531 48 561 74
rect 645 48 675 74
rect 731 48 761 74
<< polycont >>
rect 128 286 162 320
rect 196 286 230 320
rect 264 286 298 320
rect 332 286 366 320
rect 400 286 434 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 23 580 73 649
rect 23 546 39 580
rect 23 497 73 546
rect 23 463 39 497
rect 23 414 73 463
rect 23 380 39 414
rect 113 580 163 596
rect 113 546 129 580
rect 113 510 163 546
rect 113 476 129 510
rect 113 440 163 476
rect 203 580 269 649
rect 203 546 219 580
rect 253 546 269 580
rect 203 508 269 546
rect 203 474 219 508
rect 253 474 269 508
rect 203 458 269 474
rect 303 580 369 596
rect 303 546 319 580
rect 353 546 369 580
rect 303 510 369 546
rect 303 476 319 510
rect 353 476 369 510
rect 113 406 129 440
rect 303 440 369 476
rect 409 580 459 649
rect 443 546 459 580
rect 409 508 459 546
rect 443 474 459 508
rect 409 458 459 474
rect 499 580 533 596
rect 499 497 533 546
rect 303 424 319 440
rect 163 406 319 424
rect 353 424 369 440
rect 499 424 533 463
rect 353 414 533 424
rect 353 406 499 414
rect 113 390 499 406
rect 23 364 73 380
rect 112 320 450 356
rect 112 286 128 320
rect 162 286 196 320
rect 230 286 264 320
rect 298 286 332 320
rect 366 286 400 320
rect 434 286 450 320
rect 112 270 450 286
rect 499 324 533 380
rect 573 580 639 649
rect 573 546 589 580
rect 623 546 639 580
rect 573 497 639 546
rect 573 463 589 497
rect 623 463 639 497
rect 573 414 639 463
rect 573 380 589 414
rect 623 380 639 414
rect 573 364 639 380
rect 673 580 739 596
rect 673 546 689 580
rect 723 546 739 580
rect 673 497 739 546
rect 673 463 689 497
rect 723 463 739 497
rect 673 414 739 463
rect 673 380 689 414
rect 723 380 739 414
rect 673 324 739 380
rect 773 580 839 649
rect 773 546 789 580
rect 823 546 839 580
rect 773 497 839 546
rect 773 463 789 497
rect 823 463 839 497
rect 773 414 839 463
rect 773 380 789 414
rect 823 380 839 414
rect 773 364 839 380
rect 499 262 839 324
rect 484 236 839 262
rect 112 228 839 236
rect 26 210 76 226
rect 26 176 42 210
rect 26 120 76 176
rect 26 86 42 120
rect 26 17 76 86
rect 112 210 536 228
rect 112 176 128 210
rect 162 202 300 210
rect 112 120 162 176
rect 334 202 486 210
rect 112 86 128 120
rect 112 70 162 86
rect 198 152 264 168
rect 198 118 214 152
rect 248 118 264 152
rect 198 17 264 118
rect 300 120 334 176
rect 470 176 486 202
rect 520 176 536 210
rect 670 210 722 228
rect 300 70 334 86
rect 370 152 436 168
rect 370 118 386 152
rect 420 118 436 152
rect 370 17 436 118
rect 470 120 536 176
rect 470 86 486 120
rect 520 86 536 120
rect 470 70 536 86
rect 570 192 636 194
rect 570 158 586 192
rect 620 158 636 192
rect 570 116 636 158
rect 570 82 586 116
rect 620 82 636 116
rect 570 17 636 82
rect 670 176 686 210
rect 720 176 722 210
rect 670 120 722 176
rect 670 86 686 120
rect 720 86 722 120
rect 670 70 722 86
rect 756 160 772 194
rect 806 160 822 194
rect 756 120 822 160
rect 756 86 772 120
rect 806 86 822 120
rect 756 17 822 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew
flabel nbase s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew
rlabel comment s 0 0 0 0 4 inv_8
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 799 242 833 276 0 FreeSans 340 0 0 0 Y
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 864 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1820124
string GDS_START 1812808
<< end >>
