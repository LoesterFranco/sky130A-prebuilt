magic
tech sky130A
magscale 1 2
timestamp 1599588238
<< locali >>
rect 792 424 858 547
rect 972 424 1038 547
rect 473 390 1038 424
rect 473 364 743 390
rect 217 330 359 356
rect 89 264 359 330
rect 667 310 743 364
rect 409 236 633 310
rect 667 202 701 310
rect 793 270 1127 356
rect 456 168 701 202
rect 456 119 506 168
rect 644 119 701 168
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 23 364 73 649
rect 113 424 179 596
rect 219 458 253 649
rect 293 492 359 596
rect 399 526 449 649
rect 580 526 646 649
rect 692 581 1128 615
rect 692 492 758 581
rect 293 458 758 492
rect 293 424 359 458
rect 898 458 932 581
rect 113 390 359 424
rect 1078 390 1128 581
rect 113 364 179 390
rect 23 202 245 230
rect 23 196 420 202
rect 23 70 73 196
rect 211 168 420 196
rect 109 17 175 162
rect 211 70 245 168
rect 281 17 347 134
rect 386 85 420 168
rect 542 85 608 134
rect 735 202 1129 236
rect 735 85 769 202
rect 386 51 769 85
rect 805 17 871 168
rect 907 70 941 202
rect 977 17 1043 168
rect 1079 70 1129 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
rlabel locali s 217 330 359 356 6 A1
port 1 nsew signal input
rlabel locali s 89 264 359 330 6 A1
port 1 nsew signal input
rlabel locali s 793 270 1127 356 6 A2
port 2 nsew signal input
rlabel locali s 409 236 633 310 6 B1
port 3 nsew signal input
rlabel locali s 972 424 1038 547 6 Y
port 4 nsew signal output
rlabel locali s 792 424 858 547 6 Y
port 4 nsew signal output
rlabel locali s 667 310 743 364 6 Y
port 4 nsew signal output
rlabel locali s 667 202 701 310 6 Y
port 4 nsew signal output
rlabel locali s 644 119 701 168 6 Y
port 4 nsew signal output
rlabel locali s 473 390 1038 424 6 Y
port 4 nsew signal output
rlabel locali s 473 364 743 390 6 Y
port 4 nsew signal output
rlabel locali s 456 168 701 202 6 Y
port 4 nsew signal output
rlabel locali s 456 119 506 168 6 Y
port 4 nsew signal output
rlabel metal1 s 0 -49 1152 49 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1152 715 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1347034
string GDS_START 1336974
<< end >>
