magic
tech sky130A
magscale 1 2
timestamp 1604502710
<< nwell >>
rect -38 332 1670 704
<< pwell >>
rect 0 0 1632 49
<< scpmos >>
rect 83 368 119 592
rect 183 368 219 592
rect 273 368 309 592
rect 363 368 399 592
rect 453 368 489 592
rect 553 368 589 592
rect 643 368 679 592
rect 753 368 789 592
rect 843 368 879 592
rect 943 368 979 592
rect 1043 368 1079 592
rect 1133 368 1169 592
rect 1223 368 1259 592
rect 1313 368 1349 592
rect 1413 368 1449 592
rect 1503 368 1539 592
<< nmoslvt >>
rect 347 74 377 222
rect 447 74 477 222
rect 627 74 657 222
rect 727 74 757 222
rect 827 74 857 222
rect 1050 74 1080 222
rect 1164 74 1194 222
rect 1250 74 1280 222
<< ndiff >>
rect 134 210 347 222
rect 134 176 160 210
rect 194 176 231 210
rect 265 176 302 210
rect 336 176 347 210
rect 134 120 347 176
rect 134 86 160 120
rect 194 86 231 120
rect 265 86 302 120
rect 336 86 347 120
rect 134 74 347 86
rect 377 210 447 222
rect 377 176 388 210
rect 422 176 447 210
rect 377 120 447 176
rect 377 86 388 120
rect 422 86 447 120
rect 377 74 447 86
rect 477 152 627 222
rect 477 118 488 152
rect 522 118 582 152
rect 616 118 627 152
rect 477 74 627 118
rect 657 210 727 222
rect 657 176 668 210
rect 702 176 727 210
rect 657 120 727 176
rect 657 86 668 120
rect 702 86 727 120
rect 657 74 727 86
rect 757 152 827 222
rect 757 118 768 152
rect 802 118 827 152
rect 757 74 827 118
rect 857 210 1050 222
rect 857 176 868 210
rect 902 176 936 210
rect 970 176 1005 210
rect 1039 176 1050 210
rect 857 120 1050 176
rect 857 86 868 120
rect 902 86 936 120
rect 970 86 1005 120
rect 1039 86 1050 120
rect 857 74 1050 86
rect 1080 192 1164 222
rect 1080 158 1105 192
rect 1139 158 1164 192
rect 1080 120 1164 158
rect 1080 86 1105 120
rect 1139 86 1164 120
rect 1080 74 1164 86
rect 1194 210 1250 222
rect 1194 176 1205 210
rect 1239 176 1250 210
rect 1194 120 1250 176
rect 1194 86 1205 120
rect 1239 86 1250 120
rect 1194 74 1250 86
rect 1280 210 1351 222
rect 1280 176 1305 210
rect 1339 176 1351 210
rect 1280 120 1351 176
rect 1280 86 1305 120
rect 1339 86 1351 120
rect 1280 74 1351 86
<< pdiff >>
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 497 83 546
rect 27 463 39 497
rect 73 463 83 497
rect 27 414 83 463
rect 27 380 39 414
rect 73 380 83 414
rect 27 368 83 380
rect 119 580 183 592
rect 119 546 139 580
rect 173 546 183 580
rect 119 474 183 546
rect 119 440 139 474
rect 173 440 183 474
rect 119 368 183 440
rect 219 580 273 592
rect 219 546 229 580
rect 263 546 273 580
rect 219 504 273 546
rect 219 470 229 504
rect 263 470 273 504
rect 219 424 273 470
rect 219 390 229 424
rect 263 390 273 424
rect 219 368 273 390
rect 309 580 363 592
rect 309 546 319 580
rect 353 546 363 580
rect 309 508 363 546
rect 309 474 319 508
rect 353 474 363 508
rect 309 368 363 474
rect 399 580 453 592
rect 399 546 409 580
rect 443 546 453 580
rect 399 504 453 546
rect 399 470 409 504
rect 443 470 453 504
rect 399 424 453 470
rect 399 390 409 424
rect 443 390 453 424
rect 399 368 453 390
rect 489 580 553 592
rect 489 546 509 580
rect 543 546 553 580
rect 489 508 553 546
rect 489 474 509 508
rect 543 474 553 508
rect 489 368 553 474
rect 589 580 643 592
rect 589 546 599 580
rect 633 546 643 580
rect 589 504 643 546
rect 589 470 599 504
rect 633 470 643 504
rect 589 424 643 470
rect 589 390 599 424
rect 633 390 643 424
rect 589 368 643 390
rect 679 580 753 592
rect 679 546 699 580
rect 733 546 753 580
rect 679 508 753 546
rect 679 474 699 508
rect 733 474 753 508
rect 679 368 753 474
rect 789 580 843 592
rect 789 546 799 580
rect 833 546 843 580
rect 789 504 843 546
rect 789 470 799 504
rect 833 470 843 504
rect 789 424 843 470
rect 789 390 799 424
rect 833 390 843 424
rect 789 368 843 390
rect 879 547 943 592
rect 879 513 899 547
rect 933 513 943 547
rect 879 479 943 513
rect 879 445 899 479
rect 933 445 943 479
rect 879 411 943 445
rect 879 377 899 411
rect 933 377 943 411
rect 879 368 943 377
rect 979 580 1043 592
rect 979 546 999 580
rect 1033 546 1043 580
rect 979 510 1043 546
rect 979 476 999 510
rect 1033 476 1043 510
rect 979 440 1043 476
rect 979 406 999 440
rect 1033 406 1043 440
rect 979 368 1043 406
rect 1079 547 1133 592
rect 1079 513 1089 547
rect 1123 513 1133 547
rect 1079 479 1133 513
rect 1079 445 1089 479
rect 1123 445 1133 479
rect 1079 411 1133 445
rect 1079 377 1089 411
rect 1123 377 1133 411
rect 1079 368 1133 377
rect 1169 580 1223 592
rect 1169 546 1179 580
rect 1213 546 1223 580
rect 1169 497 1223 546
rect 1169 463 1179 497
rect 1213 463 1223 497
rect 1169 414 1223 463
rect 1169 380 1179 414
rect 1213 380 1223 414
rect 1169 368 1223 380
rect 1259 547 1313 592
rect 1259 513 1269 547
rect 1303 513 1313 547
rect 1259 479 1313 513
rect 1259 445 1269 479
rect 1303 445 1313 479
rect 1259 411 1313 445
rect 1259 377 1269 411
rect 1303 377 1313 411
rect 1259 368 1313 377
rect 1349 580 1413 592
rect 1349 546 1369 580
rect 1403 546 1413 580
rect 1349 497 1413 546
rect 1349 463 1369 497
rect 1403 463 1413 497
rect 1349 414 1413 463
rect 1349 380 1369 414
rect 1403 380 1413 414
rect 1349 368 1413 380
rect 1449 547 1503 592
rect 1449 513 1459 547
rect 1493 513 1503 547
rect 1449 479 1503 513
rect 1449 445 1459 479
rect 1493 445 1503 479
rect 1449 411 1503 445
rect 1449 377 1459 411
rect 1493 377 1503 411
rect 1449 368 1503 377
rect 1539 580 1605 592
rect 1539 546 1559 580
rect 1593 546 1605 580
rect 1539 497 1605 546
rect 1539 463 1559 497
rect 1593 463 1605 497
rect 1539 414 1605 463
rect 1539 380 1559 414
rect 1593 380 1605 414
rect 1539 368 1605 380
<< ndiffc >>
rect 160 176 194 210
rect 231 176 265 210
rect 302 176 336 210
rect 160 86 194 120
rect 231 86 265 120
rect 302 86 336 120
rect 388 176 422 210
rect 388 86 422 120
rect 488 118 522 152
rect 582 118 616 152
rect 668 176 702 210
rect 668 86 702 120
rect 768 118 802 152
rect 868 176 902 210
rect 936 176 970 210
rect 1005 176 1039 210
rect 868 86 902 120
rect 936 86 970 120
rect 1005 86 1039 120
rect 1105 158 1139 192
rect 1105 86 1139 120
rect 1205 176 1239 210
rect 1205 86 1239 120
rect 1305 176 1339 210
rect 1305 86 1339 120
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 139 546 173 580
rect 139 440 173 474
rect 229 546 263 580
rect 229 470 263 504
rect 229 390 263 424
rect 319 546 353 580
rect 319 474 353 508
rect 409 546 443 580
rect 409 470 443 504
rect 409 390 443 424
rect 509 546 543 580
rect 509 474 543 508
rect 599 546 633 580
rect 599 470 633 504
rect 599 390 633 424
rect 699 546 733 580
rect 699 474 733 508
rect 799 546 833 580
rect 799 470 833 504
rect 799 390 833 424
rect 899 513 933 547
rect 899 445 933 479
rect 899 377 933 411
rect 999 546 1033 580
rect 999 476 1033 510
rect 999 406 1033 440
rect 1089 513 1123 547
rect 1089 445 1123 479
rect 1089 377 1123 411
rect 1179 546 1213 580
rect 1179 463 1213 497
rect 1179 380 1213 414
rect 1269 513 1303 547
rect 1269 445 1303 479
rect 1269 377 1303 411
rect 1369 546 1403 580
rect 1369 463 1403 497
rect 1369 380 1403 414
rect 1459 513 1493 547
rect 1459 445 1493 479
rect 1459 377 1493 411
rect 1559 546 1593 580
rect 1559 463 1593 497
rect 1559 380 1593 414
<< poly >>
rect 83 592 119 618
rect 183 592 219 618
rect 273 592 309 618
rect 363 592 399 618
rect 453 592 489 618
rect 553 592 589 618
rect 643 592 679 618
rect 753 592 789 618
rect 843 592 879 618
rect 943 592 979 618
rect 1043 592 1079 618
rect 1133 592 1169 618
rect 1223 592 1259 618
rect 1313 592 1349 618
rect 1413 592 1449 618
rect 1503 592 1539 618
rect 83 345 119 368
rect 183 345 219 368
rect 273 345 309 368
rect 363 345 399 368
rect 453 345 489 368
rect 553 345 589 368
rect 643 345 679 368
rect 753 345 789 368
rect 83 320 789 345
rect 83 315 395 320
rect 347 286 395 315
rect 429 286 463 320
rect 497 286 531 320
rect 565 286 599 320
rect 633 286 667 320
rect 701 315 789 320
rect 701 286 757 315
rect 347 270 757 286
rect 347 222 377 270
rect 447 222 477 270
rect 627 222 657 270
rect 727 222 757 270
rect 843 267 879 368
rect 943 267 979 368
rect 1043 267 1079 368
rect 1133 267 1169 368
rect 1223 267 1259 368
rect 1313 267 1349 368
rect 1413 267 1449 368
rect 1503 267 1539 368
rect 827 246 1539 267
rect 827 237 1461 246
rect 827 222 857 237
rect 1050 222 1080 237
rect 1164 222 1194 237
rect 1250 222 1280 237
rect 1413 212 1461 237
rect 1495 212 1539 246
rect 1413 178 1539 212
rect 1413 144 1461 178
rect 1495 144 1539 178
rect 1413 110 1539 144
rect 1413 76 1461 110
rect 1495 76 1539 110
rect 347 48 377 74
rect 447 48 477 74
rect 627 48 657 74
rect 727 48 757 74
rect 827 48 857 74
rect 1050 48 1080 74
rect 1164 48 1194 74
rect 1250 48 1280 74
rect 1413 60 1539 76
<< polycont >>
rect 395 286 429 320
rect 463 286 497 320
rect 531 286 565 320
rect 599 286 633 320
rect 667 286 701 320
rect 1461 212 1495 246
rect 1461 144 1495 178
rect 1461 76 1495 110
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 23 580 89 596
rect 23 546 39 580
rect 73 546 89 580
rect 23 497 89 546
rect 23 463 39 497
rect 73 463 89 497
rect 23 414 89 463
rect 123 580 189 649
rect 123 546 139 580
rect 173 546 189 580
rect 123 474 189 546
rect 123 440 139 474
rect 173 440 189 474
rect 123 424 189 440
rect 229 580 263 596
rect 229 504 263 546
rect 229 424 263 470
rect 303 580 369 649
rect 303 546 319 580
rect 353 546 369 580
rect 303 508 369 546
rect 303 474 319 508
rect 353 474 369 508
rect 303 458 369 474
rect 409 580 459 596
rect 443 546 459 580
rect 409 504 459 546
rect 443 470 459 504
rect 409 424 459 470
rect 493 580 559 649
rect 493 546 509 580
rect 543 546 559 580
rect 493 508 559 546
rect 493 474 509 508
rect 543 474 559 508
rect 493 458 559 474
rect 599 580 649 596
rect 633 546 649 580
rect 599 504 649 546
rect 633 470 649 504
rect 599 424 649 470
rect 683 580 749 649
rect 683 546 699 580
rect 733 546 749 580
rect 683 508 749 546
rect 683 474 699 508
rect 733 474 749 508
rect 683 458 749 474
rect 783 581 1609 615
rect 783 580 849 581
rect 783 546 799 580
rect 833 546 849 580
rect 985 580 1037 581
rect 783 504 849 546
rect 783 470 799 504
rect 833 470 849 504
rect 783 424 849 470
rect 23 380 39 414
rect 73 390 89 414
rect 263 390 409 424
rect 443 390 599 424
rect 633 390 799 424
rect 833 390 849 424
rect 883 513 899 547
rect 933 513 949 547
rect 883 479 949 513
rect 883 445 899 479
rect 933 445 949 479
rect 883 411 949 445
rect 73 380 263 390
rect 23 356 263 380
rect 883 377 899 411
rect 933 377 949 411
rect 985 546 999 580
rect 1033 546 1037 580
rect 1175 580 1216 581
rect 985 510 1037 546
rect 985 476 999 510
rect 1033 476 1037 510
rect 985 440 1037 476
rect 985 406 999 440
rect 1033 406 1037 440
rect 985 390 1037 406
rect 1073 513 1089 547
rect 1123 513 1139 547
rect 1073 479 1139 513
rect 1073 445 1089 479
rect 1123 445 1139 479
rect 1073 411 1139 445
rect 883 356 949 377
rect 1073 377 1089 411
rect 1123 377 1139 411
rect 1073 356 1139 377
rect 1175 546 1179 580
rect 1213 546 1216 580
rect 1355 580 1407 581
rect 1175 497 1216 546
rect 1175 463 1179 497
rect 1213 463 1216 497
rect 1175 414 1216 463
rect 1175 380 1179 414
rect 1213 380 1216 414
rect 1175 364 1216 380
rect 1253 513 1269 547
rect 1303 513 1319 547
rect 1253 479 1319 513
rect 1253 445 1269 479
rect 1303 445 1319 479
rect 1253 411 1319 445
rect 1253 377 1269 411
rect 1303 377 1319 411
rect 313 320 743 356
rect 313 286 395 320
rect 429 286 463 320
rect 497 286 531 320
rect 565 286 599 320
rect 633 286 667 320
rect 701 286 743 320
rect 313 270 743 286
rect 883 330 1139 356
rect 1253 330 1319 377
rect 1355 546 1369 580
rect 1403 546 1407 580
rect 1543 580 1609 581
rect 1355 497 1407 546
rect 1355 463 1369 497
rect 1403 463 1407 497
rect 1355 414 1407 463
rect 1355 380 1369 414
rect 1403 380 1407 414
rect 1355 364 1407 380
rect 1443 513 1459 547
rect 1493 513 1509 547
rect 1443 479 1509 513
rect 1443 445 1459 479
rect 1493 445 1509 479
rect 1443 411 1509 445
rect 1443 377 1459 411
rect 1493 377 1509 411
rect 1443 330 1509 377
rect 1543 546 1559 580
rect 1593 546 1609 580
rect 1543 497 1609 546
rect 1543 463 1559 497
rect 1593 463 1609 497
rect 1543 414 1609 463
rect 1543 380 1559 414
rect 1593 380 1609 414
rect 1543 364 1609 380
rect 883 296 1509 330
rect 883 262 1255 296
rect 852 236 1255 262
rect 372 228 1255 236
rect 130 210 338 226
rect 130 176 160 210
rect 194 176 231 210
rect 265 176 302 210
rect 336 176 338 210
rect 130 120 338 176
rect 130 86 160 120
rect 194 86 231 120
rect 265 86 302 120
rect 336 86 338 120
rect 130 17 338 86
rect 372 210 1055 228
rect 372 176 388 210
rect 422 202 668 210
rect 422 176 438 202
rect 372 120 438 176
rect 652 176 668 202
rect 702 202 868 210
rect 702 176 718 202
rect 372 86 388 120
rect 422 86 438 120
rect 372 70 438 86
rect 472 152 618 168
rect 472 118 488 152
rect 522 118 582 152
rect 616 118 618 152
rect 472 17 618 118
rect 652 120 718 176
rect 852 176 868 202
rect 902 176 936 210
rect 970 176 1005 210
rect 1039 176 1055 210
rect 1189 210 1255 228
rect 1445 246 1511 262
rect 652 86 668 120
rect 702 86 718 120
rect 652 70 718 86
rect 752 152 818 168
rect 752 118 768 152
rect 802 118 818 152
rect 752 17 818 118
rect 852 120 1055 176
rect 852 86 868 120
rect 902 86 936 120
rect 970 86 1005 120
rect 1039 86 1055 120
rect 852 70 1055 86
rect 1089 192 1155 194
rect 1089 158 1105 192
rect 1139 158 1155 192
rect 1089 120 1155 158
rect 1089 86 1105 120
rect 1139 86 1155 120
rect 1089 17 1155 86
rect 1189 176 1205 210
rect 1239 176 1255 210
rect 1189 120 1255 176
rect 1189 86 1205 120
rect 1239 86 1255 120
rect 1189 70 1255 86
rect 1289 210 1355 226
rect 1289 176 1305 210
rect 1339 176 1355 210
rect 1289 120 1355 176
rect 1289 86 1305 120
rect 1339 86 1355 120
rect 1289 17 1355 86
rect 1445 212 1461 246
rect 1495 212 1511 246
rect 1445 178 1511 212
rect 1445 144 1461 178
rect 1495 144 1511 178
rect 1445 110 1511 144
rect 1445 76 1461 110
rect 1495 76 1511 110
rect 1445 60 1511 76
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
rlabel comment s 0 0 0 0 4 nor2_8
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 1471 94 1505 128 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 1471 168 1505 202 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 Y
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 1632 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1498920
string GDS_START 1487228
<< end >>
