magic
tech sky130A
magscale 1 2
timestamp 1601050082
<< locali >>
rect 21 236 87 310
rect 213 270 279 356
rect 313 270 455 356
rect 497 270 563 356
rect 601 270 677 356
rect 781 364 853 596
rect 819 226 853 364
rect 758 70 853 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 23 424 89 572
rect 123 458 305 649
rect 413 424 479 572
rect 681 458 747 649
rect 23 390 747 424
rect 23 364 155 390
rect 121 202 155 364
rect 713 330 747 390
rect 887 364 937 649
rect 713 264 785 330
rect 74 70 155 202
rect 189 104 223 226
rect 259 202 624 236
rect 259 160 324 202
rect 360 104 426 166
rect 189 70 426 104
rect 472 17 538 166
rect 574 70 624 202
rect 658 17 724 226
rect 887 17 937 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
rlabel locali s 601 270 677 356 6 A1
port 1 nsew signal input
rlabel locali s 497 270 563 356 6 A2
port 2 nsew signal input
rlabel locali s 213 270 279 356 6 B1
port 3 nsew signal input
rlabel locali s 313 270 455 356 6 B2
port 4 nsew signal input
rlabel locali s 21 236 87 310 6 C1
port 5 nsew signal input
rlabel locali s 819 226 853 364 6 X
port 6 nsew signal output
rlabel locali s 781 364 853 596 6 X
port 6 nsew signal output
rlabel locali s 758 70 853 226 6 X
port 6 nsew signal output
rlabel metal1 s 0 -49 960 49 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 617 960 715 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1512986
string GDS_START 1504652
<< end >>
