magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 503 425 579 459
rect 545 391 579 425
rect 85 289 433 323
rect 85 199 162 289
rect 196 215 355 255
rect 389 249 433 289
rect 545 351 719 391
rect 389 215 529 249
rect 671 165 719 351
rect 635 69 719 165
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 17 425 77 527
rect 111 391 187 493
rect 231 425 367 527
rect 623 425 683 527
rect 17 357 511 391
rect 17 165 51 357
rect 467 317 511 357
rect 467 283 619 317
rect 575 199 619 283
rect 17 56 110 165
rect 231 17 265 181
rect 299 131 579 165
rect 299 51 375 131
rect 419 17 499 95
rect 533 51 579 131
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel locali s 196 215 355 255 6 A
port 1 nsew signal input
rlabel locali s 389 249 433 289 6 B
port 2 nsew signal input
rlabel locali s 389 215 529 249 6 B
port 2 nsew signal input
rlabel locali s 85 289 433 323 6 B
port 2 nsew signal input
rlabel locali s 85 199 162 289 6 B
port 2 nsew signal input
rlabel locali s 671 165 719 351 6 Y
port 3 nsew signal output
rlabel locali s 635 69 719 165 6 Y
port 3 nsew signal output
rlabel locali s 545 391 579 425 6 Y
port 3 nsew signal output
rlabel locali s 545 351 719 391 6 Y
port 3 nsew signal output
rlabel locali s 503 425 579 459 6 Y
port 3 nsew signal output
rlabel metal1 s 0 -48 736 48 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 496 736 592 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 963308
string GDS_START 957716
<< end >>
