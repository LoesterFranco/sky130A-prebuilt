magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 183 425 299 493
rect 477 353 532 493
rect 17 127 137 204
rect 278 61 352 240
rect 498 147 532 353
rect 480 51 532 147
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 17 416 148 527
rect 382 418 433 527
rect 17 396 150 416
rect 103 391 150 396
rect 17 272 69 362
rect 103 342 179 391
rect 232 318 433 377
rect 232 308 454 318
rect 179 274 454 308
rect 179 272 215 274
rect 17 238 215 272
rect 171 93 215 238
rect 17 59 215 93
rect 408 198 454 274
rect 386 17 420 125
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
rlabel locali s 17 127 137 204 6 A
port 1 nsew signal input
rlabel locali s 183 425 299 493 6 B
port 2 nsew signal input
rlabel locali s 278 61 352 240 6 C
port 3 nsew signal input
rlabel locali s 498 147 532 353 6 X
port 4 nsew signal output
rlabel locali s 480 51 532 147 6 X
port 4 nsew signal output
rlabel locali s 477 353 532 493 6 X
port 4 nsew signal output
rlabel metal1 s 0 -48 552 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 552 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 552 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1517810
string GDS_START 1512672
<< end >>
