magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 17 364 87 596
rect 17 230 51 364
rect 317 290 367 356
rect 409 290 475 356
rect 17 196 215 230
rect 165 134 215 196
rect 601 114 647 134
rect 529 51 647 114
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 127 364 177 649
rect 249 390 321 596
rect 361 424 427 596
rect 467 458 507 649
rect 547 424 613 596
rect 361 390 613 424
rect 249 330 283 390
rect 547 388 613 390
rect 85 264 283 330
rect 249 256 283 264
rect 249 222 427 256
rect 251 17 317 188
rect 361 132 427 222
rect 542 202 608 268
rect 461 168 608 202
rect 461 17 495 168
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel locali s 409 290 475 356 6 A1
port 1 nsew signal input
rlabel locali s 601 114 647 134 6 A2
port 2 nsew signal input
rlabel locali s 529 51 647 114 6 A2
port 2 nsew signal input
rlabel locali s 317 290 367 356 6 B1
port 3 nsew signal input
rlabel locali s 165 134 215 196 6 X
port 4 nsew signal output
rlabel locali s 17 364 87 596 6 X
port 4 nsew signal output
rlabel locali s 17 230 51 364 6 X
port 4 nsew signal output
rlabel locali s 17 196 215 230 6 X
port 4 nsew signal output
rlabel metal1 s 0 -49 672 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 617 672 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 4084908
string GDS_START 4078508
<< end >>
