magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 552 561
rect 18 299 88 527
rect 18 215 88 265
rect 122 215 211 493
rect 292 265 340 481
rect 245 215 340 265
rect 35 17 69 181
rect 203 17 237 113
rect 389 165 432 493
rect 466 299 535 527
rect 466 199 535 265
rect 389 52 535 165
rect 0 -17 552 17
<< obsli1 >>
rect 103 147 340 181
rect 103 51 169 147
rect 274 51 340 147
<< metal1 >>
rect 0 496 552 592
rect 0 -48 552 48
<< labels >>
rlabel locali s 18 215 88 265 6 A1
port 1 nsew signal input
rlabel locali s 122 215 211 493 6 A2
port 2 nsew signal input
rlabel locali s 292 265 340 481 6 A3
port 3 nsew signal input
rlabel locali s 245 215 340 265 6 A3
port 3 nsew signal input
rlabel locali s 466 199 535 265 6 B1
port 4 nsew signal input
rlabel locali s 389 165 432 493 6 Y
port 5 nsew signal output
rlabel locali s 389 52 535 165 6 Y
port 5 nsew signal output
rlabel locali s 203 17 237 113 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 35 17 69 181 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 552 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 552 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 466 299 535 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 18 299 88 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 552 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 552 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 552 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 840362
string GDS_START 834088
<< end >>
