magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 92 53 122 137
rect 164 53 194 137
rect 255 53 285 137
rect 396 47 426 177
rect 494 47 524 177
<< pmoshvt >>
rect 83 311 119 395
rect 177 311 213 395
rect 282 297 318 381
rect 391 297 427 497
rect 485 297 521 497
<< ndiff >>
rect 325 137 396 177
rect 30 111 92 137
rect 30 77 38 111
rect 72 77 92 111
rect 30 53 92 77
rect 122 53 164 137
rect 194 53 255 137
rect 285 116 396 137
rect 285 82 313 116
rect 347 82 396 116
rect 285 53 396 82
rect 328 47 396 53
rect 426 123 494 177
rect 426 89 436 123
rect 470 89 494 123
rect 426 47 494 89
rect 524 120 584 177
rect 524 86 539 120
rect 573 86 584 120
rect 524 47 584 86
<< pdiff >>
rect 335 477 391 497
rect 335 443 345 477
rect 379 443 391 477
rect 335 408 391 443
rect 29 369 83 395
rect 29 335 37 369
rect 71 335 83 369
rect 29 311 83 335
rect 119 387 177 395
rect 119 353 131 387
rect 165 353 177 387
rect 119 311 177 353
rect 213 381 265 395
rect 335 381 345 408
rect 213 362 282 381
rect 213 328 236 362
rect 270 328 282 362
rect 213 311 282 328
rect 230 297 282 311
rect 318 374 345 381
rect 379 374 391 408
rect 318 297 391 374
rect 427 477 485 497
rect 427 443 439 477
rect 473 443 485 477
rect 427 409 485 443
rect 427 375 439 409
rect 473 375 485 409
rect 427 297 485 375
rect 521 477 600 497
rect 521 443 558 477
rect 592 443 600 477
rect 521 409 600 443
rect 521 375 558 409
rect 592 375 600 409
rect 521 297 600 375
<< ndiffc >>
rect 38 77 72 111
rect 313 82 347 116
rect 436 89 470 123
rect 539 86 573 120
<< pdiffc >>
rect 345 443 379 477
rect 37 335 71 369
rect 131 353 165 387
rect 236 328 270 362
rect 345 374 379 408
rect 439 443 473 477
rect 439 375 473 409
rect 558 443 592 477
rect 558 375 592 409
<< poly >>
rect 175 477 243 500
rect 391 497 427 523
rect 485 497 521 523
rect 175 443 189 477
rect 223 443 243 477
rect 175 427 243 443
rect 83 395 119 425
rect 175 421 215 427
rect 177 395 213 421
rect 282 381 318 407
rect 83 296 119 311
rect 177 296 213 311
rect 81 265 121 296
rect 164 279 213 296
rect 282 282 318 297
rect 391 282 427 297
rect 485 282 521 297
rect 28 249 122 265
rect 28 215 38 249
rect 72 215 122 249
rect 28 199 122 215
rect 92 137 122 199
rect 164 252 212 279
rect 280 265 320 282
rect 389 265 429 282
rect 483 265 523 282
rect 164 137 194 252
rect 255 249 322 265
rect 255 215 265 249
rect 299 215 322 249
rect 255 199 322 215
rect 364 249 524 265
rect 364 215 374 249
rect 408 215 524 249
rect 364 199 524 215
rect 255 137 285 199
rect 396 177 426 199
rect 494 177 524 199
rect 92 27 122 53
rect 164 27 194 53
rect 255 27 285 53
rect 396 21 426 47
rect 494 21 524 47
<< polycont >>
rect 189 443 223 477
rect 38 215 72 249
rect 265 215 299 249
rect 374 215 408 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 17 426 153 527
rect 20 369 71 392
rect 20 335 37 369
rect 105 391 153 426
rect 189 477 304 493
rect 223 443 304 477
rect 189 425 304 443
rect 341 477 384 527
rect 341 443 345 477
rect 379 443 384 477
rect 341 408 384 443
rect 105 387 181 391
rect 105 353 131 387
rect 165 353 181 387
rect 236 362 296 378
rect 20 319 71 335
rect 270 328 296 362
rect 341 374 345 408
rect 379 374 384 408
rect 341 358 384 374
rect 434 477 524 493
rect 434 443 439 477
rect 473 443 524 477
rect 434 409 524 443
rect 434 375 439 409
rect 473 375 524 409
rect 434 359 524 375
rect 236 319 296 328
rect 20 285 408 319
rect 17 215 38 249
rect 72 215 94 249
rect 17 153 94 215
rect 138 114 179 285
rect 362 249 408 285
rect 21 111 179 114
rect 21 77 38 111
rect 72 77 179 111
rect 21 61 179 77
rect 213 215 265 249
rect 299 215 325 249
rect 213 150 325 215
rect 362 215 374 249
rect 362 199 408 215
rect 452 289 524 359
rect 558 477 610 527
rect 592 443 610 477
rect 558 409 610 443
rect 592 375 610 409
rect 558 325 610 375
rect 452 185 585 289
rect 213 61 263 150
rect 452 143 486 185
rect 397 123 486 143
rect 297 82 313 116
rect 347 82 363 116
rect 297 17 363 82
rect 397 89 436 123
rect 470 89 486 123
rect 397 51 486 89
rect 539 120 594 149
rect 573 86 594 120
rect 539 17 594 86
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel corelocali s 230 442 230 442 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel corelocali s 402 85 436 119 0 FreeSans 200 0 0 0 X
port 8 nsew
flabel corelocali s 486 425 520 459 0 FreeSans 200 0 0 0 X
port 8 nsew
flabel corelocali s 29 153 63 187 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 215 153 249 187 0 FreeSans 400 0 0 0 C
port 3 nsew
flabel corelocali s 490 221 524 255 0 FreeSans 200 0 0 0 X
port 8 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 46 544 46 544 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
flabel metal1 s 46 0 46 0 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
rlabel comment s 0 0 0 0 4 and3_2
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1523932
string GDS_START 1517868
<< end >>
