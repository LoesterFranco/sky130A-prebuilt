magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 998 704
<< pwell >>
rect 0 0 960 49
<< scnmos >>
rect 97 74 127 222
rect 183 74 213 222
rect 417 74 447 222
rect 511 74 541 222
rect 597 74 627 222
rect 741 74 771 222
rect 813 74 843 222
<< pmoshvt >>
rect 94 368 124 592
rect 184 368 214 592
rect 414 368 444 592
rect 492 368 522 592
rect 600 368 630 592
rect 708 368 738 592
rect 816 368 846 592
<< ndiff >>
rect 44 210 97 222
rect 44 176 52 210
rect 86 176 97 210
rect 44 120 97 176
rect 44 86 52 120
rect 86 86 97 120
rect 44 74 97 86
rect 127 210 183 222
rect 127 176 138 210
rect 172 176 183 210
rect 127 120 183 176
rect 127 86 138 120
rect 172 86 183 120
rect 127 74 183 86
rect 213 152 266 222
rect 213 118 224 152
rect 258 118 266 152
rect 213 74 266 118
rect 364 210 417 222
rect 364 176 372 210
rect 406 176 417 210
rect 364 120 417 176
rect 364 86 372 120
rect 406 86 417 120
rect 364 74 417 86
rect 447 152 511 222
rect 447 118 462 152
rect 496 118 511 152
rect 447 74 511 118
rect 541 210 597 222
rect 541 176 552 210
rect 586 176 597 210
rect 541 120 597 176
rect 541 86 552 120
rect 586 86 597 120
rect 541 74 597 86
rect 627 152 741 222
rect 627 118 672 152
rect 706 118 741 152
rect 627 74 741 118
rect 771 74 813 222
rect 843 210 896 222
rect 843 176 854 210
rect 888 176 896 210
rect 843 120 896 176
rect 843 86 854 120
rect 888 86 896 120
rect 843 74 896 86
<< pdiff >>
rect 39 580 94 592
rect 39 546 47 580
rect 81 546 94 580
rect 39 497 94 546
rect 39 463 47 497
rect 81 463 94 497
rect 39 414 94 463
rect 39 380 47 414
rect 81 380 94 414
rect 39 368 94 380
rect 124 580 184 592
rect 124 546 137 580
rect 171 546 184 580
rect 124 497 184 546
rect 124 463 137 497
rect 171 463 184 497
rect 124 414 184 463
rect 124 380 137 414
rect 171 380 184 414
rect 124 368 184 380
rect 214 580 269 592
rect 214 546 227 580
rect 261 546 269 580
rect 214 508 269 546
rect 214 474 227 508
rect 261 474 269 508
rect 214 368 269 474
rect 359 580 414 592
rect 359 546 367 580
rect 401 546 414 580
rect 359 510 414 546
rect 359 476 367 510
rect 401 476 414 510
rect 359 440 414 476
rect 359 406 367 440
rect 401 406 414 440
rect 359 368 414 406
rect 444 368 492 592
rect 522 368 600 592
rect 630 580 708 592
rect 630 546 647 580
rect 681 546 708 580
rect 630 510 708 546
rect 630 476 647 510
rect 681 476 708 510
rect 630 440 708 476
rect 630 406 647 440
rect 681 406 708 440
rect 630 368 708 406
rect 738 580 816 592
rect 738 546 755 580
rect 789 546 816 580
rect 738 508 816 546
rect 738 474 755 508
rect 789 474 816 508
rect 738 368 816 474
rect 846 580 901 592
rect 846 546 859 580
rect 893 546 901 580
rect 846 510 901 546
rect 846 476 859 510
rect 893 476 901 510
rect 846 440 901 476
rect 846 406 859 440
rect 893 406 901 440
rect 846 368 901 406
<< ndiffc >>
rect 52 176 86 210
rect 52 86 86 120
rect 138 176 172 210
rect 138 86 172 120
rect 224 118 258 152
rect 372 176 406 210
rect 372 86 406 120
rect 462 118 496 152
rect 552 176 586 210
rect 552 86 586 120
rect 672 118 706 152
rect 854 176 888 210
rect 854 86 888 120
<< pdiffc >>
rect 47 546 81 580
rect 47 463 81 497
rect 47 380 81 414
rect 137 546 171 580
rect 137 463 171 497
rect 137 380 171 414
rect 227 546 261 580
rect 227 474 261 508
rect 367 546 401 580
rect 367 476 401 510
rect 367 406 401 440
rect 647 546 681 580
rect 647 476 681 510
rect 647 406 681 440
rect 755 546 789 580
rect 755 474 789 508
rect 859 546 893 580
rect 859 476 893 510
rect 859 406 893 440
<< poly >>
rect 94 592 124 618
rect 184 592 214 618
rect 414 592 444 618
rect 492 592 522 618
rect 600 592 630 618
rect 708 592 738 618
rect 816 592 846 618
rect 94 353 124 368
rect 184 353 214 368
rect 414 353 444 368
rect 492 353 522 368
rect 600 353 630 368
rect 708 353 738 368
rect 816 353 846 368
rect 91 310 127 353
rect 181 310 217 353
rect 411 336 447 353
rect 381 320 447 336
rect 91 294 272 310
rect 91 260 222 294
rect 256 260 272 294
rect 381 286 397 320
rect 431 286 447 320
rect 381 270 447 286
rect 489 336 525 353
rect 597 336 633 353
rect 705 336 741 353
rect 813 336 849 353
rect 489 320 555 336
rect 489 286 505 320
rect 539 286 555 320
rect 489 270 555 286
rect 597 320 663 336
rect 597 286 613 320
rect 647 286 663 320
rect 597 270 663 286
rect 705 320 771 336
rect 705 286 721 320
rect 755 286 771 320
rect 705 270 771 286
rect 91 244 272 260
rect 97 222 127 244
rect 183 222 213 244
rect 417 222 447 270
rect 511 222 541 270
rect 597 222 627 270
rect 741 222 771 270
rect 813 320 939 336
rect 813 286 889 320
rect 923 286 939 320
rect 813 270 939 286
rect 813 222 843 270
rect 97 48 127 74
rect 183 48 213 74
rect 417 48 447 74
rect 511 48 541 74
rect 597 48 627 74
rect 741 48 771 74
rect 813 48 843 74
<< polycont >>
rect 222 260 256 294
rect 397 286 431 320
rect 505 286 539 320
rect 613 286 647 320
rect 721 286 755 320
rect 889 286 923 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 31 580 81 649
rect 31 546 47 580
rect 31 497 81 546
rect 31 463 47 497
rect 31 414 81 463
rect 31 380 47 414
rect 31 364 81 380
rect 121 580 172 596
rect 121 546 137 580
rect 171 546 172 580
rect 121 497 172 546
rect 121 463 137 497
rect 171 463 172 497
rect 121 414 172 463
rect 211 580 277 649
rect 211 546 227 580
rect 261 546 277 580
rect 211 508 277 546
rect 211 474 227 508
rect 261 474 277 508
rect 211 458 277 474
rect 351 580 417 596
rect 351 546 367 580
rect 401 546 417 580
rect 627 580 701 596
rect 351 510 417 546
rect 351 476 367 510
rect 401 476 417 510
rect 351 440 417 476
rect 351 424 367 440
rect 121 380 137 414
rect 171 380 172 414
rect 121 310 172 380
rect 238 406 367 424
rect 401 406 417 440
rect 238 390 417 406
rect 238 310 272 390
rect 36 210 102 226
rect 36 176 52 210
rect 86 176 102 210
rect 36 120 102 176
rect 36 86 52 120
rect 86 86 102 120
rect 36 17 102 86
rect 138 210 172 310
rect 206 294 272 310
rect 206 260 222 294
rect 256 260 272 294
rect 313 320 455 356
rect 313 286 397 320
rect 431 286 455 320
rect 313 270 455 286
rect 489 320 555 578
rect 627 546 647 580
rect 681 546 701 580
rect 627 510 701 546
rect 627 476 647 510
rect 681 476 701 510
rect 627 440 701 476
rect 735 580 809 649
rect 735 546 755 580
rect 789 546 809 580
rect 735 508 809 546
rect 735 474 755 508
rect 789 474 809 508
rect 735 458 809 474
rect 843 580 909 596
rect 843 546 859 580
rect 893 546 909 580
rect 843 510 909 546
rect 843 476 859 510
rect 893 476 909 510
rect 627 406 647 440
rect 681 424 701 440
rect 843 440 909 476
rect 843 424 859 440
rect 681 406 859 424
rect 893 406 909 440
rect 627 390 909 406
rect 489 286 505 320
rect 539 286 555 320
rect 489 270 555 286
rect 597 320 663 356
rect 597 286 613 320
rect 647 286 663 320
rect 597 270 663 286
rect 697 320 839 356
rect 697 286 721 320
rect 755 286 839 320
rect 697 270 839 286
rect 873 320 939 356
rect 873 286 889 320
rect 923 286 939 320
rect 873 270 939 286
rect 206 244 272 260
rect 238 236 272 244
rect 238 210 904 236
rect 238 202 372 210
rect 138 120 172 176
rect 356 176 372 202
rect 406 202 552 210
rect 138 70 172 86
rect 208 152 274 168
rect 208 118 224 152
rect 258 118 274 152
rect 208 17 274 118
rect 356 120 406 176
rect 586 202 854 210
rect 586 176 602 202
rect 356 86 372 120
rect 356 70 406 86
rect 442 152 516 168
rect 442 118 462 152
rect 496 118 516 152
rect 442 17 516 118
rect 552 120 602 176
rect 838 176 854 202
rect 888 176 904 210
rect 586 86 602 120
rect 552 70 602 86
rect 636 152 746 168
rect 636 118 672 152
rect 706 118 746 152
rect 636 17 746 118
rect 838 120 904 176
rect 838 86 854 120
rect 888 86 904 120
rect 838 70 904 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a2111o_2
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 D1
port 5 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 D1
port 5 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 511 390 545 424 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 511 464 545 498 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 511 538 545 572 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 X
port 10 nsew
flabel corelocali s 127 390 161 424 0 FreeSans 340 0 0 0 X
port 10 nsew
flabel corelocali s 127 464 161 498 0 FreeSans 340 0 0 0 X
port 10 nsew
flabel corelocali s 127 538 161 572 0 FreeSans 340 0 0 0 X
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 960 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3893854
string GDS_START 3884908
<< end >>
