magic
tech sky130A
magscale 1 2
timestamp 1604502729
<< locali >>
rect 25 270 110 356
rect 212 360 845 414
rect 212 226 278 360
rect 212 192 850 226
rect 212 176 650 192
rect 212 70 278 176
rect 412 70 450 176
rect 584 70 650 176
rect 784 70 850 192
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 23 482 89 596
rect 123 516 189 649
rect 303 516 369 649
rect 483 516 549 649
rect 663 516 729 649
rect 869 516 935 649
rect 23 448 913 482
rect 23 390 89 448
rect 144 236 178 448
rect 26 202 178 236
rect 879 394 913 448
rect 969 462 1035 596
rect 1069 496 1135 649
rect 1169 462 1225 596
rect 969 428 1225 462
rect 879 360 1121 394
rect 333 260 964 326
rect 998 264 1121 360
rect 930 226 964 260
rect 1159 226 1225 428
rect 26 70 76 202
rect 112 17 178 168
rect 312 17 378 142
rect 484 17 550 142
rect 684 17 750 158
rect 930 176 1225 226
rect 884 17 950 142
rect 984 70 1025 176
rect 1059 17 1125 142
rect 1159 70 1225 176
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
<< metal1 >>
rect 0 683 1248 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 0 617 1248 649
rect 0 17 1248 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
rect 0 -49 1248 -17
<< labels >>
rlabel locali s 25 270 110 356 6 A
port 1 nsew signal input
rlabel locali s 784 70 850 192 6 Y
port 2 nsew signal output
rlabel locali s 584 70 650 176 6 Y
port 2 nsew signal output
rlabel locali s 412 70 450 176 6 Y
port 2 nsew signal output
rlabel locali s 212 360 845 414 6 Y
port 2 nsew signal output
rlabel locali s 212 226 278 360 6 Y
port 2 nsew signal output
rlabel locali s 212 192 850 226 6 Y
port 2 nsew signal output
rlabel locali s 212 176 650 192 6 Y
port 2 nsew signal output
rlabel locali s 212 70 278 176 6 Y
port 2 nsew signal output
rlabel metal1 s 0 -49 1248 49 8 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 617 1248 715 6 VPWR
port 4 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1248 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3419406
string GDS_START 3410234
<< end >>
