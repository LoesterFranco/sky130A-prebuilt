magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 920 561
rect 138 442 215 527
rect 17 199 114 340
rect 249 335 334 493
rect 457 442 534 527
rect 249 299 430 335
rect 264 199 430 299
rect 740 442 817 527
rect 264 165 334 199
rect 138 17 215 97
rect 249 51 334 165
rect 457 17 534 97
rect 740 17 817 97
rect 0 -17 920 17
<< obsli1 >>
rect 17 408 104 493
rect 17 374 215 408
rect 148 265 215 374
rect 368 408 423 493
rect 368 369 534 408
rect 148 199 230 265
rect 464 265 534 369
rect 568 335 617 493
rect 655 408 706 493
rect 655 369 817 408
rect 568 299 713 335
rect 464 199 549 265
rect 583 199 713 299
rect 747 265 817 369
rect 851 299 903 493
rect 747 199 832 265
rect 148 165 215 199
rect 464 165 534 199
rect 583 165 617 199
rect 747 165 817 199
rect 866 165 903 299
rect 17 131 215 165
rect 17 51 104 131
rect 372 131 534 165
rect 372 51 423 131
rect 568 51 617 165
rect 655 131 817 165
rect 655 51 706 131
rect 851 51 903 165
<< metal1 >>
rect 0 496 920 592
rect 0 -48 920 48
<< labels >>
rlabel locali s 17 199 114 340 6 A
port 1 nsew signal input
rlabel locali s 264 199 430 299 6 X
port 2 nsew signal output
rlabel locali s 264 165 334 199 6 X
port 2 nsew signal output
rlabel locali s 249 335 334 493 6 X
port 2 nsew signal output
rlabel locali s 249 299 430 335 6 X
port 2 nsew signal output
rlabel locali s 249 51 334 165 6 X
port 2 nsew signal output
rlabel locali s 740 17 817 97 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 457 17 534 97 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 138 17 215 97 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 0 -17 920 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 920 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 740 442 817 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 457 442 534 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 138 442 215 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 0 527 920 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 496 920 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 920 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2831352
string GDS_START 2823576
<< end >>
