magic
tech sky130A
magscale 1 2
timestamp 1601050047
<< nwell >>
rect -38 332 2054 704
<< pwell >>
rect 0 0 2016 49
<< scpmos >>
rect 86 373 116 573
rect 186 373 216 573
rect 294 373 324 541
rect 434 373 464 501
rect 524 373 554 501
rect 626 373 656 541
rect 851 368 881 592
rect 1053 398 1083 566
rect 1177 398 1207 566
rect 1389 368 1419 496
rect 1629 368 1659 592
rect 1719 368 1749 592
rect 1809 368 1839 592
rect 1899 368 1929 592
<< nmoslvt >>
rect 94 77 124 205
rect 194 77 224 205
rect 291 77 321 205
rect 386 121 416 205
rect 509 121 539 249
rect 599 121 629 249
rect 813 89 843 237
rect 1027 74 1057 202
rect 1138 74 1168 202
rect 1339 162 1369 246
rect 1644 98 1674 246
rect 1730 98 1760 246
rect 1816 98 1846 246
rect 1902 98 1932 246
<< ndiff >>
rect 431 237 509 249
rect 431 205 443 237
rect 37 140 94 205
rect 37 106 49 140
rect 83 106 94 140
rect 37 77 94 106
rect 124 140 194 205
rect 124 106 149 140
rect 183 106 194 140
rect 124 77 194 106
rect 224 193 291 205
rect 224 159 235 193
rect 269 159 291 193
rect 224 123 291 159
rect 224 89 235 123
rect 269 89 291 123
rect 224 77 291 89
rect 321 176 386 205
rect 321 142 341 176
rect 375 142 386 176
rect 321 121 386 142
rect 416 203 443 205
rect 477 203 509 237
rect 416 121 509 203
rect 539 225 599 249
rect 539 191 552 225
rect 586 191 599 225
rect 539 121 599 191
rect 629 121 702 249
rect 321 77 371 121
rect 644 89 702 121
rect 756 225 813 237
rect 756 191 768 225
rect 802 191 813 225
rect 756 89 813 191
rect 843 89 916 237
rect 1282 234 1339 246
rect 644 55 656 89
rect 690 55 702 89
rect 644 43 702 55
rect 858 55 870 89
rect 904 55 916 89
rect 970 190 1027 202
rect 970 156 982 190
rect 1016 156 1027 190
rect 970 120 1027 156
rect 970 86 982 120
rect 1016 86 1027 120
rect 970 74 1027 86
rect 1057 188 1138 202
rect 1057 154 1082 188
rect 1116 154 1138 188
rect 1057 120 1138 154
rect 1057 86 1082 120
rect 1116 86 1138 120
rect 1057 74 1138 86
rect 1168 179 1228 202
rect 1168 145 1182 179
rect 1216 145 1228 179
rect 1282 200 1294 234
rect 1328 200 1339 234
rect 1282 162 1339 200
rect 1369 218 1644 246
rect 1369 184 1599 218
rect 1633 184 1644 218
rect 1369 162 1644 184
rect 1168 74 1228 145
rect 1384 152 1644 162
rect 1384 118 1446 152
rect 1480 118 1524 152
rect 1558 150 1644 152
rect 1558 118 1599 150
rect 1384 116 1599 118
rect 1633 116 1644 150
rect 1384 98 1644 116
rect 1674 218 1730 246
rect 1674 184 1685 218
rect 1719 184 1730 218
rect 1674 144 1730 184
rect 1674 110 1685 144
rect 1719 110 1730 144
rect 1674 98 1730 110
rect 1760 234 1816 246
rect 1760 200 1771 234
rect 1805 200 1816 234
rect 1760 144 1816 200
rect 1760 110 1771 144
rect 1805 110 1816 144
rect 1760 98 1816 110
rect 1846 234 1902 246
rect 1846 200 1857 234
rect 1891 200 1902 234
rect 1846 144 1902 200
rect 1846 110 1857 144
rect 1891 110 1902 144
rect 1846 98 1902 110
rect 1932 234 1989 246
rect 1932 200 1943 234
rect 1977 200 1989 234
rect 1932 144 1989 200
rect 1932 110 1943 144
rect 1977 110 1989 144
rect 1932 98 1989 110
rect 1384 82 1629 98
rect 858 43 916 55
rect 1384 48 1396 82
rect 1430 48 1489 82
rect 1523 48 1583 82
rect 1617 48 1629 82
rect 1384 36 1629 48
<< pdiff >>
rect 27 561 86 573
rect 27 527 39 561
rect 73 527 86 561
rect 27 490 86 527
rect 27 456 39 490
rect 73 456 86 490
rect 27 419 86 456
rect 27 385 39 419
rect 73 385 86 419
rect 27 373 86 385
rect 116 560 186 573
rect 116 526 129 560
rect 163 526 186 560
rect 116 492 186 526
rect 116 458 129 492
rect 163 458 186 492
rect 116 373 186 458
rect 216 561 275 573
rect 216 527 229 561
rect 263 541 275 561
rect 263 527 294 541
rect 216 492 294 527
rect 216 458 229 492
rect 263 458 294 492
rect 216 424 294 458
rect 216 390 229 424
rect 263 390 294 424
rect 216 373 294 390
rect 324 501 377 541
rect 674 576 732 588
rect 674 542 686 576
rect 720 542 732 576
rect 674 541 732 542
rect 573 501 626 541
rect 324 415 434 501
rect 324 381 387 415
rect 421 381 434 415
rect 324 373 434 381
rect 464 493 524 501
rect 464 459 477 493
rect 511 459 524 493
rect 464 373 524 459
rect 554 493 626 501
rect 554 459 579 493
rect 613 459 626 493
rect 554 425 626 459
rect 554 391 579 425
rect 613 391 626 425
rect 554 373 626 391
rect 656 373 732 541
rect 1101 596 1159 608
rect 792 440 851 592
rect 792 406 804 440
rect 838 406 851 440
rect 792 368 851 406
rect 881 580 940 592
rect 881 546 894 580
rect 928 546 940 580
rect 1101 566 1113 596
rect 881 368 940 546
rect 994 444 1053 566
rect 994 410 1006 444
rect 1040 410 1053 444
rect 994 398 1053 410
rect 1083 562 1113 566
rect 1147 566 1159 596
rect 1466 580 1629 592
rect 1147 562 1177 566
rect 1083 398 1177 562
rect 1207 531 1266 566
rect 1207 497 1220 531
rect 1254 497 1266 531
rect 1466 546 1497 580
rect 1531 546 1582 580
rect 1616 546 1629 580
rect 1207 444 1266 497
rect 1466 508 1629 546
rect 1466 496 1497 508
rect 1207 410 1220 444
rect 1254 410 1266 444
rect 1207 398 1266 410
rect 1330 464 1389 496
rect 1330 430 1342 464
rect 1376 430 1389 464
rect 1330 368 1389 430
rect 1419 474 1497 496
rect 1531 499 1629 508
rect 1531 474 1582 499
rect 1419 465 1582 474
rect 1616 465 1629 499
rect 1419 418 1629 465
rect 1419 384 1537 418
rect 1571 384 1629 418
rect 1419 368 1629 384
rect 1659 580 1719 592
rect 1659 546 1672 580
rect 1706 546 1719 580
rect 1659 499 1719 546
rect 1659 465 1672 499
rect 1706 465 1719 499
rect 1659 418 1719 465
rect 1659 384 1672 418
rect 1706 384 1719 418
rect 1659 368 1719 384
rect 1749 580 1809 592
rect 1749 546 1762 580
rect 1796 546 1809 580
rect 1749 497 1809 546
rect 1749 463 1762 497
rect 1796 463 1809 497
rect 1749 414 1809 463
rect 1749 380 1762 414
rect 1796 380 1809 414
rect 1749 368 1809 380
rect 1839 580 1899 592
rect 1839 546 1852 580
rect 1886 546 1899 580
rect 1839 497 1899 546
rect 1839 463 1852 497
rect 1886 463 1899 497
rect 1839 414 1899 463
rect 1839 380 1852 414
rect 1886 380 1899 414
rect 1839 368 1899 380
rect 1929 580 1988 592
rect 1929 546 1942 580
rect 1976 546 1988 580
rect 1929 497 1988 546
rect 1929 463 1942 497
rect 1976 463 1988 497
rect 1929 414 1988 463
rect 1929 380 1942 414
rect 1976 380 1988 414
rect 1929 368 1988 380
<< ndiffc >>
rect 49 106 83 140
rect 149 106 183 140
rect 235 159 269 193
rect 235 89 269 123
rect 341 142 375 176
rect 443 203 477 237
rect 552 191 586 225
rect 768 191 802 225
rect 656 55 690 89
rect 870 55 904 89
rect 982 156 1016 190
rect 982 86 1016 120
rect 1082 154 1116 188
rect 1082 86 1116 120
rect 1182 145 1216 179
rect 1294 200 1328 234
rect 1599 184 1633 218
rect 1446 118 1480 152
rect 1524 118 1558 152
rect 1599 116 1633 150
rect 1685 184 1719 218
rect 1685 110 1719 144
rect 1771 200 1805 234
rect 1771 110 1805 144
rect 1857 200 1891 234
rect 1857 110 1891 144
rect 1943 200 1977 234
rect 1943 110 1977 144
rect 1396 48 1430 82
rect 1489 48 1523 82
rect 1583 48 1617 82
<< pdiffc >>
rect 39 527 73 561
rect 39 456 73 490
rect 39 385 73 419
rect 129 526 163 560
rect 129 458 163 492
rect 229 527 263 561
rect 229 458 263 492
rect 229 390 263 424
rect 686 542 720 576
rect 387 381 421 415
rect 477 459 511 493
rect 579 459 613 493
rect 579 391 613 425
rect 804 406 838 440
rect 894 546 928 580
rect 1006 410 1040 444
rect 1113 562 1147 596
rect 1220 497 1254 531
rect 1497 546 1531 580
rect 1582 546 1616 580
rect 1220 410 1254 444
rect 1342 430 1376 464
rect 1497 474 1531 508
rect 1582 465 1616 499
rect 1537 384 1571 418
rect 1672 546 1706 580
rect 1672 465 1706 499
rect 1672 384 1706 418
rect 1762 546 1796 580
rect 1762 463 1796 497
rect 1762 380 1796 414
rect 1852 546 1886 580
rect 1852 463 1886 497
rect 1852 380 1886 414
rect 1942 546 1976 580
rect 1942 463 1976 497
rect 1942 380 1976 414
<< poly >>
rect 291 615 777 645
rect 86 573 116 599
rect 186 573 216 599
rect 291 556 327 615
rect 294 541 324 556
rect 434 501 464 527
rect 521 516 557 615
rect 626 541 656 567
rect 524 501 554 516
rect 86 358 116 373
rect 186 358 216 373
rect 294 358 324 373
rect 434 358 464 373
rect 524 358 554 373
rect 626 358 656 373
rect 83 293 119 358
rect 183 341 219 358
rect 183 325 249 341
rect 75 277 141 293
rect 75 243 91 277
rect 125 243 141 277
rect 183 291 199 325
rect 233 291 249 325
rect 183 275 249 291
rect 291 328 327 358
rect 75 227 141 243
rect 94 205 124 227
rect 194 205 224 275
rect 291 205 321 328
rect 431 294 467 358
rect 386 264 467 294
rect 509 328 557 358
rect 623 341 659 358
rect 386 205 416 264
rect 509 249 539 328
rect 599 325 665 341
rect 599 291 615 325
rect 649 291 665 325
rect 747 336 777 615
rect 851 592 881 618
rect 1053 566 1083 592
rect 1629 592 1659 618
rect 1719 592 1749 618
rect 1809 592 1839 618
rect 1899 592 1929 618
rect 1177 566 1207 592
rect 1389 496 1419 522
rect 1053 383 1083 398
rect 1177 383 1207 398
rect 851 353 881 368
rect 1050 366 1086 383
rect 848 336 884 353
rect 747 320 884 336
rect 747 306 804 320
rect 599 275 665 291
rect 788 286 804 306
rect 838 286 884 320
rect 1024 350 1090 366
rect 1024 316 1040 350
rect 1074 316 1090 350
rect 1024 300 1090 316
rect 1174 300 1210 383
rect 1389 353 1419 368
rect 1629 353 1659 368
rect 1719 353 1749 368
rect 1809 353 1839 368
rect 1899 353 1929 368
rect 1386 336 1422 353
rect 1339 320 1422 336
rect 1626 334 1662 353
rect 1716 334 1752 353
rect 1806 334 1842 353
rect 1339 300 1372 320
rect 599 249 629 275
rect 788 270 884 286
rect 813 237 843 270
rect 94 51 124 77
rect 194 51 224 77
rect 291 51 321 77
rect 386 53 416 121
rect 509 95 539 121
rect 599 53 629 121
rect 386 23 629 53
rect 1027 202 1057 300
rect 1138 286 1372 300
rect 1406 286 1422 320
rect 1138 270 1422 286
rect 1464 333 1842 334
rect 1896 333 1932 353
rect 1464 318 1932 333
rect 1464 284 1480 318
rect 1514 284 1548 318
rect 1582 284 1616 318
rect 1650 284 1932 318
rect 1138 202 1168 270
rect 1339 246 1369 270
rect 1464 268 1932 284
rect 1644 246 1674 268
rect 1730 246 1760 268
rect 1816 246 1846 268
rect 1902 246 1932 268
rect 813 63 843 89
rect 1339 136 1369 162
rect 1027 48 1057 74
rect 1138 48 1168 74
rect 1644 72 1674 98
rect 1730 72 1760 98
rect 1816 72 1846 98
rect 1902 72 1932 98
<< polycont >>
rect 91 243 125 277
rect 199 291 233 325
rect 615 291 649 325
rect 804 286 838 320
rect 1040 316 1074 350
rect 1372 286 1406 320
rect 1480 284 1514 318
rect 1548 284 1582 318
rect 1616 284 1650 318
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 17 561 73 577
rect 17 527 39 561
rect 17 490 73 527
rect 17 456 39 490
rect 113 560 179 649
rect 113 526 129 560
rect 163 526 179 560
rect 113 492 179 526
rect 113 458 129 492
rect 163 458 179 492
rect 213 581 736 615
rect 213 561 279 581
rect 213 527 229 561
rect 263 527 279 561
rect 670 576 736 581
rect 213 492 279 527
rect 213 458 229 492
rect 263 458 279 492
rect 17 424 73 456
rect 213 424 279 458
rect 17 390 31 424
rect 65 419 73 424
rect 17 385 39 390
rect 17 369 73 385
rect 107 390 229 424
rect 263 390 279 424
rect 313 513 545 547
rect 670 542 686 576
rect 720 542 736 576
rect 878 580 944 649
rect 878 546 894 580
rect 928 546 944 580
rect 1097 596 1463 615
rect 1097 562 1113 596
rect 1147 581 1463 596
rect 1147 562 1163 581
rect 1097 546 1163 562
rect 313 424 353 513
rect 461 493 545 513
rect 1204 531 1254 547
rect 1204 512 1220 531
rect 461 459 477 493
rect 511 459 545 493
rect 461 458 545 459
rect 579 508 629 509
rect 888 508 1220 512
rect 579 497 1220 508
rect 579 493 1254 497
rect 613 478 1254 493
rect 613 474 922 478
rect 613 459 629 474
rect 313 390 319 424
rect 17 173 57 369
rect 107 293 141 390
rect 91 277 141 293
rect 125 243 141 277
rect 183 325 263 356
rect 183 291 199 325
rect 233 291 263 325
rect 183 275 263 291
rect 313 275 353 390
rect 387 424 427 431
rect 579 425 629 459
rect 387 415 415 424
rect 421 381 449 390
rect 387 335 449 381
rect 613 391 629 425
rect 579 375 629 391
rect 720 406 804 440
rect 838 406 854 440
rect 720 390 854 406
rect 720 341 754 390
rect 387 301 551 335
rect 91 241 141 243
rect 319 267 353 275
rect 91 207 285 241
rect 319 237 477 267
rect 319 233 443 237
rect 235 193 285 207
rect 427 203 443 233
rect 17 140 99 173
rect 17 106 49 140
rect 83 106 99 140
rect 17 73 99 106
rect 133 140 199 173
rect 133 106 149 140
rect 183 106 199 140
rect 133 17 199 106
rect 269 159 285 193
rect 235 123 285 159
rect 269 89 285 123
rect 325 176 391 199
rect 427 187 477 203
rect 511 241 551 301
rect 599 325 754 341
rect 599 291 615 325
rect 649 291 754 325
rect 599 275 754 291
rect 511 225 604 241
rect 511 191 552 225
rect 586 191 604 225
rect 720 225 754 275
rect 788 320 854 356
rect 788 286 804 320
rect 838 286 854 320
rect 788 270 854 286
rect 720 191 768 225
rect 802 191 818 225
rect 888 206 922 474
rect 1204 444 1254 478
rect 956 424 1006 444
rect 956 390 991 424
rect 1040 410 1056 444
rect 1025 390 1056 410
rect 1204 410 1220 444
rect 1204 394 1254 410
rect 1288 464 1392 500
rect 1288 430 1342 464
rect 1376 430 1392 464
rect 1288 398 1392 430
rect 1426 424 1463 581
rect 1497 580 1622 649
rect 1531 546 1582 580
rect 1616 546 1622 580
rect 1497 508 1622 546
rect 1531 499 1622 508
rect 1531 474 1582 499
rect 1497 465 1582 474
rect 1616 465 1622 499
rect 1497 458 1622 465
rect 956 276 990 390
rect 1024 350 1090 356
rect 1024 316 1040 350
rect 1074 344 1090 350
rect 1288 344 1322 398
rect 1426 390 1498 424
rect 1074 316 1322 344
rect 1024 310 1322 316
rect 956 242 1232 276
rect 1081 236 1232 242
rect 888 190 1032 206
rect 325 142 341 176
rect 375 153 391 176
rect 888 157 982 190
rect 511 156 982 157
rect 1016 156 1032 190
rect 511 153 1032 156
rect 375 142 1032 153
rect 325 123 1032 142
rect 325 119 545 123
rect 966 120 1032 123
rect 235 85 285 89
rect 640 85 656 89
rect 235 55 656 85
rect 690 55 706 89
rect 235 51 706 55
rect 854 55 870 89
rect 904 55 920 89
rect 966 86 982 120
rect 1016 86 1032 120
rect 966 70 1032 86
rect 1066 188 1132 202
rect 1066 154 1082 188
rect 1116 154 1132 188
rect 1066 120 1132 154
rect 1066 86 1082 120
rect 1116 86 1132 120
rect 1166 179 1232 236
rect 1278 234 1322 310
rect 1356 320 1422 356
rect 1356 286 1372 320
rect 1406 286 1422 320
rect 1356 270 1422 286
rect 1464 334 1498 390
rect 1537 418 1622 458
rect 1571 384 1622 418
rect 1537 368 1622 384
rect 1656 580 1728 596
rect 1656 546 1672 580
rect 1706 546 1728 580
rect 1656 499 1728 546
rect 1656 465 1672 499
rect 1706 465 1728 499
rect 1656 418 1728 465
rect 1656 384 1672 418
rect 1706 384 1728 418
rect 1656 368 1728 384
rect 1464 318 1660 334
rect 1464 284 1480 318
rect 1514 284 1548 318
rect 1582 284 1616 318
rect 1650 284 1660 318
rect 1464 268 1660 284
rect 1694 325 1728 368
rect 1762 580 1796 649
rect 1762 497 1796 546
rect 1762 414 1796 463
rect 1762 364 1796 380
rect 1836 580 1907 596
rect 1836 546 1852 580
rect 1886 546 1907 580
rect 1836 497 1907 546
rect 1836 463 1852 497
rect 1886 463 1907 497
rect 1836 414 1907 463
rect 1836 380 1852 414
rect 1886 380 1907 414
rect 1836 325 1907 380
rect 1942 580 1992 649
rect 1976 546 1992 580
rect 1942 497 1992 546
rect 1976 463 1992 497
rect 1942 414 1992 463
rect 1976 380 1992 414
rect 1942 364 1992 380
rect 1694 284 1907 325
rect 1464 236 1498 268
rect 1278 200 1294 234
rect 1328 200 1344 234
rect 1378 202 1498 236
rect 1694 234 1735 284
rect 1583 218 1633 234
rect 1166 145 1182 179
rect 1216 145 1232 179
rect 1378 166 1412 202
rect 1583 184 1599 218
rect 1583 168 1633 184
rect 1166 119 1232 145
rect 1266 132 1412 166
rect 1446 152 1633 168
rect 1066 85 1132 86
rect 1266 85 1300 132
rect 1480 118 1524 152
rect 1558 150 1633 152
rect 1558 118 1599 150
rect 1446 116 1599 118
rect 1446 98 1633 116
rect 854 17 920 55
rect 1066 51 1300 85
rect 1380 82 1633 98
rect 1669 218 1735 234
rect 1669 184 1685 218
rect 1719 184 1735 218
rect 1669 144 1735 184
rect 1669 110 1685 144
rect 1719 110 1735 144
rect 1669 94 1735 110
rect 1771 234 1805 250
rect 1771 144 1805 200
rect 1380 48 1396 82
rect 1430 48 1489 82
rect 1523 48 1583 82
rect 1617 48 1633 82
rect 1380 17 1633 48
rect 1771 17 1805 110
rect 1841 234 1907 284
rect 1841 200 1857 234
rect 1891 200 1907 234
rect 1841 144 1907 200
rect 1841 110 1857 144
rect 1891 110 1907 144
rect 1841 88 1907 110
rect 1943 234 1993 250
rect 1977 200 1993 234
rect 1943 144 1993 200
rect 1977 110 1993 144
rect 1943 17 1993 110
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 31 419 65 424
rect 31 390 39 419
rect 39 390 65 419
rect 319 390 353 424
rect 415 415 449 424
rect 415 390 421 415
rect 421 390 449 415
rect 991 410 1006 424
rect 1006 410 1025 424
rect 991 390 1025 410
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 19 424 77 430
rect 19 390 31 424
rect 65 421 77 424
rect 307 424 365 430
rect 307 421 319 424
rect 65 393 319 421
rect 65 390 77 393
rect 19 384 77 390
rect 307 390 319 393
rect 353 390 365 424
rect 307 384 365 390
rect 403 424 461 430
rect 403 390 415 424
rect 449 421 461 424
rect 979 424 1037 430
rect 979 421 991 424
rect 449 393 991 421
rect 449 390 461 393
rect 403 384 461 390
rect 979 390 991 393
rect 1025 390 1037 424
rect 979 384 1037 390
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
rlabel comment s 0 0 0 0 4 xnor3_4
flabel pwell s 0 0 2016 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 2016 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 2016 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 2016 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 1855 94 1889 128 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 1855 168 1889 202 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 1855 242 1889 276 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 1855 316 1889 350 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 1855 390 1889 424 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 1855 464 1889 498 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 1855 538 1889 572 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 1375 316 1409 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 2016 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 544552
string GDS_START 528686
<< end >>
