magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 335 496 401 596
rect 553 496 619 596
rect 335 462 619 496
rect 121 294 263 360
rect 505 424 619 462
rect 753 424 845 596
rect 505 390 845 424
rect 505 364 619 390
rect 25 51 96 134
rect 597 162 663 310
rect 697 270 777 356
rect 811 236 845 390
rect 697 202 845 236
rect 697 124 731 202
rect 344 70 731 124
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 23 394 89 570
rect 123 394 189 649
rect 223 428 289 570
rect 435 530 519 649
rect 223 394 471 428
rect 23 260 57 394
rect 437 310 471 394
rect 653 458 719 649
rect 337 260 403 310
rect 23 226 403 260
rect 437 244 549 310
rect 23 168 94 226
rect 437 192 471 244
rect 130 17 196 192
rect 230 158 471 192
rect 230 126 298 158
rect 765 17 831 168
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel locali s 25 51 96 134 6 A_N
port 1 nsew signal input
rlabel locali s 121 294 263 360 6 B_N
port 2 nsew signal input
rlabel locali s 597 162 663 310 6 C
port 3 nsew signal input
rlabel locali s 697 270 777 356 6 D
port 4 nsew signal input
rlabel locali s 811 236 845 390 6 Y
port 5 nsew signal output
rlabel locali s 753 424 845 596 6 Y
port 5 nsew signal output
rlabel locali s 697 202 845 236 6 Y
port 5 nsew signal output
rlabel locali s 697 124 731 202 6 Y
port 5 nsew signal output
rlabel locali s 553 496 619 596 6 Y
port 5 nsew signal output
rlabel locali s 505 424 619 462 6 Y
port 5 nsew signal output
rlabel locali s 505 390 845 424 6 Y
port 5 nsew signal output
rlabel locali s 505 364 619 390 6 Y
port 5 nsew signal output
rlabel locali s 344 70 731 124 6 Y
port 5 nsew signal output
rlabel locali s 335 496 401 596 6 Y
port 5 nsew signal output
rlabel locali s 335 462 619 496 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -49 864 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 864 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1484540
string GDS_START 1477012
<< end >>
