magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1564 561
rect 19 383 85 527
rect 119 349 153 493
rect 187 383 253 527
rect 287 349 321 493
rect 355 383 425 527
rect 30 315 321 349
rect 30 161 64 315
rect 715 383 781 527
rect 883 383 949 527
rect 1069 383 1207 527
rect 1323 383 1389 527
rect 427 215 629 256
rect 679 215 813 259
rect 855 215 995 257
rect 1031 215 1237 259
rect 1299 215 1501 259
rect 30 127 321 161
rect 19 17 85 93
rect 119 51 153 127
rect 187 17 253 93
rect 287 51 321 127
rect 355 17 425 93
rect 527 17 593 93
rect 1323 17 1389 93
rect 0 -17 1564 17
<< obsli1 >>
rect 475 459 681 493
rect 475 359 509 459
rect 543 391 609 425
rect 559 325 593 391
rect 355 291 593 325
rect 647 341 681 459
rect 815 341 849 493
rect 987 341 1021 493
rect 1255 341 1289 493
rect 1423 341 1457 493
rect 647 307 1474 341
rect 355 249 389 291
rect 98 215 389 249
rect 355 163 389 215
rect 355 129 781 163
rect 815 129 1033 163
rect 1071 129 1457 163
rect 459 51 493 129
rect 815 93 849 129
rect 631 59 849 93
rect 883 59 1221 93
rect 1423 51 1457 129
<< metal1 >>
rect 0 496 1564 592
rect 0 -48 1564 48
<< labels >>
rlabel locali s 679 215 813 259 6 A1
port 1 nsew signal input
rlabel locali s 855 215 995 257 6 A2
port 2 nsew signal input
rlabel locali s 1031 215 1237 259 6 A3
port 3 nsew signal input
rlabel locali s 1299 215 1501 259 6 A4
port 4 nsew signal input
rlabel locali s 427 215 629 256 6 B1
port 5 nsew signal input
rlabel locali s 287 349 321 493 6 X
port 6 nsew signal output
rlabel locali s 287 51 321 127 6 X
port 6 nsew signal output
rlabel locali s 119 349 153 493 6 X
port 6 nsew signal output
rlabel locali s 119 51 153 127 6 X
port 6 nsew signal output
rlabel locali s 30 315 321 349 6 X
port 6 nsew signal output
rlabel locali s 30 161 64 315 6 X
port 6 nsew signal output
rlabel locali s 30 127 321 161 6 X
port 6 nsew signal output
rlabel locali s 1323 17 1389 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 527 17 593 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 355 17 425 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 187 17 253 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 19 17 85 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 1564 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1564 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1323 383 1389 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1069 383 1207 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 883 383 949 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 715 383 781 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 355 383 425 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 187 383 253 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 19 383 85 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 1564 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 1564 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1564 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3703642
string GDS_START 3691176
<< end >>
