magic
tech sky130A
magscale 1 2
timestamp 1599588218
<< nwell >>
rect -38 332 2150 704
<< pwell >>
rect 0 0 2112 49
<< scpmos >>
rect 81 368 117 592
rect 171 368 207 592
rect 261 368 297 592
rect 351 368 387 592
rect 583 368 619 592
rect 673 368 709 592
rect 763 368 799 592
rect 853 368 889 592
rect 943 368 979 592
rect 1033 368 1069 592
rect 1123 368 1159 592
rect 1259 368 1295 592
rect 1349 368 1385 592
rect 1439 368 1475 592
rect 1529 368 1565 592
rect 1619 368 1655 592
rect 1709 368 1745 592
rect 1799 368 1835 592
rect 1889 368 1925 592
rect 1979 368 2015 592
<< nmoslvt >>
rect 110 74 140 222
rect 196 74 226 222
rect 282 74 312 222
rect 368 74 398 222
rect 587 74 617 222
rect 673 74 703 222
rect 759 74 789 222
rect 845 74 875 222
rect 931 74 961 222
rect 1017 74 1047 222
rect 1103 74 1133 222
rect 1189 74 1219 222
rect 1379 74 1409 222
rect 1465 74 1495 222
rect 1551 74 1581 222
rect 1637 74 1667 222
rect 1723 74 1753 222
rect 1809 74 1839 222
rect 1895 74 1925 222
rect 1981 74 2011 222
<< ndiff >>
rect 57 210 110 222
rect 57 176 65 210
rect 99 176 110 210
rect 57 120 110 176
rect 57 86 65 120
rect 99 86 110 120
rect 57 74 110 86
rect 140 152 196 222
rect 140 118 151 152
rect 185 118 196 152
rect 140 74 196 118
rect 226 210 282 222
rect 226 176 237 210
rect 271 176 282 210
rect 226 120 282 176
rect 226 86 237 120
rect 271 86 282 120
rect 226 74 282 86
rect 312 152 368 222
rect 312 118 323 152
rect 357 118 368 152
rect 312 74 368 118
rect 398 210 451 222
rect 398 176 409 210
rect 443 176 451 210
rect 398 120 451 176
rect 398 86 409 120
rect 443 86 451 120
rect 398 74 451 86
rect 534 144 587 222
rect 534 110 542 144
rect 576 110 587 144
rect 534 74 587 110
rect 617 116 673 222
rect 617 82 628 116
rect 662 82 673 116
rect 617 74 673 82
rect 703 144 759 222
rect 703 110 714 144
rect 748 110 759 144
rect 703 74 759 110
rect 789 116 845 222
rect 789 82 800 116
rect 834 82 845 116
rect 789 74 845 82
rect 875 184 931 222
rect 875 150 886 184
rect 920 150 931 184
rect 875 116 931 150
rect 875 82 886 116
rect 920 82 931 116
rect 875 74 931 82
rect 961 178 1017 222
rect 961 144 972 178
rect 1006 144 1017 178
rect 961 74 1017 144
rect 1047 184 1103 222
rect 1047 150 1058 184
rect 1092 150 1103 184
rect 1047 116 1103 150
rect 1047 82 1058 116
rect 1092 82 1103 116
rect 1047 74 1103 82
rect 1133 178 1189 222
rect 1133 144 1144 178
rect 1178 144 1189 178
rect 1133 74 1189 144
rect 1219 120 1272 222
rect 1219 86 1230 120
rect 1264 86 1272 120
rect 1219 74 1272 86
rect 1326 120 1379 222
rect 1326 86 1334 120
rect 1368 86 1379 120
rect 1326 74 1379 86
rect 1409 207 1465 222
rect 1409 173 1420 207
rect 1454 173 1465 207
rect 1409 74 1465 173
rect 1495 120 1551 222
rect 1495 86 1506 120
rect 1540 86 1551 120
rect 1495 74 1551 86
rect 1581 207 1637 222
rect 1581 173 1592 207
rect 1626 173 1637 207
rect 1581 74 1637 173
rect 1667 210 1723 222
rect 1667 176 1678 210
rect 1712 176 1723 210
rect 1667 120 1723 176
rect 1667 86 1678 120
rect 1712 86 1723 120
rect 1667 74 1723 86
rect 1753 152 1809 222
rect 1753 118 1764 152
rect 1798 118 1809 152
rect 1753 74 1809 118
rect 1839 210 1895 222
rect 1839 176 1850 210
rect 1884 176 1895 210
rect 1839 120 1895 176
rect 1839 86 1850 120
rect 1884 86 1895 120
rect 1839 74 1895 86
rect 1925 152 1981 222
rect 1925 118 1936 152
rect 1970 118 1981 152
rect 1925 74 1981 118
rect 2011 210 2064 222
rect 2011 176 2022 210
rect 2056 176 2064 210
rect 2011 120 2064 176
rect 2011 86 2022 120
rect 2056 86 2064 120
rect 2011 74 2064 86
<< pdiff >>
rect 29 580 81 592
rect 29 546 37 580
rect 71 546 81 580
rect 29 497 81 546
rect 29 463 37 497
rect 71 463 81 497
rect 29 414 81 463
rect 29 380 37 414
rect 71 380 81 414
rect 29 368 81 380
rect 117 531 171 592
rect 117 497 127 531
rect 161 497 171 531
rect 117 424 171 497
rect 117 390 127 424
rect 161 390 171 424
rect 117 368 171 390
rect 207 580 261 592
rect 207 546 217 580
rect 251 546 261 580
rect 207 499 261 546
rect 207 465 217 499
rect 251 465 261 499
rect 207 368 261 465
rect 297 531 351 592
rect 297 497 307 531
rect 341 497 351 531
rect 297 424 351 497
rect 297 390 307 424
rect 341 390 351 424
rect 297 368 351 390
rect 387 580 439 592
rect 387 546 397 580
rect 431 546 439 580
rect 387 499 439 546
rect 387 465 397 499
rect 431 465 439 499
rect 387 368 439 465
rect 531 580 583 592
rect 531 546 539 580
rect 573 546 583 580
rect 531 497 583 546
rect 531 463 539 497
rect 573 463 583 497
rect 531 368 583 463
rect 619 578 673 592
rect 619 544 629 578
rect 663 544 673 578
rect 619 368 673 544
rect 709 580 763 592
rect 709 546 719 580
rect 753 546 763 580
rect 709 497 763 546
rect 709 463 719 497
rect 753 463 763 497
rect 709 368 763 463
rect 799 578 853 592
rect 799 544 809 578
rect 843 544 853 578
rect 799 368 853 544
rect 889 580 943 592
rect 889 546 899 580
rect 933 546 943 580
rect 889 497 943 546
rect 889 463 899 497
rect 933 463 943 497
rect 889 368 943 463
rect 979 578 1033 592
rect 979 544 989 578
rect 1023 544 1033 578
rect 979 368 1033 544
rect 1069 580 1123 592
rect 1069 546 1079 580
rect 1113 546 1123 580
rect 1069 497 1123 546
rect 1069 463 1079 497
rect 1113 463 1123 497
rect 1069 368 1123 463
rect 1159 578 1259 592
rect 1159 544 1192 578
rect 1226 544 1259 578
rect 1159 368 1259 544
rect 1295 580 1349 592
rect 1295 546 1305 580
rect 1339 546 1349 580
rect 1295 508 1349 546
rect 1295 474 1305 508
rect 1339 474 1349 508
rect 1295 368 1349 474
rect 1385 541 1439 592
rect 1385 507 1395 541
rect 1429 507 1439 541
rect 1385 424 1439 507
rect 1385 390 1395 424
rect 1429 390 1439 424
rect 1385 368 1439 390
rect 1475 580 1529 592
rect 1475 546 1485 580
rect 1519 546 1529 580
rect 1475 508 1529 546
rect 1475 474 1485 508
rect 1519 474 1529 508
rect 1475 368 1529 474
rect 1565 541 1619 592
rect 1565 507 1575 541
rect 1609 507 1619 541
rect 1565 424 1619 507
rect 1565 390 1575 424
rect 1609 390 1619 424
rect 1565 368 1619 390
rect 1655 580 1709 592
rect 1655 546 1665 580
rect 1699 546 1709 580
rect 1655 508 1709 546
rect 1655 474 1665 508
rect 1699 474 1709 508
rect 1655 368 1709 474
rect 1745 541 1799 592
rect 1745 507 1755 541
rect 1789 507 1799 541
rect 1745 424 1799 507
rect 1745 390 1755 424
rect 1789 390 1799 424
rect 1745 368 1799 390
rect 1835 580 1889 592
rect 1835 546 1845 580
rect 1879 546 1889 580
rect 1835 508 1889 546
rect 1835 474 1845 508
rect 1879 474 1889 508
rect 1835 368 1889 474
rect 1925 541 1979 592
rect 1925 507 1935 541
rect 1969 507 1979 541
rect 1925 424 1979 507
rect 1925 390 1935 424
rect 1969 390 1979 424
rect 1925 368 1979 390
rect 2015 580 2067 592
rect 2015 546 2025 580
rect 2059 546 2067 580
rect 2015 497 2067 546
rect 2015 463 2025 497
rect 2059 463 2067 497
rect 2015 414 2067 463
rect 2015 380 2025 414
rect 2059 380 2067 414
rect 2015 368 2067 380
<< ndiffc >>
rect 65 176 99 210
rect 65 86 99 120
rect 151 118 185 152
rect 237 176 271 210
rect 237 86 271 120
rect 323 118 357 152
rect 409 176 443 210
rect 409 86 443 120
rect 542 110 576 144
rect 628 82 662 116
rect 714 110 748 144
rect 800 82 834 116
rect 886 150 920 184
rect 886 82 920 116
rect 972 144 1006 178
rect 1058 150 1092 184
rect 1058 82 1092 116
rect 1144 144 1178 178
rect 1230 86 1264 120
rect 1334 86 1368 120
rect 1420 173 1454 207
rect 1506 86 1540 120
rect 1592 173 1626 207
rect 1678 176 1712 210
rect 1678 86 1712 120
rect 1764 118 1798 152
rect 1850 176 1884 210
rect 1850 86 1884 120
rect 1936 118 1970 152
rect 2022 176 2056 210
rect 2022 86 2056 120
<< pdiffc >>
rect 37 546 71 580
rect 37 463 71 497
rect 37 380 71 414
rect 127 497 161 531
rect 127 390 161 424
rect 217 546 251 580
rect 217 465 251 499
rect 307 497 341 531
rect 307 390 341 424
rect 397 546 431 580
rect 397 465 431 499
rect 539 546 573 580
rect 539 463 573 497
rect 629 544 663 578
rect 719 546 753 580
rect 719 463 753 497
rect 809 544 843 578
rect 899 546 933 580
rect 899 463 933 497
rect 989 544 1023 578
rect 1079 546 1113 580
rect 1079 463 1113 497
rect 1192 544 1226 578
rect 1305 546 1339 580
rect 1305 474 1339 508
rect 1395 507 1429 541
rect 1395 390 1429 424
rect 1485 546 1519 580
rect 1485 474 1519 508
rect 1575 507 1609 541
rect 1575 390 1609 424
rect 1665 546 1699 580
rect 1665 474 1699 508
rect 1755 507 1789 541
rect 1755 390 1789 424
rect 1845 546 1879 580
rect 1845 474 1879 508
rect 1935 507 1969 541
rect 1935 390 1969 424
rect 2025 546 2059 580
rect 2025 463 2059 497
rect 2025 380 2059 414
<< poly >>
rect 81 592 117 618
rect 171 592 207 618
rect 261 592 297 618
rect 351 592 387 618
rect 583 592 619 618
rect 673 592 709 618
rect 763 592 799 618
rect 853 592 889 618
rect 943 592 979 618
rect 1033 592 1069 618
rect 1123 592 1159 618
rect 1259 592 1295 618
rect 1349 592 1385 618
rect 1439 592 1475 618
rect 1529 592 1565 618
rect 1619 592 1655 618
rect 1709 592 1745 618
rect 1799 592 1835 618
rect 1889 592 1925 618
rect 1979 592 2015 618
rect 81 336 117 368
rect 171 336 207 368
rect 261 336 297 368
rect 351 336 387 368
rect 81 320 387 336
rect 81 286 121 320
rect 155 286 189 320
rect 223 286 257 320
rect 291 286 325 320
rect 359 294 387 320
rect 583 336 619 368
rect 673 336 709 368
rect 763 336 799 368
rect 853 336 889 368
rect 943 336 979 368
rect 1033 336 1069 368
rect 1123 342 1159 368
rect 1259 342 1295 368
rect 1123 336 1295 342
rect 583 320 883 336
rect 359 286 398 294
rect 81 264 398 286
rect 583 286 599 320
rect 633 286 667 320
rect 701 286 735 320
rect 769 286 803 320
rect 837 286 883 320
rect 583 270 883 286
rect 931 320 1295 336
rect 931 286 947 320
rect 981 286 1015 320
rect 1049 286 1083 320
rect 1117 286 1173 320
rect 1207 286 1295 320
rect 110 222 140 264
rect 196 222 226 264
rect 282 222 312 264
rect 368 222 398 264
rect 587 222 617 270
rect 673 222 703 270
rect 759 222 789 270
rect 845 222 875 270
rect 931 264 1295 286
rect 1349 336 1385 368
rect 1439 336 1475 368
rect 1529 336 1565 368
rect 1619 336 1655 368
rect 1349 320 1655 336
rect 1349 286 1365 320
rect 1399 286 1433 320
rect 1467 286 1501 320
rect 1535 286 1569 320
rect 1603 300 1655 320
rect 1709 336 1745 368
rect 1799 336 1835 368
rect 1889 336 1925 368
rect 1979 336 2015 368
rect 1709 320 2011 336
rect 1603 286 1667 300
rect 1349 270 1667 286
rect 1709 286 1725 320
rect 1759 286 1793 320
rect 1827 286 1861 320
rect 1895 286 1929 320
rect 1963 286 2011 320
rect 1709 270 2011 286
rect 931 222 961 264
rect 1017 222 1047 264
rect 1103 222 1133 264
rect 1189 222 1219 264
rect 1379 222 1409 270
rect 1465 222 1495 270
rect 1551 222 1581 270
rect 1637 222 1667 270
rect 1723 222 1753 270
rect 1809 222 1839 270
rect 1895 222 1925 270
rect 1981 222 2011 270
rect 110 48 140 74
rect 196 48 226 74
rect 282 48 312 74
rect 368 48 398 74
rect 587 48 617 74
rect 673 48 703 74
rect 759 48 789 74
rect 845 48 875 74
rect 931 48 961 74
rect 1017 48 1047 74
rect 1103 48 1133 74
rect 1189 48 1219 74
rect 1379 48 1409 74
rect 1465 48 1495 74
rect 1551 48 1581 74
rect 1637 48 1667 74
rect 1723 48 1753 74
rect 1809 48 1839 74
rect 1895 48 1925 74
rect 1981 48 2011 74
<< polycont >>
rect 121 286 155 320
rect 189 286 223 320
rect 257 286 291 320
rect 325 286 359 320
rect 599 286 633 320
rect 667 286 701 320
rect 735 286 769 320
rect 803 286 837 320
rect 947 286 981 320
rect 1015 286 1049 320
rect 1083 286 1117 320
rect 1173 286 1207 320
rect 1365 286 1399 320
rect 1433 286 1467 320
rect 1501 286 1535 320
rect 1569 286 1603 320
rect 1725 286 1759 320
rect 1793 286 1827 320
rect 1861 286 1895 320
rect 1929 286 1963 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 21 581 447 615
rect 21 580 71 581
rect 21 546 37 580
rect 201 580 267 581
rect 21 497 71 546
rect 21 463 37 497
rect 21 414 71 463
rect 21 380 37 414
rect 111 531 167 547
rect 111 497 127 531
rect 161 497 167 531
rect 111 424 167 497
rect 201 546 217 580
rect 251 546 267 580
rect 381 580 447 581
rect 201 499 267 546
rect 201 465 217 499
rect 251 465 267 499
rect 201 458 267 465
rect 301 531 347 547
rect 301 497 307 531
rect 341 497 347 531
rect 301 424 347 497
rect 381 546 397 580
rect 431 546 447 580
rect 381 499 447 546
rect 381 465 397 499
rect 431 465 447 499
rect 381 458 447 465
rect 523 580 589 596
rect 523 546 539 580
rect 573 546 589 580
rect 523 497 589 546
rect 629 578 663 649
rect 629 526 663 544
rect 703 580 769 596
rect 703 546 719 580
rect 753 546 769 580
rect 523 463 539 497
rect 573 492 589 497
rect 703 497 769 546
rect 809 578 843 649
rect 809 526 843 544
rect 883 580 949 596
rect 883 546 899 580
rect 933 546 949 580
rect 703 492 719 497
rect 573 463 719 492
rect 753 492 769 497
rect 883 497 949 546
rect 989 578 1023 649
rect 989 526 1023 544
rect 1063 580 1129 596
rect 1063 546 1079 580
rect 1113 546 1129 580
rect 883 492 899 497
rect 753 463 899 492
rect 933 492 949 497
rect 1063 497 1129 546
rect 1163 578 1255 649
rect 1163 544 1192 578
rect 1226 544 1255 578
rect 1163 526 1255 544
rect 1289 581 2075 615
rect 1289 580 1345 581
rect 1289 546 1305 580
rect 1339 546 1345 580
rect 1479 580 1525 581
rect 1063 492 1079 497
rect 933 463 1079 492
rect 1113 492 1129 497
rect 1289 508 1345 546
rect 1289 492 1305 508
rect 1113 474 1305 492
rect 1339 474 1345 508
rect 1113 463 1345 474
rect 523 458 1345 463
rect 1379 541 1445 547
rect 1379 507 1395 541
rect 1429 507 1445 541
rect 1379 424 1445 507
rect 1479 546 1485 580
rect 1519 546 1525 580
rect 1659 580 1705 581
rect 1479 508 1525 546
rect 1479 474 1485 508
rect 1519 474 1525 508
rect 1479 458 1525 474
rect 1559 541 1625 547
rect 1559 507 1575 541
rect 1609 507 1625 541
rect 1559 424 1625 507
rect 1659 546 1665 580
rect 1699 546 1705 580
rect 1839 580 1885 581
rect 1659 508 1705 546
rect 1659 474 1665 508
rect 1699 474 1705 508
rect 1659 458 1705 474
rect 1739 541 1805 547
rect 1739 507 1755 541
rect 1789 507 1805 541
rect 1739 424 1805 507
rect 1839 546 1845 580
rect 1879 546 1885 580
rect 2025 580 2075 581
rect 1839 508 1885 546
rect 1839 474 1845 508
rect 1879 474 1885 508
rect 1839 458 1885 474
rect 1919 541 1985 547
rect 1919 507 1935 541
rect 1969 507 1985 541
rect 1919 424 1985 507
rect 111 390 127 424
rect 161 390 307 424
rect 341 390 1395 424
rect 1429 390 1575 424
rect 1609 390 1755 424
rect 1789 390 1935 424
rect 1969 390 1985 424
rect 2059 546 2075 580
rect 2025 497 2075 546
rect 2059 463 2075 497
rect 2025 414 2075 463
rect 21 236 71 380
rect 2059 380 2075 414
rect 2025 364 2075 380
rect 105 320 375 356
rect 105 286 121 320
rect 155 286 189 320
rect 223 286 257 320
rect 291 286 325 320
rect 359 286 375 320
rect 409 320 853 356
rect 409 286 599 320
rect 633 286 667 320
rect 701 286 735 320
rect 769 286 803 320
rect 837 286 853 320
rect 889 320 1223 356
rect 889 286 947 320
rect 981 286 1015 320
rect 1049 286 1083 320
rect 1117 286 1173 320
rect 1207 286 1223 320
rect 1273 320 1619 356
rect 1273 286 1365 320
rect 1399 286 1433 320
rect 1467 286 1501 320
rect 1535 286 1569 320
rect 1603 286 1619 320
rect 105 270 375 286
rect 1346 270 1619 286
rect 1657 320 1991 356
rect 1657 286 1725 320
rect 1759 286 1793 320
rect 1827 286 1861 320
rect 1895 286 1929 320
rect 1963 286 1991 320
rect 1657 270 1991 286
rect 409 236 1306 252
rect 21 218 1642 236
rect 21 210 459 218
rect 21 176 65 210
rect 99 202 237 210
rect 21 120 99 176
rect 271 202 409 210
rect 21 86 65 120
rect 21 70 99 86
rect 135 152 201 168
rect 135 118 151 152
rect 185 118 201 152
rect 135 17 201 118
rect 237 120 271 176
rect 443 176 459 210
rect 237 70 271 86
rect 307 152 373 168
rect 307 118 323 152
rect 357 118 373 152
rect 307 17 373 118
rect 409 120 459 176
rect 443 86 459 120
rect 409 70 459 86
rect 526 150 886 184
rect 920 150 936 184
rect 526 144 576 150
rect 526 110 542 144
rect 714 144 748 150
rect 526 70 576 110
rect 612 82 628 116
rect 662 82 678 116
rect 612 17 678 82
rect 886 116 936 150
rect 970 178 1008 218
rect 970 144 972 178
rect 1006 144 1008 178
rect 970 128 1008 144
rect 1042 150 1058 184
rect 1092 150 1108 184
rect 714 70 748 110
rect 784 82 800 116
rect 834 82 850 116
rect 784 17 850 82
rect 920 94 936 116
rect 1042 116 1108 150
rect 1142 178 1180 218
rect 1142 144 1144 178
rect 1178 144 1180 178
rect 1272 207 1642 218
rect 1272 173 1420 207
rect 1454 173 1592 207
rect 1626 173 1642 207
rect 1272 170 1642 173
rect 1583 154 1642 170
rect 1678 210 2072 236
rect 1712 202 1850 210
rect 1142 128 1180 144
rect 1042 94 1058 116
rect 920 82 1058 94
rect 1092 94 1108 116
rect 1214 120 1280 136
rect 1214 94 1230 120
rect 1092 86 1230 94
rect 1264 86 1280 120
rect 1092 82 1280 86
rect 886 60 1280 82
rect 1318 120 1384 136
rect 1490 120 1549 136
rect 1678 120 1712 176
rect 1884 202 2022 210
rect 1318 86 1334 120
rect 1368 86 1506 120
rect 1540 86 1678 120
rect 1318 70 1712 86
rect 1748 152 1814 168
rect 1748 118 1764 152
rect 1798 118 1814 152
rect 1748 17 1814 118
rect 1850 120 1884 176
rect 2056 176 2072 210
rect 1850 70 1884 86
rect 1920 152 1986 168
rect 1920 118 1936 152
rect 1970 118 1986 152
rect 1920 17 1986 118
rect 2022 120 2072 176
rect 2056 86 2072 120
rect 2022 70 2072 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
<< metal1 >>
rect 0 683 2112 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 0 617 2112 649
rect 0 17 2112 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
rect 0 -49 2112 -17
<< labels >>
flabel pwell s 0 0 2112 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nwell s 0 617 2112 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
rlabel comment s 0 0 0 0 4 a221oi_4
flabel metal1 s 0 617 2112 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 2112 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 31 94 65 128 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 31 168 65 202 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 31 390 65 424 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 31 464 65 498 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 31 538 65 572 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 C1
port 5 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 C1
port 5 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 C1
port 5 nsew
flabel corelocali s 1663 316 1697 350 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 1759 316 1793 350 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 1855 316 1889 350 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 1951 316 1985 350 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 1279 316 1313 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 1375 316 1409 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 1471 316 1505 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 1567 316 1601 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 1183 316 1217 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 2112 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3470398
string GDS_START 3453126
<< end >>
