magic
tech sky130A
magscale 1 2
timestamp 1604502705
<< nwell >>
rect -38 332 1190 704
<< pwell >>
rect 0 0 1152 49
<< scnmos >>
rect 87 74 117 222
rect 177 74 207 222
rect 263 74 293 222
rect 357 74 387 222
rect 465 74 495 222
rect 551 74 581 222
rect 645 74 675 222
rect 809 74 839 222
rect 909 74 939 222
rect 995 74 1025 222
<< pmoshvt >>
rect 84 368 114 592
rect 174 368 204 592
rect 264 368 294 592
rect 360 368 390 592
rect 450 368 480 592
rect 540 368 570 592
rect 734 368 764 592
rect 824 368 854 592
rect 914 368 944 592
rect 1004 368 1034 592
<< ndiff >>
rect 34 210 87 222
rect 34 176 42 210
rect 76 176 87 210
rect 34 120 87 176
rect 34 86 42 120
rect 76 86 87 120
rect 34 74 87 86
rect 117 152 177 222
rect 117 118 130 152
rect 164 118 177 152
rect 117 74 177 118
rect 207 210 263 222
rect 207 176 218 210
rect 252 176 263 210
rect 207 120 263 176
rect 207 86 218 120
rect 252 86 263 120
rect 207 74 263 86
rect 293 184 357 222
rect 293 150 304 184
rect 338 150 357 184
rect 293 116 357 150
rect 293 82 304 116
rect 338 82 357 116
rect 293 74 357 82
rect 387 116 465 222
rect 387 82 405 116
rect 439 82 465 116
rect 387 74 465 82
rect 495 184 551 222
rect 495 150 506 184
rect 540 150 551 184
rect 495 116 551 150
rect 495 82 506 116
rect 540 82 551 116
rect 495 74 551 82
rect 581 210 645 222
rect 581 176 592 210
rect 626 176 645 210
rect 581 120 645 176
rect 581 86 592 120
rect 626 86 645 120
rect 581 74 645 86
rect 675 184 809 222
rect 675 150 686 184
rect 720 150 764 184
rect 798 150 809 184
rect 675 116 809 150
rect 675 82 686 116
rect 720 82 764 116
rect 798 82 809 116
rect 675 74 809 82
rect 839 116 909 222
rect 839 82 856 116
rect 890 82 909 116
rect 839 74 909 82
rect 939 184 995 222
rect 939 150 950 184
rect 984 150 995 184
rect 939 116 995 150
rect 939 82 950 116
rect 984 82 995 116
rect 939 74 995 82
rect 1025 210 1078 222
rect 1025 176 1036 210
rect 1070 176 1078 210
rect 1025 120 1078 176
rect 1025 86 1036 120
rect 1070 86 1078 120
rect 1025 74 1078 86
<< pdiff >>
rect 29 580 84 592
rect 29 546 37 580
rect 71 546 84 580
rect 29 508 84 546
rect 29 474 37 508
rect 71 474 84 508
rect 29 368 84 474
rect 114 540 174 592
rect 114 506 127 540
rect 161 506 174 540
rect 114 429 174 506
rect 114 395 127 429
rect 161 395 174 429
rect 114 368 174 395
rect 204 580 264 592
rect 204 546 217 580
rect 251 546 264 580
rect 204 500 264 546
rect 204 466 217 500
rect 251 466 264 500
rect 204 420 264 466
rect 204 386 217 420
rect 251 386 264 420
rect 204 368 264 386
rect 294 519 360 592
rect 294 485 310 519
rect 344 485 360 519
rect 294 368 360 485
rect 390 578 450 592
rect 390 544 403 578
rect 437 544 450 578
rect 390 368 450 544
rect 480 492 540 592
rect 480 458 493 492
rect 527 458 540 492
rect 480 368 540 458
rect 570 578 625 592
rect 570 544 583 578
rect 617 544 625 578
rect 570 368 625 544
rect 679 578 734 592
rect 679 544 687 578
rect 721 544 734 578
rect 679 368 734 544
rect 764 580 824 592
rect 764 546 777 580
rect 811 546 824 580
rect 764 495 824 546
rect 764 461 777 495
rect 811 461 824 495
rect 764 368 824 461
rect 854 578 914 592
rect 854 544 867 578
rect 901 544 914 578
rect 854 368 914 544
rect 944 580 1004 592
rect 944 546 957 580
rect 991 546 1004 580
rect 944 495 1004 546
rect 944 461 957 495
rect 991 461 1004 495
rect 944 368 1004 461
rect 1034 580 1089 592
rect 1034 546 1047 580
rect 1081 546 1089 580
rect 1034 510 1089 546
rect 1034 476 1047 510
rect 1081 476 1089 510
rect 1034 440 1089 476
rect 1034 406 1047 440
rect 1081 406 1089 440
rect 1034 368 1089 406
<< ndiffc >>
rect 42 176 76 210
rect 42 86 76 120
rect 130 118 164 152
rect 218 176 252 210
rect 218 86 252 120
rect 304 150 338 184
rect 304 82 338 116
rect 405 82 439 116
rect 506 150 540 184
rect 506 82 540 116
rect 592 176 626 210
rect 592 86 626 120
rect 686 150 720 184
rect 764 150 798 184
rect 686 82 720 116
rect 764 82 798 116
rect 856 82 890 116
rect 950 150 984 184
rect 950 82 984 116
rect 1036 176 1070 210
rect 1036 86 1070 120
<< pdiffc >>
rect 37 546 71 580
rect 37 474 71 508
rect 127 506 161 540
rect 127 395 161 429
rect 217 546 251 580
rect 217 466 251 500
rect 217 386 251 420
rect 310 485 344 519
rect 403 544 437 578
rect 493 458 527 492
rect 583 544 617 578
rect 687 544 721 578
rect 777 546 811 580
rect 777 461 811 495
rect 867 544 901 578
rect 957 546 991 580
rect 957 461 991 495
rect 1047 546 1081 580
rect 1047 476 1081 510
rect 1047 406 1081 440
<< poly >>
rect 84 592 114 618
rect 174 592 204 618
rect 264 592 294 618
rect 360 592 390 618
rect 450 592 480 618
rect 540 592 570 618
rect 734 592 764 618
rect 824 592 854 618
rect 914 592 944 618
rect 1004 592 1034 618
rect 84 353 114 368
rect 174 353 204 368
rect 264 353 294 368
rect 360 353 390 368
rect 450 353 480 368
rect 540 353 570 368
rect 734 353 764 368
rect 824 353 854 368
rect 914 353 944 368
rect 1004 353 1034 368
rect 81 336 117 353
rect 171 336 207 353
rect 261 336 297 353
rect 357 336 393 353
rect 447 336 483 353
rect 81 320 207 336
rect 81 286 133 320
rect 167 286 207 320
rect 81 270 207 286
rect 249 320 315 336
rect 249 286 265 320
rect 299 286 315 320
rect 249 270 315 286
rect 357 320 483 336
rect 357 286 405 320
rect 439 300 483 320
rect 537 336 573 353
rect 731 336 767 353
rect 821 336 857 353
rect 911 336 947 353
rect 1001 336 1037 353
rect 537 320 603 336
rect 439 286 495 300
rect 357 270 495 286
rect 537 286 553 320
rect 587 286 603 320
rect 537 270 603 286
rect 645 320 767 336
rect 645 286 697 320
rect 731 286 767 320
rect 645 270 767 286
rect 809 320 947 336
rect 809 286 825 320
rect 859 286 947 320
rect 809 270 947 286
rect 995 320 1061 336
rect 995 286 1011 320
rect 1045 286 1061 320
rect 995 270 1061 286
rect 87 222 117 270
rect 177 222 207 270
rect 263 222 293 270
rect 357 222 387 270
rect 465 222 495 270
rect 551 222 581 270
rect 645 222 675 270
rect 809 222 839 270
rect 909 222 939 270
rect 995 222 1025 270
rect 87 48 117 74
rect 177 48 207 74
rect 263 48 293 74
rect 357 48 387 74
rect 465 48 495 74
rect 551 48 581 74
rect 645 48 675 74
rect 809 48 839 74
rect 909 48 939 74
rect 995 48 1025 74
<< polycont >>
rect 133 286 167 320
rect 265 286 299 320
rect 405 286 439 320
rect 553 286 587 320
rect 697 286 731 320
rect 825 286 859 320
rect 1011 286 1045 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 21 596 453 615
rect 21 581 633 596
rect 21 580 71 581
rect 21 546 37 580
rect 217 580 251 581
rect 21 508 71 546
rect 21 474 37 508
rect 21 458 71 474
rect 111 540 177 547
rect 111 506 127 540
rect 161 506 177 540
rect 111 429 177 506
rect 111 424 127 429
rect 25 395 127 424
rect 161 395 177 429
rect 25 390 177 395
rect 403 578 633 581
rect 217 500 251 546
rect 217 420 251 466
rect 291 519 363 547
rect 437 544 583 578
rect 617 544 633 578
rect 403 526 633 544
rect 671 578 721 649
rect 671 544 687 578
rect 671 526 721 544
rect 761 580 827 596
rect 761 546 777 580
rect 811 546 827 580
rect 291 485 310 519
rect 344 492 363 519
rect 761 495 827 546
rect 867 578 901 649
rect 867 526 901 544
rect 941 580 1007 596
rect 941 546 957 580
rect 991 546 1007 580
rect 761 492 777 495
rect 344 485 493 492
rect 291 458 493 485
rect 527 461 777 492
rect 811 492 827 495
rect 941 495 1007 546
rect 941 492 957 495
rect 811 461 957 492
rect 991 461 1007 495
rect 527 458 1007 461
rect 1047 580 1097 649
rect 1081 546 1097 580
rect 1047 510 1097 546
rect 1081 476 1097 510
rect 1047 440 1097 476
rect 25 236 76 390
rect 217 370 251 386
rect 285 390 647 424
rect 117 320 183 356
rect 285 336 319 390
rect 117 286 133 320
rect 167 286 183 320
rect 249 320 319 336
rect 249 286 265 320
rect 299 286 319 320
rect 389 320 455 356
rect 389 286 405 320
rect 439 286 455 320
rect 505 320 647 390
rect 505 310 553 320
rect 537 286 553 310
rect 587 310 647 320
rect 681 390 1013 424
rect 1081 406 1097 440
rect 1047 390 1097 406
rect 681 320 747 390
rect 979 356 1013 390
rect 587 286 603 310
rect 681 286 697 320
rect 731 286 747 320
rect 793 320 935 356
rect 793 286 825 320
rect 859 286 935 320
rect 979 320 1127 356
rect 979 286 1011 320
rect 1045 286 1127 320
rect 117 270 183 286
rect 218 236 1086 252
rect 25 218 1086 236
rect 25 210 252 218
rect 25 176 42 210
rect 76 202 218 210
rect 25 120 76 176
rect 590 210 636 218
rect 25 86 42 120
rect 25 70 76 86
rect 112 152 182 168
rect 112 118 130 152
rect 164 118 182 152
rect 112 17 182 118
rect 218 120 252 176
rect 218 70 252 86
rect 288 150 304 184
rect 338 150 506 184
rect 540 150 556 184
rect 288 116 354 150
rect 490 116 556 150
rect 288 82 304 116
rect 338 82 354 116
rect 288 70 354 82
rect 388 82 405 116
rect 439 82 456 116
rect 388 17 456 82
rect 490 82 506 116
rect 540 82 556 116
rect 490 66 556 82
rect 590 176 592 210
rect 626 176 636 210
rect 1036 210 1086 218
rect 590 120 636 176
rect 590 86 592 120
rect 626 86 636 120
rect 590 70 636 86
rect 670 150 686 184
rect 720 150 764 184
rect 798 150 950 184
rect 984 150 1000 184
rect 670 116 806 150
rect 940 116 1000 150
rect 670 82 686 116
rect 720 82 764 116
rect 798 82 806 116
rect 670 66 806 82
rect 840 82 856 116
rect 890 82 906 116
rect 840 17 906 82
rect 940 82 950 116
rect 984 82 1000 116
rect 940 66 1000 82
rect 1070 176 1086 210
rect 1036 120 1086 176
rect 1070 86 1086 120
rect 1036 70 1086 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a221oi_2
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 C1
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 1152 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 4128748
string GDS_START 4118786
<< end >>
