magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 736 561
rect 105 387 171 527
rect 440 387 526 527
rect 562 415 600 493
rect 634 451 700 527
rect 562 381 708 415
rect 17 199 72 265
rect 176 199 248 265
rect 306 199 364 265
rect 398 199 465 265
rect 669 157 708 381
rect 544 123 708 157
rect 278 17 345 93
rect 463 17 510 105
rect 544 51 610 123
rect 644 17 710 89
rect 0 -17 736 17
<< obsli1 >>
rect 18 353 71 493
rect 205 353 339 493
rect 18 302 533 353
rect 106 165 142 302
rect 499 265 533 302
rect 499 199 635 265
rect 19 85 142 165
rect 176 127 430 165
rect 19 51 86 85
<< metal1 >>
rect 0 496 736 592
rect 0 -48 736 48
<< labels >>
rlabel locali s 398 199 465 265 6 A1
port 1 nsew signal input
rlabel locali s 306 199 364 265 6 A2
port 2 nsew signal input
rlabel locali s 176 199 248 265 6 B1
port 3 nsew signal input
rlabel locali s 17 199 72 265 6 C1
port 4 nsew signal input
rlabel locali s 669 157 708 381 6 X
port 5 nsew signal output
rlabel locali s 562 415 600 493 6 X
port 5 nsew signal output
rlabel locali s 562 381 708 415 6 X
port 5 nsew signal output
rlabel locali s 544 123 708 157 6 X
port 5 nsew signal output
rlabel locali s 544 51 610 123 6 X
port 5 nsew signal output
rlabel locali s 644 17 710 89 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 463 17 510 105 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 278 17 345 93 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 736 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 736 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 634 451 700 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 440 387 526 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 105 387 171 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 736 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 736 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1292368
string GDS_START 1286044
<< end >>
