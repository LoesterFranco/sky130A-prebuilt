magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 2024 561
rect 108 439 153 527
rect 20 199 66 323
rect 118 199 195 323
rect 440 299 474 527
rect 508 333 558 493
rect 592 367 642 527
rect 676 333 742 493
rect 776 367 810 527
rect 844 333 910 493
rect 944 367 978 527
rect 1012 333 1078 493
rect 1122 367 1308 527
rect 1348 333 1414 493
rect 1448 367 1482 527
rect 1516 333 1582 493
rect 1616 367 1650 527
rect 1684 333 1750 493
rect 1784 367 1818 527
rect 1852 333 1918 493
rect 508 289 1918 333
rect 1952 289 2007 527
rect 740 181 798 289
rect 1224 215 1582 255
rect 1684 215 2003 255
rect 103 17 169 93
rect 508 131 798 181
rect 1684 17 1750 97
rect 1852 17 1918 97
rect 0 -17 2024 17
<< obsli1 >>
rect 17 396 74 488
rect 187 430 359 493
rect 17 357 291 396
rect 229 161 291 357
rect 17 127 291 161
rect 325 261 359 430
rect 325 255 442 261
rect 325 221 396 255
rect 430 221 442 255
rect 325 215 442 221
rect 508 215 657 249
rect 17 51 69 127
rect 325 93 359 215
rect 832 221 856 255
rect 890 221 1078 255
rect 832 215 1078 221
rect 203 51 359 93
rect 440 97 474 181
rect 844 147 1230 181
rect 844 131 1078 147
rect 1196 97 1230 147
rect 1264 131 2007 181
rect 440 51 1162 97
rect 1196 51 1582 97
<< obsli1c >>
rect 396 221 430 255
rect 856 221 890 255
<< metal1 >>
rect 0 496 2024 592
rect 0 -48 2024 48
<< obsm1 >>
rect 384 255 442 261
rect 384 221 396 255
rect 430 252 442 255
rect 844 255 902 261
rect 844 252 856 255
rect 430 224 856 252
rect 430 221 442 224
rect 384 215 442 221
rect 844 221 856 224
rect 890 221 902 255
rect 844 215 902 221
<< labels >>
rlabel locali s 20 199 66 323 6 A_N
port 1 nsew signal input
rlabel locali s 118 199 195 323 6 B_N
port 2 nsew signal input
rlabel locali s 1224 215 1582 255 6 C
port 3 nsew signal input
rlabel locali s 1684 215 2003 255 6 D
port 4 nsew signal input
rlabel locali s 1852 333 1918 493 6 Y
port 5 nsew signal output
rlabel locali s 1684 333 1750 493 6 Y
port 5 nsew signal output
rlabel locali s 1516 333 1582 493 6 Y
port 5 nsew signal output
rlabel locali s 1348 333 1414 493 6 Y
port 5 nsew signal output
rlabel locali s 1012 333 1078 493 6 Y
port 5 nsew signal output
rlabel locali s 844 333 910 493 6 Y
port 5 nsew signal output
rlabel locali s 740 181 798 289 6 Y
port 5 nsew signal output
rlabel locali s 676 333 742 493 6 Y
port 5 nsew signal output
rlabel locali s 508 333 558 493 6 Y
port 5 nsew signal output
rlabel locali s 508 289 1918 333 6 Y
port 5 nsew signal output
rlabel locali s 508 131 798 181 6 Y
port 5 nsew signal output
rlabel locali s 1852 17 1918 97 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1684 17 1750 97 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 103 17 169 93 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 2024 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 2024 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1952 289 2007 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1784 367 1818 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1616 367 1650 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1448 367 1482 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1122 367 1308 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 944 367 978 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 776 367 810 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 592 367 642 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 440 299 474 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 108 439 153 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 2024 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 2024 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2024 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1927300
string GDS_START 1912312
<< end >>
