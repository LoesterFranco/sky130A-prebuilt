magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 79 93 109 177
rect 186 47 216 177
rect 295 47 325 177
rect 488 47 518 177
rect 593 47 623 177
rect 677 47 707 177
<< pmoshvt >>
rect 81 297 117 381
rect 188 297 224 497
rect 287 297 323 497
rect 480 297 516 497
rect 585 297 621 497
rect 668 297 704 497
<< ndiff >>
rect 27 149 79 177
rect 27 115 35 149
rect 69 115 79 149
rect 27 93 79 115
rect 109 149 186 177
rect 109 115 129 149
rect 163 115 186 149
rect 109 93 186 115
rect 134 47 186 93
rect 216 93 295 177
rect 216 59 226 93
rect 260 59 295 93
rect 216 47 295 59
rect 325 93 377 177
rect 325 59 335 93
rect 369 59 377 93
rect 325 47 377 59
rect 436 161 488 177
rect 436 127 444 161
rect 478 127 488 161
rect 436 93 488 127
rect 436 59 444 93
rect 478 59 488 93
rect 436 47 488 59
rect 518 133 593 177
rect 518 99 539 133
rect 573 99 593 133
rect 518 47 593 99
rect 623 95 677 177
rect 623 61 633 95
rect 667 61 677 95
rect 623 47 677 61
rect 707 163 769 177
rect 707 129 727 163
rect 761 129 769 163
rect 707 95 769 129
rect 707 61 727 95
rect 761 61 769 95
rect 707 47 769 61
<< pdiff >>
rect 134 475 188 497
rect 134 441 142 475
rect 176 441 188 475
rect 134 381 188 441
rect 27 349 81 381
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 297 188 381
rect 224 339 287 497
rect 224 305 236 339
rect 270 305 287 339
rect 224 297 287 305
rect 323 475 480 497
rect 323 441 335 475
rect 369 441 426 475
rect 460 441 480 475
rect 323 297 480 441
rect 516 477 585 497
rect 516 443 539 477
rect 573 443 585 477
rect 516 409 585 443
rect 516 375 539 409
rect 573 375 585 409
rect 516 341 585 375
rect 516 307 539 341
rect 573 307 585 341
rect 516 297 585 307
rect 621 297 668 497
rect 704 477 762 497
rect 704 443 716 477
rect 750 443 762 477
rect 704 409 762 443
rect 704 375 716 409
rect 750 375 762 409
rect 704 297 762 375
<< ndiffc >>
rect 35 115 69 149
rect 129 115 163 149
rect 226 59 260 93
rect 335 59 369 93
rect 444 127 478 161
rect 444 59 478 93
rect 539 99 573 133
rect 633 61 667 95
rect 727 129 761 163
rect 727 61 761 95
<< pdiffc >>
rect 142 441 176 475
rect 35 315 69 349
rect 236 305 270 339
rect 335 441 369 475
rect 426 441 460 475
rect 539 443 573 477
rect 539 375 573 409
rect 539 307 573 341
rect 716 443 750 477
rect 716 375 750 409
<< poly >>
rect 188 497 224 523
rect 287 497 323 523
rect 480 497 516 523
rect 585 497 621 523
rect 668 497 704 523
rect 81 381 117 407
rect 81 282 117 297
rect 188 282 224 297
rect 287 282 323 297
rect 480 282 516 297
rect 585 282 621 297
rect 668 282 704 297
rect 79 265 119 282
rect 186 265 226 282
rect 285 265 325 282
rect 478 265 518 282
rect 583 265 623 282
rect 79 249 139 265
rect 79 215 89 249
rect 123 215 139 249
rect 79 199 139 215
rect 186 249 325 265
rect 186 215 281 249
rect 315 215 325 249
rect 186 199 325 215
rect 373 249 518 265
rect 373 215 383 249
rect 417 215 518 249
rect 373 199 518 215
rect 560 249 623 265
rect 560 215 570 249
rect 604 215 623 249
rect 560 199 623 215
rect 666 265 706 282
rect 666 249 746 265
rect 666 215 686 249
rect 720 215 746 249
rect 666 199 746 215
rect 79 177 109 199
rect 186 177 216 199
rect 295 177 325 199
rect 488 177 518 199
rect 593 177 623 199
rect 677 177 707 199
rect 79 67 109 93
rect 186 21 216 47
rect 295 21 325 47
rect 488 21 518 47
rect 593 21 623 47
rect 677 21 707 47
<< polycont >>
rect 89 215 123 249
rect 281 215 315 249
rect 383 215 417 249
rect 570 215 604 249
rect 686 215 720 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 104 475 192 527
rect 104 441 142 475
rect 176 441 192 475
rect 304 475 476 527
rect 304 441 335 475
rect 369 441 426 475
rect 460 441 476 475
rect 520 477 585 493
rect 520 443 539 477
rect 573 443 585 477
rect 520 409 585 443
rect 520 407 539 409
rect 17 373 417 407
rect 17 349 79 373
rect 17 315 35 349
rect 69 315 79 349
rect 17 299 79 315
rect 17 165 51 299
rect 121 265 165 339
rect 85 249 165 265
rect 85 215 89 249
rect 123 215 165 249
rect 85 199 165 215
rect 199 305 236 339
rect 270 305 291 339
rect 199 299 291 305
rect 17 149 69 165
rect 17 115 35 149
rect 17 86 69 115
rect 129 149 165 165
rect 163 115 165 149
rect 129 17 165 115
rect 199 93 247 299
rect 281 249 315 265
rect 281 165 315 215
rect 383 249 417 373
rect 383 199 417 215
rect 451 375 539 407
rect 573 375 585 409
rect 690 477 766 527
rect 690 443 716 477
rect 750 443 766 477
rect 690 409 766 443
rect 690 375 716 409
rect 750 375 766 409
rect 451 341 585 375
rect 451 307 539 341
rect 573 307 585 341
rect 451 291 585 307
rect 451 165 494 291
rect 529 249 636 257
rect 529 215 570 249
rect 604 215 636 249
rect 670 249 779 325
rect 670 215 686 249
rect 720 215 779 249
rect 281 161 494 165
rect 281 131 444 161
rect 428 127 444 131
rect 478 127 494 161
rect 428 93 494 127
rect 199 59 226 93
rect 260 59 276 93
rect 312 59 335 93
rect 369 59 385 93
rect 312 17 385 59
rect 428 59 444 93
rect 478 59 494 93
rect 539 163 778 181
rect 539 147 727 163
rect 539 133 589 147
rect 573 99 589 133
rect 711 129 727 147
rect 761 129 778 163
rect 539 73 589 99
rect 633 95 667 111
rect 428 51 494 59
rect 633 17 667 61
rect 711 95 778 129
rect 711 61 727 95
rect 761 61 778 95
rect 711 54 778 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel corelocali s 131 221 165 255 0 FreeSans 400 180 0 0 B1_N
port 3 nsew
flabel corelocali s 733 221 767 255 0 FreeSans 400 0 0 0 A1
port 1 nsew
flabel corelocali s 206 85 240 119 0 FreeSans 400 180 0 0 X
port 8 nsew
flabel corelocali s 579 238 579 238 0 FreeSans 400 0 0 0 A2
port 2 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
rlabel comment s 0 0 0 0 4 o21ba_2
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1076574
string GDS_START 1070062
<< end >>
