magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 644 561
rect 17 359 156 527
rect 17 199 156 325
rect 190 199 252 493
rect 286 333 396 493
rect 430 367 496 527
rect 530 333 627 493
rect 286 299 627 333
rect 286 199 356 265
rect 17 153 114 199
rect 17 17 114 119
rect 216 17 282 97
rect 397 52 440 265
rect 489 119 532 299
rect 566 153 627 265
rect 489 51 627 119
rect 0 -17 644 17
<< obsli1 >>
rect 148 131 350 165
rect 148 51 182 131
rect 316 51 350 131
<< metal1 >>
rect 0 496 644 592
rect 0 -48 644 48
<< labels >>
rlabel locali s 17 199 156 325 6 A1
port 1 nsew signal input
rlabel locali s 17 153 114 199 6 A1
port 1 nsew signal input
rlabel locali s 190 199 252 493 6 A2
port 2 nsew signal input
rlabel locali s 286 199 356 265 6 A3
port 3 nsew signal input
rlabel locali s 397 52 440 265 6 B1
port 4 nsew signal input
rlabel locali s 566 153 627 265 6 C1
port 5 nsew signal input
rlabel locali s 530 333 627 493 6 Y
port 6 nsew signal output
rlabel locali s 489 119 532 299 6 Y
port 6 nsew signal output
rlabel locali s 489 51 627 119 6 Y
port 6 nsew signal output
rlabel locali s 286 333 396 493 6 Y
port 6 nsew signal output
rlabel locali s 286 299 627 333 6 Y
port 6 nsew signal output
rlabel locali s 216 17 282 97 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 17 17 114 119 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 644 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 644 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 430 367 496 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 17 359 156 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 644 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 644 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 775652
string GDS_START 768226
<< end >>
