magic
tech sky130A
magscale 1 2
timestamp 1604502705
<< nwell >>
rect -38 332 1766 704
rect 170 315 586 332
rect 170 294 338 315
<< pwell >>
rect 0 0 1728 49
<< scnmos >>
rect 115 98 145 226
rect 229 78 259 226
rect 323 78 353 226
rect 441 78 471 226
rect 527 78 557 226
rect 679 119 709 247
rect 779 119 809 247
rect 907 119 937 247
rect 993 119 1023 247
rect 1327 74 1357 202
rect 1417 74 1447 202
rect 1513 74 1543 202
rect 1605 74 1635 202
<< pmoshvt >>
rect 86 368 116 568
rect 196 368 226 592
rect 320 368 350 592
rect 444 368 474 592
rect 568 368 598 592
rect 692 391 722 591
rect 782 391 812 591
rect 906 391 936 591
rect 996 391 1026 591
rect 1330 392 1360 592
rect 1420 392 1450 592
rect 1512 392 1542 592
rect 1602 392 1632 592
<< ndiff >>
rect 589 235 679 247
rect 589 226 601 235
rect 58 214 115 226
rect 58 180 70 214
rect 104 180 115 214
rect 58 144 115 180
rect 58 110 70 144
rect 104 110 115 144
rect 58 98 115 110
rect 145 214 229 226
rect 145 180 170 214
rect 204 180 229 214
rect 145 144 229 180
rect 145 110 170 144
rect 204 110 229 144
rect 145 98 229 110
rect 179 78 229 98
rect 259 214 323 226
rect 259 180 278 214
rect 312 180 323 214
rect 259 124 323 180
rect 259 90 278 124
rect 312 90 323 124
rect 259 78 323 90
rect 353 214 441 226
rect 353 180 378 214
rect 412 180 441 214
rect 353 124 441 180
rect 353 90 378 124
rect 412 90 441 124
rect 353 78 441 90
rect 471 214 527 226
rect 471 180 482 214
rect 516 180 527 214
rect 471 124 527 180
rect 471 90 482 124
rect 516 90 527 124
rect 471 78 527 90
rect 557 201 601 226
rect 635 201 679 235
rect 557 124 679 201
rect 557 90 601 124
rect 635 119 679 124
rect 709 235 779 247
rect 709 201 720 235
rect 754 201 779 235
rect 709 165 779 201
rect 709 131 720 165
rect 754 131 779 165
rect 709 119 779 131
rect 809 165 907 247
rect 809 131 834 165
rect 868 131 907 165
rect 809 119 907 131
rect 937 167 993 247
rect 937 133 948 167
rect 982 133 993 167
rect 937 119 993 133
rect 1023 119 1111 247
rect 635 90 647 119
rect 1038 117 1111 119
rect 557 78 647 90
rect 1038 83 1057 117
rect 1091 83 1111 117
rect 1038 71 1111 83
rect 1171 120 1327 202
rect 1171 86 1183 120
rect 1217 86 1268 120
rect 1302 86 1327 120
rect 1171 74 1327 86
rect 1357 170 1417 202
rect 1357 136 1368 170
rect 1402 136 1417 170
rect 1357 74 1417 136
rect 1447 184 1513 202
rect 1447 150 1468 184
rect 1502 150 1513 184
rect 1447 116 1513 150
rect 1447 82 1468 116
rect 1502 82 1513 116
rect 1447 74 1513 82
rect 1543 179 1605 202
rect 1543 145 1554 179
rect 1588 145 1605 179
rect 1543 74 1605 145
rect 1635 190 1701 202
rect 1635 156 1654 190
rect 1688 156 1701 190
rect 1635 120 1701 156
rect 1635 86 1654 120
rect 1688 86 1701 120
rect 1635 74 1701 86
<< pdiff >>
rect 368 617 426 629
rect 368 592 380 617
rect 134 580 196 592
rect 134 568 147 580
rect 27 556 86 568
rect 27 522 39 556
rect 73 522 86 556
rect 27 440 86 522
rect 27 406 39 440
rect 73 406 86 440
rect 27 368 86 406
rect 116 546 147 568
rect 181 546 196 580
rect 116 368 196 546
rect 226 376 320 592
rect 226 368 256 376
rect 244 342 256 368
rect 290 368 320 376
rect 350 583 380 592
rect 414 592 426 617
rect 616 617 674 629
rect 616 592 628 617
rect 414 583 444 592
rect 350 368 444 583
rect 474 397 568 592
rect 474 368 504 397
rect 290 342 302 368
rect 492 363 504 368
rect 538 368 568 397
rect 598 583 628 592
rect 662 591 674 617
rect 830 605 888 617
rect 830 591 842 605
rect 662 583 692 591
rect 598 391 692 583
rect 722 579 782 591
rect 722 545 735 579
rect 769 545 782 579
rect 722 505 782 545
rect 722 471 735 505
rect 769 471 782 505
rect 722 391 782 471
rect 812 571 842 591
rect 876 591 888 605
rect 1044 605 1102 617
rect 1044 591 1056 605
rect 876 571 906 591
rect 812 391 906 571
rect 936 437 996 591
rect 936 403 949 437
rect 983 403 996 437
rect 936 391 996 403
rect 1026 571 1056 591
rect 1090 571 1102 605
rect 1026 391 1102 571
rect 1264 440 1330 592
rect 1264 406 1279 440
rect 1313 406 1330 440
rect 1264 392 1330 406
rect 1360 578 1420 592
rect 1360 544 1373 578
rect 1407 544 1420 578
rect 1360 392 1420 544
rect 1450 440 1512 592
rect 1450 406 1464 440
rect 1498 406 1512 440
rect 1450 392 1512 406
rect 1542 576 1602 592
rect 1542 542 1555 576
rect 1589 542 1602 576
rect 1542 508 1602 542
rect 1542 474 1555 508
rect 1589 474 1602 508
rect 1542 392 1602 474
rect 1632 580 1701 592
rect 1632 546 1655 580
rect 1689 546 1701 580
rect 1632 510 1701 546
rect 1632 476 1655 510
rect 1689 476 1701 510
rect 1632 440 1701 476
rect 1632 406 1655 440
rect 1689 406 1701 440
rect 1632 392 1701 406
rect 598 368 651 391
rect 538 363 550 368
rect 244 330 302 342
rect 492 351 550 363
<< ndiffc >>
rect 70 180 104 214
rect 70 110 104 144
rect 170 180 204 214
rect 170 110 204 144
rect 278 180 312 214
rect 278 90 312 124
rect 378 180 412 214
rect 378 90 412 124
rect 482 180 516 214
rect 482 90 516 124
rect 601 201 635 235
rect 601 90 635 124
rect 720 201 754 235
rect 720 131 754 165
rect 834 131 868 165
rect 948 133 982 167
rect 1057 83 1091 117
rect 1183 86 1217 120
rect 1268 86 1302 120
rect 1368 136 1402 170
rect 1468 150 1502 184
rect 1468 82 1502 116
rect 1554 145 1588 179
rect 1654 156 1688 190
rect 1654 86 1688 120
<< pdiffc >>
rect 39 522 73 556
rect 39 406 73 440
rect 147 546 181 580
rect 256 342 290 376
rect 380 583 414 617
rect 504 363 538 397
rect 628 583 662 617
rect 735 545 769 579
rect 735 471 769 505
rect 842 571 876 605
rect 949 403 983 437
rect 1056 571 1090 605
rect 1279 406 1313 440
rect 1373 544 1407 578
rect 1464 406 1498 440
rect 1555 542 1589 576
rect 1555 474 1589 508
rect 1655 546 1689 580
rect 1655 476 1689 510
rect 1655 406 1689 440
<< poly >>
rect 86 568 116 594
rect 196 592 226 618
rect 320 592 350 618
rect 86 353 116 368
rect 196 353 226 368
rect 83 336 119 353
rect 83 320 151 336
rect 83 286 101 320
rect 135 286 151 320
rect 83 270 151 286
rect 193 271 229 353
rect 444 592 474 618
rect 568 592 598 618
rect 320 353 350 368
rect 444 353 474 368
rect 692 591 722 617
rect 782 591 812 617
rect 906 591 936 617
rect 996 591 1026 617
rect 1330 592 1360 618
rect 1420 592 1450 618
rect 1512 592 1542 618
rect 1602 592 1632 618
rect 692 376 722 391
rect 782 376 812 391
rect 906 376 936 391
rect 996 376 1026 391
rect 1330 377 1360 392
rect 1420 377 1450 392
rect 1512 377 1542 392
rect 1602 377 1632 392
rect 115 226 145 270
rect 193 241 259 271
rect 317 241 353 353
rect 229 226 259 241
rect 323 226 353 241
rect 441 241 477 353
rect 568 353 598 368
rect 689 353 725 376
rect 779 353 815 376
rect 903 353 939 376
rect 993 353 1029 376
rect 1327 356 1363 377
rect 1417 356 1453 377
rect 1509 356 1545 377
rect 1599 356 1635 377
rect 565 292 601 353
rect 527 262 601 292
rect 679 337 815 353
rect 679 303 699 337
rect 733 303 815 337
rect 679 287 815 303
rect 863 337 1029 353
rect 863 303 879 337
rect 913 303 947 337
rect 981 303 1029 337
rect 863 287 1029 303
rect 1077 340 1279 356
rect 1077 306 1093 340
rect 1127 306 1161 340
rect 1195 306 1229 340
rect 1263 306 1279 340
rect 1077 290 1279 306
rect 1327 340 1453 356
rect 1327 306 1344 340
rect 1378 320 1453 340
rect 1501 340 1635 356
rect 1378 306 1447 320
rect 1327 290 1447 306
rect 1501 306 1517 340
rect 1551 306 1585 340
rect 1619 306 1635 340
rect 1501 290 1635 306
rect 441 226 471 241
rect 527 226 557 262
rect 679 247 709 287
rect 779 247 809 287
rect 907 247 937 287
rect 993 247 1023 287
rect 115 72 145 98
rect 679 93 709 119
rect 779 93 809 119
rect 907 93 937 119
rect 993 93 1023 119
rect 229 51 259 78
rect 323 51 353 78
rect 441 51 471 78
rect 527 51 557 78
rect 1126 51 1156 290
rect 1327 202 1357 290
rect 1417 202 1447 290
rect 1513 202 1543 290
rect 1605 202 1635 290
rect 229 21 1156 51
rect 1327 48 1357 74
rect 1417 48 1447 74
rect 1513 48 1543 74
rect 1605 48 1635 74
<< polycont >>
rect 101 286 135 320
rect 699 303 733 337
rect 879 303 913 337
rect 947 303 981 337
rect 1093 306 1127 340
rect 1161 306 1195 340
rect 1229 306 1263 340
rect 1344 306 1378 340
rect 1517 306 1551 340
rect 1585 306 1619 340
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 130 580 199 649
rect 17 556 89 572
rect 17 522 39 556
rect 73 522 89 556
rect 130 546 147 580
rect 181 546 199 580
rect 364 617 430 649
rect 364 583 380 617
rect 414 583 430 617
rect 364 567 430 583
rect 612 617 678 649
rect 612 583 628 617
rect 662 583 678 617
rect 826 605 892 649
rect 612 567 678 583
rect 735 579 785 595
rect 769 545 785 579
rect 826 571 842 605
rect 876 571 892 605
rect 826 555 892 571
rect 1040 605 1090 649
rect 1040 571 1056 605
rect 1040 555 1090 571
rect 1124 578 1423 596
rect 17 512 89 522
rect 233 512 701 533
rect 17 499 701 512
rect 17 478 267 499
rect 17 440 89 478
rect 301 444 633 465
rect 17 406 39 440
rect 73 406 89 440
rect 17 390 89 406
rect 133 431 633 444
rect 133 410 335 431
rect 17 230 51 390
rect 133 356 167 410
rect 488 376 504 397
rect 85 320 167 356
rect 85 286 101 320
rect 135 286 167 320
rect 85 270 167 286
rect 217 342 256 376
rect 290 363 504 376
rect 538 363 554 397
rect 290 342 554 363
rect 599 353 633 431
rect 667 421 701 499
rect 735 521 785 545
rect 1124 544 1373 578
rect 1407 544 1423 578
rect 1124 542 1423 544
rect 1539 576 1605 596
rect 1539 542 1555 576
rect 1589 542 1605 576
rect 1124 521 1158 542
rect 735 505 1158 521
rect 1539 508 1605 542
rect 769 487 1158 505
rect 769 471 785 487
rect 735 455 785 471
rect 1192 474 1555 508
rect 1589 474 1605 508
rect 1639 580 1705 596
rect 1639 546 1655 580
rect 1689 546 1705 580
rect 1639 510 1705 546
rect 1639 476 1655 510
rect 1689 476 1705 510
rect 1192 453 1226 474
rect 933 437 1226 453
rect 1639 440 1705 476
rect 667 387 817 421
rect 933 403 949 437
rect 983 419 1226 437
rect 983 403 1028 419
rect 933 387 1028 403
rect 1260 406 1279 440
rect 1313 406 1464 440
rect 1498 406 1655 440
rect 1689 406 1705 440
rect 1260 390 1705 406
rect 783 353 817 387
rect 1260 356 1294 390
rect 217 274 551 342
rect 599 337 749 353
rect 599 303 699 337
rect 733 303 749 337
rect 599 287 749 303
rect 783 337 997 353
rect 783 303 879 337
rect 913 303 947 337
rect 981 303 997 337
rect 783 287 997 303
rect 1077 340 1294 356
rect 1077 306 1093 340
rect 1127 306 1161 340
rect 1195 306 1229 340
rect 1263 306 1294 340
rect 1077 290 1294 306
rect 1328 340 1415 356
rect 1328 306 1344 340
rect 1378 306 1415 340
rect 1328 290 1415 306
rect 1465 340 1635 356
rect 1465 306 1517 340
rect 1551 306 1585 340
rect 1619 306 1635 340
rect 1465 290 1635 306
rect 17 214 120 230
rect 17 180 70 214
rect 104 180 120 214
rect 17 144 120 180
rect 17 110 70 144
rect 104 110 120 144
rect 17 94 120 110
rect 154 214 220 230
rect 154 180 170 214
rect 204 180 220 214
rect 154 144 220 180
rect 154 110 170 144
rect 204 110 220 144
rect 154 17 220 110
rect 262 214 328 274
rect 466 214 551 274
rect 1031 253 1604 256
rect 262 180 278 214
rect 312 180 328 214
rect 262 124 328 180
rect 262 90 278 124
rect 312 90 328 124
rect 262 74 328 90
rect 362 180 378 214
rect 412 180 428 214
rect 362 124 428 180
rect 362 90 378 124
rect 412 90 428 124
rect 362 17 428 90
rect 466 180 482 214
rect 516 180 551 214
rect 466 124 551 180
rect 466 90 482 124
rect 516 90 551 124
rect 466 74 551 90
rect 585 235 651 251
rect 585 201 601 235
rect 635 201 651 235
rect 585 124 651 201
rect 585 90 601 124
rect 635 90 651 124
rect 704 235 1604 253
rect 704 201 720 235
rect 754 222 1604 235
rect 754 219 1065 222
rect 754 201 770 219
rect 704 165 770 201
rect 1099 185 1418 188
rect 704 131 720 165
rect 754 131 770 165
rect 704 115 770 131
rect 804 165 898 181
rect 804 131 834 165
rect 868 131 898 165
rect 585 17 651 90
rect 804 17 898 131
rect 932 170 1418 185
rect 932 167 1368 170
rect 932 133 948 167
rect 982 154 1368 167
rect 982 151 1133 154
rect 982 133 998 151
rect 932 115 998 133
rect 1352 136 1368 154
rect 1402 136 1418 170
rect 1034 83 1057 117
rect 1091 83 1115 117
rect 1034 17 1115 83
rect 1167 86 1183 120
rect 1217 86 1268 120
rect 1302 86 1318 120
rect 1352 119 1418 136
rect 1452 184 1518 188
rect 1452 150 1468 184
rect 1502 150 1518 184
rect 1167 85 1318 86
rect 1452 116 1518 150
rect 1554 179 1604 222
rect 1671 206 1705 390
rect 1588 145 1604 179
rect 1554 119 1604 145
rect 1638 190 1705 206
rect 1638 156 1654 190
rect 1688 156 1705 190
rect 1638 120 1705 156
rect 1452 85 1468 116
rect 1167 82 1468 85
rect 1502 85 1518 116
rect 1638 86 1654 120
rect 1688 86 1705 120
rect 1638 85 1705 86
rect 1502 82 1705 85
rect 1167 51 1705 82
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
<< metal1 >>
rect 0 683 1728 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 0 617 1728 649
rect 0 17 1728 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
rect 0 -49 1728 -17
<< labels >>
rlabel comment s 0 0 0 0 4 mux2_4
flabel pwell s 0 0 1728 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 1728 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 1728 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 1728 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 1375 316 1409 350 0 FreeSans 340 0 0 0 A0
port 1 nsew
flabel corelocali s 1471 316 1505 350 0 FreeSans 340 0 0 0 A1
port 2 nsew
flabel corelocali s 1567 316 1601 350 0 FreeSans 340 0 0 0 A1
port 2 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 S
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 1728 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1598978
string GDS_START 1586614
<< end >>
