magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 119 367 153 527
rect 287 367 321 527
rect 371 323 405 493
rect 439 367 505 527
rect 539 323 573 493
rect 607 367 673 527
rect 707 323 741 493
rect 775 367 841 527
rect 875 323 909 493
rect 371 289 909 323
rect 943 297 1009 527
rect 28 215 248 255
rect 858 263 909 289
rect 858 255 974 263
rect 858 221 861 255
rect 895 221 933 255
rect 967 221 974 255
rect 858 211 974 221
rect 858 181 909 211
rect 371 147 909 181
rect 103 17 169 113
rect 271 17 337 113
rect 371 51 405 147
rect 439 17 505 113
rect 539 51 573 147
rect 607 17 673 113
rect 707 51 741 147
rect 775 17 841 113
rect 875 51 909 147
rect 943 17 1009 177
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 861 221 895 255
rect 933 221 967 255
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< obsli1 >>
rect 19 323 85 493
rect 187 323 253 493
rect 19 289 319 323
rect 284 249 319 289
rect 284 215 809 249
rect 284 181 319 215
rect 35 147 319 181
rect 35 51 69 147
rect 203 52 237 147
<< metal1 >>
rect 0 570 1104 592
rect 0 561 1168 570
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 559 1168 561
rect 1087 529 1121 559
rect 1151 529 1168 559
rect 1075 527 1168 529
rect 0 518 1168 527
rect 0 496 1104 518
rect 404 253 532 264
rect 404 223 421 253
rect 451 223 485 253
rect 515 252 532 253
rect 849 255 979 261
rect 849 252 861 255
rect 515 224 861 252
rect 515 223 532 224
rect 404 212 532 223
rect 849 221 861 224
rect 895 221 933 255
rect 967 221 979 255
rect 849 215 979 221
rect 0 26 1104 48
rect 0 17 1168 26
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 15 1168 17
rect 1087 -15 1121 15
rect 1151 -15 1168 15
rect 1075 -17 1168 -15
rect 0 -26 1168 -17
rect 0 -48 1104 -26
<< via1 >>
rect 1057 529 1075 559
rect 1075 529 1087 559
rect 1121 529 1151 559
rect 421 223 451 253
rect 485 223 515 253
rect 1057 -15 1075 15
rect 1075 -15 1087 15
rect 1121 -15 1151 15
<< metal2 >>
rect 1027 564 1181 572
rect 1027 524 1044 564
rect 1084 559 1124 564
rect 1087 529 1121 559
rect 1084 524 1124 529
rect 1164 524 1181 564
rect 1027 516 1181 524
rect 378 258 532 266
rect 378 218 395 258
rect 435 253 475 258
rect 451 223 475 253
rect 435 218 475 223
rect 515 218 532 258
rect 378 210 532 218
rect 1027 20 1181 28
rect 1027 -20 1044 20
rect 1084 15 1124 20
rect 1087 -15 1121 15
rect 1084 -20 1124 -15
rect 1164 -20 1181 20
rect 1027 -28 1181 -20
<< via2 >>
rect 1044 559 1084 564
rect 1124 559 1164 564
rect 1044 529 1057 559
rect 1057 529 1084 559
rect 1124 529 1151 559
rect 1151 529 1164 559
rect 1044 524 1084 529
rect 1124 524 1164 529
rect 395 253 435 258
rect 475 253 515 258
rect 395 223 421 253
rect 421 223 435 253
rect 475 223 485 253
rect 485 223 515 253
rect 395 218 435 223
rect 475 218 515 223
rect 1044 15 1084 20
rect 1124 15 1164 20
rect 1044 -15 1057 15
rect 1057 -15 1084 15
rect 1124 -15 1151 15
rect 1151 -15 1164 15
rect 1044 -20 1084 -15
rect 1124 -20 1164 -15
<< metal3 >>
rect 1026 564 1182 577
rect 1026 524 1044 564
rect 1084 524 1124 564
rect 1164 524 1182 564
rect 1026 511 1182 524
rect -143 258 13 270
rect -143 218 -125 258
rect -85 218 -45 258
rect -5 218 13 258
rect -143 206 13 218
rect 377 258 533 271
rect 377 218 395 258
rect 435 218 475 258
rect 515 218 533 258
rect 377 205 533 218
rect 1026 20 1182 33
rect 1026 -20 1044 20
rect 1084 -20 1124 20
rect 1164 -20 1182 20
rect 1026 -33 1182 -20
<< via3 >>
rect 1044 524 1084 564
rect 1124 524 1164 564
rect -125 218 -85 258
rect -45 218 -5 258
rect 395 218 435 258
rect 475 218 515 258
rect 1044 -20 1084 20
rect 1124 -20 1164 20
<< metal4 >>
rect 986 685 1222 723
rect 986 525 1024 685
rect 1184 525 1222 685
rect 986 524 1044 525
rect 1084 524 1124 525
rect 1164 524 1222 525
rect 986 487 1222 524
rect -228 352 8 390
rect -228 192 -190 352
rect -30 258 8 352
rect -5 218 8 258
rect -30 192 8 218
rect -228 154 8 192
rect 292 352 528 390
rect 292 192 330 352
rect 490 258 528 352
rect 515 218 528 258
rect 490 192 528 218
rect 292 154 528 192
rect 986 20 1222 57
rect 986 19 1044 20
rect 1084 19 1124 20
rect 1164 19 1222 20
rect 986 -141 1024 19
rect 1184 -141 1222 19
rect 986 -179 1222 -141
<< via4 >>
rect 1024 564 1184 685
rect 1024 525 1044 564
rect 1044 525 1084 564
rect 1084 525 1124 564
rect 1124 525 1164 564
rect 1164 525 1184 564
rect -190 258 -30 352
rect -190 218 -125 258
rect -125 218 -85 258
rect -85 218 -45 258
rect -45 218 -30 258
rect -190 192 -30 218
rect 330 258 490 352
rect 330 218 395 258
rect 395 218 435 258
rect 435 218 475 258
rect 475 218 490 258
rect 330 192 490 218
rect 1024 -20 1044 19
rect 1044 -20 1084 19
rect 1084 -20 1124 19
rect 1124 -20 1164 19
rect 1164 -20 1184 19
rect 1024 -141 1184 -20
<< metal5 >>
rect 232 432 552 765
rect 872 685 1335 778
rect 872 525 1024 685
rect 1184 525 1335 685
rect 872 432 1335 525
rect -252 352 552 432
rect -252 192 -190 352
rect -30 192 330 352
rect 490 192 552 352
rect -252 112 552 192
rect 232 -221 552 112
rect 872 19 1335 112
rect 872 -141 1024 19
rect 1184 -141 1335 19
rect 872 -234 1335 -141
<< labels >>
rlabel locali s 28 215 248 255 6 A
port 1 nsew signal input
rlabel locali s 875 323 909 493 6 X
port 2 nsew signal output
rlabel locali s 875 51 909 147 6 X
port 2 nsew signal output
rlabel locali s 858 263 909 289 6 X
port 2 nsew signal output
rlabel locali s 858 211 974 263 6 X
port 2 nsew signal output
rlabel locali s 858 181 909 211 6 X
port 2 nsew signal output
rlabel locali s 707 323 741 493 6 X
port 2 nsew signal output
rlabel locali s 707 51 741 147 6 X
port 2 nsew signal output
rlabel locali s 539 323 573 493 6 X
port 2 nsew signal output
rlabel locali s 539 51 573 147 6 X
port 2 nsew signal output
rlabel locali s 371 323 405 493 6 X
port 2 nsew signal output
rlabel locali s 371 289 909 323 6 X
port 2 nsew signal output
rlabel locali s 371 147 909 181 6 X
port 2 nsew signal output
rlabel locali s 371 51 405 147 6 X
port 2 nsew signal output
rlabel via4 s 330 192 490 352 6 X
port 2 nsew signal output
rlabel via4 s -190 192 -30 352 4 X
port 2 nsew signal output
rlabel via3 s 475 218 515 258 6 X
port 2 nsew signal output
rlabel via3 s 395 218 435 258 6 X
port 2 nsew signal output
rlabel via3 s -45 218 -5 258 4 X
port 2 nsew signal output
rlabel via3 s -125 218 -85 258 4 X
port 2 nsew signal output
rlabel via2 s 475 218 515 258 6 X
port 2 nsew signal output
rlabel via2 s 395 218 435 258 6 X
port 2 nsew signal output
rlabel via1 s 485 223 515 253 6 X
port 2 nsew signal output
rlabel via1 s 421 223 451 253 6 X
port 2 nsew signal output
rlabel viali s 933 221 967 255 6 X
port 2 nsew signal output
rlabel viali s 861 221 895 255 6 X
port 2 nsew signal output
rlabel metal1 s 849 252 979 261 6 X
port 2 nsew signal output
rlabel metal1 s 849 215 979 224 6 X
port 2 nsew signal output
rlabel metal1 s 404 252 532 264 6 X
port 2 nsew signal output
rlabel metal1 s 404 224 979 252 6 X
port 2 nsew signal output
rlabel metal1 s 404 212 532 224 6 X
port 2 nsew signal output
rlabel metal2 s 378 210 532 266 6 X
port 2 nsew signal output
rlabel metal3 s -143 206 13 270 4 X
port 2 nsew signal output
rlabel metal3 s 377 205 533 271 6 X
port 2 nsew signal output
rlabel metal4 s -228 154 8 390 4 X
port 2 nsew signal output
rlabel metal4 s 292 154 528 390 6 X
port 2 nsew signal output
rlabel metal5 s 232 432 552 765 6 X
port 2 nsew signal output
rlabel metal5 s 232 -221 552 112 8 X
port 2 nsew signal output
rlabel metal5 s -252 112 552 432 6 X
port 2 nsew signal output
rlabel locali s 943 17 1009 177 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 775 17 841 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 607 17 673 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 439 17 505 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 271 17 337 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 103 17 169 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 0 -17 1104 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel via4 s 1024 -141 1184 19 8 VGND
port 3 nsew ground bidirectional abutment
rlabel via3 s 1124 -20 1164 20 8 VGND
port 3 nsew ground bidirectional abutment
rlabel via3 s 1044 -20 1084 20 8 VGND
port 3 nsew ground bidirectional abutment
rlabel via2 s 1124 -20 1164 20 8 VGND
port 3 nsew ground bidirectional abutment
rlabel via2 s 1044 -20 1084 20 8 VGND
port 3 nsew ground bidirectional abutment
rlabel via1 s 1121 -15 1151 15 8 VGND
port 3 nsew ground bidirectional abutment
rlabel via1 s 1057 -15 1087 15 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 1041 -17 1075 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 949 -17 983 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 857 -17 891 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 765 -17 799 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 673 -17 707 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 581 -17 615 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 489 -17 523 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 397 -17 431 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 305 -17 339 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 213 -17 247 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 121 -17 155 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 29 -17 63 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 26 1104 48 6 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -26 1168 26 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1104 -26 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal2 s 1027 -28 1181 28 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal3 s 1026 -33 1182 33 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal4 s 986 -179 1222 57 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal5 s 872 -234 1335 112 8 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 943 297 1009 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 775 367 841 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 607 367 673 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 439 367 505 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 287 367 321 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 119 367 153 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 0 527 1104 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel via4 s 1024 525 1184 685 6 VPWR
port 4 nsew power bidirectional abutment
rlabel via3 s 1124 524 1164 564 6 VPWR
port 4 nsew power bidirectional abutment
rlabel via3 s 1044 524 1084 564 6 VPWR
port 4 nsew power bidirectional abutment
rlabel via2 s 1124 524 1164 564 6 VPWR
port 4 nsew power bidirectional abutment
rlabel via2 s 1044 524 1084 564 6 VPWR
port 4 nsew power bidirectional abutment
rlabel via1 s 1121 529 1151 559 6 VPWR
port 4 nsew power bidirectional abutment
rlabel via1 s 1057 529 1087 559 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 1041 527 1075 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 949 527 983 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 857 527 891 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 765 527 799 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 673 527 707 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 581 527 615 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 489 527 523 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 397 527 431 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 305 527 339 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 213 527 247 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 121 527 155 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 29 527 63 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 570 1104 592 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 518 1168 570 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 496 1104 518 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal2 s 1027 516 1181 572 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal3 s 1026 511 1182 577 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal4 s 986 487 1222 723 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal5 s 872 432 1335 778 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1104 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 31774
string GDS_START 18966
<< end >>
