magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 644 561
rect 72 365 157 493
rect 17 146 87 331
rect 121 177 157 365
rect 191 211 265 472
rect 408 451 474 527
rect 299 211 369 347
rect 471 280 525 347
rect 407 214 525 280
rect 121 127 408 177
rect 471 132 525 214
rect 559 130 627 347
rect 157 123 408 127
rect 57 17 123 93
rect 157 51 208 123
rect 242 17 308 89
rect 342 56 408 123
rect 494 17 560 96
rect 0 -17 644 17
<< obsli1 >>
rect 308 417 374 493
rect 508 417 574 493
rect 308 381 574 417
<< metal1 >>
rect 0 496 644 592
rect 0 -48 644 48
<< labels >>
rlabel locali s 471 280 525 347 6 A1
port 1 nsew signal input
rlabel locali s 471 132 525 214 6 A1
port 1 nsew signal input
rlabel locali s 407 214 525 280 6 A1
port 1 nsew signal input
rlabel locali s 559 130 627 347 6 A2
port 2 nsew signal input
rlabel locali s 299 211 369 347 6 B1
port 3 nsew signal input
rlabel locali s 191 211 265 472 6 C1
port 4 nsew signal input
rlabel locali s 17 146 87 331 6 D1
port 5 nsew signal input
rlabel locali s 342 56 408 123 6 Y
port 6 nsew signal output
rlabel locali s 157 123 408 127 6 Y
port 6 nsew signal output
rlabel locali s 157 51 208 123 6 Y
port 6 nsew signal output
rlabel locali s 121 177 157 365 6 Y
port 6 nsew signal output
rlabel locali s 121 127 408 177 6 Y
port 6 nsew signal output
rlabel locali s 72 365 157 493 6 Y
port 6 nsew signal output
rlabel locali s 494 17 560 96 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 242 17 308 89 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 57 17 123 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 644 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 644 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 408 451 474 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 644 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 644 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3896730
string GDS_START 3889282
<< end >>
