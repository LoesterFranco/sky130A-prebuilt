magic
tech sky130A
magscale 1 2
timestamp 1604502697
<< nwell >>
rect -38 261 1050 582
<< pwell >>
rect 176 -17 220 17
<< scnmos >>
rect 87 47 117 151
rect 171 47 201 151
rect 307 47 337 131
rect 409 47 439 131
rect 540 47 570 131
rect 741 47 771 131
rect 865 47 895 151
<< pmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 299 309 335 497
rect 418 309 454 497
rect 655 309 691 497
rect 743 309 779 497
rect 857 309 893 497
<< ndiff >>
rect 27 115 87 151
rect 27 81 35 115
rect 69 81 87 115
rect 27 47 87 81
rect 117 112 171 151
rect 117 78 127 112
rect 161 78 171 112
rect 117 47 171 78
rect 201 131 263 151
rect 815 131 865 151
rect 201 93 307 131
rect 201 59 221 93
rect 255 59 307 93
rect 201 47 307 59
rect 337 47 409 131
rect 439 108 540 131
rect 439 74 482 108
rect 516 74 540 108
rect 439 47 540 74
rect 570 47 741 131
rect 771 89 865 131
rect 771 55 801 89
rect 835 55 865 89
rect 771 47 865 55
rect 895 108 947 151
rect 895 74 905 108
rect 939 74 947 108
rect 895 47 947 74
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 485 175 497
rect 117 451 129 485
rect 163 451 175 485
rect 117 417 175 451
rect 117 383 129 417
rect 163 383 175 417
rect 117 349 175 383
rect 117 315 129 349
rect 163 315 175 349
rect 117 297 175 315
rect 211 485 299 497
rect 211 451 223 485
rect 257 451 299 485
rect 211 417 299 451
rect 211 383 223 417
rect 257 383 299 417
rect 211 349 299 383
rect 211 315 223 349
rect 257 315 299 349
rect 211 309 299 315
rect 335 309 418 497
rect 454 425 655 497
rect 454 391 466 425
rect 500 391 541 425
rect 575 391 609 425
rect 643 391 655 425
rect 454 309 655 391
rect 691 309 743 497
rect 779 485 857 497
rect 779 451 809 485
rect 843 451 857 485
rect 779 417 857 451
rect 779 383 809 417
rect 843 383 857 417
rect 779 309 857 383
rect 893 485 951 497
rect 893 451 905 485
rect 939 451 951 485
rect 893 417 951 451
rect 893 383 905 417
rect 939 383 951 417
rect 893 309 951 383
rect 211 297 265 309
<< ndiffc >>
rect 35 81 69 115
rect 127 78 161 112
rect 221 59 255 93
rect 482 74 516 108
rect 801 55 835 89
rect 905 74 939 108
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 451 163 485
rect 129 383 163 417
rect 129 315 163 349
rect 223 451 257 485
rect 223 383 257 417
rect 223 315 257 349
rect 466 391 500 425
rect 541 391 575 425
rect 609 391 643 425
rect 809 451 843 485
rect 809 383 843 417
rect 905 451 939 485
rect 905 383 939 417
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 299 497 335 523
rect 418 497 454 523
rect 655 497 691 523
rect 743 497 779 523
rect 857 497 893 523
rect 81 282 117 297
rect 175 282 211 297
rect 299 294 335 309
rect 418 294 454 309
rect 655 294 691 309
rect 743 294 779 309
rect 857 294 893 309
rect 79 265 119 282
rect 173 265 213 282
rect 297 265 337 294
rect 79 249 239 265
rect 79 215 195 249
rect 229 215 239 249
rect 79 199 239 215
rect 281 249 337 265
rect 416 264 580 294
rect 653 277 693 294
rect 281 215 291 249
rect 325 215 337 249
rect 540 229 580 264
rect 639 261 693 277
rect 281 199 337 215
rect 87 151 117 199
rect 171 151 201 199
rect 307 131 337 199
rect 409 212 498 222
rect 409 178 448 212
rect 482 178 498 212
rect 409 168 498 178
rect 540 213 594 229
rect 540 179 550 213
rect 584 179 594 213
rect 639 227 649 261
rect 683 227 693 261
rect 639 211 693 227
rect 741 237 781 294
rect 855 277 895 294
rect 843 261 897 277
rect 741 221 801 237
rect 409 131 439 168
rect 540 163 594 179
rect 741 187 757 221
rect 791 187 801 221
rect 843 227 853 261
rect 887 227 897 261
rect 843 211 897 227
rect 741 171 801 187
rect 540 131 570 163
rect 741 131 771 171
rect 865 151 895 211
rect 87 21 117 47
rect 171 21 201 47
rect 307 21 337 47
rect 409 21 439 47
rect 540 21 570 47
rect 741 21 771 47
rect 865 21 895 47
<< polycont >>
rect 195 215 229 249
rect 291 215 325 249
rect 448 178 482 212
rect 550 179 584 213
rect 649 227 683 261
rect 757 187 791 221
rect 853 227 887 261
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 27 485 76 527
rect 27 451 35 485
rect 69 451 76 485
rect 27 417 76 451
rect 27 383 35 417
rect 69 383 76 417
rect 27 349 76 383
rect 27 315 35 349
rect 69 315 76 349
rect 27 299 76 315
rect 111 485 179 493
rect 111 451 129 485
rect 163 451 179 485
rect 111 417 179 451
rect 111 383 129 417
rect 163 383 179 417
rect 111 349 179 383
rect 111 315 129 349
rect 163 315 179 349
rect 111 299 179 315
rect 215 485 265 527
rect 215 451 223 485
rect 257 451 265 485
rect 215 417 265 451
rect 215 383 223 417
rect 257 383 265 417
rect 215 349 265 383
rect 215 315 223 349
rect 257 315 265 349
rect 215 299 265 315
rect 306 459 775 493
rect 27 115 77 131
rect 27 81 35 115
rect 69 81 77 115
rect 27 17 77 81
rect 111 112 161 299
rect 306 265 346 459
rect 195 249 229 265
rect 195 165 229 215
rect 291 249 346 265
rect 325 215 346 249
rect 291 199 346 215
rect 380 391 466 425
rect 500 391 541 425
rect 575 391 609 425
rect 643 391 669 425
rect 380 165 414 391
rect 195 131 414 165
rect 448 323 707 357
rect 448 212 482 323
rect 448 162 482 178
rect 550 213 615 283
rect 584 179 615 213
rect 111 78 127 112
rect 379 124 414 131
rect 379 108 516 124
rect 111 51 161 78
rect 195 93 271 97
rect 195 59 221 93
rect 255 59 271 93
rect 195 17 271 59
rect 379 74 482 108
rect 379 51 516 74
rect 550 51 615 179
rect 649 261 707 323
rect 741 326 775 459
rect 809 485 855 527
rect 843 451 855 485
rect 809 417 855 451
rect 843 383 855 417
rect 809 367 855 383
rect 889 485 969 493
rect 889 451 905 485
rect 939 451 969 485
rect 889 417 969 451
rect 889 383 905 417
rect 939 383 969 417
rect 889 367 969 383
rect 741 288 891 326
rect 683 227 707 261
rect 853 261 891 288
rect 649 51 707 227
rect 757 221 791 237
rect 887 227 891 261
rect 853 211 891 227
rect 757 173 791 187
rect 935 173 969 367
rect 757 139 969 173
rect 899 108 948 139
rect 742 89 845 105
rect 742 55 801 89
rect 835 55 845 89
rect 742 17 845 55
rect 899 74 905 108
rect 939 74 948 108
rect 899 51 948 74
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
flabel metal1 s 122 -17 156 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 122 527 156 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
flabel corelocali s 764 289 798 323 0 FreeSans 250 0 0 0 S
port 3 nsew
flabel corelocali s 673 153 707 187 0 FreeSans 250 0 0 0 A1
port 2 nsew
flabel corelocali s 673 221 707 255 0 FreeSans 250 0 0 0 A1
port 2 nsew
flabel corelocali s 581 221 615 255 0 FreeSans 250 0 0 0 A0
port 1 nsew
flabel corelocali s 122 85 156 119 0 FreeSans 250 0 0 0 X
port 8 nsew
flabel corelocali s 122 357 156 391 0 FreeSans 250 0 0 0 X
port 8 nsew
flabel corelocali s 122 425 156 459 0 FreeSans 250 0 0 0 X
port 8 nsew
flabel corelocali s 853 289 887 323 0 FreeSans 250 0 0 0 S
port 3 nsew
flabel nbase s 166 527 200 561 0 FreeSans 250 0 0 0 VPB
port 6 nsew
flabel pwell s 176 -17 220 17 0 FreeSans 250 0 0 0 VNB
port 5 nsew
rlabel comment s 0 0 0 0 4 clkmux2_2
<< properties >>
string FIXED_BBOX 0 0 1012 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3284060
string GDS_START 3276300
<< end >>
