magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 112 963 167 1009
rect 112 877 146 963
rect 67 823 146 877
rect 361 829 441 899
rect 479 829 559 899
rect 753 963 808 1009
rect 774 877 808 963
rect 940 963 995 1009
rect 940 877 974 963
rect 774 823 853 877
rect 895 823 974 877
rect 67 211 146 265
rect 112 125 146 211
rect 1189 829 1269 899
rect 1307 829 1387 899
rect 1581 963 1636 1009
rect 112 79 167 125
rect 361 189 441 259
rect 479 189 559 259
rect 1602 877 1636 963
rect 1768 963 1823 1009
rect 1768 877 1802 963
rect 1602 823 1681 877
rect 1723 823 1802 877
rect 774 211 853 265
rect 895 211 974 265
rect 774 125 808 211
rect 753 79 808 125
rect 940 125 974 211
rect 2017 829 2097 899
rect 2135 829 2215 899
rect 2409 963 2464 1009
rect 940 79 995 125
rect 1189 189 1269 259
rect 1307 189 1387 259
rect 2430 877 2464 963
rect 2596 963 2651 1009
rect 2596 877 2630 963
rect 2430 823 2509 877
rect 2551 823 2630 877
rect 1602 211 1681 265
rect 1723 211 1802 265
rect 1602 125 1636 211
rect 1581 79 1636 125
rect 1768 125 1802 211
rect 2845 829 2925 899
rect 2963 829 3043 899
rect 3237 963 3292 1009
rect 1768 79 1823 125
rect 2017 189 2097 259
rect 2135 189 2215 259
rect 3258 877 3292 963
rect 3258 823 3337 877
rect 2430 211 2509 265
rect 2551 211 2630 265
rect 2430 125 2464 211
rect 2409 79 2464 125
rect 2596 125 2630 211
rect 2596 79 2651 125
rect 2845 189 2925 259
rect 2963 189 3043 259
rect 3258 211 3337 265
rect 3258 125 3292 211
rect 3237 79 3292 125
<< obsli1 >>
rect 0 1071 29 1105
rect 63 1071 121 1105
rect 155 1071 213 1105
rect 247 1071 305 1105
rect 339 1071 397 1105
rect 431 1071 489 1105
rect 523 1071 581 1105
rect 615 1071 673 1105
rect 707 1071 765 1105
rect 799 1071 857 1105
rect 891 1071 949 1105
rect 983 1071 1041 1105
rect 1075 1071 1133 1105
rect 1167 1071 1225 1105
rect 1259 1071 1317 1105
rect 1351 1071 1409 1105
rect 1443 1071 1501 1105
rect 1535 1071 1593 1105
rect 1627 1071 1685 1105
rect 1719 1071 1777 1105
rect 1811 1071 1869 1105
rect 1903 1071 1961 1105
rect 1995 1071 2053 1105
rect 2087 1071 2145 1105
rect 2179 1071 2237 1105
rect 2271 1071 2329 1105
rect 2363 1071 2421 1105
rect 2455 1071 2513 1105
rect 2547 1071 2605 1105
rect 2639 1071 2697 1105
rect 2731 1071 2789 1105
rect 2823 1071 2881 1105
rect 2915 1071 2973 1105
rect 3007 1071 3065 1105
rect 3099 1071 3157 1105
rect 3191 1071 3249 1105
rect 3283 1071 3341 1105
rect 3375 1071 3404 1105
rect 26 911 78 1071
rect 209 921 258 1022
rect 330 971 380 1022
rect 180 887 258 921
rect 292 937 380 971
rect 427 956 493 1071
rect 540 971 590 1022
rect 540 937 628 971
rect 19 561 85 789
rect 180 737 214 887
rect 292 853 326 937
rect 248 795 326 853
rect 594 853 628 937
rect 662 921 711 1022
rect 662 887 740 921
rect 594 795 672 853
rect 248 787 388 795
rect 292 761 388 787
rect 180 731 259 737
rect 180 697 213 731
rect 247 727 259 731
rect 247 697 284 727
rect 180 691 284 697
rect 218 595 284 691
rect 322 595 388 761
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 184 561
rect 19 299 85 527
rect 218 493 259 595
rect 427 561 493 795
rect 532 787 672 795
rect 532 761 628 787
rect 532 595 598 761
rect 706 737 740 887
rect 842 911 906 1071
rect 1037 921 1086 1022
rect 1158 971 1208 1022
rect 1008 887 1086 921
rect 1120 937 1208 971
rect 1255 956 1321 1071
rect 1368 971 1418 1022
rect 1368 937 1456 971
rect 661 731 740 737
rect 661 727 673 731
rect 636 697 673 727
rect 707 697 740 731
rect 636 691 740 697
rect 636 595 702 691
rect 293 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 627 561
rect 218 397 284 493
rect 180 391 284 397
rect 180 357 213 391
rect 247 361 284 391
rect 247 357 259 361
rect 180 351 259 357
rect 26 17 78 177
rect 180 201 214 351
rect 322 327 388 493
rect 292 301 388 327
rect 248 293 388 301
rect 427 293 493 527
rect 661 493 702 595
rect 835 561 913 789
rect 1008 737 1042 887
rect 1120 853 1154 937
rect 1076 795 1154 853
rect 1422 853 1456 937
rect 1490 921 1539 1022
rect 1490 887 1568 921
rect 1422 795 1500 853
rect 1076 787 1216 795
rect 1120 761 1216 787
rect 1008 731 1087 737
rect 1008 697 1041 731
rect 1075 727 1087 731
rect 1075 697 1112 727
rect 1008 691 1112 697
rect 1046 595 1112 691
rect 1150 595 1216 761
rect 736 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 532 327 598 493
rect 636 397 702 493
rect 636 391 740 397
rect 636 361 673 391
rect 661 357 673 361
rect 707 357 740 391
rect 661 351 740 357
rect 532 301 628 327
rect 532 293 672 301
rect 248 235 326 293
rect 180 167 258 201
rect 209 66 258 167
rect 292 151 326 235
rect 594 235 672 293
rect 594 151 628 235
rect 706 201 740 351
rect 835 299 913 527
rect 1046 493 1087 595
rect 1255 561 1321 795
rect 1360 787 1500 795
rect 1360 761 1456 787
rect 1360 595 1426 761
rect 1534 737 1568 887
rect 1670 911 1734 1071
rect 1865 921 1914 1022
rect 1986 971 2036 1022
rect 1836 887 1914 921
rect 1948 937 2036 971
rect 2083 956 2149 1071
rect 2196 971 2246 1022
rect 2196 937 2284 971
rect 1489 731 1568 737
rect 1489 727 1501 731
rect 1464 697 1501 727
rect 1535 697 1568 731
rect 1464 691 1568 697
rect 1464 595 1530 691
rect 1121 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1455 561
rect 1046 397 1112 493
rect 1008 391 1112 397
rect 1008 357 1041 391
rect 1075 361 1112 391
rect 1075 357 1087 361
rect 1008 351 1087 357
rect 292 117 380 151
rect 330 66 380 117
rect 427 17 493 132
rect 540 117 628 151
rect 662 167 740 201
rect 540 66 590 117
rect 662 66 711 167
rect 842 17 906 177
rect 1008 201 1042 351
rect 1150 327 1216 493
rect 1120 301 1216 327
rect 1076 293 1216 301
rect 1255 293 1321 527
rect 1489 493 1530 595
rect 1663 561 1741 789
rect 1836 737 1870 887
rect 1948 853 1982 937
rect 1904 795 1982 853
rect 2250 853 2284 937
rect 2318 921 2367 1022
rect 2318 887 2396 921
rect 2250 795 2328 853
rect 1904 787 2044 795
rect 1948 761 2044 787
rect 1836 731 1915 737
rect 1836 697 1869 731
rect 1903 727 1915 731
rect 1903 697 1940 727
rect 1836 691 1940 697
rect 1874 595 1940 691
rect 1978 595 2044 761
rect 1564 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 1360 327 1426 493
rect 1464 397 1530 493
rect 1464 391 1568 397
rect 1464 361 1501 391
rect 1489 357 1501 361
rect 1535 357 1568 391
rect 1489 351 1568 357
rect 1360 301 1456 327
rect 1360 293 1500 301
rect 1076 235 1154 293
rect 1008 167 1086 201
rect 1037 66 1086 167
rect 1120 151 1154 235
rect 1422 235 1500 293
rect 1422 151 1456 235
rect 1534 201 1568 351
rect 1663 299 1741 527
rect 1874 493 1915 595
rect 2083 561 2149 795
rect 2188 787 2328 795
rect 2188 761 2284 787
rect 2188 595 2254 761
rect 2362 737 2396 887
rect 2498 911 2562 1071
rect 2693 921 2742 1022
rect 2814 971 2864 1022
rect 2664 887 2742 921
rect 2776 937 2864 971
rect 2911 956 2977 1071
rect 3024 971 3074 1022
rect 3024 937 3112 971
rect 2317 731 2396 737
rect 2317 727 2329 731
rect 2292 697 2329 727
rect 2363 697 2396 731
rect 2292 691 2396 697
rect 2292 595 2358 691
rect 1949 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2283 561
rect 1874 397 1940 493
rect 1836 391 1940 397
rect 1836 357 1869 391
rect 1903 361 1940 391
rect 1903 357 1915 361
rect 1836 351 1915 357
rect 1120 117 1208 151
rect 1158 66 1208 117
rect 1255 17 1321 132
rect 1368 117 1456 151
rect 1490 167 1568 201
rect 1368 66 1418 117
rect 1490 66 1539 167
rect 1670 17 1734 177
rect 1836 201 1870 351
rect 1978 327 2044 493
rect 1948 301 2044 327
rect 1904 293 2044 301
rect 2083 293 2149 527
rect 2317 493 2358 595
rect 2491 561 2569 789
rect 2664 737 2698 887
rect 2776 853 2810 937
rect 2732 795 2810 853
rect 3078 853 3112 937
rect 3146 921 3195 1022
rect 3146 887 3224 921
rect 3078 795 3156 853
rect 2732 787 2872 795
rect 2776 761 2872 787
rect 2664 731 2743 737
rect 2664 697 2697 731
rect 2731 727 2743 731
rect 2731 697 2768 727
rect 2664 691 2768 697
rect 2702 595 2768 691
rect 2806 595 2872 761
rect 2392 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2668 561
rect 2188 327 2254 493
rect 2292 397 2358 493
rect 2292 391 2396 397
rect 2292 361 2329 391
rect 2317 357 2329 361
rect 2363 357 2396 391
rect 2317 351 2396 357
rect 2188 301 2284 327
rect 2188 293 2328 301
rect 1904 235 1982 293
rect 1836 167 1914 201
rect 1865 66 1914 167
rect 1948 151 1982 235
rect 2250 235 2328 293
rect 2250 151 2284 235
rect 2362 201 2396 351
rect 2491 299 2569 527
rect 2702 493 2743 595
rect 2911 561 2977 795
rect 3016 787 3156 795
rect 3016 761 3112 787
rect 3016 595 3082 761
rect 3190 737 3224 887
rect 3326 911 3378 1071
rect 3145 731 3224 737
rect 3145 727 3157 731
rect 3120 697 3157 727
rect 3191 697 3224 731
rect 3120 691 3224 697
rect 3120 595 3186 691
rect 2777 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3111 561
rect 2702 397 2768 493
rect 2664 391 2768 397
rect 2664 357 2697 391
rect 2731 361 2768 391
rect 2731 357 2743 361
rect 2664 351 2743 357
rect 1948 117 2036 151
rect 1986 66 2036 117
rect 2083 17 2149 132
rect 2196 117 2284 151
rect 2318 167 2396 201
rect 2196 66 2246 117
rect 2318 66 2367 167
rect 2498 17 2562 177
rect 2664 201 2698 351
rect 2806 327 2872 493
rect 2776 301 2872 327
rect 2732 293 2872 301
rect 2911 293 2977 527
rect 3145 493 3186 595
rect 3319 561 3385 789
rect 3220 527 3249 561
rect 3283 527 3341 561
rect 3375 527 3404 561
rect 3016 327 3082 493
rect 3120 397 3186 493
rect 3120 391 3224 397
rect 3120 361 3157 391
rect 3145 357 3157 361
rect 3191 357 3224 391
rect 3145 351 3224 357
rect 3016 301 3112 327
rect 3016 293 3156 301
rect 2732 235 2810 293
rect 2664 167 2742 201
rect 2693 66 2742 167
rect 2776 151 2810 235
rect 3078 235 3156 293
rect 3078 151 3112 235
rect 3190 201 3224 351
rect 3319 299 3385 527
rect 2776 117 2864 151
rect 2814 66 2864 117
rect 2911 17 2977 132
rect 3024 117 3112 151
rect 3146 167 3224 201
rect 3024 66 3074 117
rect 3146 66 3195 167
rect 3326 17 3378 177
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3341 17
rect 3375 -17 3404 17
<< obsli1c >>
rect 29 1071 63 1105
rect 121 1071 155 1105
rect 213 1071 247 1105
rect 305 1071 339 1105
rect 397 1071 431 1105
rect 489 1071 523 1105
rect 581 1071 615 1105
rect 673 1071 707 1105
rect 765 1071 799 1105
rect 857 1071 891 1105
rect 949 1071 983 1105
rect 1041 1071 1075 1105
rect 1133 1071 1167 1105
rect 1225 1071 1259 1105
rect 1317 1071 1351 1105
rect 1409 1071 1443 1105
rect 1501 1071 1535 1105
rect 1593 1071 1627 1105
rect 1685 1071 1719 1105
rect 1777 1071 1811 1105
rect 1869 1071 1903 1105
rect 1961 1071 1995 1105
rect 2053 1071 2087 1105
rect 2145 1071 2179 1105
rect 2237 1071 2271 1105
rect 2329 1071 2363 1105
rect 2421 1071 2455 1105
rect 2513 1071 2547 1105
rect 2605 1071 2639 1105
rect 2697 1071 2731 1105
rect 2789 1071 2823 1105
rect 2881 1071 2915 1105
rect 2973 1071 3007 1105
rect 3065 1071 3099 1105
rect 3157 1071 3191 1105
rect 3249 1071 3283 1105
rect 3341 1071 3375 1105
rect 213 697 247 731
rect 29 527 63 561
rect 121 527 155 561
rect 673 697 707 731
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 213 357 247 391
rect 1041 697 1075 731
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 673 357 707 391
rect 1501 697 1535 731
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1041 357 1075 391
rect 1869 697 1903 731
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1501 357 1535 391
rect 2329 697 2363 731
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 1869 357 1903 391
rect 2697 697 2731 731
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2329 357 2363 391
rect 3157 697 3191 731
rect 2789 527 2823 561
rect 2881 527 2915 561
rect 2973 527 3007 561
rect 3065 527 3099 561
rect 2697 357 2731 391
rect 3249 527 3283 561
rect 3341 527 3375 561
rect 3157 357 3191 391
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
rect 2881 -17 2915 17
rect 2973 -17 3007 17
rect 3065 -17 3099 17
rect 3157 -17 3191 17
rect 3249 -17 3283 17
rect 3341 -17 3375 17
<< metal1 >>
rect 0 1105 3404 1136
rect 0 1071 29 1105
rect 63 1071 121 1105
rect 155 1071 213 1105
rect 247 1071 305 1105
rect 339 1071 397 1105
rect 431 1071 489 1105
rect 523 1071 581 1105
rect 615 1071 673 1105
rect 707 1071 765 1105
rect 799 1071 857 1105
rect 891 1071 949 1105
rect 983 1071 1041 1105
rect 1075 1071 1133 1105
rect 1167 1071 1225 1105
rect 1259 1071 1317 1105
rect 1351 1071 1409 1105
rect 1443 1071 1501 1105
rect 1535 1071 1593 1105
rect 1627 1071 1685 1105
rect 1719 1071 1777 1105
rect 1811 1071 1869 1105
rect 1903 1071 1961 1105
rect 1995 1071 2053 1105
rect 2087 1071 2145 1105
rect 2179 1071 2237 1105
rect 2271 1071 2329 1105
rect 2363 1071 2421 1105
rect 2455 1071 2513 1105
rect 2547 1071 2605 1105
rect 2639 1071 2697 1105
rect 2731 1071 2789 1105
rect 2823 1071 2881 1105
rect 2915 1071 2973 1105
rect 3007 1071 3065 1105
rect 3099 1071 3157 1105
rect 3191 1071 3249 1105
rect 3283 1071 3341 1105
rect 3375 1071 3404 1105
rect 0 1040 3404 1071
rect 201 731 259 737
rect 201 697 213 731
rect 247 728 259 731
rect 661 731 719 737
rect 661 728 673 731
rect 247 700 673 728
rect 247 697 259 700
rect 201 691 259 697
rect 661 697 673 700
rect 707 728 719 731
rect 1029 731 1087 737
rect 1029 728 1041 731
rect 707 700 1041 728
rect 707 697 719 700
rect 661 691 719 697
rect 1029 697 1041 700
rect 1075 728 1087 731
rect 1489 731 1547 737
rect 1489 728 1501 731
rect 1075 700 1501 728
rect 1075 697 1087 700
rect 1029 691 1087 697
rect 1489 697 1501 700
rect 1535 728 1547 731
rect 1857 731 1915 737
rect 1857 728 1869 731
rect 1535 700 1869 728
rect 1535 697 1547 700
rect 1489 691 1547 697
rect 1857 697 1869 700
rect 1903 728 1915 731
rect 2317 731 2375 737
rect 2317 728 2329 731
rect 1903 700 2329 728
rect 1903 697 1915 700
rect 1857 691 1915 697
rect 2317 697 2329 700
rect 2363 728 2375 731
rect 2685 731 2743 737
rect 2685 728 2697 731
rect 2363 700 2697 728
rect 2363 697 2375 700
rect 2317 691 2375 697
rect 2685 697 2697 700
rect 2731 728 2743 731
rect 3145 731 3203 737
rect 3145 728 3157 731
rect 2731 700 3157 728
rect 2731 697 2743 700
rect 2685 691 2743 697
rect 3145 697 3157 700
rect 3191 697 3203 731
rect 3145 691 3203 697
rect 0 561 3404 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3249 561
rect 3283 527 3341 561
rect 3375 527 3404 561
rect 0 496 3404 527
rect 201 391 259 397
rect 201 357 213 391
rect 247 388 259 391
rect 661 391 719 397
rect 661 388 673 391
rect 247 360 673 388
rect 247 357 259 360
rect 201 351 259 357
rect 661 357 673 360
rect 707 388 719 391
rect 1029 391 1087 397
rect 1029 388 1041 391
rect 707 360 1041 388
rect 707 357 719 360
rect 661 351 719 357
rect 1029 357 1041 360
rect 1075 388 1087 391
rect 1489 391 1547 397
rect 1489 388 1501 391
rect 1075 360 1501 388
rect 1075 357 1087 360
rect 1029 351 1087 357
rect 1489 357 1501 360
rect 1535 388 1547 391
rect 1857 391 1915 397
rect 1857 388 1869 391
rect 1535 360 1869 388
rect 1535 357 1547 360
rect 1489 351 1547 357
rect 1857 357 1869 360
rect 1903 388 1915 391
rect 2317 391 2375 397
rect 2317 388 2329 391
rect 1903 360 2329 388
rect 1903 357 1915 360
rect 1857 351 1915 357
rect 2317 357 2329 360
rect 2363 388 2375 391
rect 2685 391 2743 397
rect 2685 388 2697 391
rect 2363 360 2697 388
rect 2363 357 2375 360
rect 2317 351 2375 357
rect 2685 357 2697 360
rect 2731 388 2743 391
rect 3145 391 3203 397
rect 3145 388 3157 391
rect 2731 360 3157 388
rect 2731 357 2743 360
rect 2685 351 2743 357
rect 3145 357 3157 360
rect 3191 357 3203 391
rect 3145 351 3203 357
rect 0 17 3404 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3341 17
rect 3375 -17 3404 17
rect 0 -48 3404 -17
<< labels >>
rlabel locali s 112 125 146 211 6 D[0]
port 1 nsew signal input
rlabel locali s 112 79 167 125 6 D[0]
port 1 nsew signal input
rlabel locali s 67 211 146 265 6 D[0]
port 1 nsew signal input
rlabel locali s 774 211 853 265 6 D[1]
port 2 nsew signal input
rlabel locali s 774 125 808 211 6 D[1]
port 2 nsew signal input
rlabel locali s 753 79 808 125 6 D[1]
port 2 nsew signal input
rlabel locali s 940 125 974 211 6 D[2]
port 3 nsew signal input
rlabel locali s 940 79 995 125 6 D[2]
port 3 nsew signal input
rlabel locali s 895 211 974 265 6 D[2]
port 3 nsew signal input
rlabel locali s 1602 211 1681 265 6 D[3]
port 4 nsew signal input
rlabel locali s 1602 125 1636 211 6 D[3]
port 4 nsew signal input
rlabel locali s 1581 79 1636 125 6 D[3]
port 4 nsew signal input
rlabel locali s 1768 125 1802 211 6 D[4]
port 5 nsew signal input
rlabel locali s 1768 79 1823 125 6 D[4]
port 5 nsew signal input
rlabel locali s 1723 211 1802 265 6 D[4]
port 5 nsew signal input
rlabel locali s 2430 211 2509 265 6 D[5]
port 6 nsew signal input
rlabel locali s 2430 125 2464 211 6 D[5]
port 6 nsew signal input
rlabel locali s 2409 79 2464 125 6 D[5]
port 6 nsew signal input
rlabel locali s 2596 125 2630 211 6 D[6]
port 7 nsew signal input
rlabel locali s 2596 79 2651 125 6 D[6]
port 7 nsew signal input
rlabel locali s 2551 211 2630 265 6 D[6]
port 7 nsew signal input
rlabel locali s 3258 211 3337 265 6 D[7]
port 8 nsew signal input
rlabel locali s 3258 125 3292 211 6 D[7]
port 8 nsew signal input
rlabel locali s 3237 79 3292 125 6 D[7]
port 8 nsew signal input
rlabel locali s 112 963 167 1009 6 D[8]
port 9 nsew signal input
rlabel locali s 112 877 146 963 6 D[8]
port 9 nsew signal input
rlabel locali s 67 823 146 877 6 D[8]
port 9 nsew signal input
rlabel locali s 774 877 808 963 6 D[9]
port 10 nsew signal input
rlabel locali s 774 823 853 877 6 D[9]
port 10 nsew signal input
rlabel locali s 753 963 808 1009 6 D[9]
port 10 nsew signal input
rlabel locali s 940 963 995 1009 6 D[10]
port 11 nsew signal input
rlabel locali s 940 877 974 963 6 D[10]
port 11 nsew signal input
rlabel locali s 895 823 974 877 6 D[10]
port 11 nsew signal input
rlabel locali s 1602 877 1636 963 6 D[11]
port 12 nsew signal input
rlabel locali s 1602 823 1681 877 6 D[11]
port 12 nsew signal input
rlabel locali s 1581 963 1636 1009 6 D[11]
port 12 nsew signal input
rlabel locali s 1768 963 1823 1009 6 D[12]
port 13 nsew signal input
rlabel locali s 1768 877 1802 963 6 D[12]
port 13 nsew signal input
rlabel locali s 1723 823 1802 877 6 D[12]
port 13 nsew signal input
rlabel locali s 2430 877 2464 963 6 D[13]
port 14 nsew signal input
rlabel locali s 2430 823 2509 877 6 D[13]
port 14 nsew signal input
rlabel locali s 2409 963 2464 1009 6 D[13]
port 14 nsew signal input
rlabel locali s 2596 963 2651 1009 6 D[14]
port 15 nsew signal input
rlabel locali s 2596 877 2630 963 6 D[14]
port 15 nsew signal input
rlabel locali s 2551 823 2630 877 6 D[14]
port 15 nsew signal input
rlabel locali s 3258 877 3292 963 6 D[15]
port 16 nsew signal input
rlabel locali s 3258 823 3337 877 6 D[15]
port 16 nsew signal input
rlabel locali s 3237 963 3292 1009 6 D[15]
port 16 nsew signal input
rlabel locali s 361 189 441 259 6 S[0]
port 17 nsew signal input
rlabel locali s 479 189 559 259 6 S[1]
port 18 nsew signal input
rlabel locali s 1189 189 1269 259 6 S[2]
port 19 nsew signal input
rlabel locali s 1307 189 1387 259 6 S[3]
port 20 nsew signal input
rlabel locali s 2017 189 2097 259 6 S[4]
port 21 nsew signal input
rlabel locali s 2135 189 2215 259 6 S[5]
port 22 nsew signal input
rlabel locali s 2845 189 2925 259 6 S[6]
port 23 nsew signal input
rlabel locali s 2963 189 3043 259 6 S[7]
port 24 nsew signal input
rlabel locali s 361 829 441 899 6 S[8]
port 25 nsew signal input
rlabel locali s 479 829 559 899 6 S[9]
port 26 nsew signal input
rlabel locali s 1189 829 1269 899 6 S[10]
port 27 nsew signal input
rlabel locali s 1307 829 1387 899 6 S[11]
port 28 nsew signal input
rlabel locali s 2017 829 2097 899 6 S[12]
port 29 nsew signal input
rlabel locali s 2135 829 2215 899 6 S[13]
port 30 nsew signal input
rlabel locali s 2845 829 2925 899 6 S[14]
port 31 nsew signal input
rlabel locali s 2963 829 3043 899 6 S[15]
port 32 nsew signal input
rlabel metal1 s 3145 728 3203 737 6 Z
port 33 nsew signal output
rlabel metal1 s 3145 691 3203 700 6 Z
port 33 nsew signal output
rlabel metal1 s 3145 388 3203 397 6 Z
port 33 nsew signal output
rlabel metal1 s 3145 351 3203 360 6 Z
port 33 nsew signal output
rlabel metal1 s 2685 728 2743 737 6 Z
port 33 nsew signal output
rlabel metal1 s 2685 691 2743 700 6 Z
port 33 nsew signal output
rlabel metal1 s 2685 388 2743 397 6 Z
port 33 nsew signal output
rlabel metal1 s 2685 351 2743 360 6 Z
port 33 nsew signal output
rlabel metal1 s 2317 728 2375 737 6 Z
port 33 nsew signal output
rlabel metal1 s 2317 691 2375 700 6 Z
port 33 nsew signal output
rlabel metal1 s 2317 388 2375 397 6 Z
port 33 nsew signal output
rlabel metal1 s 2317 351 2375 360 6 Z
port 33 nsew signal output
rlabel metal1 s 1857 728 1915 737 6 Z
port 33 nsew signal output
rlabel metal1 s 1857 691 1915 700 6 Z
port 33 nsew signal output
rlabel metal1 s 1857 388 1915 397 6 Z
port 33 nsew signal output
rlabel metal1 s 1857 351 1915 360 6 Z
port 33 nsew signal output
rlabel metal1 s 1489 728 1547 737 6 Z
port 33 nsew signal output
rlabel metal1 s 1489 691 1547 700 6 Z
port 33 nsew signal output
rlabel metal1 s 1489 388 1547 397 6 Z
port 33 nsew signal output
rlabel metal1 s 1489 351 1547 360 6 Z
port 33 nsew signal output
rlabel metal1 s 1029 728 1087 737 6 Z
port 33 nsew signal output
rlabel metal1 s 1029 691 1087 700 6 Z
port 33 nsew signal output
rlabel metal1 s 1029 388 1087 397 6 Z
port 33 nsew signal output
rlabel metal1 s 1029 351 1087 360 6 Z
port 33 nsew signal output
rlabel metal1 s 661 728 719 737 6 Z
port 33 nsew signal output
rlabel metal1 s 661 691 719 700 6 Z
port 33 nsew signal output
rlabel metal1 s 661 388 719 397 6 Z
port 33 nsew signal output
rlabel metal1 s 661 351 719 360 6 Z
port 33 nsew signal output
rlabel metal1 s 201 728 259 737 6 Z
port 33 nsew signal output
rlabel metal1 s 201 700 3203 728 6 Z
port 33 nsew signal output
rlabel metal1 s 201 691 259 700 6 Z
port 33 nsew signal output
rlabel metal1 s 201 388 259 397 6 Z
port 33 nsew signal output
rlabel metal1 s 201 360 3203 388 6 Z
port 33 nsew signal output
rlabel metal1 s 201 351 259 360 6 Z
port 33 nsew signal output
rlabel metal1 s 0 1040 3404 1136 6 VGND
port 34 nsew ground bidirectional
rlabel metal1 s 0 -48 3404 48 8 VGND
port 34 nsew ground bidirectional
rlabel metal1 s 0 496 3404 592 6 VPWR
port 35 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 3404 1088
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3026090
string GDS_START 2964356
<< end >>
