magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 17 364 87 596
rect 17 226 51 364
rect 317 290 367 356
rect 409 290 551 356
rect 17 87 215 226
rect 165 69 215 87
rect 409 114 455 134
rect 409 51 575 114
rect 677 51 743 134
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 127 364 177 649
rect 271 424 337 596
rect 377 458 417 649
rect 457 424 523 596
rect 271 390 523 424
rect 85 280 283 330
rect 249 256 283 280
rect 625 256 708 596
rect 249 222 708 256
rect 456 216 708 222
rect 251 17 341 188
rect 456 168 522 216
rect 556 148 643 182
rect 609 17 643 148
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel locali s 409 290 551 356 6 A1
port 1 nsew signal input
rlabel locali s 317 290 367 356 6 A2
port 2 nsew signal input
rlabel locali s 409 114 455 134 6 B1
port 3 nsew signal input
rlabel locali s 409 51 575 114 6 B1
port 3 nsew signal input
rlabel locali s 677 51 743 134 6 C1
port 4 nsew signal input
rlabel locali s 165 69 215 87 6 X
port 5 nsew signal output
rlabel locali s 17 364 87 596 6 X
port 5 nsew signal output
rlabel locali s 17 226 51 364 6 X
port 5 nsew signal output
rlabel locali s 17 87 215 226 6 X
port 5 nsew signal output
rlabel metal1 s 0 -49 768 49 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 617 768 715 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3931658
string GDS_START 3924508
<< end >>
