magic
tech sky130A
magscale 1 2
timestamp 1604502697
<< nwell >>
rect -38 261 1326 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 288 47 318 131
rect 384 47 414 131
rect 480 47 510 131
rect 576 47 606 131
rect 672 47 702 131
rect 778 47 808 131
rect 884 47 914 131
rect 990 47 1020 131
<< pmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 270 297 306 497
rect 364 297 400 497
rect 458 297 494 497
rect 552 297 588 497
rect 646 297 682 497
rect 740 297 776 497
rect 844 297 880 497
rect 948 297 984 497
rect 1052 297 1088 497
rect 1146 297 1182 497
<< ndiff >>
rect 235 95 288 131
rect 235 61 243 95
rect 277 61 288 95
rect 235 47 288 61
rect 318 106 384 131
rect 318 72 339 106
rect 373 72 384 106
rect 318 47 384 72
rect 414 95 480 131
rect 414 61 435 95
rect 469 61 480 95
rect 414 47 480 61
rect 510 106 576 131
rect 510 72 531 106
rect 565 72 576 106
rect 510 47 576 72
rect 606 95 672 131
rect 606 61 627 95
rect 661 61 672 95
rect 606 47 672 61
rect 702 106 778 131
rect 702 72 723 106
rect 757 72 778 106
rect 702 47 778 72
rect 808 95 884 131
rect 808 61 829 95
rect 863 61 884 95
rect 808 47 884 61
rect 914 106 990 131
rect 914 72 935 106
rect 969 72 990 106
rect 914 47 990 72
rect 1020 95 1093 131
rect 1020 61 1041 95
rect 1075 61 1093 95
rect 1020 47 1093 61
<< pdiff >>
rect 27 478 81 497
rect 27 444 35 478
rect 69 444 81 478
rect 27 410 81 444
rect 27 376 35 410
rect 69 376 81 410
rect 27 297 81 376
rect 117 471 175 497
rect 117 437 129 471
rect 163 437 175 471
rect 117 403 175 437
rect 117 369 129 403
rect 163 369 175 403
rect 117 297 175 369
rect 211 478 270 497
rect 211 444 224 478
rect 258 444 270 478
rect 211 410 270 444
rect 211 376 224 410
rect 258 376 270 410
rect 211 297 270 376
rect 306 471 364 497
rect 306 437 318 471
rect 352 437 364 471
rect 306 383 364 437
rect 306 349 318 383
rect 352 349 364 383
rect 306 297 364 349
rect 400 478 458 497
rect 400 444 412 478
rect 446 444 458 478
rect 400 410 458 444
rect 400 376 412 410
rect 446 376 458 410
rect 400 297 458 376
rect 494 471 552 497
rect 494 437 506 471
rect 540 437 552 471
rect 494 383 552 437
rect 494 349 506 383
rect 540 349 552 383
rect 494 297 552 349
rect 588 478 646 497
rect 588 444 600 478
rect 634 444 646 478
rect 588 410 646 444
rect 588 376 600 410
rect 634 376 646 410
rect 588 297 646 376
rect 682 471 740 497
rect 682 437 694 471
rect 728 437 740 471
rect 682 383 740 437
rect 682 349 694 383
rect 728 349 740 383
rect 682 297 740 349
rect 776 478 844 497
rect 776 444 788 478
rect 822 444 844 478
rect 776 410 844 444
rect 776 376 788 410
rect 822 376 844 410
rect 776 297 844 376
rect 880 471 948 497
rect 880 437 892 471
rect 926 437 948 471
rect 880 383 948 437
rect 880 349 892 383
rect 926 349 948 383
rect 880 297 948 349
rect 984 478 1052 497
rect 984 444 996 478
rect 1030 444 1052 478
rect 984 410 1052 444
rect 984 376 996 410
rect 1030 376 1052 410
rect 984 297 1052 376
rect 1088 471 1146 497
rect 1088 437 1100 471
rect 1134 437 1146 471
rect 1088 383 1146 437
rect 1088 349 1100 383
rect 1134 349 1146 383
rect 1088 297 1146 349
rect 1182 478 1236 497
rect 1182 444 1194 478
rect 1228 444 1236 478
rect 1182 410 1236 444
rect 1182 376 1194 410
rect 1228 376 1236 410
rect 1182 297 1236 376
<< ndiffc >>
rect 243 61 277 95
rect 339 72 373 106
rect 435 61 469 95
rect 531 72 565 106
rect 627 61 661 95
rect 723 72 757 106
rect 829 61 863 95
rect 935 72 969 106
rect 1041 61 1075 95
<< pdiffc >>
rect 35 444 69 478
rect 35 376 69 410
rect 129 437 163 471
rect 129 369 163 403
rect 224 444 258 478
rect 224 376 258 410
rect 318 437 352 471
rect 318 349 352 383
rect 412 444 446 478
rect 412 376 446 410
rect 506 437 540 471
rect 506 349 540 383
rect 600 444 634 478
rect 600 376 634 410
rect 694 437 728 471
rect 694 349 728 383
rect 788 444 822 478
rect 788 376 822 410
rect 892 437 926 471
rect 892 349 926 383
rect 996 444 1030 478
rect 996 376 1030 410
rect 1100 437 1134 471
rect 1100 349 1134 383
rect 1194 444 1228 478
rect 1194 376 1228 410
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 270 497 306 523
rect 364 497 400 523
rect 458 497 494 523
rect 552 497 588 523
rect 646 497 682 523
rect 740 497 776 523
rect 844 497 880 523
rect 948 497 984 523
rect 1052 497 1088 523
rect 1146 497 1182 523
rect 81 282 117 297
rect 175 282 211 297
rect 270 282 306 297
rect 364 282 400 297
rect 458 282 494 297
rect 552 282 588 297
rect 646 282 682 297
rect 740 282 776 297
rect 844 282 880 297
rect 948 282 984 297
rect 1052 282 1088 297
rect 1146 282 1182 297
rect 79 277 119 282
rect 173 277 213 282
rect 268 277 308 282
rect 362 277 402 282
rect 456 277 496 282
rect 550 277 590 282
rect 644 277 684 282
rect 738 277 778 282
rect 842 277 882 282
rect 946 277 986 282
rect 1050 277 1090 282
rect 1144 277 1184 282
rect 79 249 1184 277
rect 79 215 107 249
rect 141 215 185 249
rect 219 215 263 249
rect 297 215 341 249
rect 375 215 419 249
rect 453 215 497 249
rect 531 215 565 249
rect 599 215 643 249
rect 677 215 721 249
rect 755 215 799 249
rect 833 215 887 249
rect 921 215 965 249
rect 999 215 1053 249
rect 1087 215 1184 249
rect 79 162 1184 215
rect 288 131 318 162
rect 384 131 414 162
rect 480 131 510 162
rect 576 131 606 162
rect 672 131 702 162
rect 778 131 808 162
rect 884 131 914 162
rect 990 131 1020 162
rect 288 21 318 47
rect 384 21 414 47
rect 480 21 510 47
rect 576 21 606 47
rect 672 21 702 47
rect 778 21 808 47
rect 884 21 914 47
rect 990 21 1020 47
<< polycont >>
rect 107 215 141 249
rect 185 215 219 249
rect 263 215 297 249
rect 341 215 375 249
rect 419 215 453 249
rect 497 215 531 249
rect 565 215 599 249
rect 643 215 677 249
rect 721 215 755 249
rect 799 215 833 249
rect 887 215 921 249
rect 965 215 999 249
rect 1053 215 1087 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 27 478 79 527
rect 27 444 35 478
rect 69 444 79 478
rect 27 410 79 444
rect 27 376 35 410
rect 69 376 79 410
rect 27 360 79 376
rect 123 471 171 487
rect 123 437 129 471
rect 163 437 171 471
rect 123 403 171 437
rect 123 369 129 403
rect 163 369 171 403
rect 123 326 171 369
rect 215 478 267 527
rect 215 444 224 478
rect 258 444 267 478
rect 215 410 267 444
rect 215 376 224 410
rect 258 376 267 410
rect 215 360 267 376
rect 311 471 359 487
rect 311 437 318 471
rect 352 437 359 471
rect 311 383 359 437
rect 311 349 318 383
rect 352 349 359 383
rect 403 478 455 527
rect 403 444 412 478
rect 446 444 455 478
rect 403 410 455 444
rect 403 376 412 410
rect 446 376 455 410
rect 403 360 455 376
rect 499 471 549 487
rect 499 437 506 471
rect 540 437 549 471
rect 499 383 549 437
rect 311 326 359 349
rect 499 349 506 383
rect 540 349 549 383
rect 593 478 642 527
rect 593 444 600 478
rect 634 444 642 478
rect 593 410 642 444
rect 593 376 600 410
rect 634 376 642 410
rect 593 360 642 376
rect 686 471 735 487
rect 686 437 694 471
rect 728 437 735 471
rect 686 383 735 437
rect 499 326 549 349
rect 686 349 694 383
rect 728 349 735 383
rect 779 478 840 527
rect 779 444 788 478
rect 822 444 840 478
rect 779 410 840 444
rect 779 376 788 410
rect 822 376 840 410
rect 779 360 840 376
rect 884 471 945 487
rect 884 437 892 471
rect 926 437 945 471
rect 884 383 945 437
rect 686 326 735 349
rect 884 349 892 383
rect 926 349 945 383
rect 989 478 1049 527
rect 989 444 996 478
rect 1030 444 1049 478
rect 989 410 1049 444
rect 989 376 996 410
rect 1030 376 1049 410
rect 989 360 1049 376
rect 1093 471 1141 487
rect 1093 437 1100 471
rect 1134 437 1141 471
rect 1093 383 1141 437
rect 884 326 945 349
rect 1093 349 1100 383
rect 1134 349 1141 383
rect 1185 478 1236 527
rect 1185 444 1194 478
rect 1228 444 1236 478
rect 1185 410 1236 444
rect 1185 376 1194 410
rect 1228 376 1236 410
rect 1185 360 1236 376
rect 1093 326 1141 349
rect 23 292 1266 326
rect 23 173 57 292
rect 91 249 1113 258
rect 91 215 107 249
rect 141 215 185 249
rect 219 215 263 249
rect 297 215 341 249
rect 375 215 419 249
rect 453 215 497 249
rect 531 215 565 249
rect 599 215 643 249
rect 677 215 721 249
rect 755 215 799 249
rect 833 215 887 249
rect 921 215 965 249
rect 999 215 1053 249
rect 1087 215 1113 249
rect 91 207 1113 215
rect 1212 173 1266 292
rect 23 139 1266 173
rect 337 106 375 139
rect 227 95 293 105
rect 227 61 243 95
rect 277 61 293 95
rect 227 17 293 61
rect 337 72 339 106
rect 373 72 375 106
rect 529 106 567 139
rect 337 56 375 72
rect 419 95 485 105
rect 419 61 435 95
rect 469 61 485 95
rect 419 17 485 61
rect 529 72 531 106
rect 565 72 567 106
rect 721 106 759 139
rect 529 56 567 72
rect 611 95 687 105
rect 611 61 627 95
rect 661 61 687 95
rect 611 17 687 61
rect 721 72 723 106
rect 757 72 759 106
rect 933 106 971 139
rect 721 56 759 72
rect 803 95 889 105
rect 803 61 829 95
rect 863 61 889 95
rect 803 17 889 61
rect 933 72 935 106
rect 969 72 971 106
rect 933 56 971 72
rect 1015 95 1101 105
rect 1015 61 1041 95
rect 1075 61 1101 95
rect 1015 17 1101 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
flabel corelocali s 1220 289 1254 323 0 FreeSans 400 0 0 0 Y
port 6 nsew
flabel corelocali s 1220 221 1254 255 0 FreeSans 400 0 0 0 Y
port 6 nsew
flabel corelocali s 1220 153 1254 187 0 FreeSans 400 0 0 0 Y
port 6 nsew
flabel corelocali s 507 238 507 238 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 415 238 415 238 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 323 238 323 238 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 231 238 231 238 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 856 221 890 255 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 762 221 796 255 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 673 221 707 255 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 599 238 599 238 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 132 221 166 255 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew
rlabel comment s 0 0 0 0 4 clkinv_8
<< properties >>
string FIXED_BBOX 0 0 1288 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1817926
string GDS_START 1808192
<< end >>
