magic
tech sky130A
magscale 1 2
timestamp 1604502729
<< locali >>
rect 112 378 178 547
rect 292 378 358 547
rect 472 378 538 547
rect 652 378 718 547
rect 112 344 839 378
rect 741 310 839 344
rect 82 236 692 310
rect 741 202 775 310
rect 125 168 775 202
rect 125 123 175 168
rect 309 123 375 168
rect 509 123 575 168
rect 709 119 775 168
rect 1687 282 1753 310
rect 1687 236 1799 282
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 22 581 792 615
rect 22 364 75 581
rect 214 412 255 581
rect 394 412 438 581
rect 575 412 615 581
rect 758 446 792 581
rect 832 480 898 649
rect 938 446 988 596
rect 758 412 988 446
rect 938 344 988 412
rect 1028 378 1062 649
rect 1102 344 1152 596
rect 1192 378 1242 649
rect 1282 344 1332 596
rect 1372 378 1422 649
rect 1462 344 1512 596
rect 1647 593 1713 596
rect 938 310 1512 344
rect 1555 364 1713 593
rect 1753 364 1803 649
rect 1555 323 1645 364
rect 23 85 89 202
rect 209 85 275 134
rect 409 85 475 134
rect 609 85 675 134
rect 811 242 1577 276
rect 811 85 845 242
rect 23 51 845 85
rect 881 17 947 208
rect 981 70 1031 242
rect 1067 17 1133 208
rect 1169 70 1203 242
rect 1239 17 1305 208
rect 1341 70 1391 242
rect 1425 17 1491 208
rect 1527 70 1577 242
rect 1611 202 1645 323
rect 1611 70 1701 202
rect 1735 17 1787 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
<< metal1 >>
rect 0 683 1824 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 0 617 1824 649
rect 0 17 1824 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
rect 0 -49 1824 -17
<< labels >>
rlabel locali s 82 236 692 310 6 A
port 1 nsew signal input
rlabel locali s 1687 282 1753 310 6 TE
port 2 nsew signal input
rlabel locali s 1687 236 1799 282 6 TE
port 2 nsew signal input
rlabel locali s 741 310 839 344 6 Z
port 3 nsew signal output
rlabel locali s 741 202 775 310 6 Z
port 3 nsew signal output
rlabel locali s 709 119 775 168 6 Z
port 3 nsew signal output
rlabel locali s 652 378 718 547 6 Z
port 3 nsew signal output
rlabel locali s 509 123 575 168 6 Z
port 3 nsew signal output
rlabel locali s 472 378 538 547 6 Z
port 3 nsew signal output
rlabel locali s 309 123 375 168 6 Z
port 3 nsew signal output
rlabel locali s 292 378 358 547 6 Z
port 3 nsew signal output
rlabel locali s 125 168 775 202 6 Z
port 3 nsew signal output
rlabel locali s 125 123 175 168 6 Z
port 3 nsew signal output
rlabel locali s 112 378 178 547 6 Z
port 3 nsew signal output
rlabel locali s 112 344 839 378 6 Z
port 3 nsew signal output
rlabel metal1 s 0 -49 1824 49 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 617 1824 715 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1824 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 2481548
string GDS_START 2467228
<< end >>
