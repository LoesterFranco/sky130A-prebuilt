magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 2054 704
<< pwell >>
rect 0 0 2016 49
<< scnmos >>
rect 84 74 114 222
rect 184 74 214 222
rect 270 74 300 222
rect 356 74 386 222
rect 442 74 472 222
rect 528 74 558 222
rect 614 74 644 222
rect 700 74 730 222
rect 898 74 928 222
rect 984 74 1014 222
rect 1070 74 1100 222
rect 1156 74 1186 222
rect 1256 74 1286 222
rect 1356 74 1386 222
rect 1442 74 1472 222
rect 1528 74 1558 222
rect 1614 74 1644 222
rect 1714 74 1744 222
rect 1816 74 1846 222
rect 1902 74 1932 222
<< pmoshvt >>
rect 237 368 267 592
rect 347 368 377 592
rect 437 368 467 592
rect 611 368 641 592
rect 701 368 731 592
rect 811 368 841 592
rect 1237 368 1267 592
rect 1330 368 1360 592
rect 1420 368 1450 592
rect 1510 368 1540 592
rect 1603 368 1633 592
rect 1700 368 1730 592
rect 1800 368 1830 592
rect 1900 368 1930 592
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 207 184 222
rect 114 173 139 207
rect 173 173 184 207
rect 114 74 184 173
rect 214 120 270 222
rect 214 86 225 120
rect 259 86 270 120
rect 214 74 270 86
rect 300 199 356 222
rect 300 165 311 199
rect 345 165 356 199
rect 300 74 356 165
rect 386 210 442 222
rect 386 176 397 210
rect 431 176 442 210
rect 386 120 442 176
rect 386 86 397 120
rect 431 86 442 120
rect 386 74 442 86
rect 472 120 528 222
rect 472 86 483 120
rect 517 86 528 120
rect 472 74 528 86
rect 558 207 614 222
rect 558 173 569 207
rect 603 173 614 207
rect 558 74 614 173
rect 644 120 700 222
rect 644 86 655 120
rect 689 86 700 120
rect 644 74 700 86
rect 730 207 787 222
rect 730 173 741 207
rect 775 173 787 207
rect 730 74 787 173
rect 841 207 898 222
rect 841 173 853 207
rect 887 173 898 207
rect 841 74 898 173
rect 928 120 984 222
rect 928 86 939 120
rect 973 86 984 120
rect 928 74 984 86
rect 1014 207 1070 222
rect 1014 173 1025 207
rect 1059 173 1070 207
rect 1014 74 1070 173
rect 1100 120 1156 222
rect 1100 86 1111 120
rect 1145 86 1156 120
rect 1100 74 1156 86
rect 1186 210 1256 222
rect 1186 176 1211 210
rect 1245 176 1256 210
rect 1186 120 1256 176
rect 1186 86 1211 120
rect 1245 86 1256 120
rect 1186 74 1256 86
rect 1286 148 1356 222
rect 1286 114 1311 148
rect 1345 114 1356 148
rect 1286 74 1356 114
rect 1386 210 1442 222
rect 1386 176 1397 210
rect 1431 176 1442 210
rect 1386 120 1442 176
rect 1386 86 1397 120
rect 1431 86 1442 120
rect 1386 74 1442 86
rect 1472 148 1528 222
rect 1472 114 1483 148
rect 1517 114 1528 148
rect 1472 74 1528 114
rect 1558 210 1614 222
rect 1558 176 1569 210
rect 1603 176 1614 210
rect 1558 120 1614 176
rect 1558 86 1569 120
rect 1603 86 1614 120
rect 1558 74 1614 86
rect 1644 148 1714 222
rect 1644 114 1669 148
rect 1703 114 1714 148
rect 1644 74 1714 114
rect 1744 210 1816 222
rect 1744 176 1755 210
rect 1789 176 1816 210
rect 1744 120 1816 176
rect 1744 86 1755 120
rect 1789 86 1816 120
rect 1744 74 1816 86
rect 1846 148 1902 222
rect 1846 114 1857 148
rect 1891 114 1902 148
rect 1846 74 1902 114
rect 1932 210 1989 222
rect 1932 176 1943 210
rect 1977 176 1989 210
rect 1932 120 1989 176
rect 1932 86 1943 120
rect 1977 86 1989 120
rect 1932 74 1989 86
<< pdiff >>
rect 27 580 237 592
rect 27 546 39 580
rect 73 546 114 580
rect 148 546 190 580
rect 224 546 237 580
rect 27 497 237 546
rect 27 463 39 497
rect 73 463 114 497
rect 148 463 190 497
rect 224 463 237 497
rect 27 424 237 463
rect 27 390 39 424
rect 73 390 114 424
rect 148 390 190 424
rect 224 390 237 424
rect 27 368 237 390
rect 267 580 347 592
rect 267 546 290 580
rect 324 546 347 580
rect 267 508 347 546
rect 267 474 290 508
rect 324 474 347 508
rect 267 368 347 474
rect 377 580 437 592
rect 377 546 390 580
rect 424 546 437 580
rect 377 497 437 546
rect 377 463 390 497
rect 424 463 437 497
rect 377 414 437 463
rect 377 380 390 414
rect 424 380 437 414
rect 377 368 437 380
rect 467 580 611 592
rect 467 546 480 580
rect 514 546 564 580
rect 598 546 611 580
rect 467 478 611 546
rect 467 444 480 478
rect 514 444 564 478
rect 598 444 611 478
rect 467 368 611 444
rect 641 580 701 592
rect 641 546 654 580
rect 688 546 701 580
rect 641 497 701 546
rect 641 463 654 497
rect 688 463 701 497
rect 641 414 701 463
rect 641 380 654 414
rect 688 380 701 414
rect 641 368 701 380
rect 731 580 811 592
rect 731 546 754 580
rect 788 546 811 580
rect 731 508 811 546
rect 731 474 754 508
rect 788 474 811 508
rect 731 368 811 474
rect 841 580 900 592
rect 841 546 854 580
rect 888 546 900 580
rect 841 510 900 546
rect 841 476 854 510
rect 888 476 900 510
rect 841 440 900 476
rect 841 406 854 440
rect 888 406 900 440
rect 841 368 900 406
rect 954 580 1237 592
rect 954 546 972 580
rect 1006 546 1044 580
rect 1078 546 1117 580
rect 1151 546 1189 580
rect 1223 546 1237 580
rect 954 492 1237 546
rect 954 458 972 492
rect 1006 458 1044 492
rect 1078 458 1117 492
rect 1151 458 1189 492
rect 1223 458 1237 492
rect 954 368 1237 458
rect 1267 578 1330 592
rect 1267 544 1283 578
rect 1317 544 1330 578
rect 1267 368 1330 544
rect 1360 580 1420 592
rect 1360 546 1373 580
rect 1407 546 1420 580
rect 1360 508 1420 546
rect 1360 474 1373 508
rect 1407 474 1420 508
rect 1360 368 1420 474
rect 1450 578 1510 592
rect 1450 544 1463 578
rect 1497 544 1510 578
rect 1450 368 1510 544
rect 1540 580 1603 592
rect 1540 546 1553 580
rect 1587 546 1603 580
rect 1540 508 1603 546
rect 1540 474 1553 508
rect 1587 474 1603 508
rect 1540 368 1603 474
rect 1633 531 1700 592
rect 1633 497 1653 531
rect 1687 497 1700 531
rect 1633 440 1700 497
rect 1633 406 1653 440
rect 1687 406 1700 440
rect 1633 368 1700 406
rect 1730 580 1800 592
rect 1730 546 1753 580
rect 1787 546 1800 580
rect 1730 508 1800 546
rect 1730 474 1753 508
rect 1787 474 1800 508
rect 1730 368 1800 474
rect 1830 531 1900 592
rect 1830 497 1853 531
rect 1887 497 1900 531
rect 1830 440 1900 497
rect 1830 406 1853 440
rect 1887 406 1900 440
rect 1830 368 1900 406
rect 1930 580 1989 592
rect 1930 546 1943 580
rect 1977 546 1989 580
rect 1930 497 1989 546
rect 1930 463 1943 497
rect 1977 463 1989 497
rect 1930 414 1989 463
rect 1930 380 1943 414
rect 1977 380 1989 414
rect 1930 368 1989 380
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 139 173 173 207
rect 225 86 259 120
rect 311 165 345 199
rect 397 176 431 210
rect 397 86 431 120
rect 483 86 517 120
rect 569 173 603 207
rect 655 86 689 120
rect 741 173 775 207
rect 853 173 887 207
rect 939 86 973 120
rect 1025 173 1059 207
rect 1111 86 1145 120
rect 1211 176 1245 210
rect 1211 86 1245 120
rect 1311 114 1345 148
rect 1397 176 1431 210
rect 1397 86 1431 120
rect 1483 114 1517 148
rect 1569 176 1603 210
rect 1569 86 1603 120
rect 1669 114 1703 148
rect 1755 176 1789 210
rect 1755 86 1789 120
rect 1857 114 1891 148
rect 1943 176 1977 210
rect 1943 86 1977 120
<< pdiffc >>
rect 39 546 73 580
rect 114 546 148 580
rect 190 546 224 580
rect 39 463 73 497
rect 114 463 148 497
rect 190 463 224 497
rect 39 390 73 424
rect 114 390 148 424
rect 190 390 224 424
rect 290 546 324 580
rect 290 474 324 508
rect 390 546 424 580
rect 390 463 424 497
rect 390 380 424 414
rect 480 546 514 580
rect 564 546 598 580
rect 480 444 514 478
rect 564 444 598 478
rect 654 546 688 580
rect 654 463 688 497
rect 654 380 688 414
rect 754 546 788 580
rect 754 474 788 508
rect 854 546 888 580
rect 854 476 888 510
rect 854 406 888 440
rect 972 546 1006 580
rect 1044 546 1078 580
rect 1117 546 1151 580
rect 1189 546 1223 580
rect 972 458 1006 492
rect 1044 458 1078 492
rect 1117 458 1151 492
rect 1189 458 1223 492
rect 1283 544 1317 578
rect 1373 546 1407 580
rect 1373 474 1407 508
rect 1463 544 1497 578
rect 1553 546 1587 580
rect 1553 474 1587 508
rect 1653 497 1687 531
rect 1653 406 1687 440
rect 1753 546 1787 580
rect 1753 474 1787 508
rect 1853 497 1887 531
rect 1853 406 1887 440
rect 1943 546 1977 580
rect 1943 463 1977 497
rect 1943 380 1977 414
<< poly >>
rect 237 592 267 618
rect 347 592 377 618
rect 437 592 467 618
rect 611 592 641 618
rect 701 592 731 618
rect 811 592 841 618
rect 1237 592 1267 618
rect 1330 592 1360 618
rect 1420 592 1450 618
rect 1510 592 1540 618
rect 1603 592 1633 618
rect 1700 592 1730 618
rect 1800 592 1830 618
rect 1900 592 1930 618
rect 237 353 267 368
rect 347 353 377 368
rect 437 353 467 368
rect 611 353 641 368
rect 701 353 731 368
rect 811 353 841 368
rect 1237 353 1267 368
rect 1330 353 1360 368
rect 1420 353 1450 368
rect 1510 353 1540 368
rect 1603 353 1633 368
rect 1700 353 1730 368
rect 1800 353 1830 368
rect 1900 353 1930 368
rect 234 336 270 353
rect 68 331 270 336
rect 344 331 380 353
rect 68 320 380 331
rect 68 286 84 320
rect 118 286 152 320
rect 186 286 220 320
rect 254 286 380 320
rect 434 345 470 353
rect 608 345 644 353
rect 434 315 644 345
rect 698 345 734 353
rect 808 345 844 353
rect 698 320 1186 345
rect 698 315 914 320
rect 68 267 380 286
rect 442 310 644 315
rect 442 276 458 310
rect 492 276 526 310
rect 560 276 594 310
rect 628 276 644 310
rect 442 267 644 276
rect 898 286 914 315
rect 948 286 982 320
rect 1016 286 1050 320
rect 1084 286 1118 320
rect 1152 286 1186 320
rect 898 270 1186 286
rect 68 237 386 267
rect 84 222 114 237
rect 184 222 214 237
rect 270 222 300 237
rect 356 222 386 237
rect 442 237 730 267
rect 442 222 472 237
rect 528 222 558 237
rect 614 222 644 237
rect 700 222 730 237
rect 898 222 928 270
rect 984 222 1014 270
rect 1070 222 1100 270
rect 1156 222 1186 270
rect 1234 336 1270 353
rect 1327 336 1363 353
rect 1417 336 1453 353
rect 1507 336 1543 353
rect 1234 320 1543 336
rect 1234 286 1273 320
rect 1307 286 1341 320
rect 1375 286 1409 320
rect 1443 286 1477 320
rect 1511 294 1543 320
rect 1600 336 1636 353
rect 1697 336 1733 353
rect 1797 336 1933 353
rect 1600 320 1933 336
rect 1511 286 1558 294
rect 1234 264 1558 286
rect 1256 222 1286 264
rect 1356 222 1386 264
rect 1442 222 1472 264
rect 1528 222 1558 264
rect 1600 286 1660 320
rect 1694 286 1728 320
rect 1762 286 1796 320
rect 1830 286 1864 320
rect 1898 286 1933 320
rect 1600 275 1933 286
rect 1600 245 1932 275
rect 1614 222 1644 245
rect 1714 222 1744 245
rect 1816 222 1846 245
rect 1902 222 1932 245
rect 84 48 114 74
rect 184 48 214 74
rect 270 48 300 74
rect 356 48 386 74
rect 442 48 472 74
rect 528 48 558 74
rect 614 48 644 74
rect 700 48 730 74
rect 898 48 928 74
rect 984 48 1014 74
rect 1070 48 1100 74
rect 1156 48 1186 74
rect 1256 48 1286 74
rect 1356 48 1386 74
rect 1442 48 1472 74
rect 1528 48 1558 74
rect 1614 48 1644 74
rect 1714 48 1744 74
rect 1816 48 1846 74
rect 1902 48 1932 74
<< polycont >>
rect 84 286 118 320
rect 152 286 186 320
rect 220 286 254 320
rect 458 276 492 310
rect 526 276 560 310
rect 594 276 628 310
rect 914 286 948 320
rect 982 286 1016 320
rect 1050 286 1084 320
rect 1118 286 1152 320
rect 1273 286 1307 320
rect 1341 286 1375 320
rect 1409 286 1443 320
rect 1477 286 1511 320
rect 1660 286 1694 320
rect 1728 286 1762 320
rect 1796 286 1830 320
rect 1864 286 1898 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 23 580 240 596
rect 23 546 39 580
rect 73 546 114 580
rect 148 546 190 580
rect 224 546 240 580
rect 23 497 240 546
rect 23 463 39 497
rect 73 463 114 497
rect 148 463 190 497
rect 224 463 240 497
rect 23 424 240 463
rect 274 580 340 649
rect 274 546 290 580
rect 324 546 340 580
rect 274 508 340 546
rect 274 474 290 508
rect 324 474 340 508
rect 274 458 340 474
rect 374 580 440 596
rect 374 546 390 580
rect 424 546 440 580
rect 374 497 440 546
rect 374 463 390 497
rect 424 463 440 497
rect 374 424 440 463
rect 474 580 604 649
rect 474 546 480 580
rect 514 546 564 580
rect 598 546 604 580
rect 474 478 604 546
rect 474 444 480 478
rect 514 444 564 478
rect 598 444 604 478
rect 474 428 604 444
rect 638 580 704 596
rect 638 546 654 580
rect 688 546 704 580
rect 638 497 704 546
rect 638 463 654 497
rect 688 463 704 497
rect 23 390 39 424
rect 73 390 114 424
rect 148 390 190 424
rect 224 414 440 424
rect 224 390 390 414
rect 374 380 390 390
rect 424 394 440 414
rect 638 424 704 463
rect 738 580 804 649
rect 738 546 754 580
rect 788 546 804 580
rect 738 508 804 546
rect 738 474 754 508
rect 788 474 804 508
rect 738 458 804 474
rect 838 580 904 596
rect 838 546 854 580
rect 888 546 904 580
rect 838 510 904 546
rect 838 476 854 510
rect 888 476 904 510
rect 838 440 904 476
rect 950 580 1233 596
rect 950 546 972 580
rect 1006 546 1044 580
rect 1078 546 1117 580
rect 1151 546 1189 580
rect 1223 546 1233 580
rect 950 492 1233 546
rect 1267 578 1317 649
rect 1267 544 1283 578
rect 1267 526 1317 544
rect 1357 580 1423 596
rect 1357 546 1373 580
rect 1407 546 1423 580
rect 1357 508 1423 546
rect 1463 578 1497 649
rect 1463 526 1497 544
rect 1537 581 1993 615
rect 1537 580 1603 581
rect 1537 546 1553 580
rect 1587 546 1603 580
rect 1737 580 1803 581
rect 1357 492 1373 508
rect 950 458 972 492
rect 1006 458 1044 492
rect 1078 458 1117 492
rect 1151 458 1189 492
rect 1223 474 1373 492
rect 1407 492 1423 508
rect 1537 508 1603 546
rect 1537 492 1553 508
rect 1407 474 1553 492
rect 1587 474 1603 508
rect 1223 458 1603 474
rect 1637 531 1703 547
rect 1637 497 1653 531
rect 1687 497 1703 531
rect 838 424 854 440
rect 638 414 854 424
rect 638 394 654 414
rect 424 380 654 394
rect 688 406 854 414
rect 888 424 904 440
rect 1637 440 1703 497
rect 1737 546 1753 580
rect 1787 546 1803 580
rect 1943 580 1993 581
rect 1737 508 1803 546
rect 1737 474 1753 508
rect 1787 474 1803 508
rect 1737 458 1803 474
rect 1837 531 1903 547
rect 1837 497 1853 531
rect 1887 497 1903 531
rect 1637 424 1653 440
rect 888 406 1653 424
rect 1687 424 1703 440
rect 1837 440 1903 497
rect 1837 424 1853 440
rect 1687 406 1853 424
rect 1887 406 1903 440
rect 688 390 1903 406
rect 1977 546 1993 580
rect 1943 497 1993 546
rect 1977 463 1993 497
rect 1943 414 1993 463
rect 688 380 704 390
rect 374 360 704 380
rect 1977 380 1993 414
rect 1943 364 1993 380
rect 374 356 408 360
rect 25 320 270 356
rect 25 286 84 320
rect 118 286 152 320
rect 186 286 220 320
rect 254 286 270 320
rect 25 270 270 286
rect 313 310 408 356
rect 793 326 839 356
rect 442 310 839 326
rect 313 226 361 310
rect 442 276 458 310
rect 492 276 526 310
rect 560 276 594 310
rect 628 276 839 310
rect 442 260 839 276
rect 889 320 1223 356
rect 889 286 914 320
rect 948 286 982 320
rect 1016 286 1050 320
rect 1084 286 1118 320
rect 1152 286 1223 320
rect 889 270 1223 286
rect 1257 320 1527 356
rect 1257 286 1273 320
rect 1307 286 1341 320
rect 1375 286 1409 320
rect 1443 286 1477 320
rect 1511 286 1527 320
rect 1257 270 1527 286
rect 1561 320 1898 356
rect 1561 286 1660 320
rect 1694 286 1728 320
rect 1762 286 1796 320
rect 1830 286 1864 320
rect 1561 270 1898 286
rect 1009 226 1993 236
rect 23 210 89 226
rect 23 176 39 210
rect 73 176 89 210
rect 23 120 89 176
rect 123 207 361 226
rect 123 173 139 207
rect 173 199 361 207
rect 173 173 311 199
rect 123 165 311 173
rect 345 165 361 199
rect 123 154 361 165
rect 397 210 791 226
rect 431 207 791 210
rect 431 176 569 207
rect 397 173 569 176
rect 603 173 741 207
rect 775 173 791 207
rect 397 163 791 173
rect 837 210 1993 226
rect 837 207 1211 210
rect 837 173 853 207
rect 887 173 1025 207
rect 1059 176 1211 207
rect 1245 202 1397 210
rect 1245 176 1261 202
rect 1059 173 1261 176
rect 837 170 1261 173
rect 837 163 903 170
rect 397 120 431 163
rect 1095 129 1161 136
rect 23 86 39 120
rect 73 86 225 120
rect 259 86 397 120
rect 23 70 431 86
rect 467 120 1161 129
rect 467 86 483 120
rect 517 86 655 120
rect 689 86 939 120
rect 973 86 1111 120
rect 1145 86 1161 120
rect 467 70 1161 86
rect 1195 120 1261 170
rect 1431 202 1569 210
rect 1195 86 1211 120
rect 1245 86 1261 120
rect 1195 70 1261 86
rect 1295 148 1361 164
rect 1295 114 1311 148
rect 1345 114 1361 148
rect 1295 17 1361 114
rect 1397 120 1431 176
rect 1603 202 1755 210
rect 1603 176 1619 202
rect 1397 70 1431 86
rect 1467 148 1533 164
rect 1467 114 1483 148
rect 1517 114 1533 148
rect 1467 17 1533 114
rect 1569 120 1619 176
rect 1789 202 1943 210
rect 1789 176 1805 202
rect 1603 86 1619 120
rect 1569 70 1619 86
rect 1653 148 1719 164
rect 1653 114 1669 148
rect 1703 114 1719 148
rect 1653 17 1719 114
rect 1755 120 1805 176
rect 1977 176 1993 210
rect 1789 86 1805 120
rect 1755 70 1805 86
rect 1841 148 1907 164
rect 1841 114 1857 148
rect 1891 114 1907 148
rect 1841 17 1907 114
rect 1943 120 1993 176
rect 1977 86 1993 120
rect 1943 70 1993 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o2111ai_4
flabel pwell s 0 0 2016 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nwell s 0 617 2016 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 0 617 2016 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 2016 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 1087 316 1121 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 1183 316 1217 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 1279 316 1313 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 1375 316 1409 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 1471 316 1505 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 1567 316 1601 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 1663 316 1697 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 1759 316 1793 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 1855 316 1889 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 D1
port 5 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 D1
port 5 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 D1
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 2016 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1319026
string GDS_START 1303266
<< end >>
