magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1104 561
rect 103 427 169 527
rect 18 197 66 325
rect 103 17 169 93
rect 391 367 454 527
rect 292 191 358 265
rect 755 427 789 527
rect 939 314 980 527
rect 1030 334 1087 491
rect 1053 149 1087 334
rect 375 17 441 89
rect 737 17 803 106
rect 939 17 980 143
rect 1030 83 1087 149
rect 0 -17 1104 17
<< obsli1 >>
rect 35 393 69 493
rect 35 359 156 393
rect 122 323 156 359
rect 122 280 156 289
rect 203 391 248 493
rect 203 357 214 391
rect 203 337 248 357
rect 122 214 168 280
rect 122 161 156 214
rect 35 127 156 161
rect 35 69 69 127
rect 203 69 237 337
rect 291 333 357 483
rect 554 451 721 485
rect 585 391 653 399
rect 585 357 586 391
rect 620 357 653 391
rect 291 299 428 333
rect 394 219 428 299
rect 494 323 551 337
rect 528 289 551 323
rect 494 271 551 289
rect 585 315 653 357
rect 394 157 468 219
rect 585 207 619 315
rect 687 265 721 451
rect 859 373 903 487
rect 768 307 903 373
rect 869 265 903 307
rect 687 233 835 265
rect 307 153 468 157
rect 307 123 428 153
rect 543 141 619 207
rect 666 199 835 233
rect 869 199 1019 265
rect 307 69 341 123
rect 666 107 700 199
rect 869 149 903 199
rect 568 73 700 107
rect 859 83 903 149
<< obsli1c >>
rect 122 289 156 323
rect 214 357 248 391
rect 586 357 620 391
rect 494 289 528 323
<< metal1 >>
rect 0 496 1104 592
rect 0 -48 1104 48
<< obsm1 >>
rect 202 391 260 397
rect 202 357 214 391
rect 248 388 260 391
rect 574 391 632 397
rect 574 388 586 391
rect 248 360 586 388
rect 248 357 260 360
rect 202 351 260 357
rect 574 357 586 360
rect 620 357 632 391
rect 574 351 632 357
rect 110 323 168 329
rect 110 289 122 323
rect 156 320 168 323
rect 482 323 540 329
rect 482 320 494 323
rect 156 292 494 320
rect 156 289 168 292
rect 110 283 168 289
rect 482 289 494 292
rect 528 289 540 323
rect 482 283 540 289
<< labels >>
rlabel locali s 292 191 358 265 6 D
port 1 nsew signal input
rlabel locali s 1053 149 1087 334 6 Q
port 2 nsew signal output
rlabel locali s 1030 334 1087 491 6 Q
port 2 nsew signal output
rlabel locali s 1030 83 1087 149 6 Q
port 2 nsew signal output
rlabel locali s 18 197 66 325 6 GATE
port 3 nsew clock input
rlabel locali s 939 17 980 143 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 737 17 803 106 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 375 17 441 89 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 103 17 169 93 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 1104 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1104 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 939 314 980 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 755 427 789 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 391 367 454 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 103 427 169 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 1104 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 1104 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1104 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2806144
string GDS_START 2795994
<< end >>
