magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 920 561
rect 17 299 69 527
rect 103 299 169 493
rect 203 367 305 527
rect 203 299 237 367
rect 17 17 69 177
rect 103 176 158 299
rect 355 215 431 265
rect 465 215 531 468
rect 565 215 631 468
rect 665 215 731 467
rect 813 299 879 527
rect 765 215 903 265
rect 103 51 169 176
rect 203 17 252 177
rect 497 17 550 109
rect 701 17 755 109
rect 0 -17 920 17
<< obsli1 >>
rect 339 333 429 493
rect 271 299 429 333
rect 271 265 320 299
rect 192 215 320 265
rect 286 170 320 215
rect 286 51 357 170
rect 397 143 879 181
rect 397 51 463 143
rect 591 51 657 143
rect 813 51 879 143
<< metal1 >>
rect 0 496 920 592
rect 0 -48 920 48
<< labels >>
rlabel locali s 765 215 903 265 6 A1
port 1 nsew signal input
rlabel locali s 665 215 731 467 6 A2
port 2 nsew signal input
rlabel locali s 565 215 631 468 6 A3
port 3 nsew signal input
rlabel locali s 465 215 531 468 6 A4
port 4 nsew signal input
rlabel locali s 355 215 431 265 6 B1
port 5 nsew signal input
rlabel locali s 103 299 169 493 6 X
port 6 nsew signal output
rlabel locali s 103 176 158 299 6 X
port 6 nsew signal output
rlabel locali s 103 51 169 176 6 X
port 6 nsew signal output
rlabel locali s 701 17 755 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 497 17 550 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 203 17 252 177 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 17 17 69 177 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 920 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 920 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 813 299 879 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 203 367 305 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 203 299 237 367 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 17 299 69 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 920 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 920 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 920 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 871642
string GDS_START 862562
<< end >>
