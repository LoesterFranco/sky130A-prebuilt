magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 2430 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 79 47 109 131
rect 173 47 203 131
rect 375 47 405 131
rect 487 47 517 131
rect 585 47 615 131
rect 691 47 721 131
rect 767 47 797 131
rect 981 47 1011 119
rect 1097 47 1127 119
rect 1205 47 1235 131
rect 1361 47 1391 175
rect 1462 47 1492 119
rect 1595 47 1625 119
rect 1690 47 1720 131
rect 1898 47 1928 177
rect 1982 47 2012 177
rect 2076 47 2106 177
rect 2172 47 2202 177
rect 2276 47 2306 177
<< pmoshvt >>
rect 82 363 118 491
rect 176 363 212 491
rect 374 369 410 497
rect 468 369 504 497
rect 572 369 608 497
rect 666 369 702 497
rect 769 369 805 497
rect 982 413 1018 497
rect 1085 413 1121 497
rect 1191 413 1227 497
rect 1333 347 1369 497
rect 1438 413 1474 497
rect 1532 413 1568 497
rect 1669 413 1705 497
rect 1890 297 1926 497
rect 1984 297 2020 497
rect 2078 297 2114 497
rect 2174 297 2210 497
rect 2268 297 2304 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 173 131
rect 109 59 129 93
rect 163 59 173 93
rect 109 47 173 59
rect 203 119 265 131
rect 203 85 223 119
rect 257 85 265 119
rect 203 47 265 85
rect 319 89 375 131
rect 319 55 331 89
rect 365 55 375 89
rect 319 47 375 55
rect 405 89 487 131
rect 405 55 441 89
rect 475 55 487 89
rect 405 47 487 55
rect 517 47 585 131
rect 615 89 691 131
rect 615 55 636 89
rect 670 55 691 89
rect 615 47 691 55
rect 721 47 767 131
rect 797 89 869 131
rect 1301 131 1361 175
rect 1145 119 1205 131
rect 797 55 823 89
rect 857 55 869 89
rect 797 47 869 55
rect 925 107 981 119
rect 925 73 933 107
rect 967 73 981 107
rect 925 47 981 73
rect 1011 107 1097 119
rect 1011 73 1043 107
rect 1077 73 1097 107
rect 1011 47 1097 73
rect 1127 47 1205 119
rect 1235 101 1361 131
rect 1235 67 1279 101
rect 1313 67 1361 101
rect 1235 47 1361 67
rect 1391 119 1441 175
rect 1836 162 1898 177
rect 1640 119 1690 131
rect 1391 107 1462 119
rect 1391 73 1407 107
rect 1441 73 1462 107
rect 1391 47 1462 73
rect 1492 107 1595 119
rect 1492 73 1529 107
rect 1563 73 1595 107
rect 1492 47 1595 73
rect 1625 47 1690 119
rect 1720 107 1782 131
rect 1720 73 1740 107
rect 1774 73 1782 107
rect 1720 47 1782 73
rect 1836 128 1844 162
rect 1878 128 1898 162
rect 1836 94 1898 128
rect 1836 60 1844 94
rect 1878 60 1898 94
rect 1836 47 1898 60
rect 1928 123 1982 177
rect 1928 89 1938 123
rect 1972 89 1982 123
rect 1928 47 1982 89
rect 2012 164 2076 177
rect 2012 130 2032 164
rect 2066 130 2076 164
rect 2012 96 2076 130
rect 2012 62 2032 96
rect 2066 62 2076 96
rect 2012 47 2076 62
rect 2106 96 2172 177
rect 2106 62 2128 96
rect 2162 62 2172 96
rect 2106 47 2172 62
rect 2202 164 2276 177
rect 2202 130 2222 164
rect 2256 130 2276 164
rect 2202 96 2276 130
rect 2202 62 2222 96
rect 2256 62 2276 96
rect 2202 47 2276 62
rect 2306 96 2359 177
rect 2306 62 2316 96
rect 2350 62 2359 96
rect 2306 47 2359 62
<< pdiff >>
rect 28 477 82 491
rect 28 443 36 477
rect 70 443 82 477
rect 28 409 82 443
rect 28 375 36 409
rect 70 375 82 409
rect 28 363 82 375
rect 118 461 176 491
rect 118 427 130 461
rect 164 427 176 461
rect 118 363 176 427
rect 212 477 266 491
rect 212 443 224 477
rect 258 443 266 477
rect 212 409 266 443
rect 212 375 224 409
rect 258 375 266 409
rect 212 363 266 375
rect 320 452 374 497
rect 320 418 328 452
rect 362 418 374 452
rect 320 369 374 418
rect 410 483 468 497
rect 410 449 422 483
rect 456 449 468 483
rect 410 369 468 449
rect 504 369 572 497
rect 608 483 666 497
rect 608 449 620 483
rect 654 449 666 483
rect 608 369 666 449
rect 702 369 769 497
rect 805 483 864 497
rect 805 449 822 483
rect 856 449 864 483
rect 805 369 864 449
rect 918 472 982 497
rect 918 438 926 472
rect 960 438 982 472
rect 918 413 982 438
rect 1018 472 1085 497
rect 1018 438 1035 472
rect 1069 438 1085 472
rect 1018 413 1085 438
rect 1121 413 1191 497
rect 1227 485 1333 497
rect 1227 451 1287 485
rect 1321 451 1333 485
rect 1227 417 1333 451
rect 1227 413 1287 417
rect 1244 383 1287 413
rect 1321 383 1333 417
rect 1244 347 1333 383
rect 1369 477 1438 497
rect 1369 443 1381 477
rect 1415 443 1438 477
rect 1369 413 1438 443
rect 1474 467 1532 497
rect 1474 433 1486 467
rect 1520 433 1532 467
rect 1474 413 1532 433
rect 1568 413 1669 497
rect 1705 477 1782 497
rect 1705 443 1739 477
rect 1773 443 1782 477
rect 1705 413 1782 443
rect 1836 475 1890 497
rect 1836 441 1844 475
rect 1878 441 1890 475
rect 1369 347 1421 413
rect 1836 407 1890 441
rect 1836 373 1844 407
rect 1878 373 1890 407
rect 1836 297 1890 373
rect 1926 455 1984 497
rect 1926 421 1938 455
rect 1972 421 1984 455
rect 1926 375 1984 421
rect 1926 341 1938 375
rect 1972 341 1984 375
rect 1926 297 1984 341
rect 2020 479 2078 497
rect 2020 445 2032 479
rect 2066 445 2078 479
rect 2020 411 2078 445
rect 2020 377 2032 411
rect 2066 377 2078 411
rect 2020 343 2078 377
rect 2020 309 2032 343
rect 2066 309 2078 343
rect 2020 297 2078 309
rect 2114 487 2174 497
rect 2114 453 2128 487
rect 2162 453 2174 487
rect 2114 419 2174 453
rect 2114 385 2128 419
rect 2162 385 2174 419
rect 2114 297 2174 385
rect 2210 479 2268 497
rect 2210 445 2222 479
rect 2256 445 2268 479
rect 2210 411 2268 445
rect 2210 377 2222 411
rect 2256 377 2268 411
rect 2210 343 2268 377
rect 2210 309 2222 343
rect 2256 309 2268 343
rect 2210 297 2268 309
rect 2304 487 2364 497
rect 2304 453 2316 487
rect 2350 453 2364 487
rect 2304 419 2364 453
rect 2304 385 2316 419
rect 2350 385 2364 419
rect 2304 297 2364 385
<< ndiffc >>
rect 35 85 69 119
rect 129 59 163 93
rect 223 85 257 119
rect 331 55 365 89
rect 441 55 475 89
rect 636 55 670 89
rect 823 55 857 89
rect 933 73 967 107
rect 1043 73 1077 107
rect 1279 67 1313 101
rect 1407 73 1441 107
rect 1529 73 1563 107
rect 1740 73 1774 107
rect 1844 128 1878 162
rect 1844 60 1878 94
rect 1938 89 1972 123
rect 2032 130 2066 164
rect 2032 62 2066 96
rect 2128 62 2162 96
rect 2222 130 2256 164
rect 2222 62 2256 96
rect 2316 62 2350 96
<< pdiffc >>
rect 36 443 70 477
rect 36 375 70 409
rect 130 427 164 461
rect 224 443 258 477
rect 224 375 258 409
rect 328 418 362 452
rect 422 449 456 483
rect 620 449 654 483
rect 822 449 856 483
rect 926 438 960 472
rect 1035 438 1069 472
rect 1287 451 1321 485
rect 1287 383 1321 417
rect 1381 443 1415 477
rect 1486 433 1520 467
rect 1739 443 1773 477
rect 1844 441 1878 475
rect 1844 373 1878 407
rect 1938 421 1972 455
rect 1938 341 1972 375
rect 2032 445 2066 479
rect 2032 377 2066 411
rect 2032 309 2066 343
rect 2128 453 2162 487
rect 2128 385 2162 419
rect 2222 445 2256 479
rect 2222 377 2256 411
rect 2222 309 2256 343
rect 2316 453 2350 487
rect 2316 385 2350 419
<< poly >>
rect 82 491 118 517
rect 176 491 212 517
rect 374 497 410 523
rect 468 497 504 523
rect 572 497 608 523
rect 666 497 702 523
rect 769 497 805 523
rect 982 497 1018 523
rect 1085 497 1121 523
rect 1191 497 1227 523
rect 1333 497 1369 523
rect 1438 497 1474 523
rect 1532 497 1568 523
rect 1669 497 1705 523
rect 1890 497 1926 523
rect 1984 497 2020 523
rect 2078 497 2114 523
rect 2174 497 2210 523
rect 2268 497 2304 523
rect 982 398 1018 413
rect 1085 398 1121 413
rect 1191 398 1227 413
rect 980 375 1020 398
rect 1083 381 1123 398
rect 82 348 118 363
rect 176 348 212 363
rect 374 354 410 369
rect 468 354 504 369
rect 572 354 608 369
rect 666 354 702 369
rect 769 354 805 369
rect 965 365 1041 375
rect 47 318 120 348
rect 47 265 77 318
rect 174 274 214 348
rect 372 331 412 354
rect 466 331 506 354
rect 570 337 610 354
rect 664 337 704 354
rect 360 321 506 331
rect 360 287 376 321
rect 410 301 506 321
rect 549 321 619 337
rect 410 287 436 301
rect 360 277 436 287
rect 549 287 565 321
rect 599 287 619 321
rect 549 277 619 287
rect 23 249 77 265
rect 23 215 33 249
rect 67 215 77 249
rect 129 264 214 274
rect 129 230 145 264
rect 179 230 214 264
rect 129 220 214 230
rect 23 199 77 215
rect 47 176 77 199
rect 47 146 109 176
rect 79 131 109 146
rect 173 131 203 220
rect 375 131 405 277
rect 585 271 619 277
rect 661 321 725 337
rect 661 287 671 321
rect 705 287 725 321
rect 661 271 725 287
rect 767 304 807 354
rect 965 331 981 365
rect 1015 331 1041 365
rect 965 321 1041 331
rect 1083 365 1147 381
rect 1083 331 1093 365
rect 1127 331 1147 365
rect 1083 315 1147 331
rect 767 288 831 304
rect 467 225 543 235
rect 467 191 493 225
rect 527 191 543 225
rect 467 175 543 191
rect 487 131 517 175
rect 585 131 615 271
rect 767 254 777 288
rect 811 254 831 288
rect 1083 279 1123 315
rect 767 238 831 254
rect 981 249 1123 279
rect 657 207 721 223
rect 657 173 667 207
rect 701 173 721 207
rect 657 157 721 173
rect 691 131 721 157
rect 767 131 797 238
rect 981 119 1011 249
rect 1189 213 1229 398
rect 1438 398 1474 413
rect 1532 398 1568 413
rect 1669 398 1705 413
rect 1333 332 1369 347
rect 1331 309 1371 332
rect 1436 315 1476 398
rect 1530 375 1570 398
rect 1667 381 1707 398
rect 1529 365 1605 375
rect 1529 331 1545 365
rect 1579 331 1605 365
rect 1529 321 1605 331
rect 1667 365 1755 381
rect 1667 331 1711 365
rect 1745 331 1755 365
rect 1667 315 1755 331
rect 1271 299 1371 309
rect 1271 265 1287 299
rect 1321 265 1371 299
rect 1271 255 1371 265
rect 1331 220 1371 255
rect 1423 299 1487 315
rect 1423 265 1433 299
rect 1467 279 1487 299
rect 1467 265 1625 279
rect 1423 249 1625 265
rect 1063 191 1127 207
rect 1063 157 1073 191
rect 1107 157 1127 191
rect 1189 203 1279 213
rect 1189 183 1229 203
rect 1063 141 1127 157
rect 1097 119 1127 141
rect 1205 169 1229 183
rect 1263 169 1279 203
rect 1331 190 1391 220
rect 1361 175 1391 190
rect 1462 191 1533 207
rect 1205 159 1279 169
rect 1205 131 1235 159
rect 1462 157 1489 191
rect 1523 157 1533 191
rect 1462 141 1533 157
rect 1462 119 1492 141
rect 1595 119 1625 249
rect 1690 131 1720 315
rect 1890 282 1926 297
rect 1984 282 2020 297
rect 2078 282 2114 297
rect 2174 282 2210 297
rect 2268 282 2304 297
rect 1888 265 1928 282
rect 1786 249 1928 265
rect 1786 215 1796 249
rect 1830 215 1928 249
rect 1786 199 1928 215
rect 1898 177 1928 199
rect 1982 265 2022 282
rect 2076 265 2116 282
rect 2172 265 2212 282
rect 2266 265 2306 282
rect 1982 249 2306 265
rect 1982 215 1992 249
rect 2026 215 2070 249
rect 2104 215 2148 249
rect 2182 215 2226 249
rect 2260 215 2306 249
rect 1982 199 2306 215
rect 1982 177 2012 199
rect 2076 177 2106 199
rect 2172 177 2202 199
rect 2276 177 2306 199
rect 79 21 109 47
rect 173 21 203 47
rect 375 21 405 47
rect 487 21 517 47
rect 585 21 615 47
rect 691 21 721 47
rect 767 21 797 47
rect 981 21 1011 47
rect 1097 21 1127 47
rect 1205 21 1235 47
rect 1361 21 1391 47
rect 1462 21 1492 47
rect 1595 21 1625 47
rect 1690 21 1720 47
rect 1898 21 1928 47
rect 1982 21 2012 47
rect 2076 21 2106 47
rect 2172 21 2202 47
rect 2276 21 2306 47
<< polycont >>
rect 376 287 410 321
rect 565 287 599 321
rect 33 215 67 249
rect 145 230 179 264
rect 671 287 705 321
rect 981 331 1015 365
rect 1093 331 1127 365
rect 493 191 527 225
rect 777 254 811 288
rect 667 173 701 207
rect 1545 331 1579 365
rect 1711 331 1745 365
rect 1287 265 1321 299
rect 1433 265 1467 299
rect 1073 157 1107 191
rect 1229 169 1263 203
rect 1489 157 1523 191
rect 1796 215 1830 249
rect 1992 215 2026 249
rect 2070 215 2104 249
rect 2148 215 2182 249
rect 2226 215 2260 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2392 561
rect 36 477 70 493
rect 36 409 70 443
rect 104 461 180 527
rect 104 427 130 461
rect 164 427 180 461
rect 223 477 269 493
rect 223 443 224 477
rect 258 443 269 477
rect 223 409 269 443
rect 70 382 179 393
rect 70 375 133 382
rect 36 359 133 375
rect 167 348 179 382
rect 19 249 89 325
rect 19 215 33 249
rect 67 215 89 249
rect 19 195 89 215
rect 133 264 179 348
rect 133 230 145 264
rect 133 161 179 230
rect 35 127 179 161
rect 223 375 224 409
rect 258 375 269 409
rect 223 178 269 375
rect 223 144 231 178
rect 265 144 269 178
rect 35 119 69 127
rect 223 119 269 144
rect 35 69 69 85
rect 103 59 129 93
rect 163 59 179 93
rect 257 85 269 119
rect 223 69 269 85
rect 307 452 362 489
rect 307 418 328 452
rect 396 483 472 527
rect 822 483 856 527
rect 396 449 422 483
rect 456 449 472 483
rect 579 449 620 483
rect 654 449 778 483
rect 307 415 362 418
rect 307 372 705 415
rect 307 89 341 372
rect 376 321 443 337
rect 410 287 443 321
rect 376 157 443 287
rect 477 225 511 372
rect 549 321 630 337
rect 549 287 565 321
rect 599 287 630 321
rect 549 271 630 287
rect 666 321 705 372
rect 744 399 778 449
rect 822 433 856 449
rect 913 472 960 488
rect 1287 485 1321 527
rect 913 438 926 472
rect 1009 438 1035 472
rect 1069 438 1253 472
rect 913 413 960 438
rect 913 399 947 413
rect 744 365 947 399
rect 1077 382 1175 402
rect 666 287 671 321
rect 666 271 705 287
rect 745 288 819 331
rect 745 254 777 288
rect 811 254 819 288
rect 477 191 493 225
rect 527 191 543 225
rect 667 207 701 223
rect 745 207 819 254
rect 913 173 947 365
rect 667 157 701 173
rect 376 123 701 157
rect 745 139 947 173
rect 981 365 1039 381
rect 1015 331 1039 365
rect 1077 365 1133 382
rect 1077 331 1093 365
rect 1127 348 1133 365
rect 1167 348 1175 382
rect 1127 331 1175 348
rect 981 207 1039 331
rect 1209 315 1253 438
rect 1287 417 1321 451
rect 1287 367 1321 383
rect 1355 477 1415 493
rect 1355 443 1381 477
rect 1713 477 1774 527
rect 1355 427 1415 443
rect 1460 433 1486 467
rect 1520 433 1667 467
rect 1209 299 1321 315
rect 1209 297 1287 299
rect 1145 265 1287 297
rect 1145 249 1321 265
rect 981 191 1107 207
rect 981 178 1073 191
rect 981 144 1031 178
rect 1065 157 1073 178
rect 1065 144 1107 157
rect 981 141 1107 144
rect 745 89 779 139
rect 913 107 947 139
rect 1145 107 1179 249
rect 1355 213 1399 427
rect 1433 382 1481 393
rect 1433 348 1445 382
rect 1479 348 1481 382
rect 1433 299 1481 348
rect 1467 265 1481 299
rect 1433 249 1481 265
rect 1515 365 1589 381
rect 1515 331 1545 365
rect 1579 331 1589 365
rect 1515 315 1589 331
rect 1213 203 1399 213
rect 1515 207 1553 315
rect 1633 281 1667 433
rect 1713 443 1739 477
rect 1773 443 1774 477
rect 1713 427 1774 443
rect 1844 475 1901 491
rect 1878 441 1901 475
rect 1844 407 1901 441
rect 1711 373 1844 381
rect 1878 373 1901 407
rect 1711 365 1901 373
rect 1745 331 1901 365
rect 1711 315 1901 331
rect 1938 455 1972 527
rect 2128 487 2162 527
rect 1938 375 1972 421
rect 1938 325 1972 341
rect 2006 445 2032 479
rect 2066 445 2082 479
rect 2006 411 2082 445
rect 2006 377 2032 411
rect 2066 377 2082 411
rect 2006 343 2082 377
rect 2316 487 2350 527
rect 2128 419 2162 453
rect 2128 369 2162 385
rect 2196 445 2222 479
rect 2256 445 2272 479
rect 2196 411 2272 445
rect 2196 377 2222 411
rect 2256 377 2272 411
rect 1213 169 1229 203
rect 1263 169 1399 203
rect 1213 153 1399 169
rect 103 17 179 59
rect 307 55 331 89
rect 365 55 381 89
rect 425 55 441 89
rect 475 55 491 89
rect 614 55 636 89
rect 670 55 779 89
rect 823 89 863 105
rect 857 55 863 89
rect 913 73 933 107
rect 967 73 983 107
rect 1027 73 1043 107
rect 1077 73 1179 107
rect 1245 101 1319 117
rect 425 17 491 55
rect 823 17 863 55
rect 1245 67 1279 101
rect 1313 67 1319 101
rect 1355 107 1399 153
rect 1433 191 1553 207
rect 1433 178 1489 191
rect 1433 144 1445 178
rect 1479 157 1489 178
rect 1523 157 1553 191
rect 1479 144 1553 157
rect 1433 141 1553 144
rect 1597 265 1667 281
rect 1864 265 1901 315
rect 2006 309 2032 343
rect 2066 335 2082 343
rect 2196 343 2272 377
rect 2316 419 2350 453
rect 2316 369 2350 385
rect 2196 335 2222 343
rect 2066 309 2222 335
rect 2256 335 2272 343
rect 2256 309 2370 335
rect 2006 301 2370 309
rect 1597 249 1830 265
rect 1597 215 1796 249
rect 1597 199 1830 215
rect 1864 249 2276 265
rect 1864 215 1992 249
rect 2026 215 2070 249
rect 2104 215 2148 249
rect 2182 215 2226 249
rect 2260 215 2276 249
rect 1597 107 1641 199
rect 1864 165 1900 215
rect 2310 181 2370 301
rect 1828 162 1900 165
rect 1828 128 1844 162
rect 1878 128 1900 162
rect 2006 164 2370 181
rect 1355 73 1407 107
rect 1441 73 1457 107
rect 1513 73 1529 107
rect 1563 73 1641 107
rect 1690 107 1774 123
rect 1690 73 1740 107
rect 1245 17 1319 67
rect 1690 17 1774 73
rect 1828 94 1900 128
rect 1828 60 1844 94
rect 1878 60 1900 94
rect 1938 123 1972 139
rect 1938 17 1972 89
rect 2006 130 2032 164
rect 2066 147 2222 164
rect 2066 130 2082 147
rect 2006 96 2082 130
rect 2196 130 2222 147
rect 2256 147 2370 164
rect 2256 130 2272 147
rect 2006 62 2032 96
rect 2066 62 2082 96
rect 2006 61 2082 62
rect 2128 96 2162 113
rect 2128 17 2162 62
rect 2196 96 2272 130
rect 2196 62 2222 96
rect 2256 62 2272 96
rect 2196 61 2272 62
rect 2316 96 2350 113
rect 2316 17 2350 62
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2392 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 133 348 167 382
rect 231 144 265 178
rect 1133 348 1167 382
rect 1031 144 1065 178
rect 1445 348 1479 382
rect 1445 144 1479 178
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
<< metal1 >>
rect 0 561 2392 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2392 561
rect 0 496 2392 527
rect 121 382 1491 388
rect 121 348 133 382
rect 167 360 1133 382
rect 167 348 179 360
rect 121 342 179 348
rect 1111 348 1133 360
rect 1167 360 1445 382
rect 1167 348 1179 360
rect 1111 342 1179 348
rect 1423 348 1445 360
rect 1479 348 1491 382
rect 1423 342 1491 348
rect 219 178 1491 184
rect 219 144 231 178
rect 265 156 1031 178
rect 265 144 277 156
rect 219 138 277 144
rect 1009 144 1031 156
rect 1065 156 1445 178
rect 1065 144 1077 156
rect 1009 138 1077 144
rect 1423 144 1445 156
rect 1479 144 1491 178
rect 1423 138 1491 144
rect 0 17 2392 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2392 17
rect 0 -48 2392 -17
<< labels >>
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
flabel corelocali s 764 221 798 255 0 FreeSans 300 0 0 0 SCD
port 3 nsew
flabel corelocali s 581 289 615 323 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel corelocali s 397 152 431 186 0 FreeSans 300 0 0 0 SCE
port 4 nsew
flabel corelocali s 29 221 63 255 0 FreeSans 400 0 0 0 CLK
port 1 nsew
flabel corelocali s 2324 221 2358 255 0 FreeSans 300 0 0 0 Q
port 9 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel nbase s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
port 7 nsew
rlabel comment s 0 0 0 0 4 sdfxtp_4
<< properties >>
string FIXED_BBOX 0 0 2392 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 369710
string GDS_START 352612
<< end >>
