magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 1173 391 1215 493
rect 1173 357 1300 391
rect 18 215 88 255
rect 1266 323 1300 357
rect 1353 323 1403 493
rect 213 289 609 323
rect 213 215 346 289
rect 390 215 499 255
rect 533 215 609 289
rect 661 289 1045 323
rect 1266 289 1542 323
rect 661 215 791 289
rect 995 255 1045 289
rect 825 215 951 255
rect 995 215 1107 255
rect 1473 181 1542 289
rect 1147 147 1542 181
rect 1147 145 1411 147
rect 1147 51 1223 145
rect 1335 51 1411 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 29 291 79 527
rect 123 391 173 493
rect 217 425 267 527
rect 311 459 549 493
rect 311 425 361 459
rect 499 425 549 459
rect 593 425 745 527
rect 789 459 1027 493
rect 789 425 839 459
rect 977 425 1027 459
rect 1071 425 1121 527
rect 1259 425 1309 527
rect 123 357 1129 391
rect 17 95 69 179
rect 123 173 179 357
rect 1095 323 1129 357
rect 1447 359 1497 527
rect 1095 289 1185 323
rect 1141 255 1185 289
rect 1141 215 1411 255
rect 103 129 179 173
rect 223 95 257 181
rect 291 145 1035 181
rect 291 129 847 145
rect 17 51 651 95
rect 687 17 753 93
rect 797 51 847 129
rect 891 17 925 111
rect 959 51 1035 145
rect 1079 17 1113 181
rect 1267 17 1301 111
rect 1455 17 1506 113
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
<< metal1 >>
rect 0 561 1564 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 0 496 1564 527
rect 0 17 1564 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
rect 0 -48 1564 -17
<< labels >>
rlabel locali s 995 255 1045 289 6 A1
port 1 nsew signal input
rlabel locali s 995 215 1107 255 6 A1
port 1 nsew signal input
rlabel locali s 661 289 1045 323 6 A1
port 1 nsew signal input
rlabel locali s 661 215 791 289 6 A1
port 1 nsew signal input
rlabel locali s 825 215 951 255 6 A2
port 2 nsew signal input
rlabel locali s 533 215 609 289 6 B1
port 3 nsew signal input
rlabel locali s 213 289 609 323 6 B1
port 3 nsew signal input
rlabel locali s 213 215 346 289 6 B1
port 3 nsew signal input
rlabel locali s 390 215 499 255 6 B2
port 4 nsew signal input
rlabel locali s 18 215 88 255 6 C1
port 5 nsew signal input
rlabel locali s 1473 181 1542 289 6 X
port 6 nsew signal output
rlabel locali s 1353 323 1403 493 6 X
port 6 nsew signal output
rlabel locali s 1335 51 1411 145 6 X
port 6 nsew signal output
rlabel locali s 1266 323 1300 357 6 X
port 6 nsew signal output
rlabel locali s 1266 289 1542 323 6 X
port 6 nsew signal output
rlabel locali s 1173 391 1215 493 6 X
port 6 nsew signal output
rlabel locali s 1173 357 1300 391 6 X
port 6 nsew signal output
rlabel locali s 1147 147 1542 181 6 X
port 6 nsew signal output
rlabel locali s 1147 145 1411 147 6 X
port 6 nsew signal output
rlabel locali s 1147 51 1223 145 6 X
port 6 nsew signal output
rlabel metal1 s 0 -48 1564 48 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 496 1564 592 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1564 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 847230
string GDS_START 835908
<< end >>
