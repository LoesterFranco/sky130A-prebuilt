magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 460 561
rect 26 299 79 527
rect 113 333 179 493
rect 213 367 247 527
rect 281 337 347 493
rect 381 435 423 527
rect 281 333 434 337
rect 113 299 434 333
rect 21 215 347 265
rect 381 181 434 299
rect 113 145 434 181
rect 26 17 79 109
rect 113 51 179 145
rect 213 17 247 109
rect 281 51 347 145
rect 381 17 431 110
rect 0 -17 460 17
<< metal1 >>
rect 0 496 460 592
rect 0 -48 460 48
<< labels >>
rlabel locali s 21 215 347 265 6 A
port 1 nsew signal input
rlabel locali s 381 181 434 299 6 Y
port 2 nsew signal output
rlabel locali s 281 337 347 493 6 Y
port 2 nsew signal output
rlabel locali s 281 333 434 337 6 Y
port 2 nsew signal output
rlabel locali s 281 51 347 145 6 Y
port 2 nsew signal output
rlabel locali s 113 333 179 493 6 Y
port 2 nsew signal output
rlabel locali s 113 299 434 333 6 Y
port 2 nsew signal output
rlabel locali s 113 145 434 181 6 Y
port 2 nsew signal output
rlabel locali s 113 51 179 145 6 Y
port 2 nsew signal output
rlabel locali s 381 17 431 110 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 213 17 247 109 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 26 17 79 109 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 0 -17 460 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 460 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 381 435 423 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 213 367 247 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 26 299 79 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 0 527 460 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 496 460 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 460 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2235240
string GDS_START 2230250
<< end >>
