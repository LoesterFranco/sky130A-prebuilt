magic
tech sky130A
magscale 1 2
timestamp 1601050088
<< locali >>
rect 217 290 314 356
rect 505 282 556 547
rect 21 57 87 134
rect 505 230 647 282
rect 681 264 747 356
rect 793 270 935 356
rect 416 196 759 230
rect 416 78 450 196
rect 693 154 759 196
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 116 388 182 649
rect 284 390 382 596
rect 348 330 382 390
rect 416 581 646 615
rect 416 364 466 581
rect 348 264 441 330
rect 596 424 646 581
rect 686 458 752 649
rect 792 424 826 596
rect 866 458 932 649
rect 972 424 1022 596
rect 596 390 1022 424
rect 596 364 646 390
rect 972 364 1022 390
rect 348 256 382 264
rect 121 17 171 234
rect 207 222 382 256
rect 207 98 266 222
rect 314 17 380 188
rect 486 17 552 162
rect 795 202 1017 236
rect 795 120 829 202
rect 607 70 829 120
rect 865 17 915 168
rect 951 70 1017 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 683 1056 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 0 617 1056 649
rect 0 17 1056 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -49 1056 -17
<< labels >>
rlabel locali s 21 57 87 134 6 A1_N
port 1 nsew signal input
rlabel locali s 217 290 314 356 6 A2_N
port 2 nsew signal input
rlabel locali s 793 270 935 356 6 B1
port 3 nsew signal input
rlabel locali s 681 264 747 356 6 B2
port 4 nsew signal input
rlabel locali s 693 154 759 196 6 Y
port 5 nsew signal output
rlabel locali s 505 282 556 547 6 Y
port 5 nsew signal output
rlabel locali s 505 230 647 282 6 Y
port 5 nsew signal output
rlabel locali s 416 196 759 230 6 Y
port 5 nsew signal output
rlabel locali s 416 78 450 196 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -49 1056 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 1056 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1056 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3657914
string GDS_START 3649220
<< end >>
