magic
tech sky130A
magscale 1 2
timestamp 1599588232
<< locali >>
rect 261 424 327 596
rect 461 424 559 596
rect 261 390 559 424
rect 461 364 559 390
rect 89 270 167 356
rect 203 270 269 356
rect 313 270 383 356
rect 525 230 559 364
rect 485 158 559 230
rect 450 74 559 158
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 21 390 120 540
rect 161 390 227 649
rect 361 458 427 649
rect 21 230 55 390
rect 417 264 491 330
rect 417 230 451 264
rect 21 196 451 230
rect 21 112 75 196
rect 109 17 244 162
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
rlabel locali s 89 270 167 356 6 A_N
port 1 nsew signal input
rlabel locali s 313 270 383 356 6 B
port 2 nsew signal input
rlabel locali s 203 270 269 356 6 C
port 3 nsew signal input
rlabel locali s 525 230 559 364 6 Y
port 4 nsew signal output
rlabel locali s 485 158 559 230 6 Y
port 4 nsew signal output
rlabel locali s 461 424 559 596 6 Y
port 4 nsew signal output
rlabel locali s 461 364 559 390 6 Y
port 4 nsew signal output
rlabel locali s 450 74 559 158 6 Y
port 4 nsew signal output
rlabel locali s 261 424 327 596 6 Y
port 4 nsew signal output
rlabel locali s 261 390 559 424 6 Y
port 4 nsew signal output
rlabel metal1 s 0 -49 576 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 6 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 617 576 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 576 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 2088790
string GDS_START 2083154
<< end >>
