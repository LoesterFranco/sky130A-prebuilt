magic
tech sky130A
magscale 1 2
timestamp 1604502701
<< nwell >>
rect -38 332 1670 704
<< pwell >>
rect 0 0 1632 49
<< scpmos >>
rect 86 368 116 592
rect 176 368 206 592
rect 276 368 306 592
rect 366 368 396 592
rect 466 368 496 592
rect 556 368 586 592
rect 656 368 686 592
rect 746 368 776 592
rect 836 368 866 592
rect 926 368 956 592
rect 1020 368 1050 592
rect 1116 368 1146 592
rect 1226 368 1256 592
rect 1316 368 1346 592
rect 1426 368 1456 592
rect 1516 368 1546 592
<< nmoslvt >>
rect 98 74 128 222
rect 184 74 214 222
rect 284 74 314 222
rect 370 74 400 222
rect 470 74 500 222
rect 556 74 586 222
rect 656 74 686 222
rect 742 74 772 222
rect 828 74 858 222
rect 914 74 944 222
rect 1014 74 1044 222
rect 1100 74 1130 222
rect 1214 74 1244 222
rect 1300 74 1330 222
rect 1418 74 1448 222
rect 1504 74 1534 222
<< ndiff >>
rect 45 210 98 222
rect 45 176 53 210
rect 87 176 98 210
rect 45 120 98 176
rect 45 86 53 120
rect 87 86 98 120
rect 45 74 98 86
rect 128 210 184 222
rect 128 176 139 210
rect 173 176 184 210
rect 128 120 184 176
rect 128 86 139 120
rect 173 86 184 120
rect 128 74 184 86
rect 214 210 284 222
rect 214 176 239 210
rect 273 176 284 210
rect 214 120 284 176
rect 214 86 239 120
rect 273 86 284 120
rect 214 74 284 86
rect 314 210 370 222
rect 314 176 325 210
rect 359 176 370 210
rect 314 120 370 176
rect 314 86 325 120
rect 359 86 370 120
rect 314 74 370 86
rect 400 210 470 222
rect 400 176 411 210
rect 445 176 470 210
rect 400 120 470 176
rect 400 86 411 120
rect 445 86 470 120
rect 400 74 470 86
rect 500 210 556 222
rect 500 176 511 210
rect 545 176 556 210
rect 500 120 556 176
rect 500 86 511 120
rect 545 86 556 120
rect 500 74 556 86
rect 586 210 656 222
rect 586 176 607 210
rect 641 176 656 210
rect 586 120 656 176
rect 586 86 607 120
rect 641 86 656 120
rect 586 74 656 86
rect 686 210 742 222
rect 686 176 697 210
rect 731 176 742 210
rect 686 120 742 176
rect 686 86 697 120
rect 731 86 742 120
rect 686 74 742 86
rect 772 210 828 222
rect 772 176 783 210
rect 817 176 828 210
rect 772 120 828 176
rect 772 86 783 120
rect 817 86 828 120
rect 772 74 828 86
rect 858 210 914 222
rect 858 176 869 210
rect 903 176 914 210
rect 858 120 914 176
rect 858 86 869 120
rect 903 86 914 120
rect 858 74 914 86
rect 944 210 1014 222
rect 944 176 962 210
rect 996 176 1014 210
rect 944 123 1014 176
rect 944 89 962 123
rect 996 89 1014 123
rect 944 74 1014 89
rect 1044 210 1100 222
rect 1044 176 1055 210
rect 1089 176 1100 210
rect 1044 120 1100 176
rect 1044 86 1055 120
rect 1089 86 1100 120
rect 1044 74 1100 86
rect 1130 210 1214 222
rect 1130 176 1155 210
rect 1189 176 1214 210
rect 1130 123 1214 176
rect 1130 89 1155 123
rect 1189 89 1214 123
rect 1130 74 1214 89
rect 1244 210 1300 222
rect 1244 176 1255 210
rect 1289 176 1300 210
rect 1244 120 1300 176
rect 1244 86 1255 120
rect 1289 86 1300 120
rect 1244 74 1300 86
rect 1330 210 1418 222
rect 1330 176 1357 210
rect 1391 176 1418 210
rect 1330 123 1418 176
rect 1330 89 1357 123
rect 1391 89 1418 123
rect 1330 74 1418 89
rect 1448 210 1504 222
rect 1448 176 1459 210
rect 1493 176 1504 210
rect 1448 120 1504 176
rect 1448 86 1459 120
rect 1493 86 1504 120
rect 1448 74 1504 86
rect 1534 210 1587 222
rect 1534 176 1545 210
rect 1579 176 1587 210
rect 1534 120 1587 176
rect 1534 86 1545 120
rect 1579 86 1587 120
rect 1534 74 1587 86
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 497 86 546
rect 27 463 39 497
rect 73 463 86 497
rect 27 414 86 463
rect 27 380 39 414
rect 73 380 86 414
rect 27 368 86 380
rect 116 580 176 592
rect 116 546 129 580
rect 163 546 176 580
rect 116 497 176 546
rect 116 463 129 497
rect 163 463 176 497
rect 116 414 176 463
rect 116 380 129 414
rect 163 380 176 414
rect 116 368 176 380
rect 206 580 276 592
rect 206 546 219 580
rect 253 546 276 580
rect 206 506 276 546
rect 206 472 219 506
rect 253 472 276 506
rect 206 438 276 472
rect 206 404 219 438
rect 253 404 276 438
rect 206 368 276 404
rect 306 580 366 592
rect 306 546 319 580
rect 353 546 366 580
rect 306 501 366 546
rect 306 467 319 501
rect 353 467 366 501
rect 306 422 366 467
rect 306 388 319 422
rect 353 388 366 422
rect 306 368 366 388
rect 396 580 466 592
rect 396 546 409 580
rect 443 546 466 580
rect 396 506 466 546
rect 396 472 409 506
rect 443 472 466 506
rect 396 438 466 472
rect 396 404 409 438
rect 443 404 466 438
rect 396 368 466 404
rect 496 580 556 592
rect 496 546 509 580
rect 543 546 556 580
rect 496 497 556 546
rect 496 463 509 497
rect 543 463 556 497
rect 496 414 556 463
rect 496 380 509 414
rect 543 380 556 414
rect 496 368 556 380
rect 586 580 656 592
rect 586 546 599 580
rect 633 546 656 580
rect 586 506 656 546
rect 586 472 599 506
rect 633 472 656 506
rect 586 438 656 472
rect 586 404 599 438
rect 633 404 656 438
rect 586 368 656 404
rect 686 580 746 592
rect 686 546 699 580
rect 733 546 746 580
rect 686 497 746 546
rect 686 463 699 497
rect 733 463 746 497
rect 686 414 746 463
rect 686 380 699 414
rect 733 380 746 414
rect 686 368 746 380
rect 776 580 836 592
rect 776 546 789 580
rect 823 546 836 580
rect 776 506 836 546
rect 776 472 789 506
rect 823 472 836 506
rect 776 438 836 472
rect 776 404 789 438
rect 823 404 836 438
rect 776 368 836 404
rect 866 580 926 592
rect 866 546 879 580
rect 913 546 926 580
rect 866 497 926 546
rect 866 463 879 497
rect 913 463 926 497
rect 866 414 926 463
rect 866 380 879 414
rect 913 380 926 414
rect 866 368 926 380
rect 956 580 1020 592
rect 956 546 969 580
rect 1003 546 1020 580
rect 956 506 1020 546
rect 956 472 969 506
rect 1003 472 1020 506
rect 956 438 1020 472
rect 956 404 969 438
rect 1003 404 1020 438
rect 956 368 1020 404
rect 1050 580 1116 592
rect 1050 546 1069 580
rect 1103 546 1116 580
rect 1050 497 1116 546
rect 1050 463 1069 497
rect 1103 463 1116 497
rect 1050 414 1116 463
rect 1050 380 1069 414
rect 1103 380 1116 414
rect 1050 368 1116 380
rect 1146 580 1226 592
rect 1146 546 1169 580
rect 1203 546 1226 580
rect 1146 506 1226 546
rect 1146 472 1169 506
rect 1203 472 1226 506
rect 1146 438 1226 472
rect 1146 404 1169 438
rect 1203 404 1226 438
rect 1146 368 1226 404
rect 1256 580 1316 592
rect 1256 546 1269 580
rect 1303 546 1316 580
rect 1256 497 1316 546
rect 1256 463 1269 497
rect 1303 463 1316 497
rect 1256 414 1316 463
rect 1256 380 1269 414
rect 1303 380 1316 414
rect 1256 368 1316 380
rect 1346 580 1426 592
rect 1346 546 1369 580
rect 1403 546 1426 580
rect 1346 506 1426 546
rect 1346 472 1369 506
rect 1403 472 1426 506
rect 1346 438 1426 472
rect 1346 404 1369 438
rect 1403 404 1426 438
rect 1346 368 1426 404
rect 1456 580 1516 592
rect 1456 546 1469 580
rect 1503 546 1516 580
rect 1456 497 1516 546
rect 1456 463 1469 497
rect 1503 463 1516 497
rect 1456 414 1516 463
rect 1456 380 1469 414
rect 1503 380 1516 414
rect 1456 368 1516 380
rect 1546 580 1605 592
rect 1546 546 1559 580
rect 1593 546 1605 580
rect 1546 497 1605 546
rect 1546 463 1559 497
rect 1593 463 1605 497
rect 1546 414 1605 463
rect 1546 380 1559 414
rect 1593 380 1605 414
rect 1546 368 1605 380
<< ndiffc >>
rect 53 176 87 210
rect 53 86 87 120
rect 139 176 173 210
rect 139 86 173 120
rect 239 176 273 210
rect 239 86 273 120
rect 325 176 359 210
rect 325 86 359 120
rect 411 176 445 210
rect 411 86 445 120
rect 511 176 545 210
rect 511 86 545 120
rect 607 176 641 210
rect 607 86 641 120
rect 697 176 731 210
rect 697 86 731 120
rect 783 176 817 210
rect 783 86 817 120
rect 869 176 903 210
rect 869 86 903 120
rect 962 176 996 210
rect 962 89 996 123
rect 1055 176 1089 210
rect 1055 86 1089 120
rect 1155 176 1189 210
rect 1155 89 1189 123
rect 1255 176 1289 210
rect 1255 86 1289 120
rect 1357 176 1391 210
rect 1357 89 1391 123
rect 1459 176 1493 210
rect 1459 86 1493 120
rect 1545 176 1579 210
rect 1545 86 1579 120
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 129 546 163 580
rect 129 463 163 497
rect 129 380 163 414
rect 219 546 253 580
rect 219 472 253 506
rect 219 404 253 438
rect 319 546 353 580
rect 319 467 353 501
rect 319 388 353 422
rect 409 546 443 580
rect 409 472 443 506
rect 409 404 443 438
rect 509 546 543 580
rect 509 463 543 497
rect 509 380 543 414
rect 599 546 633 580
rect 599 472 633 506
rect 599 404 633 438
rect 699 546 733 580
rect 699 463 733 497
rect 699 380 733 414
rect 789 546 823 580
rect 789 472 823 506
rect 789 404 823 438
rect 879 546 913 580
rect 879 463 913 497
rect 879 380 913 414
rect 969 546 1003 580
rect 969 472 1003 506
rect 969 404 1003 438
rect 1069 546 1103 580
rect 1069 463 1103 497
rect 1069 380 1103 414
rect 1169 546 1203 580
rect 1169 472 1203 506
rect 1169 404 1203 438
rect 1269 546 1303 580
rect 1269 463 1303 497
rect 1269 380 1303 414
rect 1369 546 1403 580
rect 1369 472 1403 506
rect 1369 404 1403 438
rect 1469 546 1503 580
rect 1469 463 1503 497
rect 1469 380 1503 414
rect 1559 546 1593 580
rect 1559 463 1593 497
rect 1559 380 1593 414
<< poly >>
rect 86 592 116 618
rect 176 592 206 618
rect 276 592 306 618
rect 366 592 396 618
rect 466 592 496 618
rect 556 592 586 618
rect 656 592 686 618
rect 746 592 776 618
rect 836 592 866 618
rect 926 592 956 618
rect 1020 592 1050 618
rect 1116 592 1146 618
rect 1226 592 1256 618
rect 1316 592 1346 618
rect 1426 592 1456 618
rect 1516 592 1546 618
rect 86 353 116 368
rect 176 353 206 368
rect 276 353 306 368
rect 366 353 396 368
rect 466 353 496 368
rect 556 353 586 368
rect 656 353 686 368
rect 746 353 776 368
rect 836 353 866 368
rect 926 353 956 368
rect 1020 353 1050 368
rect 1116 353 1146 368
rect 1226 353 1256 368
rect 1316 353 1346 368
rect 1426 353 1456 368
rect 1516 353 1546 368
rect 83 336 119 353
rect 173 336 209 353
rect 273 336 309 353
rect 363 336 399 353
rect 463 336 499 353
rect 553 336 589 353
rect 653 336 689 353
rect 743 336 779 353
rect 833 336 869 353
rect 923 336 959 353
rect 1017 336 1053 353
rect 1113 336 1149 353
rect 1223 336 1259 353
rect 1313 336 1349 353
rect 1423 336 1459 353
rect 1513 336 1549 353
rect 83 320 1549 336
rect 83 286 229 320
rect 263 286 417 320
rect 451 286 605 320
rect 639 286 788 320
rect 822 286 970 320
rect 1004 286 1169 320
rect 1203 286 1368 320
rect 1402 286 1549 320
rect 83 270 1549 286
rect 98 222 128 270
rect 184 222 214 270
rect 284 222 314 270
rect 370 222 400 270
rect 470 222 500 270
rect 556 222 586 270
rect 656 222 686 270
rect 742 222 772 270
rect 828 222 858 270
rect 914 222 944 270
rect 1014 222 1044 270
rect 1100 222 1130 270
rect 1214 222 1244 270
rect 1300 222 1330 270
rect 1418 222 1448 270
rect 1504 222 1534 270
rect 98 48 128 74
rect 184 48 214 74
rect 284 48 314 74
rect 370 48 400 74
rect 470 48 500 74
rect 556 48 586 74
rect 656 48 686 74
rect 742 48 772 74
rect 828 48 858 74
rect 914 48 944 74
rect 1014 48 1044 74
rect 1100 48 1130 74
rect 1214 48 1244 74
rect 1300 48 1330 74
rect 1418 48 1448 74
rect 1504 48 1534 74
<< polycont >>
rect 229 286 263 320
rect 417 286 451 320
rect 605 286 639 320
rect 788 286 822 320
rect 970 286 1004 320
rect 1169 286 1203 320
rect 1368 286 1402 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 23 580 73 649
rect 23 546 39 580
rect 23 497 73 546
rect 23 463 39 497
rect 23 414 73 463
rect 23 380 39 414
rect 23 364 73 380
rect 113 580 177 599
rect 113 546 129 580
rect 163 546 177 580
rect 113 497 177 546
rect 113 463 129 497
rect 163 463 177 497
rect 113 424 177 463
rect 113 380 129 424
rect 163 380 177 424
rect 211 580 269 649
rect 211 546 219 580
rect 253 546 269 580
rect 211 506 269 546
rect 211 472 219 506
rect 253 472 269 506
rect 211 438 269 472
rect 211 404 219 438
rect 253 404 269 438
rect 211 388 269 404
rect 303 580 369 596
rect 303 546 319 580
rect 353 546 369 580
rect 303 501 369 546
rect 303 467 319 501
rect 353 467 369 501
rect 303 424 369 467
rect 303 388 319 424
rect 353 388 369 424
rect 409 580 459 649
rect 443 546 459 580
rect 409 506 459 546
rect 443 472 459 506
rect 409 438 459 472
rect 443 404 459 438
rect 409 388 459 404
rect 493 580 559 596
rect 493 546 509 580
rect 543 546 559 580
rect 493 497 559 546
rect 493 463 509 497
rect 543 463 559 497
rect 493 424 559 463
rect 493 388 509 424
rect 113 266 177 380
rect 214 350 276 354
rect 214 286 229 350
rect 263 286 276 350
rect 214 270 276 286
rect 123 226 177 266
rect 37 210 89 226
rect 37 176 53 210
rect 87 176 89 210
rect 37 120 89 176
rect 37 86 53 120
rect 87 86 89 120
rect 37 17 89 86
rect 123 210 189 226
rect 123 176 139 210
rect 173 176 189 210
rect 123 120 189 176
rect 123 86 139 120
rect 173 86 189 120
rect 123 70 189 86
rect 223 210 275 226
rect 223 176 239 210
rect 273 176 275 210
rect 223 120 275 176
rect 223 86 239 120
rect 273 86 275 120
rect 223 17 275 86
rect 311 210 369 388
rect 497 380 509 388
rect 543 380 559 424
rect 599 580 649 649
rect 633 546 649 580
rect 599 506 649 546
rect 633 472 649 506
rect 599 438 649 472
rect 633 404 649 438
rect 599 388 649 404
rect 683 580 742 596
rect 683 546 699 580
rect 733 546 742 580
rect 683 497 742 546
rect 683 463 699 497
rect 733 463 742 497
rect 683 424 742 463
rect 404 350 462 354
rect 404 286 417 350
rect 451 286 462 350
rect 404 270 462 286
rect 311 176 325 210
rect 359 176 369 210
rect 311 120 369 176
rect 311 86 325 120
rect 359 86 369 120
rect 311 70 369 86
rect 405 210 461 226
rect 405 176 411 210
rect 445 176 461 210
rect 405 120 461 176
rect 405 86 411 120
rect 445 86 461 120
rect 405 17 461 86
rect 497 210 559 380
rect 683 380 699 424
rect 733 380 742 424
rect 783 580 830 649
rect 783 546 789 580
rect 823 546 830 580
rect 783 506 830 546
rect 783 472 789 506
rect 823 472 830 506
rect 783 438 830 472
rect 783 404 789 438
rect 823 404 830 438
rect 783 388 830 404
rect 868 580 926 596
rect 868 546 879 580
rect 913 546 926 580
rect 868 497 926 546
rect 868 463 879 497
rect 913 463 926 497
rect 868 424 926 463
rect 594 350 649 354
rect 594 286 605 350
rect 639 286 649 350
rect 594 270 649 286
rect 497 176 511 210
rect 545 176 559 210
rect 497 120 559 176
rect 497 86 511 120
rect 545 86 559 120
rect 497 70 559 86
rect 595 210 649 226
rect 595 176 607 210
rect 641 176 649 210
rect 595 120 649 176
rect 595 86 607 120
rect 641 86 649 120
rect 595 17 649 86
rect 683 210 742 380
rect 868 380 879 424
rect 913 388 926 424
rect 962 580 1019 649
rect 962 546 969 580
rect 1003 546 1019 580
rect 962 506 1019 546
rect 962 472 969 506
rect 1003 472 1019 506
rect 962 438 1019 472
rect 962 404 969 438
rect 1003 404 1019 438
rect 962 388 1019 404
rect 1053 580 1116 596
rect 1053 546 1069 580
rect 1103 546 1116 580
rect 1053 497 1116 546
rect 1053 463 1069 497
rect 1103 463 1116 497
rect 1053 424 1116 463
rect 913 380 919 388
rect 777 350 833 354
rect 777 286 788 350
rect 822 286 833 350
rect 777 270 833 286
rect 683 176 697 210
rect 731 176 742 210
rect 683 120 742 176
rect 683 86 697 120
rect 731 86 742 120
rect 683 70 742 86
rect 778 210 830 226
rect 778 176 783 210
rect 817 176 830 210
rect 778 120 830 176
rect 778 86 783 120
rect 817 86 830 120
rect 778 17 830 86
rect 868 210 919 380
rect 1053 380 1069 424
rect 1103 380 1116 424
rect 1153 580 1219 649
rect 1153 546 1169 580
rect 1203 546 1219 580
rect 1153 506 1219 546
rect 1153 472 1169 506
rect 1203 472 1219 506
rect 1153 438 1219 472
rect 1153 404 1169 438
rect 1203 404 1219 438
rect 1153 388 1219 404
rect 1253 580 1319 596
rect 1253 546 1269 580
rect 1303 546 1319 580
rect 1253 497 1319 546
rect 1253 463 1269 497
rect 1303 463 1319 497
rect 1253 424 1319 463
rect 954 350 1017 354
rect 954 286 970 350
rect 1004 286 1017 350
rect 954 270 1017 286
rect 1053 257 1116 380
rect 1253 380 1269 424
rect 1303 380 1319 424
rect 1353 580 1419 649
rect 1353 546 1369 580
rect 1403 546 1419 580
rect 1353 506 1419 546
rect 1353 472 1369 506
rect 1403 472 1419 506
rect 1353 438 1419 472
rect 1353 404 1369 438
rect 1403 404 1419 438
rect 1353 388 1419 404
rect 1453 580 1509 596
rect 1453 546 1469 580
rect 1503 546 1509 580
rect 1453 497 1509 546
rect 1453 463 1469 497
rect 1503 463 1509 497
rect 1453 424 1509 463
rect 1151 350 1218 354
rect 1151 286 1169 350
rect 1203 286 1218 350
rect 1151 270 1218 286
rect 1253 257 1319 380
rect 1453 380 1469 424
rect 1503 380 1509 424
rect 1354 350 1418 354
rect 1354 286 1368 350
rect 1402 286 1418 350
rect 1354 270 1418 286
rect 1053 236 1105 257
rect 1253 236 1305 257
rect 868 176 869 210
rect 903 176 919 210
rect 868 120 919 176
rect 868 86 869 120
rect 903 86 919 120
rect 868 70 919 86
rect 953 210 1005 226
rect 953 176 962 210
rect 996 176 1005 210
rect 953 123 1005 176
rect 953 89 962 123
rect 996 89 1005 123
rect 953 17 1005 89
rect 1043 210 1105 236
rect 1043 176 1055 210
rect 1089 176 1105 210
rect 1043 120 1105 176
rect 1043 86 1055 120
rect 1089 86 1105 120
rect 1043 70 1105 86
rect 1141 210 1205 226
rect 1141 176 1155 210
rect 1189 176 1205 210
rect 1141 123 1205 176
rect 1141 89 1155 123
rect 1189 89 1205 123
rect 1141 17 1205 89
rect 1239 210 1305 236
rect 1453 226 1509 380
rect 1547 580 1609 649
rect 1547 546 1559 580
rect 1593 546 1609 580
rect 1547 497 1609 546
rect 1547 463 1559 497
rect 1593 463 1609 497
rect 1547 414 1609 463
rect 1547 380 1559 414
rect 1593 380 1609 414
rect 1547 364 1609 380
rect 1239 176 1255 210
rect 1289 176 1305 210
rect 1239 120 1305 176
rect 1239 86 1255 120
rect 1289 86 1305 120
rect 1239 70 1305 86
rect 1341 210 1409 226
rect 1341 176 1357 210
rect 1391 176 1409 210
rect 1341 123 1409 176
rect 1341 89 1357 123
rect 1391 89 1409 123
rect 1341 17 1409 89
rect 1443 210 1509 226
rect 1443 176 1459 210
rect 1493 176 1509 210
rect 1443 120 1509 176
rect 1443 86 1459 120
rect 1493 86 1509 120
rect 1443 70 1509 86
rect 1543 210 1609 226
rect 1543 176 1545 210
rect 1579 176 1609 210
rect 1543 120 1609 176
rect 1543 86 1545 120
rect 1579 86 1609 120
rect 1543 17 1609 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 129 414 163 424
rect 129 390 163 414
rect 319 422 353 424
rect 319 390 353 422
rect 509 414 543 424
rect 509 390 543 414
rect 229 320 263 350
rect 229 316 263 320
rect 417 320 451 350
rect 417 316 451 320
rect 699 414 733 424
rect 699 390 733 414
rect 605 320 639 350
rect 605 316 639 320
rect 879 414 913 424
rect 879 390 913 414
rect 788 320 822 350
rect 788 316 822 320
rect 1069 414 1103 424
rect 1069 390 1103 414
rect 970 320 1004 350
rect 970 316 1004 320
rect 1269 414 1303 424
rect 1269 390 1303 414
rect 1169 320 1203 350
rect 1169 316 1203 320
rect 1469 414 1503 424
rect 1469 390 1503 414
rect 1368 320 1402 350
rect 1368 316 1402 320
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 117 424 1515 430
rect 117 390 129 424
rect 163 390 319 424
rect 353 390 509 424
rect 543 390 699 424
rect 733 390 879 424
rect 913 390 1069 424
rect 1103 390 1269 424
rect 1303 390 1469 424
rect 1503 390 1515 424
rect 117 384 1515 390
rect 217 350 1414 356
rect 217 316 229 350
rect 263 316 417 350
rect 451 316 605 350
rect 639 316 788 350
rect 822 316 970 350
rect 1004 316 1169 350
rect 1203 316 1368 350
rect 1402 316 1414 350
rect 217 310 1414 316
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
rlabel comment s 0 0 0 0 4 inv_16
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew
flabel nbase s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew
flabel metal1 s 117 384 1515 430 0 FreeSans 400 0 0 0 Y
port 6 nsew
flabel metal1 s 217 310 1414 356 0 FreeSans 400 0 0 0 A
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 1632 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1851672
string GDS_START 1837552
<< end >>
