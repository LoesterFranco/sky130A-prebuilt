magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 113 378 179 596
rect 313 378 379 596
rect 113 344 379 378
rect 113 310 179 344
rect 123 200 173 310
rect 513 294 647 360
rect 793 290 935 356
rect 985 290 1173 356
rect 1223 290 1415 356
rect 123 166 345 200
rect 123 70 173 166
rect 311 66 345 166
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 23 364 73 649
rect 213 412 279 649
rect 413 364 479 649
rect 525 562 815 596
rect 525 394 591 562
rect 625 394 715 528
rect 23 17 89 226
rect 213 260 467 310
rect 681 260 715 394
rect 749 424 815 562
rect 849 458 915 649
rect 949 424 1015 596
rect 1049 458 1115 649
rect 1151 424 1217 596
rect 1251 458 1317 649
rect 1351 424 1417 596
rect 749 390 1417 424
rect 213 256 718 260
rect 213 244 950 256
rect 379 226 950 244
rect 209 17 275 132
rect 386 17 452 192
rect 498 70 548 226
rect 684 222 950 226
rect 584 17 650 192
rect 684 70 750 222
rect 784 85 850 188
rect 884 119 950 222
rect 996 222 1406 256
rect 996 119 1046 222
rect 1082 85 1148 188
rect 784 51 1148 85
rect 1184 70 1218 222
rect 1254 17 1320 188
rect 1356 70 1406 222
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 683 1440 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 0 617 1440 649
rect 0 17 1440 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -49 1440 -17
<< labels >>
rlabel locali s 793 290 935 356 6 A1
port 1 nsew signal input
rlabel locali s 985 290 1173 356 6 A2
port 2 nsew signal input
rlabel locali s 1223 290 1415 356 6 A3
port 3 nsew signal input
rlabel locali s 513 294 647 360 6 B1
port 4 nsew signal input
rlabel locali s 313 378 379 596 6 X
port 5 nsew signal output
rlabel locali s 311 66 345 166 6 X
port 5 nsew signal output
rlabel locali s 123 200 173 310 6 X
port 5 nsew signal output
rlabel locali s 123 166 345 200 6 X
port 5 nsew signal output
rlabel locali s 123 70 173 166 6 X
port 5 nsew signal output
rlabel locali s 113 378 179 596 6 X
port 5 nsew signal output
rlabel locali s 113 344 379 378 6 X
port 5 nsew signal output
rlabel locali s 113 310 179 344 6 X
port 5 nsew signal output
rlabel metal1 s 0 -49 1440 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 1440 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1440 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3802782
string GDS_START 3789944
<< end >>
