magic
tech sky130A
magscale 1 2
timestamp 1604502710
<< nwell >>
rect -38 332 998 704
<< pwell >>
rect 0 0 960 49
<< scpmos >>
rect 83 368 119 592
rect 173 368 209 592
rect 313 368 349 568
rect 397 368 433 568
rect 505 368 541 568
rect 619 368 655 568
rect 733 368 769 568
<< nmoslvt >>
rect 119 74 149 222
rect 205 74 235 222
rect 319 74 349 222
rect 405 74 435 222
rect 519 74 549 222
rect 619 74 649 222
rect 832 74 862 222
<< ndiff >>
rect 27 206 119 222
rect 27 172 39 206
rect 73 172 119 206
rect 27 120 119 172
rect 27 86 74 120
rect 108 86 119 120
rect 27 74 119 86
rect 149 210 205 222
rect 149 176 160 210
rect 194 176 205 210
rect 149 120 205 176
rect 149 86 160 120
rect 194 86 205 120
rect 149 74 205 86
rect 235 210 319 222
rect 235 176 260 210
rect 294 176 319 210
rect 235 120 319 176
rect 235 86 260 120
rect 294 86 319 120
rect 235 74 319 86
rect 349 210 405 222
rect 349 176 360 210
rect 394 176 405 210
rect 349 120 405 176
rect 349 86 360 120
rect 394 86 405 120
rect 349 74 405 86
rect 435 152 519 222
rect 435 118 460 152
rect 494 118 519 152
rect 435 74 519 118
rect 549 210 619 222
rect 549 176 560 210
rect 594 176 619 210
rect 549 120 619 176
rect 549 86 560 120
rect 594 86 619 120
rect 549 74 619 86
rect 649 193 832 222
rect 649 159 660 193
rect 694 159 787 193
rect 821 159 832 193
rect 649 74 832 159
rect 862 186 933 222
rect 862 152 873 186
rect 907 152 933 186
rect 862 116 933 152
rect 862 82 873 116
rect 907 82 933 116
rect 862 74 933 82
<< pdiff >>
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 497 83 546
rect 27 463 39 497
rect 73 463 83 497
rect 27 414 83 463
rect 27 380 39 414
rect 73 380 83 414
rect 27 368 83 380
rect 119 580 173 592
rect 119 546 129 580
rect 163 546 173 580
rect 119 497 173 546
rect 119 463 129 497
rect 163 463 173 497
rect 119 414 173 463
rect 119 380 129 414
rect 163 380 173 414
rect 119 368 173 380
rect 209 568 259 592
rect 209 562 313 568
rect 209 528 219 562
rect 253 528 313 562
rect 209 494 313 528
rect 209 460 268 494
rect 302 460 313 494
rect 209 368 313 460
rect 349 368 397 568
rect 433 368 505 568
rect 541 560 619 568
rect 541 526 563 560
rect 597 526 619 560
rect 541 492 619 526
rect 541 458 563 492
rect 597 458 619 492
rect 541 424 619 458
rect 541 390 563 424
rect 597 390 619 424
rect 541 368 619 390
rect 655 368 733 568
rect 769 560 825 568
rect 769 526 779 560
rect 813 526 825 560
rect 769 492 825 526
rect 769 458 779 492
rect 813 458 825 492
rect 769 368 825 458
<< ndiffc >>
rect 39 172 73 206
rect 74 86 108 120
rect 160 176 194 210
rect 160 86 194 120
rect 260 176 294 210
rect 260 86 294 120
rect 360 176 394 210
rect 360 86 394 120
rect 460 118 494 152
rect 560 176 594 210
rect 560 86 594 120
rect 660 159 694 193
rect 787 159 821 193
rect 873 152 907 186
rect 873 82 907 116
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 129 546 163 580
rect 129 463 163 497
rect 129 380 163 414
rect 219 528 253 562
rect 268 460 302 494
rect 563 526 597 560
rect 563 458 597 492
rect 563 390 597 424
rect 779 526 813 560
rect 779 458 813 492
<< poly >>
rect 83 592 119 618
rect 173 592 209 618
rect 313 568 349 594
rect 397 568 433 594
rect 505 568 541 594
rect 619 568 655 594
rect 733 568 769 594
rect 83 294 119 368
rect 173 330 209 368
rect 313 345 349 368
rect 173 314 241 330
rect 173 294 191 314
rect 83 280 191 294
rect 225 280 241 314
rect 83 264 241 280
rect 283 320 349 345
rect 283 286 299 320
rect 333 286 349 320
rect 283 270 349 286
rect 397 336 433 368
rect 505 336 541 368
rect 619 336 655 368
rect 397 320 463 336
rect 397 286 413 320
rect 447 286 463 320
rect 397 270 463 286
rect 505 320 571 336
rect 505 286 521 320
rect 555 286 571 320
rect 505 270 571 286
rect 619 320 685 336
rect 619 286 635 320
rect 669 286 685 320
rect 619 270 685 286
rect 733 310 769 368
rect 733 294 937 310
rect 733 280 887 294
rect 119 222 149 264
rect 205 222 235 264
rect 319 222 349 270
rect 405 222 435 270
rect 519 222 549 270
rect 619 222 649 270
rect 832 260 887 280
rect 921 260 937 294
rect 832 244 937 260
rect 832 222 862 244
rect 119 48 149 74
rect 205 48 235 74
rect 319 48 349 74
rect 405 48 435 74
rect 519 48 549 74
rect 619 48 649 74
rect 832 48 862 74
<< polycont >>
rect 191 280 225 314
rect 299 286 333 320
rect 413 286 447 320
rect 521 286 555 320
rect 635 286 669 320
rect 887 260 921 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 23 580 73 649
rect 23 546 39 580
rect 23 497 73 546
rect 23 463 39 497
rect 23 414 73 463
rect 23 380 39 414
rect 23 364 73 380
rect 107 580 179 596
rect 107 546 129 580
rect 163 546 179 580
rect 107 497 179 546
rect 107 463 129 497
rect 163 463 179 497
rect 107 414 179 463
rect 213 562 320 649
rect 213 528 219 562
rect 253 528 320 562
rect 213 494 320 528
rect 213 460 268 494
rect 302 460 320 494
rect 213 458 320 460
rect 535 560 622 576
rect 535 526 563 560
rect 597 526 622 560
rect 535 492 622 526
rect 535 458 563 492
rect 597 458 622 492
rect 763 560 829 649
rect 763 526 779 560
rect 813 526 829 560
rect 763 492 829 526
rect 763 458 779 492
rect 813 458 829 492
rect 535 424 622 458
rect 107 380 129 414
rect 163 380 179 414
rect 107 364 179 380
rect 213 390 563 424
rect 597 390 837 424
rect 23 206 73 228
rect 23 172 39 206
rect 107 226 141 364
rect 213 330 247 390
rect 175 314 247 330
rect 175 280 191 314
rect 225 280 247 314
rect 175 264 247 280
rect 283 320 359 356
rect 283 286 299 320
rect 333 286 359 320
rect 283 270 359 286
rect 397 320 463 356
rect 397 286 413 320
rect 447 286 463 320
rect 397 270 463 286
rect 505 320 571 356
rect 505 286 521 320
rect 555 286 571 320
rect 505 270 571 286
rect 619 320 743 356
rect 619 286 635 320
rect 669 286 743 320
rect 619 270 743 286
rect 107 210 210 226
rect 107 192 160 210
rect 23 158 73 172
rect 144 176 160 192
rect 194 176 210 210
rect 23 120 108 158
rect 23 86 74 120
rect 23 17 108 86
rect 144 120 210 176
rect 144 86 160 120
rect 194 86 210 120
rect 144 70 210 86
rect 244 210 310 226
rect 244 176 260 210
rect 294 176 310 210
rect 244 120 310 176
rect 244 86 260 120
rect 294 86 310 120
rect 244 17 310 86
rect 344 210 610 236
rect 344 176 360 210
rect 394 202 560 210
rect 394 176 410 202
rect 344 120 410 176
rect 544 176 560 202
rect 594 176 610 210
rect 803 209 837 390
rect 871 294 937 578
rect 871 260 887 294
rect 921 260 937 294
rect 871 236 937 260
rect 344 86 360 120
rect 394 86 410 120
rect 344 70 410 86
rect 444 152 510 168
rect 444 118 460 152
rect 494 118 510 152
rect 444 17 510 118
rect 544 120 610 176
rect 644 193 837 209
rect 644 159 660 193
rect 694 159 787 193
rect 821 159 837 193
rect 644 143 837 159
rect 871 186 923 202
rect 871 152 873 186
rect 907 152 923 186
rect 544 86 560 120
rect 594 104 610 120
rect 871 116 923 152
rect 871 104 873 116
rect 594 86 873 104
rect 544 82 873 86
rect 907 82 923 116
rect 544 70 923 82
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
rlabel comment s 0 0 0 0 4 o32a_2
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 895 242 929 276 0 FreeSans 340 0 0 0 B1
port 4 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 B1
port 4 nsew
flabel corelocali s 895 390 929 424 0 FreeSans 340 0 0 0 B1
port 4 nsew
flabel corelocali s 895 464 929 498 0 FreeSans 340 0 0 0 B1
port 4 nsew
flabel corelocali s 895 538 929 572 0 FreeSans 340 0 0 0 B1
port 4 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 B2
port 5 nsew
flabel corelocali s 127 390 161 424 0 FreeSans 340 0 0 0 X
port 10 nsew
flabel corelocali s 127 464 161 498 0 FreeSans 340 0 0 0 X
port 10 nsew
flabel corelocali s 127 538 161 572 0 FreeSans 340 0 0 0 X
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 960 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 665538
string GDS_START 657422
<< end >>
