magic
tech sky130A
magscale 1 2
timestamp 1599588218
<< nwell >>
rect -38 332 1190 704
<< pwell >>
rect 0 0 1152 49
<< scpmos >>
rect 82 392 118 592
rect 184 392 220 592
rect 274 392 310 592
rect 376 392 412 592
rect 471 392 507 592
rect 561 392 597 592
rect 663 392 699 592
rect 765 368 801 592
rect 855 368 891 592
rect 945 368 981 592
rect 1035 368 1071 592
<< nmoslvt >>
rect 88 136 118 264
rect 477 74 507 222
rect 577 74 607 222
rect 663 74 693 222
rect 765 74 795 222
rect 856 74 886 222
rect 952 74 982 222
rect 1038 74 1068 222
<< ndiff >>
rect 31 232 88 264
rect 31 198 43 232
rect 77 198 88 232
rect 31 136 88 198
rect 118 136 278 264
rect 193 112 278 136
rect 193 78 218 112
rect 252 78 278 112
rect 193 66 278 78
rect 421 196 477 222
rect 421 162 432 196
rect 466 162 477 196
rect 421 120 477 162
rect 421 86 432 120
rect 466 86 477 120
rect 421 74 477 86
rect 507 124 577 222
rect 507 90 532 124
rect 566 90 577 124
rect 507 74 577 90
rect 607 196 663 222
rect 607 162 618 196
rect 652 162 663 196
rect 607 120 663 162
rect 607 86 618 120
rect 652 86 663 120
rect 607 74 663 86
rect 693 120 765 222
rect 693 86 719 120
rect 753 86 765 120
rect 693 74 765 86
rect 795 210 856 222
rect 795 176 811 210
rect 845 176 856 210
rect 795 120 856 176
rect 795 86 811 120
rect 845 86 856 120
rect 795 74 856 86
rect 886 136 952 222
rect 886 102 897 136
rect 931 102 952 136
rect 886 74 952 102
rect 982 210 1038 222
rect 982 176 993 210
rect 1027 176 1038 210
rect 982 120 1038 176
rect 982 86 993 120
rect 1027 86 1038 120
rect 982 74 1038 86
rect 1068 142 1125 222
rect 1068 108 1079 142
rect 1113 108 1125 142
rect 1068 74 1125 108
<< pdiff >>
rect 27 580 82 592
rect 27 546 38 580
rect 72 546 82 580
rect 27 509 82 546
rect 27 475 38 509
rect 72 475 82 509
rect 27 438 82 475
rect 27 404 38 438
rect 72 404 82 438
rect 27 392 82 404
rect 118 580 184 592
rect 118 546 128 580
rect 162 546 184 580
rect 118 509 184 546
rect 118 475 128 509
rect 162 475 184 509
rect 118 438 184 475
rect 118 404 128 438
rect 162 404 184 438
rect 118 392 184 404
rect 220 580 274 592
rect 220 546 230 580
rect 264 546 274 580
rect 220 512 274 546
rect 220 478 230 512
rect 264 478 274 512
rect 220 444 274 478
rect 220 410 230 444
rect 264 410 274 444
rect 220 392 274 410
rect 310 577 376 592
rect 310 543 332 577
rect 366 543 376 577
rect 310 392 376 543
rect 412 438 471 592
rect 412 404 424 438
rect 458 404 471 438
rect 412 392 471 404
rect 507 577 561 592
rect 507 543 517 577
rect 551 543 561 577
rect 507 392 561 543
rect 597 580 663 592
rect 597 546 617 580
rect 651 546 663 580
rect 597 512 663 546
rect 597 478 617 512
rect 651 478 663 512
rect 597 392 663 478
rect 699 580 765 592
rect 699 546 717 580
rect 751 546 765 580
rect 699 512 765 546
rect 699 478 717 512
rect 751 478 765 512
rect 699 392 765 478
rect 715 368 765 392
rect 801 580 855 592
rect 801 546 811 580
rect 845 546 855 580
rect 801 497 855 546
rect 801 463 811 497
rect 845 463 855 497
rect 801 414 855 463
rect 801 380 811 414
rect 845 380 855 414
rect 801 368 855 380
rect 891 580 945 592
rect 891 546 901 580
rect 935 546 945 580
rect 891 478 945 546
rect 891 444 901 478
rect 935 444 945 478
rect 891 368 945 444
rect 981 580 1035 592
rect 981 546 991 580
rect 1025 546 1035 580
rect 981 497 1035 546
rect 981 463 991 497
rect 1025 463 1035 497
rect 981 414 1035 463
rect 981 380 991 414
rect 1025 380 1035 414
rect 981 368 1035 380
rect 1071 580 1125 592
rect 1071 546 1081 580
rect 1115 546 1125 580
rect 1071 478 1125 546
rect 1071 444 1081 478
rect 1115 444 1125 478
rect 1071 368 1125 444
<< ndiffc >>
rect 43 198 77 232
rect 218 78 252 112
rect 432 162 466 196
rect 432 86 466 120
rect 532 90 566 124
rect 618 162 652 196
rect 618 86 652 120
rect 719 86 753 120
rect 811 176 845 210
rect 811 86 845 120
rect 897 102 931 136
rect 993 176 1027 210
rect 993 86 1027 120
rect 1079 108 1113 142
<< pdiffc >>
rect 38 546 72 580
rect 38 475 72 509
rect 38 404 72 438
rect 128 546 162 580
rect 128 475 162 509
rect 128 404 162 438
rect 230 546 264 580
rect 230 478 264 512
rect 230 410 264 444
rect 332 543 366 577
rect 424 404 458 438
rect 517 543 551 577
rect 617 546 651 580
rect 617 478 651 512
rect 717 546 751 580
rect 717 478 751 512
rect 811 546 845 580
rect 811 463 845 497
rect 811 380 845 414
rect 901 546 935 580
rect 901 444 935 478
rect 991 546 1025 580
rect 991 463 1025 497
rect 991 380 1025 414
rect 1081 546 1115 580
rect 1081 444 1115 478
<< poly >>
rect 82 592 118 618
rect 184 592 220 618
rect 274 592 310 618
rect 376 592 412 618
rect 471 592 507 618
rect 561 592 597 618
rect 663 592 699 618
rect 765 592 801 618
rect 855 592 891 618
rect 945 592 981 618
rect 1035 592 1071 618
rect 82 279 118 392
rect 184 352 220 392
rect 274 360 310 392
rect 160 336 226 352
rect 160 302 176 336
rect 210 302 226 336
rect 160 286 226 302
rect 268 344 334 360
rect 268 310 284 344
rect 318 310 334 344
rect 268 294 334 310
rect 88 264 118 279
rect 376 267 412 392
rect 471 267 507 392
rect 561 360 597 392
rect 549 344 615 360
rect 549 310 565 344
rect 599 310 615 344
rect 663 310 699 392
rect 765 326 801 368
rect 855 326 891 368
rect 945 326 981 368
rect 1035 326 1071 368
rect 765 310 1071 326
rect 549 294 615 310
rect 657 294 723 310
rect 376 237 507 267
rect 376 196 406 237
rect 477 222 507 237
rect 577 222 607 294
rect 657 260 673 294
rect 707 260 723 294
rect 657 244 723 260
rect 765 276 781 310
rect 815 276 849 310
rect 883 276 917 310
rect 951 276 985 310
rect 1019 276 1071 310
rect 765 260 1071 276
rect 663 222 693 244
rect 765 222 795 260
rect 856 222 886 260
rect 952 222 982 260
rect 1038 222 1068 260
rect 88 114 118 136
rect 21 98 155 114
rect 21 64 37 98
rect 71 64 105 98
rect 139 64 155 98
rect 316 180 406 196
rect 316 146 332 180
rect 366 146 406 180
rect 316 112 406 146
rect 316 78 332 112
rect 366 78 406 112
rect 21 48 155 64
rect 316 62 406 78
rect 477 48 507 74
rect 577 48 607 74
rect 663 48 693 74
rect 765 48 795 74
rect 856 48 886 74
rect 952 48 982 74
rect 1038 48 1068 74
<< polycont >>
rect 176 302 210 336
rect 284 310 318 344
rect 565 310 599 344
rect 673 260 707 294
rect 781 276 815 310
rect 849 276 883 310
rect 917 276 951 310
rect 985 276 1019 310
rect 37 64 71 98
rect 105 64 139 98
rect 332 146 366 180
rect 332 78 366 112
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 22 580 72 596
rect 22 546 38 580
rect 22 509 72 546
rect 22 475 38 509
rect 22 438 72 475
rect 22 404 38 438
rect 22 268 72 404
rect 112 580 178 649
rect 112 546 128 580
rect 162 546 178 580
rect 112 509 178 546
rect 112 475 128 509
rect 162 475 178 509
rect 112 438 178 475
rect 112 404 128 438
rect 162 404 178 438
rect 112 388 178 404
rect 214 580 280 596
rect 214 546 230 580
rect 264 546 280 580
rect 214 512 280 546
rect 316 577 567 596
rect 316 543 332 577
rect 366 543 517 577
rect 551 543 567 577
rect 316 540 567 543
rect 601 580 667 596
rect 601 546 617 580
rect 651 546 667 580
rect 214 478 230 512
rect 264 506 280 512
rect 601 512 667 546
rect 601 506 617 512
rect 264 478 617 506
rect 651 478 667 512
rect 214 472 667 478
rect 214 444 280 472
rect 601 462 667 472
rect 701 580 767 649
rect 701 546 717 580
rect 751 546 767 580
rect 701 512 767 546
rect 701 478 717 512
rect 751 478 767 512
rect 701 462 767 478
rect 811 580 845 596
rect 811 497 845 546
rect 214 410 230 444
rect 264 410 280 444
rect 214 394 280 410
rect 406 404 424 438
rect 458 428 477 438
rect 458 404 777 428
rect 406 394 777 404
rect 160 336 226 352
rect 160 302 176 336
rect 210 302 226 336
rect 22 232 93 268
rect 22 198 43 232
rect 77 198 93 232
rect 160 264 226 302
rect 268 344 615 360
rect 268 310 284 344
rect 318 310 565 344
rect 599 310 615 344
rect 743 326 777 394
rect 811 414 845 463
rect 885 580 935 649
rect 885 546 901 580
rect 885 478 935 546
rect 885 444 901 478
rect 885 428 935 444
rect 975 580 1041 596
rect 975 546 991 580
rect 1025 546 1041 580
rect 975 497 1041 546
rect 975 463 991 497
rect 1025 463 1041 497
rect 975 414 1041 463
rect 1081 580 1131 649
rect 1115 546 1131 580
rect 1081 478 1131 546
rect 1115 444 1131 478
rect 1081 428 1131 444
rect 975 394 991 414
rect 845 380 991 394
rect 1025 394 1041 414
rect 1025 380 1127 394
rect 811 360 1127 380
rect 743 310 1035 326
rect 268 298 334 310
rect 657 294 709 310
rect 657 276 673 294
rect 601 264 673 276
rect 160 260 673 264
rect 707 260 709 294
rect 160 230 709 260
rect 743 276 781 310
rect 815 276 849 310
rect 883 276 917 310
rect 951 276 985 310
rect 1019 276 1035 310
rect 743 260 1035 276
rect 22 196 93 198
rect 743 196 777 260
rect 1081 226 1127 360
rect 22 180 382 196
rect 22 162 332 180
rect 316 146 332 162
rect 366 146 382 180
rect 21 98 155 128
rect 21 64 37 98
rect 71 64 105 98
rect 139 64 155 98
rect 21 51 155 64
rect 189 112 282 128
rect 189 78 218 112
rect 252 78 282 112
rect 189 17 282 78
rect 316 112 382 146
rect 316 78 332 112
rect 366 78 382 112
rect 316 62 382 78
rect 416 162 432 196
rect 466 162 618 196
rect 652 162 777 196
rect 811 210 1127 226
rect 845 192 993 210
rect 416 120 482 162
rect 416 86 432 120
rect 466 86 482 120
rect 416 70 482 86
rect 516 124 582 128
rect 516 90 532 124
rect 566 90 582 124
rect 516 17 582 90
rect 618 120 668 162
rect 811 120 845 176
rect 977 176 993 192
rect 1027 192 1127 210
rect 652 86 668 120
rect 618 70 668 86
rect 702 86 719 120
rect 753 86 770 120
rect 702 17 770 86
rect 811 70 845 86
rect 881 136 931 158
rect 881 102 897 136
rect 881 17 931 102
rect 977 120 1027 176
rect 977 86 993 120
rect 977 70 1027 86
rect 1063 142 1129 158
rect 1063 108 1079 142
rect 1113 108 1129 142
rect 1063 17 1129 108
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
rlabel comment s 0 0 0 0 4 or3b_4
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 607 242 641 276 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 31 94 65 128 0 FreeSans 340 0 0 0 C_N
port 3 nsew
flabel corelocali s 1087 242 1121 276 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 1087 316 1121 350 0 FreeSans 340 0 0 0 X
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 1152 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 823870
string GDS_START 814030
<< end >>
