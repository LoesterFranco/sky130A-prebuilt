magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 644 561
rect 58 439 124 527
rect 158 405 205 493
rect 242 451 308 527
rect 350 405 419 493
rect 17 357 419 405
rect 17 177 63 357
rect 454 323 523 474
rect 557 359 623 527
rect 97 215 163 323
rect 17 51 138 177
rect 205 51 271 323
rect 305 199 363 323
rect 397 199 523 323
rect 557 201 623 323
rect 457 17 523 91
rect 0 -17 644 17
<< obsli1 >>
rect 350 125 623 165
rect 350 51 419 125
rect 557 51 623 125
<< metal1 >>
rect 0 496 644 592
rect 0 -48 644 48
<< labels >>
rlabel locali s 557 201 623 323 6 A1
port 1 nsew signal input
rlabel locali s 454 323 523 474 6 A2
port 2 nsew signal input
rlabel locali s 397 199 523 323 6 A2
port 2 nsew signal input
rlabel locali s 305 199 363 323 6 B1
port 3 nsew signal input
rlabel locali s 205 51 271 323 6 C1
port 4 nsew signal input
rlabel locali s 97 215 163 323 6 D1
port 5 nsew signal input
rlabel locali s 350 405 419 493 6 Y
port 6 nsew signal output
rlabel locali s 158 405 205 493 6 Y
port 6 nsew signal output
rlabel locali s 17 357 419 405 6 Y
port 6 nsew signal output
rlabel locali s 17 177 63 357 6 Y
port 6 nsew signal output
rlabel locali s 17 51 138 177 6 Y
port 6 nsew signal output
rlabel locali s 457 17 523 91 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 644 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 644 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 557 359 623 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 242 451 308 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 58 439 124 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 644 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 644 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1254158
string GDS_START 1248122
<< end >>
