magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 132 425 572 483
rect 17 151 85 265
rect 324 199 482 323
rect 724 299 799 493
rect 526 199 615 265
rect 745 152 799 299
rect 724 83 799 152
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 17 312 85 527
rect 129 265 177 384
rect 216 357 572 391
rect 616 367 672 527
rect 216 299 280 357
rect 538 333 572 357
rect 129 199 260 265
rect 538 299 683 333
rect 649 265 683 299
rect 649 199 701 265
rect 17 17 85 117
rect 129 61 178 199
rect 649 165 683 199
rect 333 131 683 165
rect 217 17 283 117
rect 333 61 367 131
rect 402 17 478 97
rect 522 61 556 131
rect 590 17 676 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
rlabel locali s 526 199 615 265 6 A
port 1 nsew signal input
rlabel locali s 132 425 572 483 6 B
port 2 nsew signal input
rlabel locali s 324 199 482 323 6 C
port 3 nsew signal input
rlabel locali s 17 151 85 265 6 D_N
port 4 nsew signal input
rlabel locali s 745 152 799 299 6 X
port 5 nsew signal output
rlabel locali s 724 299 799 493 6 X
port 5 nsew signal output
rlabel locali s 724 83 799 152 6 X
port 5 nsew signal output
rlabel metal1 s 0 -48 828 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 828 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 520464
string GDS_START 513080
<< end >>
