magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1012 561
rect 103 451 169 527
rect 271 451 337 527
rect 455 435 505 527
rect 543 451 995 485
rect 950 357 995 451
rect 86 199 156 265
rect 494 215 712 255
rect 862 199 927 323
rect 116 145 156 199
rect 103 17 167 109
rect 287 17 337 177
rect 455 17 489 109
rect 961 93 995 357
rect 543 59 995 93
rect 0 -17 1012 17
<< obsli1 >>
rect 17 427 69 493
rect 371 427 416 493
rect 17 333 52 427
rect 382 401 416 427
rect 543 401 870 417
rect 187 367 347 401
rect 382 383 870 401
rect 382 367 577 383
rect 313 333 347 367
rect 627 333 693 343
rect 17 299 279 333
rect 313 299 693 333
rect 17 135 52 299
rect 245 265 279 299
rect 245 231 397 265
rect 331 215 397 231
rect 203 153 214 187
rect 248 153 251 187
rect 17 69 69 135
rect 203 115 251 153
rect 371 147 693 181
rect 371 59 405 147
rect 627 131 693 147
rect 804 165 821 187
rect 804 153 869 165
rect 770 131 869 153
<< obsli1c >>
rect 214 153 248 187
rect 770 153 804 187
<< metal1 >>
rect 0 496 1012 592
rect 0 -48 1012 48
<< obsm1 >>
rect 202 187 260 193
rect 202 153 214 187
rect 248 184 260 187
rect 758 187 816 193
rect 758 184 770 187
rect 248 156 770 184
rect 248 153 260 156
rect 202 147 260 153
rect 758 153 770 156
rect 804 153 816 187
rect 758 147 816 153
<< labels >>
rlabel locali s 494 215 712 255 6 A0
port 1 nsew signal input
rlabel locali s 862 199 927 323 6 A1
port 2 nsew signal input
rlabel locali s 116 145 156 199 6 S
port 3 nsew signal input
rlabel locali s 86 199 156 265 6 S
port 3 nsew signal input
rlabel locali s 961 93 995 357 6 Y
port 4 nsew signal output
rlabel locali s 950 357 995 451 6 Y
port 4 nsew signal output
rlabel locali s 543 451 995 485 6 Y
port 4 nsew signal output
rlabel locali s 543 59 995 93 6 Y
port 4 nsew signal output
rlabel locali s 455 17 489 109 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 287 17 337 177 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 103 17 167 109 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 1012 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1012 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 455 435 505 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 271 451 337 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 103 451 169 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 1012 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 1012 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1012 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1686858
string GDS_START 1678844
<< end >>
