magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 19 53 71 491
rect 213 203 322 265
rect 356 203 443 265
rect 397 75 443 203
rect 482 199 532 265
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 105 381 183 527
rect 219 345 273 491
rect 109 301 273 345
rect 319 349 365 491
rect 401 385 477 527
rect 521 349 573 491
rect 319 301 573 349
rect 109 167 177 301
rect 109 127 363 167
rect 133 17 267 91
rect 303 53 363 127
rect 515 17 573 163
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 397 75 443 203 6 A1
port 1 nsew signal input
rlabel locali s 356 203 443 265 6 A1
port 1 nsew signal input
rlabel locali s 482 199 532 265 6 A2
port 2 nsew signal input
rlabel locali s 213 203 322 265 6 B1
port 3 nsew signal input
rlabel locali s 19 53 71 491 6 X
port 4 nsew signal output
rlabel metal1 s 0 -48 644 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1180152
string GDS_START 1173906
<< end >>
