magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 17 199 90 335
rect 335 84 431 339
rect 465 84 523 339
rect 557 133 615 339
rect 727 299 799 493
rect 745 161 799 299
rect 704 59 799 161
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 34 403 69 493
rect 103 439 179 527
rect 240 409 274 493
rect 331 445 475 527
rect 526 409 560 493
rect 612 445 678 527
rect 34 369 170 403
rect 136 265 170 369
rect 240 375 683 409
rect 136 199 205 265
rect 136 165 170 199
rect 34 131 170 165
rect 34 51 69 131
rect 240 117 274 375
rect 103 17 179 93
rect 228 51 274 117
rect 649 265 683 375
rect 649 199 707 265
rect 591 17 670 93
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
rlabel locali s 17 199 90 335 6 A_N
port 1 nsew signal input
rlabel locali s 335 84 431 339 6 B
port 2 nsew signal input
rlabel locali s 465 84 523 339 6 C
port 3 nsew signal input
rlabel locali s 557 133 615 339 6 D
port 4 nsew signal input
rlabel locali s 745 161 799 299 6 X
port 5 nsew signal output
rlabel locali s 727 299 799 493 6 X
port 5 nsew signal output
rlabel locali s 704 59 799 161 6 X
port 5 nsew signal output
rlabel metal1 s 0 -48 828 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 828 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1581260
string GDS_START 1573514
<< end >>
