magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 736 561
rect 18 383 85 485
rect 18 112 69 383
rect 135 367 201 527
rect 358 443 424 527
rect 665 265 706 323
rect 214 199 264 265
rect 306 133 360 265
rect 398 133 456 265
rect 490 132 574 265
rect 636 199 706 265
rect 18 60 85 112
rect 119 17 185 97
rect 651 17 717 161
rect 0 -17 736 17
<< obsli1 >>
rect 250 409 307 493
rect 469 459 701 493
rect 469 409 535 459
rect 250 375 535 409
rect 581 333 615 425
rect 667 359 701 459
rect 141 299 615 333
rect 141 265 175 299
rect 114 199 175 265
rect 141 165 175 199
rect 141 131 253 165
rect 219 97 253 131
rect 219 63 542 97
<< metal1 >>
rect 0 496 736 592
rect 0 -48 736 48
<< labels >>
rlabel locali s 398 133 456 265 6 A1
port 1 nsew signal input
rlabel locali s 306 133 360 265 6 A2
port 2 nsew signal input
rlabel locali s 214 199 264 265 6 A3
port 3 nsew signal input
rlabel locali s 490 132 574 265 6 B1
port 4 nsew signal input
rlabel locali s 665 265 706 323 6 B2
port 5 nsew signal input
rlabel locali s 636 199 706 265 6 B2
port 5 nsew signal input
rlabel locali s 18 383 85 485 6 X
port 6 nsew signal output
rlabel locali s 18 112 69 383 6 X
port 6 nsew signal output
rlabel locali s 18 60 85 112 6 X
port 6 nsew signal output
rlabel locali s 651 17 717 161 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 119 17 185 97 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 736 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 736 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 358 443 424 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 135 367 201 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 736 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 736 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3620700
string GDS_START 3613326
<< end >>
