magic
tech sky130A
magscale 1 2
timestamp 1604502710
<< nwell >>
rect -38 332 1958 704
rect 277 330 1074 332
rect 854 315 1074 330
<< pwell >>
rect 0 0 1920 49
<< scpmos >>
rect 83 395 119 563
rect 167 395 203 563
rect 426 424 462 592
rect 645 379 681 547
rect 752 455 788 539
rect 836 455 872 539
rect 946 351 982 575
rect 1149 368 1185 536
rect 1256 368 1292 592
rect 1385 368 1421 592
rect 1485 368 1521 592
rect 1601 368 1637 592
rect 1701 368 1737 592
rect 1800 368 1836 592
<< nmoslvt >>
rect 89 143 119 253
rect 184 143 214 253
rect 324 105 354 253
rect 604 74 634 184
rect 714 74 744 158
rect 792 74 822 158
rect 964 74 994 222
rect 1162 74 1192 222
rect 1262 74 1292 222
rect 1340 74 1370 222
rect 1538 74 1568 222
rect 1634 74 1664 222
rect 1720 74 1750 222
rect 1806 74 1836 222
<< ndiff >>
rect 27 215 89 253
rect 27 181 39 215
rect 73 181 89 215
rect 27 143 89 181
rect 119 215 184 253
rect 119 181 139 215
rect 173 181 184 215
rect 119 143 184 181
rect 214 143 324 253
rect 229 105 324 143
rect 354 241 411 253
rect 354 207 365 241
rect 399 207 411 241
rect 354 105 411 207
rect 465 141 604 184
rect 465 107 488 141
rect 522 107 604 141
rect 229 73 309 105
rect 465 74 604 107
rect 634 172 699 184
rect 634 138 649 172
rect 683 158 699 172
rect 914 158 964 222
rect 683 138 714 158
rect 634 74 714 138
rect 744 74 792 158
rect 822 124 964 158
rect 822 90 837 124
rect 871 90 964 124
rect 822 74 964 90
rect 994 183 1051 222
rect 994 149 1005 183
rect 1039 149 1051 183
rect 994 74 1051 149
rect 1105 202 1162 222
rect 1105 168 1117 202
rect 1151 168 1162 202
rect 1105 120 1162 168
rect 1105 86 1117 120
rect 1151 86 1162 120
rect 1105 74 1162 86
rect 1192 202 1262 222
rect 1192 168 1217 202
rect 1251 168 1262 202
rect 1192 120 1262 168
rect 1192 86 1217 120
rect 1251 86 1262 120
rect 1192 74 1262 86
rect 1292 74 1340 222
rect 1370 210 1427 222
rect 1370 176 1381 210
rect 1415 176 1427 210
rect 1370 120 1427 176
rect 1370 86 1381 120
rect 1415 86 1427 120
rect 1370 74 1427 86
rect 1481 131 1538 222
rect 1481 97 1493 131
rect 1527 97 1538 131
rect 1481 74 1538 97
rect 1568 210 1634 222
rect 1568 176 1589 210
rect 1623 176 1634 210
rect 1568 120 1634 176
rect 1568 86 1589 120
rect 1623 86 1634 120
rect 1568 74 1634 86
rect 1664 131 1720 222
rect 1664 97 1675 131
rect 1709 97 1720 131
rect 1664 74 1720 97
rect 1750 210 1806 222
rect 1750 176 1761 210
rect 1795 176 1806 210
rect 1750 120 1806 176
rect 1750 86 1761 120
rect 1795 86 1806 120
rect 1750 74 1806 86
rect 1836 210 1893 222
rect 1836 176 1847 210
rect 1881 176 1893 210
rect 1836 120 1893 176
rect 1836 86 1847 120
rect 1881 86 1893 120
rect 1836 74 1893 86
rect 229 39 252 73
rect 286 39 309 73
rect 229 27 309 39
<< pdiff >>
rect 313 572 426 592
rect 27 551 83 563
rect 27 517 39 551
rect 73 517 83 551
rect 27 441 83 517
rect 27 407 39 441
rect 73 407 83 441
rect 27 395 83 407
rect 119 395 167 563
rect 203 551 259 563
rect 203 517 213 551
rect 247 517 259 551
rect 203 441 259 517
rect 203 407 213 441
rect 247 407 259 441
rect 313 538 381 572
rect 415 538 426 572
rect 313 424 426 538
rect 462 424 535 592
rect 203 395 259 407
rect 477 412 535 424
rect 477 378 489 412
rect 523 378 535 412
rect 589 535 645 547
rect 589 501 601 535
rect 635 501 645 535
rect 589 431 645 501
rect 589 397 601 431
rect 635 397 645 431
rect 589 379 645 397
rect 681 539 737 547
rect 890 563 946 575
rect 890 539 902 563
rect 681 535 752 539
rect 681 501 691 535
rect 725 501 752 535
rect 681 455 752 501
rect 788 455 836 539
rect 872 529 902 539
rect 936 529 946 563
rect 872 465 946 529
rect 872 455 902 465
rect 681 431 737 455
rect 681 397 691 431
rect 725 397 737 431
rect 681 379 737 397
rect 477 366 535 378
rect 890 431 902 455
rect 936 431 946 465
rect 890 351 946 431
rect 982 563 1038 575
rect 982 529 992 563
rect 1026 529 1038 563
rect 1200 566 1256 592
rect 1200 536 1212 566
rect 982 480 1038 529
rect 982 446 992 480
rect 1026 446 1038 480
rect 982 397 1038 446
rect 982 363 992 397
rect 1026 363 1038 397
rect 1092 414 1149 536
rect 1092 380 1104 414
rect 1138 380 1149 414
rect 1092 368 1149 380
rect 1185 532 1212 536
rect 1246 532 1256 566
rect 1185 368 1256 532
rect 1292 580 1385 592
rect 1292 546 1341 580
rect 1375 546 1385 580
rect 1292 497 1385 546
rect 1292 463 1341 497
rect 1375 463 1385 497
rect 1292 414 1385 463
rect 1292 380 1341 414
rect 1375 380 1385 414
rect 1292 368 1385 380
rect 1421 580 1485 592
rect 1421 546 1441 580
rect 1475 546 1485 580
rect 1421 478 1485 546
rect 1421 444 1441 478
rect 1475 444 1485 478
rect 1421 368 1485 444
rect 1521 580 1601 592
rect 1521 546 1557 580
rect 1591 546 1601 580
rect 1521 497 1601 546
rect 1521 463 1557 497
rect 1591 463 1601 497
rect 1521 414 1601 463
rect 1521 380 1557 414
rect 1591 380 1601 414
rect 1521 368 1601 380
rect 1637 580 1701 592
rect 1637 546 1647 580
rect 1681 546 1701 580
rect 1637 478 1701 546
rect 1637 444 1647 478
rect 1681 444 1701 478
rect 1637 368 1701 444
rect 1737 580 1800 592
rect 1737 546 1747 580
rect 1781 546 1800 580
rect 1737 497 1800 546
rect 1737 463 1747 497
rect 1781 463 1800 497
rect 1737 414 1800 463
rect 1737 380 1747 414
rect 1781 380 1800 414
rect 1737 368 1800 380
rect 1836 580 1893 592
rect 1836 546 1847 580
rect 1881 546 1893 580
rect 1836 497 1893 546
rect 1836 463 1847 497
rect 1881 463 1893 497
rect 1836 414 1893 463
rect 1836 380 1847 414
rect 1881 380 1893 414
rect 1836 368 1893 380
rect 982 351 1038 363
<< ndiffc >>
rect 39 181 73 215
rect 139 181 173 215
rect 365 207 399 241
rect 488 107 522 141
rect 649 138 683 172
rect 837 90 871 124
rect 1005 149 1039 183
rect 1117 168 1151 202
rect 1117 86 1151 120
rect 1217 168 1251 202
rect 1217 86 1251 120
rect 1381 176 1415 210
rect 1381 86 1415 120
rect 1493 97 1527 131
rect 1589 176 1623 210
rect 1589 86 1623 120
rect 1675 97 1709 131
rect 1761 176 1795 210
rect 1761 86 1795 120
rect 1847 176 1881 210
rect 1847 86 1881 120
rect 252 39 286 73
<< pdiffc >>
rect 39 517 73 551
rect 39 407 73 441
rect 213 517 247 551
rect 213 407 247 441
rect 381 538 415 572
rect 489 378 523 412
rect 601 501 635 535
rect 601 397 635 431
rect 691 501 725 535
rect 902 529 936 563
rect 691 397 725 431
rect 902 431 936 465
rect 992 529 1026 563
rect 992 446 1026 480
rect 992 363 1026 397
rect 1104 380 1138 414
rect 1212 532 1246 566
rect 1341 546 1375 580
rect 1341 463 1375 497
rect 1341 380 1375 414
rect 1441 546 1475 580
rect 1441 444 1475 478
rect 1557 546 1591 580
rect 1557 463 1591 497
rect 1557 380 1591 414
rect 1647 546 1681 580
rect 1647 444 1681 478
rect 1747 546 1781 580
rect 1747 463 1781 497
rect 1747 380 1781 414
rect 1847 546 1881 580
rect 1847 463 1881 497
rect 1847 380 1881 414
<< poly >>
rect 426 615 788 645
rect 426 592 462 615
rect 83 563 119 589
rect 167 563 203 589
rect 645 547 681 573
rect 83 357 119 395
rect 44 341 119 357
rect 44 307 60 341
rect 94 307 119 341
rect 44 291 119 307
rect 167 357 203 395
rect 167 341 233 357
rect 167 307 183 341
rect 217 307 233 341
rect 167 291 233 307
rect 426 298 462 424
rect 752 539 788 615
rect 946 575 982 601
rect 1256 592 1292 618
rect 1385 592 1421 618
rect 1485 592 1521 618
rect 1601 592 1637 618
rect 1701 592 1737 618
rect 1800 592 1836 618
rect 836 539 872 565
rect 752 429 788 455
rect 836 381 872 455
rect 645 347 681 379
rect 585 331 681 347
rect 89 253 119 291
rect 184 253 214 291
rect 324 268 515 298
rect 585 297 601 331
rect 635 311 681 331
rect 792 365 872 381
rect 792 331 808 365
rect 842 331 872 365
rect 1149 536 1185 562
rect 792 315 872 331
rect 635 297 744 311
rect 585 281 744 297
rect 324 253 354 268
rect 426 263 515 268
rect 89 117 119 143
rect 184 117 214 143
rect 426 229 465 263
rect 499 239 515 263
rect 499 229 634 239
rect 426 209 634 229
rect 604 184 634 209
rect 324 79 354 105
rect 714 158 744 281
rect 792 158 822 315
rect 946 313 982 351
rect 920 297 994 313
rect 920 263 936 297
rect 970 263 994 297
rect 920 247 994 263
rect 964 222 994 247
rect 1149 310 1185 368
rect 1256 310 1292 368
rect 1385 326 1421 368
rect 1149 294 1292 310
rect 1149 260 1173 294
rect 1207 260 1292 294
rect 1149 244 1292 260
rect 1162 222 1192 244
rect 1262 222 1292 244
rect 1340 310 1421 326
rect 1340 276 1356 310
rect 1390 276 1421 310
rect 1340 260 1421 276
rect 1485 326 1521 368
rect 1601 326 1637 368
rect 1701 326 1737 368
rect 1800 326 1836 368
rect 1485 310 1836 326
rect 1485 276 1501 310
rect 1535 276 1569 310
rect 1603 276 1637 310
rect 1671 276 1836 310
rect 1485 260 1836 276
rect 1340 222 1370 260
rect 1538 222 1568 260
rect 1634 222 1664 260
rect 1720 222 1750 260
rect 1806 222 1836 260
rect 604 48 634 74
rect 714 48 744 74
rect 792 48 822 74
rect 964 48 994 74
rect 1162 48 1192 74
rect 1262 48 1292 74
rect 1340 48 1370 74
rect 1538 48 1568 74
rect 1634 48 1664 74
rect 1720 48 1750 74
rect 1806 48 1836 74
<< polycont >>
rect 60 307 94 341
rect 183 307 217 341
rect 601 297 635 331
rect 808 331 842 365
rect 465 229 499 263
rect 936 263 970 297
rect 1173 260 1207 294
rect 1356 276 1390 310
rect 1501 276 1535 310
rect 1569 276 1603 310
rect 1637 276 1671 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 23 551 89 649
rect 309 572 432 649
rect 23 517 39 551
rect 73 517 89 551
rect 23 441 89 517
rect 23 407 39 441
rect 73 407 89 441
rect 23 391 89 407
rect 197 551 263 567
rect 197 517 213 551
rect 247 517 263 551
rect 309 538 381 572
rect 415 538 432 572
rect 886 563 936 649
rect 309 530 432 538
rect 585 535 651 551
rect 197 496 263 517
rect 585 501 601 535
rect 635 501 651 535
rect 585 496 651 501
rect 197 462 651 496
rect 197 441 331 462
rect 197 407 213 441
rect 247 407 331 441
rect 585 431 651 462
rect 197 391 331 407
rect 25 341 110 357
rect 25 307 60 341
rect 94 307 110 341
rect 25 291 110 307
rect 167 341 263 357
rect 167 307 183 341
rect 217 307 263 341
rect 167 291 263 307
rect 23 215 89 257
rect 23 181 39 215
rect 73 181 89 215
rect 23 17 89 181
rect 123 215 189 257
rect 123 181 139 215
rect 173 181 189 215
rect 123 157 189 181
rect 297 157 331 391
rect 473 412 539 428
rect 473 378 489 412
rect 523 378 539 412
rect 585 397 601 431
rect 635 397 651 431
rect 585 381 651 397
rect 685 535 741 551
rect 685 501 691 535
rect 725 501 741 535
rect 685 431 741 501
rect 685 397 691 431
rect 725 397 741 431
rect 886 529 902 563
rect 886 465 936 529
rect 886 431 902 465
rect 886 415 936 431
rect 976 563 1054 579
rect 976 529 992 563
rect 1026 529 1054 563
rect 976 482 1054 529
rect 1196 566 1262 649
rect 1196 532 1212 566
rect 1246 532 1262 566
rect 1196 516 1262 532
rect 1325 580 1391 596
rect 1325 546 1341 580
rect 1375 546 1391 580
rect 1325 497 1391 546
rect 976 480 1291 482
rect 976 446 992 480
rect 1026 448 1291 480
rect 1026 446 1054 448
rect 473 347 539 378
rect 365 331 651 347
rect 365 313 601 331
rect 365 241 415 313
rect 585 297 601 313
rect 635 297 651 331
rect 585 281 651 297
rect 685 281 741 397
rect 976 397 1054 446
rect 976 381 992 397
rect 792 365 992 381
rect 792 331 808 365
rect 842 363 992 365
rect 1026 363 1054 397
rect 1088 380 1104 414
rect 1138 380 1155 414
rect 1088 364 1155 380
rect 842 347 1054 363
rect 842 331 858 347
rect 792 315 858 331
rect 920 297 986 313
rect 920 281 936 297
rect 399 207 415 241
rect 449 263 515 279
rect 449 229 465 263
rect 499 247 515 263
rect 685 263 936 281
rect 970 263 986 297
rect 685 247 986 263
rect 499 229 595 247
rect 449 213 595 229
rect 365 191 415 207
rect 461 157 527 179
rect 123 141 527 157
rect 123 123 488 141
rect 461 107 488 123
rect 522 107 527 141
rect 225 73 313 89
rect 225 39 252 73
rect 286 39 313 73
rect 461 70 527 107
rect 561 88 595 213
rect 685 188 719 247
rect 1020 213 1054 347
rect 629 172 719 188
rect 629 138 649 172
rect 683 138 719 172
rect 629 122 719 138
rect 753 179 955 213
rect 753 88 787 179
rect 561 54 787 88
rect 821 124 887 145
rect 821 90 837 124
rect 871 90 887 124
rect 225 17 313 39
rect 821 17 887 90
rect 921 85 955 179
rect 989 183 1055 213
rect 989 149 1005 183
rect 1039 149 1055 183
rect 989 119 1055 149
rect 1089 202 1123 364
rect 1257 326 1291 448
rect 1325 463 1341 497
rect 1375 463 1391 497
rect 1325 414 1391 463
rect 1425 580 1491 649
rect 1425 546 1441 580
rect 1475 546 1491 580
rect 1425 478 1491 546
rect 1425 444 1441 478
rect 1475 444 1491 478
rect 1425 428 1491 444
rect 1541 580 1607 596
rect 1541 546 1557 580
rect 1591 546 1607 580
rect 1541 497 1607 546
rect 1541 463 1557 497
rect 1591 463 1607 497
rect 1325 380 1341 414
rect 1375 394 1391 414
rect 1541 414 1607 463
rect 1647 580 1697 649
rect 1681 546 1697 580
rect 1647 478 1697 546
rect 1681 444 1697 478
rect 1647 428 1697 444
rect 1731 580 1797 596
rect 1731 546 1747 580
rect 1781 546 1797 580
rect 1731 497 1797 546
rect 1731 463 1747 497
rect 1781 463 1797 497
rect 1375 380 1507 394
rect 1325 360 1507 380
rect 1541 380 1557 414
rect 1591 394 1607 414
rect 1731 414 1797 463
rect 1731 394 1747 414
rect 1591 380 1747 394
rect 1781 380 1797 414
rect 1541 360 1797 380
rect 1831 580 1897 649
rect 1831 546 1847 580
rect 1881 546 1897 580
rect 1831 497 1897 546
rect 1831 463 1847 497
rect 1881 463 1897 497
rect 1831 414 1897 463
rect 1831 380 1847 414
rect 1881 380 1897 414
rect 1831 364 1897 380
rect 1473 326 1507 360
rect 1257 310 1406 326
rect 1157 294 1223 310
rect 1157 260 1173 294
rect 1207 260 1223 294
rect 1257 276 1356 310
rect 1390 276 1406 310
rect 1257 260 1406 276
rect 1473 310 1687 326
rect 1473 276 1501 310
rect 1535 276 1569 310
rect 1603 276 1637 310
rect 1671 276 1687 310
rect 1473 260 1687 276
rect 1745 282 1797 360
rect 1157 236 1223 260
rect 1473 226 1507 260
rect 1745 226 1811 282
rect 1365 210 1507 226
rect 1089 168 1117 202
rect 1151 168 1167 202
rect 1089 120 1167 168
rect 1089 86 1117 120
rect 1151 86 1167 120
rect 1089 85 1167 86
rect 921 51 1167 85
rect 1201 168 1217 202
rect 1251 168 1267 202
rect 1201 120 1267 168
rect 1201 86 1217 120
rect 1251 86 1267 120
rect 1201 17 1267 86
rect 1365 176 1381 210
rect 1415 192 1507 210
rect 1573 210 1811 226
rect 1415 176 1431 192
rect 1365 120 1431 176
rect 1573 176 1589 210
rect 1623 192 1761 210
rect 1365 86 1381 120
rect 1415 86 1431 120
rect 1365 70 1431 86
rect 1477 131 1527 158
rect 1477 97 1493 131
rect 1477 17 1527 97
rect 1573 120 1623 176
rect 1745 176 1761 192
rect 1795 176 1811 210
rect 1573 86 1589 120
rect 1573 70 1623 86
rect 1659 131 1709 158
rect 1659 97 1675 131
rect 1659 17 1709 97
rect 1745 120 1811 176
rect 1745 86 1761 120
rect 1795 86 1811 120
rect 1745 70 1811 86
rect 1847 210 1897 226
rect 1881 176 1897 210
rect 1847 120 1897 176
rect 1881 86 1897 120
rect 1847 17 1897 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
<< metal1 >>
rect 0 683 1920 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 0 617 1920 649
rect 0 17 1920 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
rect 0 -49 1920 -17
<< labels >>
flabel pwell s 0 0 1920 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 1920 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
rlabel comment s 0 0 0 0 4 sdlclkp_4
flabel metal1 s 0 617 1920 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 1920 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 SCE
port 3 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 GATE
port 2 nsew
flabel corelocali s 1183 242 1217 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 1759 242 1793 276 0 FreeSans 340 0 0 0 GCLK
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 1920 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 338952
string GDS_START 326072
<< end >>
