magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 17 299 85 493
rect 17 177 52 299
rect 270 215 363 255
rect 397 215 474 255
rect 508 215 616 255
rect 17 51 85 177
rect 563 87 616 215
rect 728 215 801 265
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 129 299 163 527
rect 217 367 267 527
rect 417 333 493 493
rect 552 367 618 527
rect 694 333 760 493
rect 201 299 760 333
rect 201 249 235 299
rect 86 215 235 249
rect 129 17 179 177
rect 217 147 482 181
rect 217 51 283 147
rect 327 17 372 109
rect 406 51 482 147
rect 650 173 694 299
rect 650 51 760 173
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
rlabel locali s 270 215 363 255 6 A1
port 1 nsew signal input
rlabel locali s 397 215 474 255 6 A2
port 2 nsew signal input
rlabel locali s 563 87 616 215 6 B1
port 3 nsew signal input
rlabel locali s 508 215 616 255 6 B1
port 3 nsew signal input
rlabel locali s 728 215 801 265 6 C1
port 4 nsew signal input
rlabel locali s 17 299 85 493 6 X
port 5 nsew signal output
rlabel locali s 17 177 52 299 6 X
port 5 nsew signal output
rlabel locali s 17 51 85 177 6 X
port 5 nsew signal output
rlabel metal1 s 0 -48 828 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 828 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2568290
string GDS_START 2561202
<< end >>
