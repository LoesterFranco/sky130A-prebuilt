magic
tech sky130A
magscale 1 2
timestamp 1604502697
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 89 47 119 177
rect 183 47 213 177
rect 277 47 307 177
rect 371 47 401 177
rect 465 47 495 177
<< pmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 457 297 493 497
<< ndiff >>
rect 27 129 89 177
rect 27 95 35 129
rect 69 95 89 129
rect 27 47 89 95
rect 119 97 183 177
rect 119 63 129 97
rect 163 63 183 97
rect 119 47 183 63
rect 213 129 277 177
rect 213 95 223 129
rect 257 95 277 129
rect 213 47 277 95
rect 307 97 371 177
rect 307 63 317 97
rect 351 63 371 97
rect 307 47 371 63
rect 401 129 465 177
rect 401 95 411 129
rect 445 95 465 129
rect 401 47 465 95
rect 495 161 547 177
rect 495 127 505 161
rect 539 127 547 161
rect 495 93 547 127
rect 495 59 505 93
rect 539 59 547 93
rect 495 47 547 59
<< pdiff >>
rect 27 479 81 497
rect 27 445 35 479
rect 69 445 81 479
rect 27 411 81 445
rect 27 377 35 411
rect 69 377 81 411
rect 27 343 81 377
rect 27 309 35 343
rect 69 309 81 343
rect 27 297 81 309
rect 117 485 175 497
rect 117 451 129 485
rect 163 451 175 485
rect 117 417 175 451
rect 117 383 129 417
rect 163 383 175 417
rect 117 297 175 383
rect 211 463 269 497
rect 211 429 223 463
rect 257 429 269 463
rect 211 368 269 429
rect 211 334 223 368
rect 257 334 269 368
rect 211 297 269 334
rect 305 485 363 497
rect 305 451 317 485
rect 351 451 363 485
rect 305 417 363 451
rect 305 383 317 417
rect 351 383 363 417
rect 305 297 363 383
rect 399 463 457 497
rect 399 429 411 463
rect 445 429 457 463
rect 399 368 457 429
rect 399 334 411 368
rect 445 334 457 368
rect 399 297 457 334
rect 493 485 547 497
rect 493 451 505 485
rect 539 451 547 485
rect 493 417 547 451
rect 493 383 505 417
rect 539 383 547 417
rect 493 349 547 383
rect 493 315 505 349
rect 539 315 547 349
rect 493 297 547 315
<< ndiffc >>
rect 35 95 69 129
rect 129 63 163 97
rect 223 95 257 129
rect 317 63 351 97
rect 411 95 445 129
rect 505 127 539 161
rect 505 59 539 93
<< pdiffc >>
rect 35 445 69 479
rect 35 377 69 411
rect 35 309 69 343
rect 129 451 163 485
rect 129 383 163 417
rect 223 429 257 463
rect 223 334 257 368
rect 317 451 351 485
rect 317 383 351 417
rect 411 429 445 463
rect 411 334 445 368
rect 505 451 539 485
rect 505 383 539 417
rect 505 315 539 349
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 457 497 493 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 457 282 493 297
rect 79 261 119 282
rect 28 249 119 261
rect 173 259 213 282
rect 267 259 307 282
rect 361 259 401 282
rect 455 259 495 282
rect 28 215 44 249
rect 78 215 119 249
rect 28 203 119 215
rect 172 249 495 259
rect 172 215 188 249
rect 222 215 495 249
rect 172 205 495 215
rect 89 177 119 203
rect 183 177 213 205
rect 277 177 307 205
rect 371 177 401 205
rect 465 177 495 205
rect 89 21 119 47
rect 183 21 213 47
rect 277 21 307 47
rect 371 21 401 47
rect 465 21 495 47
<< polycont >>
rect 44 215 78 249
rect 188 215 222 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 19 479 85 493
rect 19 445 35 479
rect 69 445 85 479
rect 19 411 85 445
rect 19 377 35 411
rect 69 377 85 411
rect 19 343 85 377
rect 129 485 177 527
rect 163 451 177 485
rect 129 417 177 451
rect 163 383 177 417
rect 129 367 177 383
rect 223 463 257 493
rect 223 368 257 429
rect 19 309 35 343
rect 69 331 85 343
rect 291 485 367 527
rect 291 451 317 485
rect 351 451 367 485
rect 291 417 367 451
rect 291 383 317 417
rect 351 383 367 417
rect 291 367 367 383
rect 411 463 445 493
rect 411 368 445 429
rect 69 309 172 331
rect 19 297 172 309
rect 18 249 94 263
rect 18 215 44 249
rect 78 215 94 249
rect 138 249 172 297
rect 223 323 257 334
rect 411 323 445 334
rect 223 289 445 323
rect 479 485 555 527
rect 479 451 505 485
rect 539 451 555 485
rect 479 417 555 451
rect 479 383 505 417
rect 539 383 555 417
rect 479 349 555 383
rect 479 315 505 349
rect 539 315 555 349
rect 479 297 555 315
rect 138 215 188 249
rect 222 215 248 249
rect 138 181 172 215
rect 384 181 445 289
rect 35 147 172 181
rect 223 147 445 181
rect 35 129 69 147
rect 223 129 257 147
rect 35 51 69 95
rect 105 97 163 113
rect 105 63 129 97
rect 105 17 163 63
rect 411 129 445 147
rect 223 51 257 95
rect 291 97 367 113
rect 291 63 317 97
rect 351 63 367 97
rect 291 17 367 63
rect 411 51 445 95
rect 479 161 555 177
rect 479 127 505 161
rect 539 127 555 161
rect 479 93 555 127
rect 479 59 505 93
rect 539 59 555 93
rect 479 17 555 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel corelocali s 395 221 429 255 0 FreeSans 200 0 0 0 X
port 6 nsew
flabel corelocali s 395 289 429 323 0 FreeSans 200 0 0 0 X
port 6 nsew
flabel corelocali s 395 153 429 187 0 FreeSans 200 0 0 0 X
port 6 nsew
flabel corelocali s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew
flabel corelocali s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew
rlabel comment s 0 0 0 0 4 buf_4
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1666920
string GDS_START 1661252
<< end >>
