magic
tech sky130A
magscale 1 2
timestamp 1604502729
<< locali >>
rect 125 390 310 596
rect 23 236 89 310
rect 125 226 159 390
rect 193 270 263 356
rect 307 270 373 356
rect 409 260 555 356
rect 123 131 213 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 25 364 91 649
rect 451 390 517 649
rect 23 97 89 202
rect 268 192 534 226
rect 268 97 334 192
rect 23 63 334 97
rect 368 17 434 158
rect 468 70 534 192
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
rlabel locali s 409 260 555 356 6 A1
port 1 nsew signal input
rlabel locali s 307 270 373 356 6 A2
port 2 nsew signal input
rlabel locali s 23 236 89 310 6 B1
port 3 nsew signal input
rlabel locali s 193 270 263 356 6 B2
port 4 nsew signal input
rlabel locali s 125 390 310 596 6 Y
port 5 nsew signal output
rlabel locali s 125 226 159 390 6 Y
port 5 nsew signal output
rlabel locali s 123 131 213 226 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -49 576 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 576 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 576 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1297950
string GDS_START 1292270
<< end >>
