magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1196 561
rect 127 443 193 527
rect 295 443 361 527
rect 463 443 529 527
rect 121 257 177 341
rect 85 215 177 257
rect 211 289 445 341
rect 640 427 690 527
rect 211 181 291 289
rect 143 17 177 181
rect 211 145 445 181
rect 987 367 1053 527
rect 756 215 964 255
rect 998 215 1179 255
rect 211 51 277 145
rect 311 17 345 111
rect 379 51 445 145
rect 479 17 513 111
rect 835 17 869 111
rect 1003 17 1037 111
rect 0 -17 1196 17
<< obsli1 >>
rect 17 409 87 493
rect 17 375 513 409
rect 17 291 87 375
rect 17 171 51 291
rect 479 323 513 375
rect 563 393 597 493
rect 737 459 953 493
rect 737 427 785 459
rect 827 393 876 425
rect 563 359 876 393
rect 479 289 581 323
rect 325 215 513 255
rect 547 249 581 289
rect 547 215 627 249
rect 17 53 109 171
rect 479 179 513 215
rect 679 179 717 359
rect 827 289 876 359
rect 919 333 953 459
rect 1087 333 1142 493
rect 919 291 1142 333
rect 479 145 717 179
rect 647 129 717 145
rect 751 145 1142 181
rect 751 95 801 145
rect 561 51 801 95
rect 903 51 969 145
rect 1071 53 1142 145
<< metal1 >>
rect 0 496 1196 592
rect 0 -48 1196 48
<< labels >>
rlabel locali s 998 215 1179 255 6 A1
port 1 nsew signal input
rlabel locali s 756 215 964 255 6 A2
port 2 nsew signal input
rlabel locali s 121 257 177 341 6 B1_N
port 3 nsew signal input
rlabel locali s 85 215 177 257 6 B1_N
port 3 nsew signal input
rlabel locali s 379 51 445 145 6 X
port 4 nsew signal output
rlabel locali s 211 289 445 341 6 X
port 4 nsew signal output
rlabel locali s 211 181 291 289 6 X
port 4 nsew signal output
rlabel locali s 211 145 445 181 6 X
port 4 nsew signal output
rlabel locali s 211 51 277 145 6 X
port 4 nsew signal output
rlabel locali s 1003 17 1037 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 835 17 869 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 479 17 513 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 311 17 345 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 143 17 177 181 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 1196 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1196 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 987 367 1053 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 640 427 690 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 463 443 529 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 295 443 361 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 127 443 193 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 1196 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 1196 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1388840
string GDS_START 1379840
<< end >>
