magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 301 444 633 465
rect 133 431 633 444
rect 133 410 335 431
rect 133 356 167 410
rect 488 376 554 397
rect 85 270 167 356
rect 217 342 554 376
rect 599 353 633 431
rect 217 274 551 342
rect 599 287 749 353
rect 1328 290 1415 356
rect 1465 290 1635 356
rect 262 74 328 274
rect 466 74 551 274
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 17 512 89 572
rect 130 546 199 649
rect 364 567 430 649
rect 612 567 678 649
rect 233 512 701 533
rect 17 499 701 512
rect 17 478 267 499
rect 17 390 89 478
rect 17 230 51 390
rect 667 421 701 499
rect 735 521 785 595
rect 826 555 892 649
rect 1040 555 1090 649
rect 1124 542 1423 596
rect 1124 521 1158 542
rect 735 487 1158 521
rect 1539 508 1605 596
rect 735 455 785 487
rect 1192 474 1605 508
rect 1192 453 1226 474
rect 667 387 817 421
rect 933 419 1226 453
rect 1639 440 1705 596
rect 933 387 1028 419
rect 1260 390 1705 440
rect 783 353 817 387
rect 1260 356 1294 390
rect 783 287 997 353
rect 1077 290 1294 356
rect 17 94 120 230
rect 154 17 220 230
rect 362 17 428 214
rect 1031 253 1604 256
rect 585 17 651 251
rect 704 222 1604 253
rect 704 219 1065 222
rect 704 115 770 219
rect 1099 185 1418 188
rect 804 17 898 181
rect 932 154 1418 185
rect 932 151 1133 154
rect 932 115 998 151
rect 1034 17 1115 117
rect 1167 85 1318 120
rect 1352 119 1418 154
rect 1452 85 1518 188
rect 1554 119 1604 222
rect 1671 206 1705 390
rect 1638 85 1705 206
rect 1167 51 1705 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
<< metal1 >>
rect 0 683 1728 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 0 617 1728 649
rect 0 17 1728 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
rect 0 -49 1728 -17
<< labels >>
rlabel locali s 1328 290 1415 356 6 A0
port 1 nsew signal input
rlabel locali s 1465 290 1635 356 6 A1
port 2 nsew signal input
rlabel locali s 599 353 633 431 6 S
port 3 nsew signal input
rlabel locali s 599 287 749 353 6 S
port 3 nsew signal input
rlabel locali s 301 444 633 465 6 S
port 3 nsew signal input
rlabel locali s 133 431 633 444 6 S
port 3 nsew signal input
rlabel locali s 133 410 335 431 6 S
port 3 nsew signal input
rlabel locali s 133 356 167 410 6 S
port 3 nsew signal input
rlabel locali s 85 270 167 356 6 S
port 3 nsew signal input
rlabel locali s 488 376 554 397 6 X
port 4 nsew signal output
rlabel locali s 466 74 551 274 6 X
port 4 nsew signal output
rlabel locali s 262 74 328 274 6 X
port 4 nsew signal output
rlabel locali s 217 342 554 376 6 X
port 4 nsew signal output
rlabel locali s 217 274 551 342 6 X
port 4 nsew signal output
rlabel metal1 s 0 -49 1728 49 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1728 715 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1728 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1598978
string GDS_START 1586614
<< end >>
