magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 155 47 185 177
rect 284 47 314 177
rect 356 47 386 177
rect 481 47 511 177
rect 577 47 607 177
rect 673 47 703 177
rect 779 47 809 177
<< pmoshvt >>
rect 147 297 183 497
rect 276 297 312 497
rect 372 297 408 497
rect 483 297 519 497
rect 579 297 615 497
rect 675 297 711 497
rect 771 297 807 497
<< ndiff >>
rect 94 161 155 177
rect 94 127 110 161
rect 144 127 155 161
rect 94 93 155 127
rect 94 59 110 93
rect 144 59 155 93
rect 94 47 155 59
rect 185 47 284 177
rect 314 47 356 177
rect 386 89 481 177
rect 386 55 427 89
rect 461 55 481 89
rect 386 47 481 55
rect 511 153 577 177
rect 511 119 532 153
rect 566 119 577 153
rect 511 47 577 119
rect 607 89 673 177
rect 607 55 628 89
rect 662 55 673 89
rect 607 47 673 55
rect 703 169 779 177
rect 703 135 724 169
rect 758 135 779 169
rect 703 101 779 135
rect 703 67 724 101
rect 758 67 779 101
rect 703 47 779 67
rect 809 89 866 177
rect 809 55 820 89
rect 854 55 866 89
rect 809 47 866 55
<< pdiff >>
rect 85 477 147 497
rect 85 443 101 477
rect 135 443 147 477
rect 85 409 147 443
rect 85 375 101 409
rect 135 375 147 409
rect 85 297 147 375
rect 183 489 276 497
rect 183 455 219 489
rect 253 455 276 489
rect 183 421 276 455
rect 183 387 219 421
rect 253 387 276 421
rect 183 297 276 387
rect 312 477 372 497
rect 312 443 325 477
rect 359 443 372 477
rect 312 409 372 443
rect 312 375 325 409
rect 359 375 372 409
rect 312 297 372 375
rect 408 489 483 497
rect 408 455 428 489
rect 462 455 483 489
rect 408 421 483 455
rect 408 387 428 421
rect 462 387 483 421
rect 408 297 483 387
rect 519 477 579 497
rect 519 443 532 477
rect 566 443 579 477
rect 519 409 579 443
rect 519 375 532 409
rect 566 375 579 409
rect 519 297 579 375
rect 615 489 675 497
rect 615 455 628 489
rect 662 455 675 489
rect 615 421 675 455
rect 615 387 628 421
rect 662 387 675 421
rect 615 297 675 387
rect 711 477 771 497
rect 711 443 724 477
rect 758 443 771 477
rect 711 409 771 443
rect 711 375 724 409
rect 758 375 771 409
rect 711 341 771 375
rect 711 307 724 341
rect 758 307 771 341
rect 711 297 771 307
rect 807 489 866 497
rect 807 455 820 489
rect 854 455 866 489
rect 807 421 866 455
rect 807 387 820 421
rect 854 387 866 421
rect 807 297 866 387
<< ndiffc >>
rect 110 127 144 161
rect 110 59 144 93
rect 427 55 461 89
rect 532 119 566 153
rect 628 55 662 89
rect 724 135 758 169
rect 724 67 758 101
rect 820 55 854 89
<< pdiffc >>
rect 101 443 135 477
rect 101 375 135 409
rect 219 455 253 489
rect 219 387 253 421
rect 325 443 359 477
rect 325 375 359 409
rect 428 455 462 489
rect 428 387 462 421
rect 532 443 566 477
rect 532 375 566 409
rect 628 455 662 489
rect 628 387 662 421
rect 724 443 758 477
rect 724 375 758 409
rect 724 307 758 341
rect 820 455 854 489
rect 820 387 854 421
<< poly >>
rect 147 497 183 523
rect 276 497 312 523
rect 372 497 408 523
rect 483 497 519 523
rect 579 497 615 523
rect 675 497 711 523
rect 771 497 807 523
rect 147 282 183 297
rect 276 282 312 297
rect 372 282 408 297
rect 483 282 519 297
rect 579 282 615 297
rect 675 282 711 297
rect 771 282 807 297
rect 145 265 185 282
rect 274 265 314 282
rect 370 265 410 282
rect 481 265 521 282
rect 577 265 617 282
rect 673 265 713 282
rect 769 265 809 282
rect 121 249 185 265
rect 121 215 131 249
rect 165 215 185 249
rect 121 199 185 215
rect 227 249 314 265
rect 227 215 237 249
rect 271 215 314 249
rect 227 199 314 215
rect 155 177 185 199
rect 284 177 314 199
rect 356 249 420 265
rect 356 215 366 249
rect 400 215 420 249
rect 356 199 420 215
rect 481 249 809 265
rect 481 215 497 249
rect 531 215 575 249
rect 609 215 653 249
rect 687 215 731 249
rect 765 215 809 249
rect 481 199 809 215
rect 356 177 386 199
rect 481 177 511 199
rect 577 177 607 199
rect 673 177 703 199
rect 779 177 809 199
rect 155 21 185 47
rect 284 21 314 47
rect 356 21 386 47
rect 481 21 511 47
rect 577 21 607 47
rect 673 21 703 47
rect 779 21 809 47
<< polycont >>
rect 131 215 165 249
rect 237 215 271 249
rect 366 215 400 249
rect 497 215 531 249
rect 575 215 609 249
rect 653 215 687 249
rect 731 215 765 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 100 477 136 493
rect 23 268 66 467
rect 100 443 101 477
rect 135 443 136 477
rect 100 409 136 443
rect 100 375 101 409
rect 135 375 136 409
rect 179 489 279 527
rect 179 455 219 489
rect 253 455 279 489
rect 179 421 279 455
rect 179 387 219 421
rect 253 387 279 421
rect 324 477 360 493
rect 324 443 325 477
rect 359 443 360 477
rect 324 409 360 443
rect 100 350 136 375
rect 324 375 325 409
rect 359 375 360 409
rect 412 489 478 527
rect 412 455 428 489
rect 462 455 478 489
rect 412 421 478 455
rect 412 387 428 421
rect 462 387 478 421
rect 530 477 568 493
rect 530 443 532 477
rect 566 443 568 477
rect 530 409 568 443
rect 324 350 360 375
rect 530 375 532 409
rect 566 375 568 409
rect 602 489 678 527
rect 602 455 628 489
rect 662 455 678 489
rect 602 421 678 455
rect 602 387 628 421
rect 662 387 678 421
rect 722 477 760 493
rect 722 443 724 477
rect 758 443 760 477
rect 722 409 760 443
rect 530 352 568 375
rect 722 375 724 409
rect 758 375 760 409
rect 794 489 870 527
rect 794 455 820 489
rect 854 455 870 489
rect 794 421 870 455
rect 794 387 820 421
rect 854 387 870 421
rect 722 353 760 375
rect 722 352 898 353
rect 100 316 486 350
rect 444 271 486 316
rect 530 341 898 352
rect 530 307 724 341
rect 758 307 898 341
rect 23 249 175 268
rect 23 215 131 249
rect 165 215 175 249
rect 23 199 175 215
rect 209 249 271 268
rect 209 215 237 249
rect 93 127 110 161
rect 144 127 160 161
rect 209 149 271 215
rect 305 249 410 265
rect 305 215 366 249
rect 400 215 410 249
rect 305 199 410 215
rect 444 249 781 271
rect 444 215 497 249
rect 531 215 575 249
rect 609 215 653 249
rect 687 215 731 249
rect 765 215 781 249
rect 444 204 781 215
rect 444 161 486 204
rect 842 169 898 307
rect 93 93 160 127
rect 93 59 110 93
rect 144 89 160 93
rect 327 123 486 161
rect 530 153 724 169
rect 327 89 365 123
rect 530 119 532 153
rect 566 135 724 153
rect 758 135 898 169
rect 566 123 898 135
rect 566 119 568 123
rect 530 103 568 119
rect 722 101 760 123
rect 144 59 365 89
rect 93 51 365 59
rect 411 55 427 89
rect 461 55 477 89
rect 411 17 477 55
rect 602 55 628 89
rect 662 55 678 89
rect 602 17 678 55
rect 722 67 724 101
rect 758 67 760 101
rect 722 51 760 67
rect 794 55 820 89
rect 854 55 870 89
rect 794 17 870 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel corelocali s 111 221 145 255 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 223 221 257 255 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 322 238 322 238 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 852 153 886 187 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
rlabel comment s 0 0 0 0 4 and3_4
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1531194
string GDS_START 1523990
<< end >>
