magic
tech sky130A
magscale 1 2
timestamp 1599588238
<< locali >>
rect 25 294 243 360
rect 285 294 359 360
rect 393 270 459 356
rect 25 101 71 134
rect 25 51 112 101
rect 585 70 651 596
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 39 394 89 649
rect 129 581 399 615
rect 129 394 179 581
rect 219 428 285 547
rect 319 462 399 581
rect 433 462 545 649
rect 219 394 551 428
rect 44 226 257 260
rect 501 236 551 394
rect 44 168 110 226
rect 146 17 189 192
rect 223 125 257 226
rect 297 202 551 236
rect 297 159 363 202
rect 223 75 449 125
rect 499 17 549 168
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel locali s 393 270 459 356 6 A1
port 1 nsew signal input
rlabel locali s 25 101 71 134 6 A2
port 2 nsew signal input
rlabel locali s 25 51 112 101 6 A2
port 2 nsew signal input
rlabel locali s 285 294 359 360 6 B1
port 3 nsew signal input
rlabel locali s 25 294 243 360 6 B2
port 4 nsew signal input
rlabel locali s 585 70 651 596 6 X
port 5 nsew signal output
rlabel metal1 s 0 -49 672 49 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 617 672 715 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3463794
string GDS_START 3456366
<< end >>
