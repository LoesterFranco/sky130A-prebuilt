magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 1050 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 94 47 124 177
rect 190 47 220 177
rect 286 47 316 177
rect 382 47 412 177
rect 590 47 620 177
rect 691 47 721 177
rect 782 47 812 177
rect 879 47 909 177
<< pmoshvt >>
rect 86 297 122 497
rect 182 297 218 497
rect 278 297 314 497
rect 374 297 410 497
rect 582 297 618 497
rect 678 297 714 497
rect 774 297 810 497
rect 870 297 906 497
<< ndiff >>
rect 27 89 94 177
rect 27 55 39 89
rect 73 55 94 89
rect 27 47 94 55
rect 124 169 190 177
rect 124 135 135 169
rect 169 135 190 169
rect 124 47 190 135
rect 220 158 286 177
rect 220 124 231 158
rect 265 124 286 158
rect 220 89 286 124
rect 220 55 231 89
rect 265 55 286 89
rect 220 47 286 55
rect 316 165 382 177
rect 316 131 327 165
rect 361 131 382 165
rect 316 47 382 131
rect 412 89 469 177
rect 412 55 423 89
rect 457 55 469 89
rect 412 47 469 55
rect 523 89 590 177
rect 523 55 535 89
rect 569 55 590 89
rect 523 47 590 55
rect 620 165 691 177
rect 620 131 631 165
rect 665 131 691 165
rect 620 47 691 131
rect 721 89 782 177
rect 721 55 731 89
rect 765 55 782 89
rect 721 47 782 55
rect 812 153 879 177
rect 812 119 823 153
rect 857 119 879 153
rect 812 47 879 119
rect 909 89 970 177
rect 909 55 924 89
rect 958 55 970 89
rect 909 47 970 55
<< pdiff >>
rect 31 485 86 497
rect 31 451 39 485
rect 73 451 86 485
rect 31 297 86 451
rect 122 477 182 497
rect 122 443 135 477
rect 169 443 182 477
rect 122 381 182 443
rect 122 347 135 381
rect 169 347 182 381
rect 122 297 182 347
rect 218 485 278 497
rect 218 451 231 485
rect 265 451 278 485
rect 218 417 278 451
rect 218 383 231 417
rect 265 383 278 417
rect 218 297 278 383
rect 314 477 374 497
rect 314 443 327 477
rect 361 443 374 477
rect 314 386 374 443
rect 314 352 327 386
rect 361 352 374 386
rect 314 297 374 352
rect 410 485 465 497
rect 410 451 423 485
rect 457 451 465 485
rect 410 417 465 451
rect 410 383 423 417
rect 457 383 465 417
rect 410 297 465 383
rect 527 477 582 497
rect 527 443 535 477
rect 569 443 582 477
rect 527 297 582 443
rect 618 425 678 497
rect 618 391 631 425
rect 665 391 678 425
rect 618 357 678 391
rect 618 323 631 357
rect 665 323 678 357
rect 618 297 678 323
rect 714 477 774 497
rect 714 443 727 477
rect 761 443 774 477
rect 714 382 774 443
rect 714 348 727 382
rect 761 348 774 382
rect 714 297 774 348
rect 810 485 870 497
rect 810 451 823 485
rect 857 451 870 485
rect 810 407 870 451
rect 810 373 823 407
rect 857 373 870 407
rect 810 297 870 373
rect 906 477 961 497
rect 906 443 919 477
rect 953 443 961 477
rect 906 409 961 443
rect 906 375 919 409
rect 953 375 961 409
rect 906 297 961 375
<< ndiffc >>
rect 39 55 73 89
rect 135 135 169 169
rect 231 124 265 158
rect 231 55 265 89
rect 327 131 361 165
rect 423 55 457 89
rect 535 55 569 89
rect 631 131 665 165
rect 731 55 765 89
rect 823 119 857 153
rect 924 55 958 89
<< pdiffc >>
rect 39 451 73 485
rect 135 443 169 477
rect 135 347 169 381
rect 231 451 265 485
rect 231 383 265 417
rect 327 443 361 477
rect 327 352 361 386
rect 423 451 457 485
rect 423 383 457 417
rect 535 443 569 477
rect 631 391 665 425
rect 631 323 665 357
rect 727 443 761 477
rect 727 348 761 382
rect 823 451 857 485
rect 823 373 857 407
rect 919 443 953 477
rect 919 375 953 409
<< poly >>
rect 86 497 122 523
rect 182 497 218 523
rect 278 497 314 523
rect 374 497 410 523
rect 582 497 618 523
rect 678 497 714 523
rect 774 497 810 523
rect 870 497 906 523
rect 86 282 122 297
rect 182 282 218 297
rect 278 282 314 297
rect 374 282 410 297
rect 582 282 618 297
rect 678 282 714 297
rect 774 282 810 297
rect 870 282 906 297
rect 84 265 124 282
rect 180 265 220 282
rect 276 265 316 282
rect 372 265 412 282
rect 580 265 620 282
rect 676 265 716 282
rect 772 265 812 282
rect 868 265 908 282
rect 21 249 220 265
rect 21 215 31 249
rect 65 215 220 249
rect 21 199 220 215
rect 262 249 412 265
rect 262 215 272 249
rect 306 215 350 249
rect 384 215 412 249
rect 262 199 412 215
rect 579 249 721 265
rect 579 215 589 249
rect 623 215 667 249
rect 701 215 721 249
rect 579 199 721 215
rect 767 249 909 265
rect 767 215 777 249
rect 811 215 855 249
rect 889 215 909 249
rect 767 199 909 215
rect 94 177 124 199
rect 190 177 220 199
rect 286 177 316 199
rect 382 177 412 199
rect 590 177 620 199
rect 691 177 721 199
rect 782 177 812 199
rect 879 177 909 199
rect 94 21 124 47
rect 190 21 220 47
rect 286 21 316 47
rect 382 21 412 47
rect 590 21 620 47
rect 691 21 721 47
rect 782 21 812 47
rect 879 21 909 47
<< polycont >>
rect 31 215 65 249
rect 272 215 306 249
rect 350 215 384 249
rect 589 215 623 249
rect 667 215 701 249
rect 777 215 811 249
rect 855 215 889 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 23 485 75 527
rect 23 451 39 485
rect 73 451 75 485
rect 23 435 75 451
rect 109 477 171 493
rect 109 443 135 477
rect 169 443 171 477
rect 17 249 75 394
rect 17 215 31 249
rect 65 215 75 249
rect 17 199 75 215
rect 109 381 171 443
rect 205 485 281 527
rect 205 451 231 485
rect 265 451 281 485
rect 205 417 281 451
rect 205 383 231 417
rect 265 383 281 417
rect 325 477 363 493
rect 325 443 327 477
rect 361 443 363 477
rect 325 386 363 443
rect 109 347 135 381
rect 169 347 171 381
rect 109 342 171 347
rect 325 352 327 386
rect 361 352 363 386
rect 397 485 473 527
rect 397 451 423 485
rect 457 451 473 485
rect 397 417 473 451
rect 519 477 763 493
rect 519 443 535 477
rect 569 459 727 477
rect 569 443 571 459
rect 519 420 571 443
rect 725 443 727 459
rect 761 443 763 477
rect 397 383 423 417
rect 457 383 473 417
rect 605 391 631 425
rect 665 391 681 425
rect 325 342 363 352
rect 605 357 681 391
rect 605 342 631 357
rect 109 323 631 342
rect 665 323 681 357
rect 109 308 681 323
rect 725 382 763 443
rect 725 348 727 382
rect 761 348 763 382
rect 797 485 873 527
rect 797 451 823 485
rect 857 451 873 485
rect 797 407 873 451
rect 797 373 823 407
rect 857 373 873 407
rect 917 477 969 493
rect 917 443 919 477
rect 953 443 969 477
rect 917 409 969 443
rect 917 375 919 409
rect 953 375 969 409
rect 725 339 763 348
rect 917 339 969 375
rect 109 169 185 308
rect 725 305 969 339
rect 243 249 442 273
rect 243 215 272 249
rect 306 215 350 249
rect 384 215 442 249
rect 534 249 727 271
rect 534 215 589 249
rect 623 215 667 249
rect 701 215 727 249
rect 761 249 983 259
rect 761 215 777 249
rect 811 215 855 249
rect 889 215 983 249
rect 109 135 135 169
rect 169 135 185 169
rect 109 134 185 135
rect 229 158 267 178
rect 229 124 231 158
rect 265 124 267 158
rect 301 165 859 169
rect 301 131 327 165
rect 361 131 631 165
rect 665 153 859 165
rect 893 153 983 215
rect 665 131 823 153
rect 301 127 823 131
rect 229 93 267 124
rect 821 119 823 127
rect 857 119 859 153
rect 821 103 859 119
rect 229 89 473 93
rect 19 55 39 89
rect 73 55 231 89
rect 265 55 423 89
rect 457 55 473 89
rect 19 51 473 55
rect 519 55 535 89
rect 569 55 585 89
rect 519 17 585 55
rect 705 55 731 89
rect 765 55 781 89
rect 705 17 781 55
rect 893 55 924 89
rect 958 55 974 89
rect 893 17 974 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
flabel corelocali s 937 153 971 187 0 FreeSans 400 0 0 0 A1
port 1 nsew
flabel corelocali s 581 221 615 255 0 FreeSans 400 0 0 0 A2
port 2 nsew
flabel corelocali s 302 221 336 255 0 FreeSans 400 0 0 0 B1
port 3 nsew
flabel corelocali s 131 153 165 187 0 FreeSans 400 0 0 0 Y
port 9 nsew
flabel corelocali s 29 289 63 323 0 FreeSans 400 0 0 0 C1
port 4 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
rlabel comment s 0 0 0 0 4 o211ai_2
<< properties >>
string FIXED_BBOX 0 0 1012 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 987786
string GDS_START 980022
<< end >>
