magic
tech sky130A
magscale 1 2
timestamp 1599588232
<< locali >>
rect 148 424 214 596
rect 348 424 414 596
rect 937 424 1003 547
rect 1137 424 1203 547
rect 148 390 1319 424
rect 348 364 414 390
rect 937 364 1003 390
rect 25 260 248 356
rect 449 286 839 356
rect 1037 328 1239 356
rect 897 286 1239 328
rect 1273 252 1319 390
rect 1353 270 1555 356
rect 282 220 1319 252
rect 1833 270 2087 356
rect 109 218 1319 220
rect 109 154 348 218
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 23 390 89 649
rect 248 458 314 649
rect 448 458 781 649
rect 837 581 1713 615
rect 837 458 903 581
rect 1037 458 1103 581
rect 1257 458 1323 581
rect 1357 424 1423 547
rect 1457 458 1523 581
rect 1557 430 1613 547
rect 1647 466 1713 581
rect 1759 466 1825 649
rect 1859 430 1905 596
rect 1939 466 2005 649
rect 2039 430 2095 596
rect 1557 424 2095 430
rect 1357 390 2095 424
rect 2135 364 2185 649
rect 23 120 73 226
rect 1589 260 1795 294
rect 1589 236 1623 260
rect 1378 202 1623 236
rect 1745 226 1795 260
rect 1378 184 1428 202
rect 384 150 780 184
rect 814 150 1428 184
rect 384 120 418 150
rect 23 70 418 120
rect 814 116 848 150
rect 454 66 848 116
rect 882 17 948 116
rect 984 70 1034 150
rect 1070 17 1136 116
rect 1172 70 1238 150
rect 1274 17 1342 116
rect 1378 70 1428 150
rect 1464 17 1530 165
rect 1589 70 1623 202
rect 1659 17 1709 226
rect 1745 192 2083 226
rect 1745 70 1795 192
rect 1831 17 1999 158
rect 2033 70 2083 192
rect 2119 17 2185 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
<< metal1 >>
rect 0 683 2208 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 0 617 2208 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 2208 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
rect 0 -49 2208 -17
<< labels >>
rlabel locali s 1833 270 2087 356 6 A1
port 1 nsew signal input
rlabel locali s 1353 270 1555 356 6 A2
port 2 nsew signal input
rlabel locali s 1037 328 1239 356 6 A3
port 3 nsew signal input
rlabel locali s 897 286 1239 328 6 A3
port 3 nsew signal input
rlabel locali s 449 286 839 356 6 B1
port 4 nsew signal input
rlabel locali s 25 260 248 356 6 C1
port 5 nsew signal input
rlabel locali s 1273 252 1319 390 6 Y
port 6 nsew signal output
rlabel locali s 1137 424 1203 547 6 Y
port 6 nsew signal output
rlabel locali s 937 424 1003 547 6 Y
port 6 nsew signal output
rlabel locali s 937 364 1003 390 6 Y
port 6 nsew signal output
rlabel locali s 348 424 414 596 6 Y
port 6 nsew signal output
rlabel locali s 348 364 414 390 6 Y
port 6 nsew signal output
rlabel locali s 282 220 1319 252 6 Y
port 6 nsew signal output
rlabel locali s 148 424 214 596 6 Y
port 6 nsew signal output
rlabel locali s 148 390 1319 424 6 Y
port 6 nsew signal output
rlabel locali s 109 218 1319 220 6 Y
port 6 nsew signal output
rlabel locali s 109 154 348 218 6 Y
port 6 nsew signal output
rlabel metal1 s 0 -49 2208 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 8 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 9 nsew power bidirectional
rlabel metal1 s 0 617 2208 715 6 VPWR
port 10 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2208 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1423308
string GDS_START 1406396
<< end >>
