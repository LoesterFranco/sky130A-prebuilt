magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 18 215 84 323
rect 121 181 181 425
rect 346 289 713 323
rect 346 215 438 289
rect 472 215 603 255
rect 637 215 713 289
rect 747 289 1054 323
rect 747 215 813 289
rect 1020 255 1054 289
rect 847 215 983 255
rect 1020 215 1177 255
rect 121 173 959 181
rect 105 145 959 173
rect 105 61 181 145
rect 487 129 567 145
rect 883 129 959 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 18 459 275 493
rect 18 359 87 459
rect 225 391 275 459
rect 321 459 755 493
rect 321 425 371 459
rect 509 425 559 459
rect 415 391 465 425
rect 603 391 653 425
rect 225 357 653 391
rect 705 391 755 459
rect 807 425 857 527
rect 901 391 951 493
rect 995 425 1045 527
rect 1098 391 1139 493
rect 705 357 1139 391
rect 225 299 275 357
rect 1098 291 1139 357
rect 21 17 71 179
rect 225 17 363 111
rect 397 51 661 95
rect 714 17 748 111
rect 1003 95 1053 181
rect 789 51 1053 95
rect 1097 17 1131 181
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
rlabel locali s 847 215 983 255 6 A1
port 1 nsew signal input
rlabel locali s 1020 255 1054 289 6 A2
port 2 nsew signal input
rlabel locali s 1020 215 1177 255 6 A2
port 2 nsew signal input
rlabel locali s 747 289 1054 323 6 A2
port 2 nsew signal input
rlabel locali s 747 215 813 289 6 A2
port 2 nsew signal input
rlabel locali s 472 215 603 255 6 B1
port 3 nsew signal input
rlabel locali s 637 215 713 289 6 B2
port 4 nsew signal input
rlabel locali s 346 289 713 323 6 B2
port 4 nsew signal input
rlabel locali s 346 215 438 289 6 B2
port 4 nsew signal input
rlabel locali s 18 215 84 323 6 C1
port 5 nsew signal input
rlabel locali s 883 129 959 145 6 Y
port 6 nsew signal output
rlabel locali s 487 129 567 145 6 Y
port 6 nsew signal output
rlabel locali s 121 181 181 425 6 Y
port 6 nsew signal output
rlabel locali s 121 173 959 181 6 Y
port 6 nsew signal output
rlabel locali s 105 145 959 173 6 Y
port 6 nsew signal output
rlabel locali s 105 61 181 145 6 Y
port 6 nsew signal output
rlabel metal1 s 0 -48 1196 48 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 496 1196 592 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1231362
string GDS_START 1221708
<< end >>
