magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 2392 561
rect 103 427 169 527
rect 17 195 88 325
rect 287 427 357 527
rect 103 17 169 93
rect 350 201 432 325
rect 682 441 758 527
rect 976 383 1042 527
rect 1465 451 1541 527
rect 287 17 357 93
rect 718 193 784 213
rect 718 147 800 193
rect 1729 451 2006 527
rect 714 17 748 105
rect 1492 147 1567 213
rect 2040 326 2097 493
rect 1863 219 1938 265
rect 1070 17 1136 93
rect 1453 17 1505 105
rect 1940 17 2006 161
rect 2056 143 2097 326
rect 2040 51 2097 143
rect 2230 353 2289 527
rect 2323 289 2375 493
rect 2332 165 2375 289
rect 2230 17 2289 109
rect 2323 51 2375 165
rect 0 -17 2392 17
<< obsli1 >>
rect 17 393 69 493
rect 17 391 168 393
rect 17 359 122 391
rect 156 357 168 391
rect 122 161 168 357
rect 17 127 168 161
rect 203 187 248 493
rect 391 393 425 493
rect 468 450 634 484
rect 203 153 214 187
rect 17 69 69 127
rect 203 69 248 153
rect 282 359 425 393
rect 282 165 316 359
rect 466 357 490 391
rect 524 357 566 391
rect 466 315 566 357
rect 282 127 425 165
rect 466 141 510 315
rect 600 281 634 450
rect 818 407 852 475
rect 668 357 938 407
rect 1251 450 1417 484
rect 1213 391 1260 397
rect 668 315 718 357
rect 820 281 870 297
rect 600 247 870 281
rect 600 239 680 247
rect 546 187 612 203
rect 546 153 578 187
rect 546 129 612 153
rect 391 61 425 127
rect 646 93 680 239
rect 826 231 870 247
rect 904 213 938 357
rect 1213 357 1226 391
rect 972 323 1173 331
rect 972 289 1134 323
rect 1168 289 1173 323
rect 1213 315 1260 357
rect 972 283 1173 289
rect 972 247 1038 283
rect 1308 261 1349 381
rect 1225 255 1349 261
rect 1100 213 1166 247
rect 904 179 1166 213
rect 1225 221 1226 255
rect 1260 225 1349 255
rect 1383 281 1417 450
rect 1589 417 1623 475
rect 1451 383 2006 417
rect 1451 315 1501 383
rect 1383 247 1653 281
rect 1260 221 1282 225
rect 904 153 948 179
rect 882 119 948 153
rect 481 53 680 93
rect 782 85 848 109
rect 982 85 1016 143
rect 1225 141 1282 221
rect 1383 93 1417 247
rect 1609 215 1653 247
rect 1687 156 1723 383
rect 1657 119 1723 156
rect 1757 323 1909 349
rect 1757 289 1778 323
rect 1812 315 1909 323
rect 1757 185 1812 289
rect 1972 265 2006 383
rect 1972 199 2022 265
rect 1757 151 1895 185
rect 782 51 1016 85
rect 1264 53 1417 93
rect 1557 85 1623 109
rect 1757 85 1791 117
rect 1557 51 1791 85
rect 1848 53 1895 151
rect 2131 265 2194 483
rect 2131 199 2298 265
rect 2131 51 2194 199
<< obsli1c >>
rect 122 357 156 391
rect 214 153 248 187
rect 490 357 524 391
rect 578 153 612 187
rect 1226 357 1260 391
rect 1134 289 1168 323
rect 1226 221 1260 255
rect 1778 289 1812 323
<< metal1 >>
rect 0 496 2392 592
rect 754 184 812 193
rect 1490 184 1548 193
rect 754 156 1548 184
rect 754 147 812 156
rect 1490 147 1548 156
rect 0 -48 2392 48
<< obsm1 >>
rect 110 391 168 397
rect 110 357 122 391
rect 156 388 168 391
rect 478 391 536 397
rect 478 388 490 391
rect 156 360 490 388
rect 156 357 168 360
rect 110 351 168 357
rect 478 357 490 360
rect 524 388 536 391
rect 1214 391 1272 397
rect 1214 388 1226 391
rect 524 360 1226 388
rect 524 357 536 360
rect 478 351 536 357
rect 1214 357 1226 360
rect 1260 357 1272 391
rect 1214 351 1272 357
rect 1122 323 1180 329
rect 1122 289 1134 323
rect 1168 320 1180 323
rect 1766 323 1824 329
rect 1766 320 1778 323
rect 1168 292 1778 320
rect 1168 289 1180 292
rect 1122 283 1180 289
rect 1766 289 1778 292
rect 1812 289 1824 323
rect 1766 283 1824 289
rect 1214 255 1272 261
rect 1214 252 1226 255
rect 585 224 1226 252
rect 585 193 624 224
rect 1214 221 1226 224
rect 1260 221 1272 255
rect 1214 215 1272 221
rect 202 187 260 193
rect 202 153 214 187
rect 248 184 260 187
rect 566 187 624 193
rect 566 184 578 187
rect 248 156 578 184
rect 248 153 260 156
rect 202 147 260 153
rect 566 153 578 156
rect 612 153 624 187
rect 566 147 624 153
<< labels >>
rlabel locali s 350 201 432 325 6 D
port 1 nsew signal input
rlabel locali s 2332 165 2375 289 6 Q
port 2 nsew signal output
rlabel locali s 2323 289 2375 493 6 Q
port 2 nsew signal output
rlabel locali s 2323 51 2375 165 6 Q
port 2 nsew signal output
rlabel locali s 2056 143 2097 326 6 Q_N
port 3 nsew signal output
rlabel locali s 2040 326 2097 493 6 Q_N
port 3 nsew signal output
rlabel locali s 2040 51 2097 143 6 Q_N
port 3 nsew signal output
rlabel locali s 1863 219 1938 265 6 RESET_B
port 4 nsew signal input
rlabel locali s 718 193 784 213 6 SET_B
port 5 nsew signal input
rlabel locali s 718 147 800 193 6 SET_B
port 5 nsew signal input
rlabel locali s 1492 147 1567 213 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1490 184 1548 193 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1490 147 1548 156 6 SET_B
port 5 nsew signal input
rlabel metal1 s 754 184 812 193 6 SET_B
port 5 nsew signal input
rlabel metal1 s 754 156 1548 184 6 SET_B
port 5 nsew signal input
rlabel metal1 s 754 147 812 156 6 SET_B
port 5 nsew signal input
rlabel locali s 17 195 88 325 6 CLK
port 6 nsew clock input
rlabel locali s 2230 17 2289 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1940 17 2006 161 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1453 17 1505 105 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1070 17 1136 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 714 17 748 105 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 287 17 357 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 103 17 169 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 2392 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 2392 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 2230 353 2289 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1729 451 2006 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1465 451 1541 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 976 383 1042 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 682 441 758 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 287 427 357 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 103 427 169 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 2392 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 2392 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2392 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3280032
string GDS_START 3261014
<< end >>
