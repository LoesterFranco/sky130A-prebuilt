magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 552 561
rect 105 435 171 527
rect 94 240 179 391
rect 213 331 261 493
rect 395 435 433 527
rect 213 240 322 331
rect 110 17 229 122
rect 263 51 322 240
rect 356 153 434 323
rect 468 153 523 287
rect 467 17 533 119
rect 0 -17 552 17
<< obsli1 >>
rect 19 417 71 493
rect 19 206 60 417
rect 295 401 361 493
rect 467 401 533 493
rect 295 365 533 401
rect 19 156 229 206
rect 19 56 76 156
<< metal1 >>
rect 0 496 552 592
rect 0 -48 552 48
<< labels >>
rlabel locali s 356 153 434 323 6 A1
port 1 nsew signal input
rlabel locali s 468 153 523 287 6 A2
port 2 nsew signal input
rlabel locali s 94 240 179 391 6 B1_N
port 3 nsew signal input
rlabel locali s 263 51 322 240 6 Y
port 4 nsew signal output
rlabel locali s 213 331 261 493 6 Y
port 4 nsew signal output
rlabel locali s 213 240 322 331 6 Y
port 4 nsew signal output
rlabel locali s 467 17 533 119 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 110 17 229 122 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 552 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 552 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 395 435 433 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 105 435 171 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 552 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 552 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 552 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 4003052
string GDS_START 3997876
<< end >>
