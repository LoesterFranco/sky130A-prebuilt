magic
tech sky130A
magscale 1 2
timestamp 1599588244
<< locali >>
rect 25 162 103 314
rect 1341 236 1409 334
rect 2179 308 2213 580
rect 2595 364 2661 596
rect 2179 282 2345 308
rect 2179 264 2375 282
rect 2239 154 2375 264
rect 2239 70 2291 154
rect 2627 226 2661 364
rect 2612 66 2678 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 23 593 287 649
rect 23 388 102 593
rect 321 581 555 615
rect 321 559 355 581
rect 136 525 355 559
rect 136 390 202 525
rect 297 457 394 491
rect 137 128 171 390
rect 205 350 263 356
rect 205 316 223 350
rect 257 316 263 350
rect 205 290 263 316
rect 297 237 331 457
rect 437 423 487 547
rect 521 491 555 581
rect 589 525 639 649
rect 673 581 892 615
rect 673 491 707 581
rect 858 563 892 581
rect 521 457 707 491
rect 758 423 824 547
rect 858 497 992 563
rect 1085 519 1157 596
rect 1198 553 1300 649
rect 1463 581 1644 615
rect 1463 519 1501 581
rect 858 482 895 497
rect 365 389 824 423
rect 365 294 431 389
rect 477 350 551 355
rect 477 316 511 350
rect 545 316 551 350
rect 477 289 551 316
rect 585 311 651 355
rect 777 322 824 389
rect 585 237 619 311
rect 297 203 619 237
rect 669 221 743 277
rect 777 255 827 322
rect 861 221 895 482
rect 1085 485 1501 519
rect 1085 448 1157 485
rect 929 382 1157 448
rect 1341 434 1407 451
rect 1019 368 1157 382
rect 1219 368 1501 434
rect 65 78 171 128
rect 229 17 295 162
rect 329 93 395 203
rect 441 17 507 156
rect 541 85 575 203
rect 669 187 895 221
rect 929 153 979 320
rect 1019 200 1085 368
rect 1219 334 1253 368
rect 1119 268 1307 334
rect 1273 193 1307 268
rect 1542 305 1576 547
rect 1443 271 1576 305
rect 1610 321 1644 581
rect 1678 419 1728 477
rect 1853 458 1925 649
rect 1966 424 2032 477
rect 2073 458 2139 649
rect 1678 385 1779 419
rect 609 119 979 153
rect 1013 132 1239 166
rect 1013 85 1047 132
rect 541 51 1047 85
rect 1121 17 1171 98
rect 1205 85 1239 132
rect 1273 127 1392 193
rect 1443 85 1477 271
rect 1610 255 1711 321
rect 1745 253 1779 385
rect 1813 390 2135 424
rect 1813 291 1866 390
rect 1908 350 1991 356
rect 1908 316 1951 350
rect 1985 316 1991 350
rect 1908 290 1991 316
rect 1511 153 1545 237
rect 1745 221 2067 253
rect 1581 187 2067 221
rect 2101 153 2135 390
rect 2253 348 2319 649
rect 2379 348 2461 556
rect 2495 364 2561 649
rect 2695 364 2761 649
rect 2427 326 2461 348
rect 1511 119 1847 153
rect 1205 51 1756 85
rect 1797 70 1847 119
rect 1883 17 1949 144
rect 2041 70 2135 153
rect 2169 17 2203 220
rect 2427 260 2593 326
rect 2325 17 2393 120
rect 2427 70 2486 260
rect 2526 17 2576 226
rect 2712 17 2764 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 223 316 257 350
rect 511 316 545 350
rect 1951 316 1985 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
<< metal1 >>
rect 0 683 2784 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 0 617 2784 649
rect 0 616 50 617
rect 211 350 269 356
rect 211 316 223 350
rect 257 347 269 350
rect 499 350 557 356
rect 499 347 511 350
rect 257 319 511 347
rect 257 316 269 319
rect 211 310 269 316
rect 499 316 511 319
rect 545 347 557 350
rect 1939 350 1997 356
rect 1939 347 1951 350
rect 545 319 1951 347
rect 545 316 557 319
rect 499 310 557 316
rect 1939 316 1951 319
rect 1985 316 1997 350
rect 1939 310 1997 316
rect 0 49 50 50
rect 0 17 2784 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
rect 0 -49 2784 -17
<< labels >>
rlabel locali s 25 162 103 314 6 D
port 1 nsew signal input
rlabel locali s 2627 226 2661 364 6 Q
port 2 nsew signal output
rlabel locali s 2612 66 2678 226 6 Q
port 2 nsew signal output
rlabel locali s 2595 364 2661 596 6 Q
port 2 nsew signal output
rlabel locali s 2239 154 2375 264 6 Q_N
port 3 nsew signal output
rlabel locali s 2239 70 2291 154 6 Q_N
port 3 nsew signal output
rlabel locali s 2179 308 2213 580 6 Q_N
port 3 nsew signal output
rlabel locali s 2179 282 2345 308 6 Q_N
port 3 nsew signal output
rlabel locali s 2179 264 2375 282 6 Q_N
port 3 nsew signal output
rlabel metal1 s 1939 347 1997 356 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 1939 310 1997 319 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 499 347 557 356 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 499 310 557 319 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 211 347 269 356 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 211 319 1997 347 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 211 310 269 319 6 RESET_B
port 4 nsew signal input
rlabel locali s 1341 236 1409 334 6 CLK
port 5 nsew clock input
rlabel metal1 s 0 -49 2784 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 7 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 617 2784 715 6 VPWR
port 9 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2784 666
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 2623448
string GDS_START 2603700
<< end >>
