magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1104 561
rect 103 367 164 527
rect 683 451 749 527
rect 86 199 148 265
rect 296 199 350 323
rect 393 199 487 265
rect 536 199 679 265
rect 783 349 817 493
rect 851 383 917 527
rect 951 349 985 493
rect 1019 383 1085 527
rect 783 315 1086 349
rect 114 161 148 199
rect 536 161 570 199
rect 114 127 570 161
rect 1040 161 1086 315
rect 783 127 1086 161
rect 103 17 169 93
rect 683 17 749 93
rect 783 51 817 127
rect 851 17 917 93
rect 951 51 985 127
rect 1019 17 1085 93
rect 0 -17 1104 17
<< obsli1 >>
rect 18 333 69 493
rect 198 455 554 489
rect 198 387 268 455
rect 615 421 649 493
rect 306 387 649 421
rect 713 353 747 357
rect 18 299 216 333
rect 18 125 52 299
rect 182 199 216 299
rect 396 319 747 353
rect 713 249 747 319
rect 713 215 1006 249
rect 713 165 747 215
rect 612 131 747 165
rect 18 59 69 125
rect 612 93 646 131
rect 395 59 646 93
<< metal1 >>
rect 0 496 1104 592
rect 0 -48 1104 48
<< labels >>
rlabel locali s 296 199 350 323 6 A0
port 1 nsew signal input
rlabel locali s 393 199 487 265 6 A1
port 2 nsew signal input
rlabel locali s 536 199 679 265 6 S
port 3 nsew signal input
rlabel locali s 536 161 570 199 6 S
port 3 nsew signal input
rlabel locali s 114 161 148 199 6 S
port 3 nsew signal input
rlabel locali s 114 127 570 161 6 S
port 3 nsew signal input
rlabel locali s 86 199 148 265 6 S
port 3 nsew signal input
rlabel locali s 1040 161 1086 315 6 X
port 4 nsew signal output
rlabel locali s 951 349 985 493 6 X
port 4 nsew signal output
rlabel locali s 951 51 985 127 6 X
port 4 nsew signal output
rlabel locali s 783 349 817 493 6 X
port 4 nsew signal output
rlabel locali s 783 315 1086 349 6 X
port 4 nsew signal output
rlabel locali s 783 127 1086 161 6 X
port 4 nsew signal output
rlabel locali s 783 51 817 127 6 X
port 4 nsew signal output
rlabel locali s 1019 17 1085 93 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 851 17 917 93 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 683 17 749 93 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 103 17 169 93 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 1104 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1104 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 1019 383 1085 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 851 383 917 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 683 451 749 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 103 367 164 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 1104 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 1104 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1104 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1659120
string GDS_START 1650786
<< end >>
