magic
tech sky130A
magscale 1 2
timestamp 1604502705
<< nwell >>
rect -38 332 2726 704
<< pwell >>
rect 0 0 2688 49
<< scnmos >>
rect 93 74 123 158
rect 193 74 223 158
rect 271 74 301 158
rect 420 74 450 158
rect 498 74 528 158
rect 600 74 630 222
rect 798 74 828 222
rect 991 97 1021 181
rect 1143 97 1173 181
rect 1243 74 1273 158
rect 1395 74 1425 184
rect 1481 74 1511 184
rect 1633 74 1663 158
rect 1711 74 1741 158
rect 1887 74 1917 222
rect 2099 74 2129 222
rect 2185 74 2215 222
rect 2383 98 2413 226
rect 2485 78 2515 226
rect 2574 78 2604 226
<< pmoshvt >>
rect 118 453 148 581
rect 208 453 238 581
rect 292 453 322 581
rect 393 453 423 581
rect 490 453 520 581
rect 632 368 662 592
rect 878 368 908 592
rect 1080 499 1110 583
rect 1187 499 1217 583
rect 1271 499 1301 583
rect 1395 424 1425 592
rect 1554 424 1584 592
rect 1661 508 1691 592
rect 1745 508 1775 592
rect 1893 392 1923 592
rect 2091 368 2121 592
rect 2181 368 2211 592
rect 2379 368 2409 568
rect 2484 368 2514 592
rect 2574 368 2604 592
<< ndiff >>
rect 543 210 600 222
rect 543 176 555 210
rect 589 176 600 210
rect 543 158 600 176
rect 36 125 93 158
rect 36 91 48 125
rect 82 91 93 125
rect 36 74 93 91
rect 123 125 193 158
rect 123 91 148 125
rect 182 91 193 125
rect 123 74 193 91
rect 223 74 271 158
rect 301 128 420 158
rect 301 94 343 128
rect 377 94 420 128
rect 301 74 420 94
rect 450 74 498 158
rect 528 120 600 158
rect 528 86 555 120
rect 589 86 600 120
rect 528 74 600 86
rect 630 210 687 222
rect 630 176 641 210
rect 675 176 687 210
rect 630 120 687 176
rect 630 86 641 120
rect 675 86 687 120
rect 630 74 687 86
rect 741 136 798 222
rect 741 102 753 136
rect 787 102 798 136
rect 741 74 798 102
rect 828 210 882 222
rect 828 176 839 210
rect 873 176 882 210
rect 828 120 882 176
rect 828 86 839 120
rect 873 86 882 120
rect 936 169 991 181
rect 936 135 946 169
rect 980 135 991 169
rect 936 97 991 135
rect 1021 156 1143 181
rect 1021 122 1098 156
rect 1132 122 1143 156
rect 1021 97 1143 122
rect 1173 158 1223 181
rect 1345 158 1395 184
rect 1173 97 1243 158
rect 828 74 882 86
rect 1193 74 1243 97
rect 1273 120 1395 158
rect 1273 86 1284 120
rect 1318 86 1395 120
rect 1273 74 1395 86
rect 1425 170 1481 184
rect 1425 136 1436 170
rect 1470 136 1481 170
rect 1425 74 1481 136
rect 1511 158 1561 184
rect 1837 158 1887 222
rect 1511 133 1633 158
rect 1511 99 1588 133
rect 1622 99 1633 133
rect 1511 74 1633 99
rect 1663 74 1711 158
rect 1741 127 1887 158
rect 1741 93 1752 127
rect 1786 124 1887 127
rect 1786 93 1842 124
rect 1741 90 1842 93
rect 1876 90 1887 124
rect 1741 74 1887 90
rect 1917 141 1974 222
rect 1917 107 1928 141
rect 1962 107 1974 141
rect 1917 74 1974 107
rect 2028 210 2099 222
rect 2028 176 2040 210
rect 2074 176 2099 210
rect 2028 120 2099 176
rect 2028 86 2040 120
rect 2074 86 2099 120
rect 2028 74 2099 86
rect 2129 210 2185 222
rect 2129 176 2140 210
rect 2174 176 2185 210
rect 2129 120 2185 176
rect 2129 86 2140 120
rect 2174 86 2185 120
rect 2129 74 2185 86
rect 2215 210 2272 222
rect 2215 176 2226 210
rect 2260 176 2272 210
rect 2215 120 2272 176
rect 2215 86 2226 120
rect 2260 86 2272 120
rect 2326 218 2383 226
rect 2326 184 2338 218
rect 2372 184 2383 218
rect 2326 150 2383 184
rect 2326 116 2338 150
rect 2372 116 2383 150
rect 2326 98 2383 116
rect 2413 214 2485 226
rect 2413 180 2434 214
rect 2468 180 2485 214
rect 2413 127 2485 180
rect 2413 98 2440 127
rect 2215 74 2272 86
rect 2428 93 2440 98
rect 2474 93 2485 127
rect 2428 78 2485 93
rect 2515 214 2574 226
rect 2515 180 2527 214
rect 2561 180 2574 214
rect 2515 78 2574 180
rect 2604 142 2654 226
rect 2604 127 2661 142
rect 2604 93 2615 127
rect 2649 93 2661 127
rect 2604 78 2661 93
<< pdiff >>
rect 1319 625 1377 637
rect 538 592 614 604
rect 538 581 559 592
rect 42 569 118 581
rect 42 535 54 569
rect 88 535 118 569
rect 42 499 118 535
rect 42 465 54 499
rect 88 465 118 499
rect 42 453 118 465
rect 148 569 208 581
rect 148 535 161 569
rect 195 535 208 569
rect 148 499 208 535
rect 148 465 161 499
rect 195 465 208 499
rect 148 453 208 465
rect 238 453 292 581
rect 322 569 393 581
rect 322 535 346 569
rect 380 535 393 569
rect 322 499 393 535
rect 322 465 346 499
rect 380 465 393 499
rect 322 453 393 465
rect 423 453 490 581
rect 520 558 559 581
rect 593 558 632 592
rect 520 453 632 558
rect 579 368 632 453
rect 662 440 763 592
rect 662 406 676 440
rect 710 406 763 440
rect 662 368 763 406
rect 819 578 878 592
rect 819 544 831 578
rect 865 544 878 578
rect 819 368 878 544
rect 908 419 967 592
rect 1319 591 1331 625
rect 1365 592 1377 625
rect 1365 591 1395 592
rect 1319 583 1395 591
rect 1021 560 1080 583
rect 1021 526 1033 560
rect 1067 526 1080 560
rect 1021 499 1080 526
rect 1110 558 1187 583
rect 1110 524 1123 558
rect 1157 524 1187 558
rect 1110 499 1187 524
rect 1217 499 1271 583
rect 1301 499 1395 583
rect 908 385 921 419
rect 955 385 967 419
rect 908 368 967 385
rect 1342 424 1395 499
rect 1425 473 1554 592
rect 1425 439 1441 473
rect 1475 439 1554 473
rect 1425 424 1554 439
rect 1584 580 1661 592
rect 1584 546 1597 580
rect 1631 546 1661 580
rect 1584 508 1661 546
rect 1691 508 1745 592
rect 1775 580 1893 592
rect 1775 546 1812 580
rect 1846 546 1893 580
rect 1775 508 1893 546
rect 1584 470 1643 508
rect 1584 436 1597 470
rect 1631 436 1643 470
rect 1584 424 1643 436
rect 1840 392 1893 508
rect 1923 580 1980 592
rect 1923 546 1936 580
rect 1970 546 1980 580
rect 1923 509 1980 546
rect 1923 475 1936 509
rect 1970 475 1980 509
rect 1923 438 1980 475
rect 1923 404 1936 438
rect 1970 404 1980 438
rect 1923 392 1980 404
rect 2034 580 2091 592
rect 2034 546 2044 580
rect 2078 546 2091 580
rect 2034 497 2091 546
rect 2034 463 2044 497
rect 2078 463 2091 497
rect 2034 414 2091 463
rect 2034 380 2044 414
rect 2078 380 2091 414
rect 2034 368 2091 380
rect 2121 580 2181 592
rect 2121 546 2134 580
rect 2168 546 2181 580
rect 2121 497 2181 546
rect 2121 463 2134 497
rect 2168 463 2181 497
rect 2121 414 2181 463
rect 2121 380 2134 414
rect 2168 380 2181 414
rect 2121 368 2181 380
rect 2211 580 2268 592
rect 2211 546 2224 580
rect 2258 546 2268 580
rect 2427 580 2484 592
rect 2427 568 2437 580
rect 2211 497 2268 546
rect 2211 463 2224 497
rect 2258 463 2268 497
rect 2211 414 2268 463
rect 2211 380 2224 414
rect 2258 380 2268 414
rect 2211 368 2268 380
rect 2322 556 2379 568
rect 2322 522 2332 556
rect 2366 522 2379 556
rect 2322 485 2379 522
rect 2322 451 2332 485
rect 2366 451 2379 485
rect 2322 414 2379 451
rect 2322 380 2332 414
rect 2366 380 2379 414
rect 2322 368 2379 380
rect 2409 546 2437 568
rect 2471 546 2484 580
rect 2409 497 2484 546
rect 2409 463 2437 497
rect 2471 463 2484 497
rect 2409 414 2484 463
rect 2409 380 2437 414
rect 2471 380 2484 414
rect 2409 368 2484 380
rect 2514 580 2574 592
rect 2514 546 2527 580
rect 2561 546 2574 580
rect 2514 497 2574 546
rect 2514 463 2527 497
rect 2561 463 2574 497
rect 2514 414 2574 463
rect 2514 380 2527 414
rect 2561 380 2574 414
rect 2514 368 2574 380
rect 2604 580 2661 592
rect 2604 546 2617 580
rect 2651 546 2661 580
rect 2604 498 2661 546
rect 2604 464 2617 498
rect 2651 464 2661 498
rect 2604 368 2661 464
<< ndiffc >>
rect 555 176 589 210
rect 48 91 82 125
rect 148 91 182 125
rect 343 94 377 128
rect 555 86 589 120
rect 641 176 675 210
rect 641 86 675 120
rect 753 102 787 136
rect 839 176 873 210
rect 839 86 873 120
rect 946 135 980 169
rect 1098 122 1132 156
rect 1284 86 1318 120
rect 1436 136 1470 170
rect 1588 99 1622 133
rect 1752 93 1786 127
rect 1842 90 1876 124
rect 1928 107 1962 141
rect 2040 176 2074 210
rect 2040 86 2074 120
rect 2140 176 2174 210
rect 2140 86 2174 120
rect 2226 176 2260 210
rect 2226 86 2260 120
rect 2338 184 2372 218
rect 2338 116 2372 150
rect 2434 180 2468 214
rect 2440 93 2474 127
rect 2527 180 2561 214
rect 2615 93 2649 127
<< pdiffc >>
rect 54 535 88 569
rect 54 465 88 499
rect 161 535 195 569
rect 161 465 195 499
rect 346 535 380 569
rect 346 465 380 499
rect 559 558 593 592
rect 676 406 710 440
rect 831 544 865 578
rect 1331 591 1365 625
rect 1033 526 1067 560
rect 1123 524 1157 558
rect 921 385 955 419
rect 1441 439 1475 473
rect 1597 546 1631 580
rect 1812 546 1846 580
rect 1597 436 1631 470
rect 1936 546 1970 580
rect 1936 475 1970 509
rect 1936 404 1970 438
rect 2044 546 2078 580
rect 2044 463 2078 497
rect 2044 380 2078 414
rect 2134 546 2168 580
rect 2134 463 2168 497
rect 2134 380 2168 414
rect 2224 546 2258 580
rect 2224 463 2258 497
rect 2224 380 2258 414
rect 2332 522 2366 556
rect 2332 451 2366 485
rect 2332 380 2366 414
rect 2437 546 2471 580
rect 2437 463 2471 497
rect 2437 380 2471 414
rect 2527 546 2561 580
rect 2527 463 2561 497
rect 2527 380 2561 414
rect 2617 546 2651 580
rect 2617 464 2651 498
<< poly >>
rect 118 581 148 607
rect 208 581 238 607
rect 292 581 322 607
rect 393 581 423 607
rect 490 581 520 607
rect 632 592 662 618
rect 878 592 908 618
rect 118 438 148 453
rect 208 438 238 453
rect 292 438 322 453
rect 393 438 423 453
rect 490 438 520 453
rect 39 408 241 438
rect 39 246 69 408
rect 289 360 325 438
rect 390 411 426 438
rect 487 421 523 438
rect 373 395 439 411
rect 373 361 389 395
rect 423 361 439 395
rect 117 344 223 360
rect 117 310 133 344
rect 167 310 223 344
rect 117 294 223 310
rect 265 344 331 360
rect 373 345 439 361
rect 481 405 547 421
rect 481 371 497 405
rect 531 371 547 405
rect 481 355 547 371
rect 1080 583 1110 609
rect 1187 583 1217 609
rect 1271 583 1301 609
rect 1395 592 1425 618
rect 1554 592 1584 618
rect 1661 592 1691 618
rect 1745 592 1775 618
rect 1893 592 1923 618
rect 2091 592 2121 618
rect 2181 592 2211 618
rect 1080 484 1110 499
rect 1187 484 1217 499
rect 1271 484 1301 499
rect 1077 467 1113 484
rect 1001 451 1113 467
rect 1001 417 1017 451
rect 1051 437 1113 451
rect 1184 449 1220 484
rect 1051 417 1067 437
rect 1001 401 1067 417
rect 1160 433 1226 449
rect 1160 399 1176 433
rect 1210 399 1226 433
rect 265 310 281 344
rect 315 310 331 344
rect 265 294 331 310
rect 39 230 151 246
rect 39 196 101 230
rect 135 196 151 230
rect 39 180 151 196
rect 93 158 123 180
rect 193 158 223 294
rect 271 158 301 294
rect 349 230 450 246
rect 349 196 365 230
rect 399 196 450 230
rect 349 180 450 196
rect 420 158 450 180
rect 498 158 528 355
rect 632 353 662 368
rect 878 353 908 368
rect 1160 353 1226 399
rect 629 336 665 353
rect 629 320 719 336
rect 629 300 669 320
rect 600 286 669 300
rect 703 286 719 320
rect 600 270 719 286
rect 762 323 1226 353
rect 762 320 828 323
rect 762 286 778 320
rect 812 286 828 320
rect 762 270 828 286
rect 600 222 630 270
rect 798 222 828 270
rect 991 181 1021 323
rect 1268 281 1304 484
rect 1661 493 1691 508
rect 1745 493 1775 508
rect 1658 428 1694 493
rect 1742 476 1778 493
rect 1742 460 1808 476
rect 1395 409 1425 424
rect 1554 409 1584 424
rect 1392 389 1428 409
rect 1346 373 1428 389
rect 1551 386 1587 409
rect 1658 398 1700 428
rect 1742 426 1758 460
rect 1792 426 1808 460
rect 1742 410 1808 426
rect 1346 339 1362 373
rect 1396 339 1428 373
rect 1346 323 1428 339
rect 1513 370 1587 386
rect 1513 336 1529 370
rect 1563 350 1587 370
rect 1563 336 1628 350
rect 1135 259 1201 275
rect 1135 225 1151 259
rect 1185 225 1201 259
rect 1135 209 1201 225
rect 1243 265 1316 281
rect 1243 231 1266 265
rect 1300 231 1316 265
rect 1243 215 1316 231
rect 1143 181 1173 209
rect 1243 158 1273 215
rect 1395 184 1425 323
rect 1513 320 1628 336
rect 1481 256 1556 272
rect 1481 222 1506 256
rect 1540 222 1556 256
rect 1481 206 1556 222
rect 1481 184 1511 206
rect 1598 203 1628 320
rect 1670 311 1700 398
rect 1670 295 1736 311
rect 1670 261 1686 295
rect 1720 261 1736 295
rect 1670 245 1736 261
rect 1778 203 1808 410
rect 1893 377 1923 392
rect 1890 310 1926 377
rect 2379 568 2409 594
rect 2484 592 2514 618
rect 2574 592 2604 618
rect 2091 353 2121 368
rect 2181 353 2211 368
rect 2379 353 2409 368
rect 2484 353 2514 368
rect 2574 353 2604 368
rect 2088 326 2124 353
rect 1856 294 1926 310
rect 1856 260 1872 294
rect 1906 260 1926 294
rect 1988 310 2129 326
rect 1988 276 2004 310
rect 2038 276 2072 310
rect 2106 290 2129 310
rect 2178 290 2214 353
rect 2376 290 2412 353
rect 2481 330 2517 353
rect 2571 330 2607 353
rect 2481 314 2607 330
rect 2106 276 2413 290
rect 1988 260 2413 276
rect 2481 280 2497 314
rect 2531 280 2607 314
rect 2481 264 2607 280
rect 1856 244 1926 260
rect 1887 222 1917 244
rect 2099 222 2129 260
rect 2185 222 2215 260
rect 2383 226 2413 260
rect 2485 226 2515 264
rect 2574 226 2604 264
rect 93 48 123 74
rect 193 48 223 74
rect 271 48 301 74
rect 420 48 450 74
rect 498 48 528 74
rect 600 48 630 74
rect 798 48 828 74
rect 991 71 1021 97
rect 1143 71 1173 97
rect 1598 173 1663 203
rect 1633 158 1663 173
rect 1711 173 1808 203
rect 1711 158 1741 173
rect 1243 48 1273 74
rect 1395 48 1425 74
rect 1481 48 1511 74
rect 1633 48 1663 74
rect 1711 48 1741 74
rect 1887 48 1917 74
rect 2099 48 2129 74
rect 2185 48 2215 74
rect 2383 72 2413 98
rect 2485 52 2515 78
rect 2574 52 2604 78
<< polycont >>
rect 389 361 423 395
rect 133 310 167 344
rect 497 371 531 405
rect 1017 417 1051 451
rect 1176 399 1210 433
rect 281 310 315 344
rect 101 196 135 230
rect 365 196 399 230
rect 669 286 703 320
rect 778 286 812 320
rect 1758 426 1792 460
rect 1362 339 1396 373
rect 1529 336 1563 370
rect 1151 225 1185 259
rect 1266 231 1300 265
rect 1506 222 1540 256
rect 1686 261 1720 295
rect 1872 260 1906 294
rect 2004 276 2038 310
rect 2072 276 2106 310
rect 2497 280 2531 314
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2688 683
rect 17 569 104 585
rect 17 535 54 569
rect 88 535 104 569
rect 17 499 104 535
rect 17 465 54 499
rect 88 465 104 499
rect 17 360 104 465
rect 145 569 211 649
rect 534 592 618 649
rect 145 535 161 569
rect 195 535 211 569
rect 145 499 211 535
rect 145 465 161 499
rect 195 465 211 499
rect 145 462 211 465
rect 330 569 396 585
rect 330 535 346 569
rect 380 535 396 569
rect 534 558 559 592
rect 593 558 618 592
rect 534 542 618 558
rect 815 578 881 649
rect 1315 625 1381 649
rect 1315 591 1331 625
rect 1365 591 1381 625
rect 815 544 831 578
rect 865 544 881 578
rect 815 542 881 544
rect 1017 560 1067 587
rect 330 508 396 535
rect 1017 533 1033 560
rect 915 526 1033 533
rect 915 508 1067 526
rect 330 499 1067 508
rect 1101 558 1173 587
rect 1101 524 1123 558
rect 1157 524 1173 558
rect 1581 580 1647 596
rect 330 465 346 499
rect 380 474 949 499
rect 1101 495 1173 524
rect 1207 523 1547 557
rect 380 465 396 474
rect 330 462 396 465
rect 149 395 439 428
rect 149 394 389 395
rect 149 360 183 394
rect 373 361 389 394
rect 423 361 439 395
rect 17 344 183 360
rect 17 310 133 344
rect 167 310 183 344
rect 17 294 183 310
rect 217 344 331 360
rect 373 345 439 361
rect 481 405 551 430
rect 481 371 497 405
rect 531 371 551 405
rect 481 355 551 371
rect 217 310 281 344
rect 315 310 331 344
rect 217 294 331 310
rect 585 304 619 474
rect 659 406 676 440
rect 710 406 819 440
rect 659 390 819 406
rect 17 146 51 294
rect 449 270 619 304
rect 653 320 737 356
rect 653 286 669 320
rect 703 286 737 320
rect 653 270 737 286
rect 771 320 819 390
rect 771 286 778 320
rect 812 286 819 320
rect 853 330 887 474
rect 1001 451 1067 465
rect 1001 440 1017 451
rect 921 419 1017 440
rect 955 417 1017 419
rect 1051 417 1067 451
rect 955 401 1067 417
rect 955 385 971 401
rect 921 364 971 385
rect 853 296 980 330
rect 771 270 819 286
rect 85 230 415 246
rect 85 196 101 230
rect 135 196 365 230
rect 399 196 415 230
rect 85 180 415 196
rect 313 162 415 180
rect 17 125 98 146
rect 17 91 48 125
rect 82 91 98 125
rect 17 70 98 91
rect 132 125 198 146
rect 449 128 483 270
rect 771 236 805 270
rect 132 91 148 125
rect 182 91 198 125
rect 132 17 198 91
rect 296 94 343 128
rect 377 94 483 128
rect 296 78 483 94
rect 539 210 589 226
rect 539 176 555 210
rect 539 120 589 176
rect 539 86 555 120
rect 539 17 589 86
rect 625 210 805 236
rect 625 176 641 210
rect 675 202 805 210
rect 839 210 889 226
rect 675 176 691 202
rect 625 120 691 176
rect 873 176 889 210
rect 625 86 641 120
rect 675 86 691 120
rect 625 70 691 86
rect 737 136 803 168
rect 737 102 753 136
rect 787 102 803 136
rect 737 17 803 102
rect 839 120 889 176
rect 873 86 889 120
rect 930 169 980 296
rect 930 135 946 169
rect 930 119 980 135
rect 839 85 889 86
rect 1014 85 1048 401
rect 1101 349 1135 495
rect 1207 449 1241 523
rect 1169 433 1241 449
rect 1169 399 1176 433
rect 1210 399 1241 433
rect 1422 473 1479 489
rect 1422 439 1441 473
rect 1475 439 1479 473
rect 1422 423 1479 439
rect 1169 383 1241 399
rect 1346 373 1402 389
rect 1346 349 1362 373
rect 1082 339 1362 349
rect 1396 339 1402 373
rect 1082 315 1402 339
rect 1082 175 1116 315
rect 1436 281 1470 423
rect 1513 386 1547 523
rect 1581 546 1597 580
rect 1631 546 1647 580
rect 1581 470 1647 546
rect 1772 580 1886 649
rect 1772 546 1812 580
rect 1846 546 1886 580
rect 1772 530 1886 546
rect 1920 580 1990 596
rect 1920 546 1936 580
rect 1970 546 1990 580
rect 1920 509 1990 546
rect 1920 476 1936 509
rect 1581 436 1597 470
rect 1631 436 1647 470
rect 1581 420 1647 436
rect 1513 370 1579 386
rect 1513 336 1529 370
rect 1563 336 1579 370
rect 1613 378 1647 420
rect 1742 475 1936 476
rect 1970 475 1990 509
rect 1742 460 1990 475
rect 1742 426 1758 460
rect 1792 438 1990 460
rect 1792 426 1936 438
rect 1742 412 1936 426
rect 1920 404 1936 412
rect 1970 404 1990 438
rect 1920 388 1990 404
rect 1613 344 1804 378
rect 1513 320 1579 336
rect 1150 259 1216 275
rect 1150 225 1151 259
rect 1185 225 1216 259
rect 1150 209 1216 225
rect 1250 265 1470 281
rect 1670 295 1736 310
rect 1670 279 1686 295
rect 1250 231 1266 265
rect 1300 231 1470 265
rect 1250 222 1470 231
rect 1182 188 1216 209
rect 1082 156 1148 175
rect 1082 122 1098 156
rect 1132 122 1148 156
rect 1082 119 1148 122
rect 1182 154 1402 188
rect 1182 85 1216 154
rect 839 51 1216 85
rect 1268 86 1284 120
rect 1318 86 1334 120
rect 1268 17 1334 86
rect 1368 85 1402 154
rect 1436 170 1470 222
rect 1436 119 1470 136
rect 1504 261 1686 279
rect 1720 261 1736 295
rect 1504 256 1736 261
rect 1504 222 1506 256
rect 1540 245 1736 256
rect 1770 245 1804 344
rect 1956 326 1990 388
rect 2028 580 2078 649
rect 2028 546 2044 580
rect 2028 497 2078 546
rect 2028 463 2044 497
rect 2028 414 2078 463
rect 2028 380 2044 414
rect 2028 364 2078 380
rect 2118 580 2168 596
rect 2118 546 2134 580
rect 2118 497 2168 546
rect 2118 463 2134 497
rect 2118 414 2168 463
rect 2208 580 2274 649
rect 2208 546 2224 580
rect 2258 546 2274 580
rect 2421 580 2471 649
rect 2208 497 2274 546
rect 2208 463 2224 497
rect 2258 463 2274 497
rect 2208 428 2274 463
rect 2118 380 2134 414
rect 2224 414 2274 428
rect 2168 380 2190 394
rect 2118 360 2190 380
rect 2258 380 2274 414
rect 2224 364 2274 380
rect 2316 556 2382 572
rect 2316 522 2332 556
rect 2366 522 2382 556
rect 2316 485 2382 522
rect 2316 451 2332 485
rect 2366 451 2382 485
rect 2316 414 2382 451
rect 2316 380 2332 414
rect 2366 380 2382 414
rect 1956 310 2122 326
rect 1856 294 1922 310
rect 1856 260 1872 294
rect 1906 260 1922 294
rect 1856 245 1922 260
rect 1540 222 1556 245
rect 1504 206 1556 222
rect 1770 211 1922 245
rect 1956 276 2004 310
rect 2038 276 2072 310
rect 2106 276 2122 310
rect 1956 260 2122 276
rect 1504 85 1538 206
rect 1604 177 1804 211
rect 1956 177 1990 260
rect 2156 226 2190 360
rect 2316 330 2382 380
rect 2421 546 2437 580
rect 2421 497 2471 546
rect 2421 463 2437 497
rect 2421 414 2471 463
rect 2421 380 2437 414
rect 2421 364 2471 380
rect 2511 580 2567 596
rect 2511 546 2527 580
rect 2561 546 2567 580
rect 2511 497 2567 546
rect 2511 463 2527 497
rect 2561 463 2567 497
rect 2601 580 2667 649
rect 2601 546 2617 580
rect 2651 546 2667 580
rect 2601 498 2667 546
rect 2601 464 2617 498
rect 2651 464 2667 498
rect 2511 430 2567 463
rect 2511 414 2663 430
rect 2511 380 2527 414
rect 2561 380 2663 414
rect 2511 364 2663 380
rect 2316 314 2547 330
rect 2316 280 2497 314
rect 2531 280 2547 314
rect 2316 264 2547 280
rect 1604 162 1638 177
rect 1368 51 1538 85
rect 1572 133 1638 162
rect 1572 99 1588 133
rect 1622 99 1638 133
rect 1572 70 1638 99
rect 1736 127 1878 143
rect 1736 93 1752 127
rect 1786 124 1878 127
rect 1786 93 1842 124
rect 1736 90 1842 93
rect 1876 90 1878 124
rect 1736 17 1878 90
rect 1912 141 1990 177
rect 1912 107 1928 141
rect 1962 107 1990 141
rect 1912 70 1990 107
rect 2024 210 2090 226
rect 2024 176 2040 210
rect 2074 176 2090 210
rect 2024 120 2090 176
rect 2024 86 2040 120
rect 2074 86 2090 120
rect 2024 17 2090 86
rect 2124 210 2190 226
rect 2124 176 2140 210
rect 2174 176 2190 210
rect 2124 120 2190 176
rect 2124 86 2140 120
rect 2174 86 2190 120
rect 2124 70 2190 86
rect 2226 210 2276 226
rect 2260 176 2276 210
rect 2226 120 2276 176
rect 2260 86 2276 120
rect 2316 218 2388 264
rect 2615 230 2663 364
rect 2316 184 2338 218
rect 2372 184 2388 218
rect 2316 150 2388 184
rect 2316 116 2338 150
rect 2372 116 2388 150
rect 2316 112 2388 116
rect 2424 214 2476 230
rect 2424 180 2434 214
rect 2468 180 2476 214
rect 2510 214 2663 230
rect 2510 180 2527 214
rect 2561 180 2663 214
rect 2424 146 2476 180
rect 2424 127 2490 146
rect 2226 17 2276 86
rect 2424 93 2440 127
rect 2474 93 2490 127
rect 2424 17 2490 93
rect 2599 127 2665 146
rect 2599 93 2615 127
rect 2649 93 2665 127
rect 2599 17 2665 93
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2688 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
<< metal1 >>
rect 0 683 2688 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2688 683
rect 0 617 2688 649
rect 0 17 2688 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2688 17
rect 0 -49 2688 -17
<< labels >>
rlabel comment s 0 0 0 0 4 sdfxbp_2
flabel comment s 1004 343 1004 343 0 FreeSans 200 0 0 0 no_jumper_check
flabel pwell s 0 0 2688 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 2688 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 2688 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 2688 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 319 168 353 202 0 FreeSans 340 0 0 0 SCE
port 4 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 511 390 545 424 0 FreeSans 340 0 0 0 SCD
port 3 nsew
flabel corelocali s 2143 94 2177 128 0 FreeSans 340 0 0 0 Q
port 9 nsew
flabel corelocali s 2143 168 2177 202 0 FreeSans 340 0 0 0 Q
port 9 nsew
flabel corelocali s 2623 242 2657 276 0 FreeSans 340 0 0 0 Q_N
port 10 nsew
flabel corelocali s 2623 316 2657 350 0 FreeSans 340 0 0 0 Q_N
port 10 nsew
flabel corelocali s 2623 390 2657 424 0 FreeSans 340 0 0 0 Q_N
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 2688 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 277842
string GDS_START 258190
<< end >>
