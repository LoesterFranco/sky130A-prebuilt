magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 93 47 123 177
rect 177 47 207 177
rect 281 47 311 177
rect 367 47 397 177
rect 565 47 595 177
rect 659 47 689 177
rect 760 47 790 177
rect 844 47 874 177
rect 948 47 978 177
rect 1032 47 1062 177
<< pmoshvt >>
rect 85 297 121 497
rect 179 297 215 497
rect 273 297 309 497
rect 369 297 405 497
rect 557 297 593 497
rect 651 297 687 497
rect 752 297 788 497
rect 846 297 882 497
rect 940 297 976 497
rect 1034 297 1070 497
<< ndiff >>
rect 27 163 93 177
rect 27 129 39 163
rect 73 129 93 163
rect 27 95 93 129
rect 27 61 39 95
rect 73 61 93 95
rect 27 47 93 61
rect 123 163 177 177
rect 123 129 133 163
rect 167 129 177 163
rect 123 95 177 129
rect 123 61 133 95
rect 167 61 177 95
rect 123 47 177 61
rect 207 163 281 177
rect 207 129 227 163
rect 261 129 281 163
rect 207 47 281 129
rect 311 95 367 177
rect 311 61 321 95
rect 355 61 367 95
rect 311 47 367 61
rect 397 95 449 177
rect 397 61 407 95
rect 441 61 449 95
rect 397 47 449 61
rect 503 95 565 177
rect 503 61 511 95
rect 545 61 565 95
rect 503 47 565 61
rect 595 163 659 177
rect 595 129 605 163
rect 639 129 659 163
rect 595 47 659 129
rect 689 163 760 177
rect 689 129 699 163
rect 733 129 760 163
rect 689 95 760 129
rect 689 61 699 95
rect 733 61 760 95
rect 689 47 760 61
rect 790 95 844 177
rect 790 61 800 95
rect 834 61 844 95
rect 790 47 844 61
rect 874 163 948 177
rect 874 129 894 163
rect 928 129 948 163
rect 874 95 948 129
rect 874 61 894 95
rect 928 61 948 95
rect 874 47 948 61
rect 978 95 1032 177
rect 978 61 988 95
rect 1022 61 1032 95
rect 978 47 1032 61
rect 1062 163 1124 177
rect 1062 129 1082 163
rect 1116 129 1124 163
rect 1062 95 1124 129
rect 1062 61 1082 95
rect 1116 61 1124 95
rect 1062 47 1124 61
<< pdiff >>
rect 27 477 85 497
rect 27 443 39 477
rect 73 443 85 477
rect 27 409 85 443
rect 27 375 39 409
rect 73 375 85 409
rect 27 297 85 375
rect 121 477 179 497
rect 121 443 133 477
rect 167 443 179 477
rect 121 409 179 443
rect 121 375 133 409
rect 167 375 179 409
rect 121 297 179 375
rect 215 477 273 497
rect 215 443 227 477
rect 261 443 273 477
rect 215 297 273 443
rect 309 391 369 497
rect 309 357 321 391
rect 355 357 369 391
rect 309 297 369 357
rect 405 477 557 497
rect 405 443 417 477
rect 451 443 511 477
rect 545 443 557 477
rect 405 297 557 443
rect 593 477 651 497
rect 593 443 605 477
rect 639 443 651 477
rect 593 409 651 443
rect 593 375 605 409
rect 639 375 651 409
rect 593 341 651 375
rect 593 307 605 341
rect 639 307 651 341
rect 593 297 651 307
rect 687 477 752 497
rect 687 443 699 477
rect 733 443 752 477
rect 687 297 752 443
rect 788 477 846 497
rect 788 443 800 477
rect 834 443 846 477
rect 788 297 846 443
rect 882 409 940 497
rect 882 375 894 409
rect 928 375 940 409
rect 882 297 940 375
rect 976 477 1034 497
rect 976 443 988 477
rect 1022 443 1034 477
rect 976 409 1034 443
rect 976 375 988 409
rect 1022 375 1034 409
rect 976 297 1034 375
rect 1070 477 1129 497
rect 1070 443 1083 477
rect 1117 443 1129 477
rect 1070 409 1129 443
rect 1070 375 1083 409
rect 1117 375 1129 409
rect 1070 297 1129 375
<< ndiffc >>
rect 39 129 73 163
rect 39 61 73 95
rect 133 129 167 163
rect 133 61 167 95
rect 227 129 261 163
rect 321 61 355 95
rect 407 61 441 95
rect 511 61 545 95
rect 605 129 639 163
rect 699 129 733 163
rect 699 61 733 95
rect 800 61 834 95
rect 894 129 928 163
rect 894 61 928 95
rect 988 61 1022 95
rect 1082 129 1116 163
rect 1082 61 1116 95
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 133 443 167 477
rect 133 375 167 409
rect 227 443 261 477
rect 321 357 355 391
rect 417 443 451 477
rect 511 443 545 477
rect 605 443 639 477
rect 605 375 639 409
rect 605 307 639 341
rect 699 443 733 477
rect 800 443 834 477
rect 894 375 928 409
rect 988 443 1022 477
rect 988 375 1022 409
rect 1083 443 1117 477
rect 1083 375 1117 409
<< poly >>
rect 85 497 121 523
rect 179 497 215 523
rect 273 497 309 523
rect 369 497 405 523
rect 557 497 593 523
rect 651 497 687 523
rect 752 497 788 523
rect 846 497 882 523
rect 940 497 976 523
rect 1034 497 1070 523
rect 85 282 121 297
rect 179 282 215 297
rect 273 282 309 297
rect 369 282 405 297
rect 557 282 593 297
rect 651 282 687 297
rect 752 282 788 297
rect 846 282 882 297
rect 940 282 976 297
rect 1034 282 1070 297
rect 83 265 123 282
rect 69 249 123 265
rect 69 215 79 249
rect 113 215 123 249
rect 69 199 123 215
rect 93 177 123 199
rect 177 265 217 282
rect 271 265 311 282
rect 177 249 311 265
rect 177 215 226 249
rect 260 215 311 249
rect 177 199 311 215
rect 177 177 207 199
rect 281 177 311 199
rect 367 265 407 282
rect 555 265 595 282
rect 649 265 689 282
rect 750 265 790 282
rect 367 249 421 265
rect 367 215 377 249
rect 411 215 421 249
rect 367 199 421 215
rect 495 249 689 265
rect 495 215 511 249
rect 545 215 689 249
rect 495 199 689 215
rect 736 249 790 265
rect 736 215 746 249
rect 780 215 790 249
rect 736 199 790 215
rect 367 177 397 199
rect 565 177 595 199
rect 659 177 689 199
rect 760 177 790 199
rect 844 265 884 282
rect 938 265 978 282
rect 844 249 978 265
rect 844 215 894 249
rect 928 215 978 249
rect 844 199 978 215
rect 844 177 874 199
rect 948 177 978 199
rect 1032 265 1072 282
rect 1032 249 1096 265
rect 1032 215 1042 249
rect 1076 215 1096 249
rect 1032 199 1096 215
rect 1032 177 1062 199
rect 93 21 123 47
rect 177 21 207 47
rect 281 21 311 47
rect 367 21 397 47
rect 565 21 595 47
rect 659 21 689 47
rect 760 21 790 47
rect 844 21 874 47
rect 948 21 978 47
rect 1032 21 1062 47
<< polycont >>
rect 79 215 113 249
rect 226 215 260 249
rect 377 215 411 249
rect 511 215 545 249
rect 746 215 780 249
rect 894 215 928 249
rect 1042 215 1076 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 30 477 80 527
rect 30 443 39 477
rect 73 443 80 477
rect 30 409 80 443
rect 30 375 39 409
rect 73 375 80 409
rect 30 359 80 375
rect 125 477 175 493
rect 125 443 133 477
rect 167 443 175 477
rect 125 409 175 443
rect 219 477 269 527
rect 219 443 227 477
rect 261 443 269 477
rect 219 427 269 443
rect 407 477 545 527
rect 407 443 417 477
rect 451 443 511 477
rect 407 427 545 443
rect 579 477 647 493
rect 579 443 605 477
rect 639 443 647 477
rect 125 375 133 409
rect 167 393 175 409
rect 579 409 647 443
rect 691 477 748 527
rect 691 443 699 477
rect 733 443 748 477
rect 691 425 748 443
rect 792 477 1030 493
rect 792 443 800 477
rect 834 459 988 477
rect 834 443 842 459
rect 792 425 842 443
rect 980 443 988 459
rect 1022 443 1030 477
rect 167 391 497 393
rect 167 375 321 391
rect 125 357 321 375
rect 355 357 497 391
rect 18 289 429 323
rect 18 249 135 289
rect 18 215 79 249
rect 113 215 135 249
rect 169 249 300 255
rect 169 215 226 249
rect 260 215 300 249
rect 353 249 429 289
rect 353 215 377 249
rect 411 215 429 249
rect 463 265 497 357
rect 579 375 605 409
rect 639 391 647 409
rect 886 409 936 425
rect 886 391 894 409
rect 639 375 894 391
rect 928 375 936 409
rect 579 357 936 375
rect 980 409 1030 443
rect 980 375 988 409
rect 1022 375 1030 409
rect 980 357 1030 375
rect 1083 477 1124 527
rect 1117 443 1124 477
rect 1083 409 1124 443
rect 1117 375 1124 409
rect 1083 359 1124 375
rect 579 341 693 357
rect 579 307 605 341
rect 639 307 693 341
rect 463 249 545 265
rect 463 215 511 249
rect 463 199 545 215
rect 579 215 693 307
rect 730 289 1092 323
rect 730 249 808 289
rect 730 215 746 249
rect 780 215 808 249
rect 852 249 980 255
rect 852 215 894 249
rect 928 215 980 249
rect 1026 249 1092 289
rect 1026 215 1042 249
rect 1076 215 1092 249
rect 463 181 497 199
rect 39 163 73 179
rect 39 95 73 129
rect 107 163 167 179
rect 107 129 133 163
rect 201 163 497 181
rect 201 129 227 163
rect 261 145 497 163
rect 579 163 655 215
rect 261 129 277 145
rect 579 129 605 163
rect 639 129 655 163
rect 699 163 1132 181
rect 733 147 894 163
rect 733 129 756 147
rect 107 95 167 129
rect 407 95 441 111
rect 107 61 133 95
rect 167 61 321 95
rect 355 61 371 95
rect 39 17 73 61
rect 407 17 441 61
rect 495 95 545 111
rect 699 95 756 129
rect 868 129 894 147
rect 928 145 1082 163
rect 928 129 944 145
rect 495 61 511 95
rect 545 61 699 95
rect 733 61 756 95
rect 495 51 756 61
rect 800 95 834 111
rect 800 17 834 61
rect 868 95 944 129
rect 1056 129 1082 145
rect 1116 129 1132 163
rect 868 61 894 95
rect 928 61 944 95
rect 868 51 944 61
rect 988 95 1022 111
rect 988 17 1022 61
rect 1056 95 1132 129
rect 1056 61 1082 95
rect 1116 61 1132 95
rect 1056 51 1132 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
flabel corelocali s 926 238 926 238 0 FreeSans 400 180 0 0 B2
port 4 nsew
flabel corelocali s 626 289 660 323 0 FreeSans 400 0 0 0 Y
port 9 nsew
flabel corelocali s 79 238 79 238 0 FreeSans 400 0 0 0 A1_N
port 1 nsew
flabel corelocali s 231 238 231 238 0 FreeSans 400 0 0 0 A2_N
port 2 nsew
flabel corelocali s 1039 221 1073 255 0 FreeSans 400 180 0 0 B1
port 3 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
rlabel comment s 0 0 0 0 4 o2bb2ai_2
<< properties >>
string FIXED_BBOX 0 0 1196 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 670776
string GDS_START 661926
<< end >>
