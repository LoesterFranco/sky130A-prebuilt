magic
tech sky130A
magscale 1 2
timestamp 1601050056
<< nwell >>
rect -38 356 2822 704
rect -38 332 1166 356
rect 1945 332 2822 356
rect 823 311 1166 332
<< pwell >>
rect 0 0 2784 49
<< scpmos >>
rect 83 464 119 592
rect 173 464 209 592
rect 251 464 287 592
rect 438 464 474 592
rect 516 464 552 592
rect 640 464 676 592
rect 924 347 960 547
rect 1041 347 1077 547
rect 1253 457 1289 541
rect 1345 457 1381 541
rect 1429 457 1465 541
rect 1525 457 1561 541
rect 1719 392 1755 592
rect 1906 392 1942 592
rect 2009 508 2045 592
rect 2091 508 2127 592
rect 2246 508 2282 592
rect 2336 508 2372 592
rect 2548 424 2584 592
rect 2664 368 2700 592
<< nmoslvt >>
rect 84 88 114 172
rect 294 81 324 165
rect 366 81 396 165
rect 508 81 538 165
rect 586 81 616 165
rect 674 81 704 165
rect 930 74 960 222
rect 1039 74 1069 222
rect 1243 131 1273 215
rect 1379 131 1409 215
rect 1453 131 1483 215
rect 1525 131 1555 215
rect 1655 144 1685 272
rect 1797 144 1827 272
rect 2043 74 2073 158
rect 2123 74 2153 158
rect 2235 74 2265 158
rect 2313 74 2343 158
rect 2554 74 2584 184
rect 2670 74 2700 222
<< ndiff >>
rect 27 147 84 172
rect 27 113 39 147
rect 73 113 84 147
rect 27 88 84 113
rect 114 147 185 172
rect 864 202 930 222
rect 864 168 881 202
rect 915 168 930 202
rect 114 113 139 147
rect 173 113 185 147
rect 114 88 185 113
rect 239 132 294 165
rect 239 98 249 132
rect 283 98 294 132
rect 239 81 294 98
rect 324 81 366 165
rect 396 153 508 165
rect 396 119 435 153
rect 469 119 508 153
rect 396 81 508 119
rect 538 81 586 165
rect 616 140 674 165
rect 616 106 628 140
rect 662 106 674 140
rect 616 81 674 106
rect 704 140 810 165
rect 704 106 747 140
rect 781 106 810 140
rect 704 81 810 106
rect 864 129 930 168
rect 864 95 881 129
rect 915 95 930 129
rect 864 74 930 95
rect 960 124 1039 222
rect 960 90 983 124
rect 1017 90 1039 124
rect 960 74 1039 90
rect 1069 202 1130 222
rect 1069 168 1088 202
rect 1122 168 1130 202
rect 1069 129 1130 168
rect 1069 95 1088 129
rect 1122 95 1130 129
rect 1069 74 1130 95
rect 1605 215 1655 272
rect 1190 190 1243 215
rect 1190 156 1198 190
rect 1232 156 1243 190
rect 1190 131 1243 156
rect 1273 203 1379 215
rect 1273 169 1334 203
rect 1368 169 1379 203
rect 1273 131 1379 169
rect 1409 131 1453 215
rect 1483 131 1525 215
rect 1555 144 1655 215
rect 1685 260 1797 272
rect 1685 226 1746 260
rect 1780 226 1797 260
rect 1685 190 1797 226
rect 1685 156 1746 190
rect 1780 156 1797 190
rect 1685 144 1797 156
rect 1827 179 1877 272
rect 1827 175 1885 179
rect 1827 168 1888 175
rect 1827 158 2016 168
rect 2599 210 2670 222
rect 2599 184 2625 210
rect 1827 156 2043 158
rect 1827 144 1882 156
rect 1555 131 1640 144
rect 1582 124 1640 131
rect 1582 90 1594 124
rect 1628 90 1640 124
rect 1582 78 1640 90
rect 1844 122 1882 144
rect 1916 140 2043 156
rect 1916 122 1998 140
rect 1844 106 1998 122
rect 2032 106 2043 140
rect 1844 74 2043 106
rect 2073 74 2123 158
rect 2153 120 2235 158
rect 2153 86 2176 120
rect 2210 86 2235 120
rect 2153 74 2235 86
rect 2265 74 2313 158
rect 2343 140 2443 158
rect 2343 106 2375 140
rect 2409 106 2443 140
rect 2343 74 2443 106
rect 2497 146 2554 184
rect 2497 112 2509 146
rect 2543 112 2554 146
rect 2497 74 2554 112
rect 2584 176 2625 184
rect 2659 176 2670 210
rect 2584 128 2670 176
rect 2584 94 2611 128
rect 2645 94 2670 128
rect 2584 74 2670 94
rect 2700 210 2757 222
rect 2700 176 2711 210
rect 2745 176 2757 210
rect 2700 120 2757 176
rect 2700 86 2711 120
rect 2745 86 2757 120
rect 2700 74 2757 86
rect 1844 62 2028 74
<< pdiff >>
rect 567 628 625 639
rect 567 594 579 628
rect 613 594 625 628
rect 567 592 625 594
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 510 83 546
rect 27 476 39 510
rect 73 476 83 510
rect 27 464 83 476
rect 119 578 173 592
rect 119 544 129 578
rect 163 544 173 578
rect 119 464 173 544
rect 209 464 251 592
rect 287 576 438 592
rect 287 542 297 576
rect 331 542 394 576
rect 428 542 438 576
rect 287 464 438 542
rect 474 464 516 592
rect 552 464 640 592
rect 676 580 732 592
rect 676 546 686 580
rect 720 546 732 580
rect 975 547 1026 560
rect 676 510 732 546
rect 676 476 686 510
rect 720 476 732 510
rect 676 464 732 476
rect 859 400 924 547
rect 859 366 878 400
rect 912 366 924 400
rect 859 347 924 366
rect 960 544 1041 547
rect 960 510 984 544
rect 1018 510 1041 544
rect 960 347 1041 510
rect 1077 400 1130 547
rect 1667 580 1719 592
rect 1667 546 1675 580
rect 1709 546 1719 580
rect 1197 522 1253 541
rect 1197 488 1208 522
rect 1242 488 1253 522
rect 1197 457 1253 488
rect 1289 522 1345 541
rect 1289 488 1300 522
rect 1334 488 1345 522
rect 1289 457 1345 488
rect 1381 457 1429 541
rect 1465 522 1525 541
rect 1465 488 1475 522
rect 1509 488 1525 522
rect 1465 457 1525 488
rect 1561 522 1613 541
rect 1561 488 1571 522
rect 1605 488 1613 522
rect 1561 457 1613 488
rect 1667 496 1719 546
rect 1667 462 1675 496
rect 1709 462 1719 496
rect 1077 366 1088 400
rect 1122 366 1130 400
rect 1077 347 1130 366
rect 1667 392 1719 462
rect 1755 580 1906 592
rect 1755 546 1775 580
rect 1809 546 1862 580
rect 1896 546 1906 580
rect 1755 512 1906 546
rect 1755 478 1775 512
rect 1809 478 1862 512
rect 1896 478 1906 512
rect 1755 444 1906 478
rect 1755 410 1775 444
rect 1809 410 1862 444
rect 1896 410 1906 444
rect 1755 392 1906 410
rect 1942 580 2009 592
rect 1942 546 1963 580
rect 1997 546 2009 580
rect 1942 512 2009 546
rect 1942 478 1952 512
rect 1986 508 2009 512
rect 2045 508 2091 592
rect 2127 580 2246 592
rect 2127 546 2164 580
rect 2198 546 2246 580
rect 2127 508 2246 546
rect 2282 567 2336 592
rect 2282 533 2292 567
rect 2326 533 2336 567
rect 2282 508 2336 533
rect 2372 578 2438 592
rect 2372 544 2392 578
rect 2426 544 2438 578
rect 2372 508 2438 544
rect 2492 580 2548 592
rect 2492 546 2504 580
rect 2538 546 2548 580
rect 1986 478 1994 508
rect 1942 444 1994 478
rect 1942 410 1952 444
rect 1986 410 1994 444
rect 1942 392 1994 410
rect 2492 470 2548 546
rect 2492 436 2504 470
rect 2538 436 2548 470
rect 2492 424 2548 436
rect 2584 580 2664 592
rect 2584 546 2611 580
rect 2645 546 2664 580
rect 2584 497 2664 546
rect 2584 463 2611 497
rect 2645 463 2664 497
rect 2584 424 2664 463
rect 2599 414 2664 424
rect 2599 380 2611 414
rect 2645 380 2664 414
rect 2599 368 2664 380
rect 2700 580 2757 592
rect 2700 546 2711 580
rect 2745 546 2757 580
rect 2700 497 2757 546
rect 2700 463 2711 497
rect 2745 463 2757 497
rect 2700 414 2757 463
rect 2700 380 2711 414
rect 2745 380 2757 414
rect 2700 368 2757 380
<< ndiffc >>
rect 39 113 73 147
rect 881 168 915 202
rect 139 113 173 147
rect 249 98 283 132
rect 435 119 469 153
rect 628 106 662 140
rect 747 106 781 140
rect 881 95 915 129
rect 983 90 1017 124
rect 1088 168 1122 202
rect 1088 95 1122 129
rect 1198 156 1232 190
rect 1334 169 1368 203
rect 1746 226 1780 260
rect 1746 156 1780 190
rect 1594 90 1628 124
rect 1882 122 1916 156
rect 1998 106 2032 140
rect 2176 86 2210 120
rect 2375 106 2409 140
rect 2509 112 2543 146
rect 2625 176 2659 210
rect 2611 94 2645 128
rect 2711 176 2745 210
rect 2711 86 2745 120
<< pdiffc >>
rect 579 594 613 628
rect 39 546 73 580
rect 39 476 73 510
rect 129 544 163 578
rect 297 542 331 576
rect 394 542 428 576
rect 686 546 720 580
rect 686 476 720 510
rect 878 366 912 400
rect 984 510 1018 544
rect 1675 546 1709 580
rect 1208 488 1242 522
rect 1300 488 1334 522
rect 1475 488 1509 522
rect 1571 488 1605 522
rect 1675 462 1709 496
rect 1088 366 1122 400
rect 1775 546 1809 580
rect 1862 546 1896 580
rect 1775 478 1809 512
rect 1862 478 1896 512
rect 1775 410 1809 444
rect 1862 410 1896 444
rect 1963 546 1997 580
rect 1952 478 1986 512
rect 2164 546 2198 580
rect 2292 533 2326 567
rect 2392 544 2426 578
rect 2504 546 2538 580
rect 1952 410 1986 444
rect 2504 436 2538 470
rect 2611 546 2645 580
rect 2611 463 2645 497
rect 2611 380 2645 414
rect 2711 546 2745 580
rect 2711 463 2745 497
rect 2711 380 2745 414
<< poly >>
rect 83 592 119 618
rect 173 592 209 618
rect 251 592 287 618
rect 438 592 474 618
rect 516 592 552 618
rect 640 615 1561 645
rect 640 592 676 615
rect 924 547 960 573
rect 1041 547 1077 573
rect 83 416 119 464
rect 173 416 209 464
rect 84 400 209 416
rect 84 366 123 400
rect 157 386 209 400
rect 251 422 287 464
rect 251 406 396 422
rect 251 392 346 406
rect 157 366 173 386
rect 84 332 173 366
rect 330 372 346 392
rect 380 372 396 406
rect 330 356 396 372
rect 84 298 123 332
rect 157 298 173 332
rect 84 282 173 298
rect 84 172 114 282
rect 258 237 324 253
rect 258 203 274 237
rect 308 203 324 237
rect 258 187 324 203
rect 294 165 324 187
rect 366 165 396 356
rect 438 377 474 464
rect 516 449 552 464
rect 640 449 676 464
rect 516 419 590 449
rect 640 419 704 449
rect 438 361 509 377
rect 438 327 459 361
rect 493 327 509 361
rect 438 311 509 327
rect 560 371 590 419
rect 674 405 704 419
rect 674 389 747 405
rect 560 355 626 371
rect 560 321 576 355
rect 610 321 626 355
rect 560 305 626 321
rect 674 355 697 389
rect 731 355 747 389
rect 674 321 747 355
rect 1253 541 1289 567
rect 1345 541 1381 567
rect 1429 541 1465 567
rect 1525 541 1561 615
rect 1719 592 1755 618
rect 1906 592 1942 618
rect 2009 592 2045 618
rect 2091 592 2127 618
rect 2246 592 2282 618
rect 2336 592 2372 618
rect 2548 592 2584 618
rect 2664 592 2700 618
rect 1253 442 1289 457
rect 1145 412 1289 442
rect 924 332 960 347
rect 1041 332 1077 347
rect 1145 332 1175 412
rect 444 241 538 257
rect 444 207 460 241
rect 494 207 538 241
rect 444 191 538 207
rect 508 165 538 191
rect 586 165 616 305
rect 674 287 697 321
rect 731 287 747 321
rect 674 271 747 287
rect 829 294 960 332
rect 674 165 704 271
rect 829 260 871 294
rect 905 260 960 294
rect 829 242 960 260
rect 1010 299 1175 332
rect 1345 393 1381 457
rect 1345 319 1375 393
rect 1429 360 1465 457
rect 1525 360 1561 457
rect 1719 360 1755 392
rect 1010 265 1026 299
rect 1060 265 1175 299
rect 1010 242 1175 265
rect 930 222 960 242
rect 1039 222 1069 242
rect 84 62 114 88
rect 294 55 324 81
rect 366 55 396 81
rect 508 55 538 81
rect 586 55 616 81
rect 674 55 704 81
rect 930 48 960 74
rect 1039 48 1069 74
rect 1145 51 1175 242
rect 1243 303 1375 319
rect 1243 269 1266 303
rect 1300 283 1375 303
rect 1417 344 1483 360
rect 1417 310 1433 344
rect 1467 310 1483 344
rect 1417 294 1483 310
rect 1300 269 1316 283
rect 1243 253 1316 269
rect 1243 215 1273 253
rect 1379 215 1409 241
rect 1453 215 1483 294
rect 1525 344 1603 360
rect 1525 310 1547 344
rect 1581 310 1603 344
rect 1525 294 1603 310
rect 1645 344 1755 360
rect 1645 310 1661 344
rect 1695 310 1755 344
rect 1645 294 1755 310
rect 1797 344 1864 360
rect 1797 310 1814 344
rect 1848 310 1864 344
rect 1797 294 1864 310
rect 1525 215 1555 294
rect 1655 272 1685 294
rect 1797 272 1827 294
rect 1906 256 1942 392
rect 2009 324 2045 508
rect 2091 476 2127 508
rect 2246 487 2282 508
rect 2087 460 2153 476
rect 2087 426 2103 460
rect 2137 426 2153 460
rect 2087 410 2153 426
rect 2009 308 2079 324
rect 2009 274 2029 308
rect 2063 274 2079 308
rect 2009 258 2079 274
rect 1899 240 1965 256
rect 1899 206 1915 240
rect 1949 216 1965 240
rect 1949 206 2073 216
rect 1899 186 2073 206
rect 2043 158 2073 186
rect 2123 158 2153 410
rect 2235 457 2282 487
rect 2235 308 2265 457
rect 2336 409 2372 508
rect 2548 409 2584 424
rect 2336 379 2584 409
rect 2336 314 2366 379
rect 2664 337 2700 368
rect 2496 321 2700 337
rect 2199 292 2265 308
rect 2199 258 2215 292
rect 2249 258 2265 292
rect 2199 242 2265 258
rect 2235 158 2265 242
rect 2313 298 2379 314
rect 2313 264 2329 298
rect 2363 264 2379 298
rect 2496 287 2512 321
rect 2546 287 2700 321
rect 2496 271 2700 287
rect 2313 230 2379 264
rect 2313 196 2329 230
rect 2363 229 2379 230
rect 2363 199 2584 229
rect 2670 222 2700 271
rect 2363 196 2379 199
rect 2313 180 2379 196
rect 2554 184 2584 199
rect 2313 158 2343 180
rect 1243 93 1273 131
rect 1379 51 1409 131
rect 1453 93 1483 131
rect 1525 93 1555 131
rect 1655 118 1685 144
rect 1797 51 1827 144
rect 1145 21 1827 51
rect 2043 48 2073 74
rect 2123 48 2153 74
rect 2235 48 2265 74
rect 2313 48 2343 74
rect 2554 48 2584 74
rect 2670 48 2700 74
<< polycont >>
rect 123 366 157 400
rect 346 372 380 406
rect 123 298 157 332
rect 274 203 308 237
rect 459 327 493 361
rect 576 321 610 355
rect 697 355 731 389
rect 460 207 494 241
rect 697 287 731 321
rect 871 260 905 294
rect 1026 265 1060 299
rect 1266 269 1300 303
rect 1433 310 1467 344
rect 1547 310 1581 344
rect 1661 310 1695 344
rect 1814 310 1848 344
rect 2103 426 2137 460
rect 2029 274 2063 308
rect 1915 206 1949 240
rect 2215 258 2249 292
rect 2329 264 2363 298
rect 2512 287 2546 321
rect 2329 196 2363 230
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 23 580 73 596
rect 23 546 39 580
rect 23 510 73 546
rect 113 578 179 649
rect 563 628 629 649
rect 563 594 579 628
rect 613 594 629 628
rect 113 544 129 578
rect 163 544 179 578
rect 113 526 179 544
rect 281 576 444 592
rect 281 542 297 576
rect 331 542 394 576
rect 428 560 444 576
rect 686 580 736 596
rect 428 546 686 560
rect 720 546 736 580
rect 428 542 736 546
rect 281 526 736 542
rect 23 476 39 510
rect 686 520 736 526
rect 968 544 1034 649
rect 686 510 903 520
rect 968 510 984 544
rect 1018 510 1034 544
rect 1193 522 1247 541
rect 73 476 509 492
rect 23 458 509 476
rect 720 476 903 510
rect 1193 488 1208 522
rect 1242 488 1247 522
rect 1193 476 1247 488
rect 686 460 1247 476
rect 23 248 73 458
rect 107 400 173 416
rect 107 366 123 400
rect 157 366 173 400
rect 107 332 173 366
rect 217 406 396 424
rect 217 372 346 406
rect 380 372 396 406
rect 217 356 396 372
rect 443 361 509 458
rect 781 436 1247 460
rect 1283 522 1370 541
rect 1283 488 1300 522
rect 1334 488 1370 522
rect 1283 455 1370 488
rect 1459 522 1509 649
rect 1659 580 1725 649
rect 1659 546 1675 580
rect 1709 546 1725 580
rect 1459 488 1475 522
rect 1459 472 1509 488
rect 1557 522 1625 541
rect 1557 488 1571 522
rect 1605 488 1625 522
rect 107 298 123 332
rect 157 316 173 332
rect 443 327 459 361
rect 493 327 509 361
rect 443 316 509 327
rect 560 355 647 430
rect 560 321 576 355
rect 610 321 647 355
rect 157 298 409 316
rect 560 305 647 321
rect 681 389 747 405
rect 681 355 697 389
rect 731 355 747 389
rect 681 350 747 355
rect 681 321 703 350
rect 107 282 409 298
rect 681 287 697 321
rect 737 316 747 350
rect 731 287 747 316
rect 23 237 324 248
rect 23 210 274 237
rect 23 147 89 210
rect 258 203 274 210
rect 308 203 324 237
rect 258 187 324 203
rect 375 241 510 282
rect 681 271 747 287
rect 375 207 460 241
rect 494 207 510 241
rect 781 237 815 436
rect 862 400 1038 402
rect 862 366 878 400
rect 912 366 1038 400
rect 862 364 1038 366
rect 988 315 1038 364
rect 1072 400 1147 402
rect 1072 366 1088 400
rect 1122 366 1147 400
rect 1072 349 1147 366
rect 855 294 935 310
rect 855 260 871 294
rect 905 260 935 294
rect 855 242 935 260
rect 988 299 1060 315
rect 988 265 1026 299
rect 988 244 1060 265
rect 375 191 510 207
rect 544 192 815 237
rect 988 202 1054 244
rect 1094 218 1147 349
rect 23 113 39 147
rect 73 113 89 147
rect 23 84 89 113
rect 123 147 189 176
rect 544 153 578 192
rect 865 168 881 202
rect 915 168 1054 202
rect 865 162 1054 168
rect 1088 202 1147 218
rect 1122 168 1147 202
rect 123 113 139 147
rect 173 113 189 147
rect 123 17 189 113
rect 233 132 299 153
rect 233 98 249 132
rect 283 98 299 132
rect 391 119 435 153
rect 469 119 578 153
rect 612 140 678 156
rect 233 85 299 98
rect 612 106 628 140
rect 662 106 678 140
rect 612 85 678 106
rect 233 51 678 85
rect 731 140 797 156
rect 731 106 747 140
rect 781 106 797 140
rect 731 17 797 106
rect 865 129 932 162
rect 865 95 881 129
rect 915 95 932 129
rect 1088 129 1147 168
rect 865 79 932 95
rect 967 124 1033 128
rect 967 90 983 124
rect 1017 90 1033 124
rect 967 17 1033 90
rect 1122 95 1147 129
rect 1182 368 1247 436
rect 1334 438 1370 455
rect 1557 438 1625 488
rect 1659 496 1725 546
rect 1659 462 1675 496
rect 1709 462 1725 496
rect 1759 580 1899 596
rect 1759 546 1775 580
rect 1809 546 1862 580
rect 1896 546 1899 580
rect 1759 512 1899 546
rect 1759 478 1775 512
rect 1809 478 1862 512
rect 1896 478 1899 512
rect 1334 428 1625 438
rect 1759 444 1899 478
rect 1759 433 1775 444
rect 1334 394 1698 428
rect 1182 190 1232 368
rect 1182 156 1198 190
rect 1182 127 1232 156
rect 1266 303 1300 334
rect 1088 93 1147 95
rect 1266 93 1300 269
rect 1334 215 1370 394
rect 1415 344 1483 360
rect 1415 310 1433 344
rect 1467 310 1483 344
rect 1415 294 1483 310
rect 1531 350 1607 360
rect 1531 344 1567 350
rect 1531 310 1547 344
rect 1601 316 1607 350
rect 1581 310 1607 316
rect 1531 294 1607 310
rect 1645 344 1698 394
rect 1645 310 1661 344
rect 1695 310 1698 344
rect 1645 294 1698 310
rect 1746 410 1775 433
rect 1809 410 1862 444
rect 1896 410 1899 444
rect 1746 394 1899 410
rect 1947 580 2013 596
rect 1947 546 1963 580
rect 1997 546 2013 580
rect 1947 512 2013 546
rect 2121 580 2242 649
rect 2121 546 2164 580
rect 2198 546 2242 580
rect 2121 530 2242 546
rect 2276 567 2342 596
rect 2276 533 2292 567
rect 2326 533 2342 567
rect 1947 478 1952 512
rect 1986 478 2013 512
rect 2276 492 2342 533
rect 2376 578 2442 649
rect 2376 544 2392 578
rect 2426 544 2442 578
rect 2376 526 2442 544
rect 2488 580 2559 596
rect 2488 546 2504 580
rect 2538 546 2559 580
rect 1947 444 2013 478
rect 1947 410 1952 444
rect 1986 410 2013 444
rect 2087 460 2447 492
rect 2087 426 2103 460
rect 2137 458 2447 460
rect 2087 410 2137 426
rect 1447 260 1483 294
rect 1746 260 1780 394
rect 1947 376 2013 410
rect 2171 390 2379 424
rect 2171 376 2205 390
rect 1814 344 1870 360
rect 1848 310 1870 344
rect 1947 342 2205 376
rect 2239 350 2279 356
rect 1814 308 1870 310
rect 2273 316 2279 350
rect 2239 308 2279 316
rect 1814 274 2029 308
rect 2063 274 2079 308
rect 1447 226 1746 260
rect 2013 258 2079 274
rect 2199 292 2279 308
rect 2199 258 2215 292
rect 2249 258 2279 292
rect 2199 242 2279 258
rect 2313 298 2379 390
rect 2313 264 2329 298
rect 2363 264 2379 298
rect 1334 203 1384 215
rect 1368 169 1384 203
rect 1334 127 1384 169
rect 1418 158 1712 192
rect 1418 93 1452 158
rect 1088 51 1452 93
rect 1578 90 1594 124
rect 1628 90 1644 124
rect 1578 17 1644 90
rect 1678 106 1712 158
rect 1746 190 1780 226
rect 1746 140 1780 156
rect 1814 206 1915 240
rect 1949 206 1965 240
rect 2313 230 2379 264
rect 2313 208 2329 230
rect 1814 106 1848 206
rect 2061 196 2329 208
rect 2363 196 2379 230
rect 2061 174 2379 196
rect 2061 172 2095 174
rect 1882 156 2095 172
rect 1916 140 2095 156
rect 2413 140 2447 458
rect 1916 122 1998 140
rect 1882 106 1998 122
rect 2032 106 2095 140
rect 2146 120 2240 136
rect 1678 72 1848 106
rect 2146 86 2176 120
rect 2210 86 2240 120
rect 2338 106 2375 140
rect 2409 106 2447 140
rect 2338 90 2447 106
rect 2488 470 2559 546
rect 2488 436 2504 470
rect 2538 436 2559 470
rect 2488 337 2559 436
rect 2595 580 2661 649
rect 2595 546 2611 580
rect 2645 546 2661 580
rect 2595 497 2661 546
rect 2595 463 2611 497
rect 2645 463 2661 497
rect 2595 414 2661 463
rect 2595 380 2611 414
rect 2645 380 2661 414
rect 2595 364 2661 380
rect 2695 580 2761 596
rect 2695 546 2711 580
rect 2745 546 2761 580
rect 2695 497 2761 546
rect 2695 463 2711 497
rect 2745 463 2761 497
rect 2695 414 2761 463
rect 2695 380 2711 414
rect 2745 380 2761 414
rect 2488 321 2562 337
rect 2488 287 2512 321
rect 2546 287 2562 321
rect 2488 271 2562 287
rect 2488 146 2559 271
rect 2488 112 2509 146
rect 2543 112 2559 146
rect 2146 17 2240 86
rect 2488 70 2559 112
rect 2595 210 2661 226
rect 2595 176 2625 210
rect 2659 176 2661 210
rect 2595 128 2661 176
rect 2595 94 2611 128
rect 2645 94 2661 128
rect 2595 17 2661 94
rect 2695 210 2761 380
rect 2695 176 2711 210
rect 2745 176 2761 210
rect 2695 120 2761 176
rect 2695 86 2711 120
rect 2745 86 2761 120
rect 2695 70 2761 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 703 321 737 350
rect 703 316 731 321
rect 731 316 737 321
rect 1567 344 1601 350
rect 1567 316 1581 344
rect 1581 316 1601 344
rect 2239 316 2273 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
<< metal1 >>
rect 0 683 2784 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 0 617 2784 649
rect 691 350 749 356
rect 691 316 703 350
rect 737 347 749 350
rect 1555 350 1613 356
rect 1555 347 1567 350
rect 737 319 1567 347
rect 737 316 749 319
rect 691 310 749 316
rect 1555 316 1567 319
rect 1601 347 1613 350
rect 2227 350 2285 356
rect 2227 347 2239 350
rect 1601 319 2239 347
rect 1601 316 1613 319
rect 1555 310 1613 316
rect 2227 316 2239 319
rect 2273 316 2285 350
rect 2227 310 2285 316
rect 0 17 2784 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
rect 0 -49 2784 -17
<< labels >>
flabel pwell s 0 0 2784 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 0 617 2784 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel comment s 1150 630 1150 630 0 FreeSans 300 0 0 0 no_jumper_check
flabel comment s 1471 36 1471 36 0 FreeSans 300 0 0 0 no_jumper_check
rlabel comment s 0 0 0 0 4 sdfrtn_1
flabel metal1 s 703 316 737 350 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew
flabel metal1 s 0 617 2784 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 2784 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 2719 94 2753 128 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2719 168 2753 202 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2719 242 2753 276 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2719 316 2753 350 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2719 390 2753 424 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2719 464 2753 498 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2719 538 2753 572 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 895 242 929 276 0 FreeSans 340 0 0 0 CLK_N
port 1 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 SCD
port 4 nsew
flabel corelocali s 607 390 641 424 0 FreeSans 340 0 0 0 SCD
port 4 nsew
flabel corelocali s 415 242 449 276 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 223 390 257 424 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 319 390 353 424 0 FreeSans 340 0 0 0 D
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 2784 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 252634
string GDS_START 231904
<< end >>
