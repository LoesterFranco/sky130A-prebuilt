magic
tech sky130A
magscale 1 2
timestamp 1601050047
<< nwell >>
rect -38 332 806 704
<< pwell >>
rect 0 0 768 49
<< scpmos >>
rect 128 392 158 592
rect 212 392 242 592
rect 422 368 452 592
rect 536 368 566 592
rect 636 368 666 592
<< nmoslvt >>
rect 164 125 194 235
rect 323 125 353 235
rect 425 87 455 235
rect 503 87 533 235
rect 617 87 647 235
<< ndiff >>
rect 43 182 164 235
rect 43 148 51 182
rect 85 148 119 182
rect 153 148 164 182
rect 43 125 164 148
rect 194 192 323 235
rect 194 158 205 192
rect 239 158 278 192
rect 312 158 323 192
rect 194 125 323 158
rect 353 223 425 235
rect 353 189 380 223
rect 414 189 425 223
rect 353 133 425 189
rect 353 125 380 133
rect 368 99 380 125
rect 414 99 425 133
rect 368 87 425 99
rect 455 87 503 235
rect 533 214 617 235
rect 533 180 544 214
rect 578 180 617 214
rect 533 133 617 180
rect 533 99 544 133
rect 578 99 617 133
rect 533 87 617 99
rect 647 133 728 235
rect 647 99 658 133
rect 692 99 728 133
rect 647 87 728 99
<< pdiff >>
rect 69 580 128 592
rect 69 546 81 580
rect 115 546 128 580
rect 69 509 128 546
rect 69 475 81 509
rect 115 475 128 509
rect 69 438 128 475
rect 69 404 81 438
rect 115 404 128 438
rect 69 392 128 404
rect 158 392 212 592
rect 242 580 301 592
rect 242 546 255 580
rect 289 546 301 580
rect 242 510 301 546
rect 242 476 255 510
rect 289 476 301 510
rect 242 440 301 476
rect 242 406 255 440
rect 289 406 301 440
rect 242 392 301 406
rect 355 580 422 592
rect 355 546 367 580
rect 401 546 422 580
rect 355 508 422 546
rect 355 474 367 508
rect 401 474 422 508
rect 355 368 422 474
rect 452 580 536 592
rect 452 546 478 580
rect 512 546 536 580
rect 452 368 536 546
rect 566 580 636 592
rect 566 546 589 580
rect 623 546 636 580
rect 566 508 636 546
rect 566 474 589 508
rect 623 474 636 508
rect 566 368 636 474
rect 666 580 735 592
rect 666 546 689 580
rect 723 546 735 580
rect 666 497 735 546
rect 666 463 689 497
rect 723 463 735 497
rect 666 414 735 463
rect 666 380 689 414
rect 723 380 735 414
rect 666 368 735 380
<< ndiffc >>
rect 51 148 85 182
rect 119 148 153 182
rect 205 158 239 192
rect 278 158 312 192
rect 380 189 414 223
rect 380 99 414 133
rect 544 180 578 214
rect 544 99 578 133
rect 658 99 692 133
<< pdiffc >>
rect 81 546 115 580
rect 81 475 115 509
rect 81 404 115 438
rect 255 546 289 580
rect 255 476 289 510
rect 255 406 289 440
rect 367 546 401 580
rect 367 474 401 508
rect 478 546 512 580
rect 589 546 623 580
rect 589 474 623 508
rect 689 546 723 580
rect 689 463 723 497
rect 689 380 723 414
<< poly >>
rect 128 592 158 618
rect 212 592 242 618
rect 422 592 452 618
rect 536 592 566 618
rect 636 592 666 618
rect 128 377 158 392
rect 212 377 242 392
rect 125 335 161 377
rect 209 369 245 377
rect 209 339 287 369
rect 422 353 452 368
rect 536 353 566 368
rect 636 353 666 368
rect 125 323 155 335
rect 21 307 155 323
rect 21 273 37 307
rect 71 273 105 307
rect 139 287 155 307
rect 257 323 353 339
rect 257 289 273 323
rect 307 289 353 323
rect 139 273 194 287
rect 257 273 353 289
rect 21 257 194 273
rect 164 235 194 257
rect 323 235 353 273
rect 419 250 455 353
rect 533 336 569 353
rect 425 235 455 250
rect 503 320 569 336
rect 633 330 669 353
rect 503 286 519 320
rect 553 286 569 320
rect 503 270 569 286
rect 617 314 683 330
rect 617 280 633 314
rect 667 280 683 314
rect 503 235 533 270
rect 617 264 683 280
rect 617 235 647 264
rect 164 51 194 125
rect 323 99 353 125
rect 425 51 455 87
rect 503 61 533 87
rect 617 61 647 87
rect 164 21 455 51
<< polycont >>
rect 37 273 71 307
rect 105 273 139 307
rect 273 289 307 323
rect 519 286 553 320
rect 633 280 667 314
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 65 580 131 649
rect 65 546 81 580
rect 115 546 131 580
rect 65 509 131 546
rect 65 475 81 509
rect 115 475 131 509
rect 65 438 131 475
rect 65 404 81 438
rect 115 404 131 438
rect 65 388 131 404
rect 189 580 305 596
rect 189 546 255 580
rect 289 546 305 580
rect 189 510 305 546
rect 189 476 255 510
rect 289 476 305 510
rect 189 440 305 476
rect 351 580 417 596
rect 351 546 367 580
rect 401 546 417 580
rect 351 508 417 546
rect 451 580 539 649
rect 451 546 478 580
rect 512 546 539 580
rect 451 530 539 546
rect 573 580 639 596
rect 573 546 589 580
rect 623 546 639 580
rect 351 474 367 508
rect 401 492 417 508
rect 573 508 639 546
rect 573 492 589 508
rect 401 474 589 492
rect 623 474 639 508
rect 351 458 639 474
rect 673 580 751 596
rect 673 546 689 580
rect 723 546 751 580
rect 673 497 751 546
rect 673 463 689 497
rect 723 463 751 497
rect 189 406 255 440
rect 289 424 305 440
rect 289 406 639 424
rect 189 390 639 406
rect 21 307 155 323
rect 21 273 37 307
rect 71 273 105 307
rect 139 273 155 307
rect 21 236 155 273
rect 189 208 223 390
rect 503 339 569 356
rect 257 323 569 339
rect 257 289 273 323
rect 307 320 569 323
rect 307 289 519 320
rect 257 286 519 289
rect 553 286 569 320
rect 257 273 569 286
rect 503 270 569 273
rect 605 330 639 390
rect 673 414 751 463
rect 673 380 689 414
rect 723 380 751 414
rect 673 364 751 380
rect 605 314 683 330
rect 605 280 633 314
rect 667 280 683 314
rect 605 264 683 280
rect 364 223 430 239
rect 717 230 751 364
rect 35 182 155 198
rect 35 148 51 182
rect 85 148 119 182
rect 153 148 155 182
rect 35 17 155 148
rect 189 192 328 208
rect 189 158 205 192
rect 239 158 278 192
rect 312 158 328 192
rect 189 142 328 158
rect 364 189 380 223
rect 414 189 430 223
rect 364 133 430 189
rect 364 99 380 133
rect 414 99 430 133
rect 364 17 430 99
rect 505 214 751 230
rect 505 180 544 214
rect 578 196 751 214
rect 578 180 594 196
rect 505 133 594 180
rect 505 99 544 133
rect 578 99 594 133
rect 505 83 594 99
rect 642 133 708 149
rect 642 99 658 133
rect 692 99 708 133
rect 642 17 708 99
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel comment s 0 0 0 0 4 xor2_1
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 511 94 545 128 0 FreeSans 340 0 0 0 X
port 7 nsew
flabel corelocali s 511 168 545 202 0 FreeSans 340 0 0 0 X
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 768 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 550900
string GDS_START 544608
<< end >>
