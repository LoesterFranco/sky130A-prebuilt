magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 388 2822 704
rect -38 332 833 388
rect 1105 332 2822 388
rect 1105 321 2490 332
rect 1897 306 2490 321
<< pwell >>
rect 0 0 2784 49
<< scnmos >>
rect 83 112 113 260
rect 201 132 231 260
rect 410 84 440 232
rect 614 104 644 232
rect 951 167 981 295
rect 1052 125 1082 253
rect 1138 125 1168 253
rect 1238 107 1268 235
rect 1508 74 1538 222
rect 1738 94 1768 222
rect 1888 94 1918 222
rect 2006 94 2036 222
rect 2240 94 2270 222
rect 2342 74 2372 222
rect 2564 74 2594 202
rect 2670 74 2700 202
<< pmoshvt >>
rect 86 368 116 592
rect 222 380 252 580
rect 543 368 573 592
rect 672 377 702 577
rect 814 424 844 592
rect 1026 424 1056 592
rect 1239 373 1269 541
rect 1390 373 1420 541
rect 1497 357 1527 581
rect 1719 374 1749 542
rect 1819 374 1849 542
rect 2154 368 2184 536
rect 2244 368 2274 536
rect 2345 368 2375 592
rect 2567 392 2597 592
rect 2667 392 2697 592
<< ndiff >>
rect 27 248 83 260
rect 27 214 38 248
rect 72 214 83 248
rect 27 158 83 214
rect 27 124 38 158
rect 72 124 83 158
rect 27 112 83 124
rect 113 132 201 260
rect 231 248 294 260
rect 231 214 245 248
rect 279 214 294 248
rect 231 132 294 214
rect 113 112 186 132
rect 128 78 140 112
rect 174 78 186 112
rect 128 66 186 78
rect 659 232 717 233
rect 354 130 410 232
rect 354 96 365 130
rect 399 96 410 130
rect 354 84 410 96
rect 440 130 614 232
rect 440 96 451 130
rect 485 104 614 130
rect 644 221 717 232
rect 644 187 671 221
rect 705 187 717 221
rect 644 104 717 187
rect 901 167 951 295
rect 981 269 1037 295
rect 981 235 992 269
rect 1026 253 1037 269
rect 1026 235 1052 253
rect 981 167 1052 235
rect 901 113 931 167
rect 485 96 497 104
rect 440 84 497 96
rect 879 101 936 113
rect 879 67 891 101
rect 925 67 936 101
rect 879 55 936 67
rect 1002 125 1052 167
rect 1082 223 1138 253
rect 1082 189 1093 223
rect 1127 189 1138 223
rect 1082 125 1138 189
rect 1168 235 1218 253
rect 1168 172 1238 235
rect 1168 138 1193 172
rect 1227 138 1238 172
rect 1168 125 1238 138
rect 1188 107 1238 125
rect 1268 192 1325 235
rect 1268 158 1279 192
rect 1313 158 1325 192
rect 1268 107 1325 158
rect 1665 226 1723 238
rect 1451 210 1508 222
rect 1451 176 1463 210
rect 1497 176 1508 210
rect 1451 120 1508 176
rect 1451 86 1463 120
rect 1497 86 1508 120
rect 1451 74 1508 86
rect 1538 90 1611 222
rect 1665 192 1677 226
rect 1711 222 1723 226
rect 1933 226 1991 238
rect 1933 222 1945 226
rect 1711 192 1738 222
rect 1665 94 1738 192
rect 1768 94 1888 222
rect 1918 192 1945 222
rect 1979 222 1991 226
rect 1979 192 2006 222
rect 1918 94 2006 192
rect 2036 181 2240 222
rect 2036 147 2113 181
rect 2147 147 2240 181
rect 2036 94 2240 147
rect 2270 210 2342 222
rect 2270 176 2297 210
rect 2331 176 2342 210
rect 2270 120 2342 176
rect 2270 94 2297 120
rect 1538 74 1565 90
rect 1553 56 1565 74
rect 1599 56 1611 90
rect 1783 90 1873 94
rect 1553 44 1611 56
rect 1783 56 1811 90
rect 1845 56 1873 90
rect 2285 86 2297 94
rect 2331 86 2342 120
rect 2285 74 2342 86
rect 2372 108 2445 222
rect 2372 74 2399 108
rect 2433 74 2445 108
rect 2499 190 2564 202
rect 2499 156 2511 190
rect 2545 156 2564 190
rect 2499 120 2564 156
rect 2499 86 2511 120
rect 2545 86 2564 120
rect 2499 74 2564 86
rect 2594 190 2670 202
rect 2594 156 2611 190
rect 2645 156 2670 190
rect 2594 120 2670 156
rect 2594 86 2611 120
rect 2645 86 2670 120
rect 2594 74 2670 86
rect 2700 190 2757 202
rect 2700 156 2711 190
rect 2745 156 2757 190
rect 2700 120 2757 156
rect 2700 86 2711 120
rect 2745 86 2757 120
rect 2700 74 2757 86
rect 1783 44 1873 56
rect 2387 62 2445 74
<< pdiff >>
rect 591 627 654 639
rect 467 609 525 621
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 497 86 546
rect 27 463 39 497
rect 73 463 86 497
rect 27 414 86 463
rect 27 380 39 414
rect 73 380 86 414
rect 27 368 86 380
rect 116 580 178 592
rect 116 546 129 580
rect 163 546 222 580
rect 116 508 222 546
rect 116 474 129 508
rect 163 474 222 508
rect 116 380 222 474
rect 252 531 311 580
rect 252 497 265 531
rect 299 497 311 531
rect 252 440 311 497
rect 467 575 479 609
rect 513 592 525 609
rect 591 593 605 627
rect 639 593 654 627
rect 591 592 654 593
rect 513 575 543 592
rect 252 406 265 440
rect 299 406 311 440
rect 252 380 311 406
rect 116 368 169 380
rect 467 368 543 575
rect 573 577 654 592
rect 761 577 814 592
rect 573 377 672 577
rect 702 424 814 577
rect 844 539 1026 592
rect 844 505 857 539
rect 891 505 1026 539
rect 844 468 1026 505
rect 844 434 857 468
rect 891 434 1026 468
rect 844 424 1026 434
rect 1056 580 1221 592
rect 1056 546 1069 580
rect 1103 546 1175 580
rect 1209 546 1221 580
rect 1056 541 1221 546
rect 1438 569 1497 581
rect 1438 541 1450 569
rect 1056 424 1239 541
rect 702 423 796 424
rect 702 389 732 423
rect 766 389 796 423
rect 702 377 796 389
rect 573 368 626 377
rect 1186 373 1239 424
rect 1269 512 1390 541
rect 1269 478 1282 512
rect 1316 478 1390 512
rect 1269 373 1390 478
rect 1420 535 1450 541
rect 1484 535 1497 569
rect 1420 498 1497 535
rect 1420 464 1450 498
rect 1484 464 1497 498
rect 1420 427 1497 464
rect 1420 393 1450 427
rect 1484 393 1497 427
rect 1420 373 1497 393
rect 1444 357 1497 373
rect 1527 569 1596 581
rect 1527 535 1550 569
rect 1584 535 1596 569
rect 1527 486 1596 535
rect 1527 452 1550 486
rect 1584 452 1596 486
rect 1527 403 1596 452
rect 1527 369 1550 403
rect 1584 369 1596 403
rect 1527 357 1596 369
rect 1660 530 1719 542
rect 1660 496 1672 530
rect 1706 496 1719 530
rect 1660 426 1719 496
rect 1660 392 1672 426
rect 1706 392 1719 426
rect 1660 374 1719 392
rect 1749 531 1819 542
rect 1749 497 1772 531
rect 1806 497 1819 531
rect 1749 432 1819 497
rect 1749 398 1772 432
rect 1806 398 1819 432
rect 1749 374 1819 398
rect 1849 536 2136 542
rect 2393 608 2454 620
rect 2393 592 2406 608
rect 2292 536 2345 592
rect 1849 479 2154 536
rect 1849 445 1879 479
rect 1913 445 1962 479
rect 1996 445 2045 479
rect 2079 445 2154 479
rect 1849 411 2154 445
rect 1849 377 1879 411
rect 1913 377 1962 411
rect 1996 377 2045 411
rect 2079 377 2154 411
rect 1849 374 2154 377
rect 1867 368 2154 374
rect 2184 528 2244 536
rect 2184 494 2197 528
rect 2231 494 2244 528
rect 2184 413 2244 494
rect 2184 379 2197 413
rect 2231 379 2244 413
rect 2184 368 2244 379
rect 2274 528 2345 536
rect 2274 494 2292 528
rect 2326 494 2345 528
rect 2274 415 2345 494
rect 2274 381 2292 415
rect 2326 381 2345 415
rect 2274 368 2345 381
rect 2375 574 2406 592
rect 2440 574 2454 608
rect 2375 540 2454 574
rect 2375 506 2406 540
rect 2440 506 2454 540
rect 2375 472 2454 506
rect 2375 438 2406 472
rect 2440 438 2454 472
rect 2375 368 2454 438
rect 2508 580 2567 592
rect 2508 546 2520 580
rect 2554 546 2567 580
rect 2508 512 2567 546
rect 2508 478 2520 512
rect 2554 478 2567 512
rect 2508 444 2567 478
rect 2508 410 2520 444
rect 2554 410 2567 444
rect 2508 392 2567 410
rect 2597 580 2667 592
rect 2597 546 2610 580
rect 2644 546 2667 580
rect 2597 512 2667 546
rect 2597 478 2610 512
rect 2644 478 2667 512
rect 2597 444 2667 478
rect 2597 410 2610 444
rect 2644 410 2667 444
rect 2597 392 2667 410
rect 2697 580 2757 592
rect 2697 546 2710 580
rect 2744 546 2757 580
rect 2697 512 2757 546
rect 2697 478 2710 512
rect 2744 478 2757 512
rect 2697 444 2757 478
rect 2697 410 2710 444
rect 2744 410 2757 444
rect 2697 392 2757 410
<< ndiffc >>
rect 38 214 72 248
rect 38 124 72 158
rect 245 214 279 248
rect 140 78 174 112
rect 365 96 399 130
rect 451 96 485 130
rect 671 187 705 221
rect 992 235 1026 269
rect 891 67 925 101
rect 1093 189 1127 223
rect 1193 138 1227 172
rect 1279 158 1313 192
rect 1463 176 1497 210
rect 1463 86 1497 120
rect 1677 192 1711 226
rect 1945 192 1979 226
rect 2113 147 2147 181
rect 2297 176 2331 210
rect 1565 56 1599 90
rect 1811 56 1845 90
rect 2297 86 2331 120
rect 2399 74 2433 108
rect 2511 156 2545 190
rect 2511 86 2545 120
rect 2611 156 2645 190
rect 2611 86 2645 120
rect 2711 156 2745 190
rect 2711 86 2745 120
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 129 546 163 580
rect 129 474 163 508
rect 265 497 299 531
rect 479 575 513 609
rect 605 593 639 627
rect 265 406 299 440
rect 857 505 891 539
rect 857 434 891 468
rect 1069 546 1103 580
rect 1175 546 1209 580
rect 732 389 766 423
rect 1282 478 1316 512
rect 1450 535 1484 569
rect 1450 464 1484 498
rect 1450 393 1484 427
rect 1550 535 1584 569
rect 1550 452 1584 486
rect 1550 369 1584 403
rect 1672 496 1706 530
rect 1672 392 1706 426
rect 1772 497 1806 531
rect 1772 398 1806 432
rect 1879 445 1913 479
rect 1962 445 1996 479
rect 2045 445 2079 479
rect 1879 377 1913 411
rect 1962 377 1996 411
rect 2045 377 2079 411
rect 2197 494 2231 528
rect 2197 379 2231 413
rect 2292 494 2326 528
rect 2292 381 2326 415
rect 2406 574 2440 608
rect 2406 506 2440 540
rect 2406 438 2440 472
rect 2520 546 2554 580
rect 2520 478 2554 512
rect 2520 410 2554 444
rect 2610 546 2644 580
rect 2610 478 2644 512
rect 2610 410 2644 444
rect 2710 546 2744 580
rect 2710 478 2744 512
rect 2710 410 2744 444
<< poly >>
rect 86 592 116 618
rect 222 580 252 606
rect 543 592 573 618
rect 332 457 435 473
rect 332 423 385 457
rect 419 423 435 457
rect 332 389 435 423
rect 86 353 116 368
rect 222 365 252 380
rect 83 275 119 353
rect 219 348 255 365
rect 332 355 385 389
rect 419 355 435 389
rect 672 577 702 603
rect 814 592 844 618
rect 1023 615 1423 645
rect 1023 607 1059 615
rect 1026 592 1056 607
rect 1239 541 1269 567
rect 1387 556 1423 615
rect 1611 615 2277 645
rect 1497 581 1527 607
rect 1390 541 1420 556
rect 814 409 844 424
rect 1026 409 1056 424
rect 811 379 946 409
rect 1023 379 1082 409
rect 201 332 267 348
rect 201 298 217 332
rect 251 298 267 332
rect 201 282 267 298
rect 332 339 435 355
rect 543 353 573 368
rect 672 362 702 377
rect 540 350 576 353
rect 83 260 113 275
rect 201 260 231 282
rect 332 277 362 339
rect 500 320 576 350
rect 669 337 705 362
rect 916 340 946 379
rect 669 321 868 337
rect 500 311 566 320
rect 500 291 516 311
rect 309 247 362 277
rect 410 277 516 291
rect 550 277 566 311
rect 669 287 750 321
rect 784 287 818 321
rect 852 287 868 321
rect 916 310 981 340
rect 951 295 981 310
rect 669 278 868 287
rect 410 261 566 277
rect 83 51 113 112
rect 201 106 231 132
rect 309 51 339 247
rect 410 232 440 261
rect 614 248 868 278
rect 614 232 644 248
rect 1052 253 1082 379
rect 1239 358 1269 373
rect 1390 358 1420 373
rect 1124 328 1272 358
rect 1124 325 1190 328
rect 1124 291 1140 325
rect 1174 291 1190 325
rect 1124 275 1190 291
rect 1387 280 1423 358
rect 1497 342 1527 357
rect 1611 342 1641 615
rect 1719 542 1749 568
rect 1816 557 1852 615
rect 1819 542 1849 557
rect 2154 536 2184 563
rect 2241 552 2277 615
rect 2345 592 2375 624
rect 2244 536 2274 552
rect 1719 359 1749 374
rect 1819 359 1849 374
rect 2567 592 2597 618
rect 2667 592 2697 618
rect 2567 377 2597 392
rect 2667 377 2697 392
rect 1716 342 1752 359
rect 1494 312 1641 342
rect 1702 326 1768 342
rect 1138 253 1168 275
rect 1238 260 1423 280
rect 410 58 440 84
rect 614 78 644 104
rect 83 21 339 51
rect 951 51 981 167
rect 1238 250 1363 260
rect 1238 235 1268 250
rect 1052 99 1082 125
rect 1138 51 1168 125
rect 1347 226 1363 250
rect 1397 250 1423 260
rect 1397 226 1417 250
rect 1347 192 1417 226
rect 1508 222 1538 312
rect 1702 292 1718 326
rect 1752 292 1768 326
rect 1702 276 1768 292
rect 1347 158 1363 192
rect 1397 158 1417 192
rect 1347 142 1417 158
rect 1238 81 1268 107
rect 1738 222 1768 276
rect 1816 310 1852 359
rect 2154 353 2184 368
rect 2244 353 2274 368
rect 2345 353 2375 368
rect 2564 360 2600 377
rect 2664 360 2700 377
rect 2151 310 2187 353
rect 1816 294 1918 310
rect 1816 260 1845 294
rect 1879 260 1918 294
rect 1816 244 1918 260
rect 1888 222 1918 244
rect 2006 294 2187 310
rect 2241 300 2277 353
rect 2006 260 2045 294
rect 2079 280 2187 294
rect 2079 260 2095 280
rect 2006 244 2095 260
rect 2240 270 2277 300
rect 2342 310 2378 353
rect 2564 344 2700 360
rect 2564 310 2580 344
rect 2614 310 2648 344
rect 2682 310 2700 344
rect 2342 294 2516 310
rect 2006 222 2036 244
rect 2240 222 2270 270
rect 2342 260 2466 294
rect 2500 260 2516 294
rect 2342 244 2516 260
rect 2564 294 2700 310
rect 2342 222 2372 244
rect 951 21 1168 51
rect 1508 48 1538 74
rect 1738 68 1768 94
rect 1888 68 1918 94
rect 2006 68 2036 94
rect 2240 68 2270 94
rect 2564 202 2594 294
rect 2670 202 2700 294
rect 2342 48 2372 74
rect 2564 48 2594 74
rect 2670 48 2700 74
<< polycont >>
rect 385 423 419 457
rect 385 355 419 389
rect 217 298 251 332
rect 516 277 550 311
rect 750 287 784 321
rect 818 287 852 321
rect 1140 291 1174 325
rect 1363 226 1397 260
rect 1718 292 1752 326
rect 1363 158 1397 192
rect 1845 260 1879 294
rect 2045 260 2079 294
rect 2580 310 2614 344
rect 2648 310 2682 344
rect 2466 260 2500 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 22 580 89 596
rect 22 546 39 580
rect 73 546 89 580
rect 22 497 89 546
rect 22 463 39 497
rect 73 463 89 497
rect 22 414 89 463
rect 129 580 163 649
rect 587 627 658 649
rect 129 508 163 546
rect 129 458 163 474
rect 197 609 529 615
rect 197 581 479 609
rect 197 424 231 581
rect 463 575 479 581
rect 513 575 529 609
rect 587 593 605 627
rect 639 593 658 627
rect 692 581 1400 615
rect 692 559 726 581
rect 22 380 39 414
rect 73 380 89 414
rect 22 248 89 380
rect 22 214 38 248
rect 72 214 89 248
rect 22 158 89 214
rect 22 124 38 158
rect 72 124 89 158
rect 133 390 231 424
rect 265 541 335 547
rect 563 541 726 559
rect 941 580 1225 581
rect 265 531 726 541
rect 299 525 726 531
rect 841 539 907 547
rect 299 507 597 525
rect 299 497 335 507
rect 265 440 335 497
rect 841 505 857 539
rect 891 505 907 539
rect 841 491 907 505
rect 631 473 907 491
rect 299 406 335 440
rect 265 390 335 406
rect 133 180 167 390
rect 201 332 267 356
rect 201 298 217 332
rect 251 298 267 332
rect 201 282 267 298
rect 301 248 335 390
rect 226 214 245 248
rect 279 214 335 248
rect 369 468 907 473
rect 369 457 857 468
rect 369 423 385 457
rect 419 439 665 457
rect 419 423 435 439
rect 841 434 857 457
rect 891 434 907 468
rect 369 389 435 423
rect 699 405 732 423
rect 369 355 385 389
rect 419 355 435 389
rect 369 214 435 355
rect 601 389 732 405
rect 766 389 800 423
rect 841 420 907 434
rect 941 546 1069 580
rect 1103 546 1175 580
rect 1209 546 1225 580
rect 601 371 800 389
rect 601 350 689 371
rect 941 353 975 546
rect 1266 512 1332 528
rect 1266 498 1282 512
rect 500 311 566 327
rect 601 316 607 350
rect 641 316 689 350
rect 834 337 975 353
rect 500 277 516 311
rect 550 282 566 311
rect 550 277 621 282
rect 500 248 621 277
rect 369 180 553 214
rect 133 146 335 180
rect 22 108 89 124
rect 301 130 415 146
rect 124 78 140 112
rect 174 78 190 112
rect 301 96 365 130
rect 399 96 415 130
rect 301 80 415 96
rect 451 130 485 146
rect 124 17 190 78
rect 451 17 485 96
rect 519 85 553 180
rect 587 153 621 248
rect 655 237 689 316
rect 734 321 975 337
rect 734 287 750 321
rect 784 287 818 321
rect 852 319 975 321
rect 1009 478 1282 498
rect 1316 478 1332 512
rect 1009 464 1332 478
rect 852 287 868 319
rect 1009 285 1043 464
rect 1266 458 1332 464
rect 976 269 1043 285
rect 1081 424 1127 430
rect 1366 424 1400 581
rect 1081 390 1087 424
rect 1121 390 1127 424
rect 1081 341 1127 390
rect 1211 390 1400 424
rect 1434 569 1500 585
rect 1434 535 1450 569
rect 1484 535 1500 569
rect 1434 498 1500 535
rect 1434 464 1450 498
rect 1484 464 1500 498
rect 1434 427 1500 464
rect 1434 393 1450 427
rect 1484 393 1500 427
rect 1434 390 1500 393
rect 1081 325 1177 341
rect 1081 291 1140 325
rect 1174 291 1177 325
rect 1081 275 1177 291
rect 976 253 992 269
rect 655 221 721 237
rect 655 187 671 221
rect 705 187 721 221
rect 755 235 992 253
rect 1026 235 1043 269
rect 1211 241 1245 390
rect 755 219 1043 235
rect 1077 223 1245 241
rect 755 153 789 219
rect 1077 189 1093 223
rect 1127 207 1245 223
rect 1279 350 1319 356
rect 1313 316 1319 350
rect 1279 310 1319 316
rect 1369 350 1415 356
rect 1369 316 1375 350
rect 1409 316 1415 350
rect 1369 310 1415 316
rect 1127 189 1143 207
rect 1077 187 1143 189
rect 1279 192 1313 310
rect 1369 276 1413 310
rect 587 119 789 153
rect 823 153 1009 185
rect 1177 172 1243 173
rect 1177 153 1193 172
rect 823 151 1193 153
rect 823 85 857 151
rect 975 138 1193 151
rect 1227 138 1243 172
rect 975 119 1243 138
rect 1279 134 1313 158
rect 1347 260 1413 276
rect 1347 226 1363 260
rect 1397 226 1413 260
rect 1466 226 1500 390
rect 1534 569 1600 649
rect 1534 535 1550 569
rect 1584 535 1600 569
rect 1534 486 1600 535
rect 1534 452 1550 486
rect 1584 452 1600 486
rect 1534 403 1600 452
rect 1534 369 1550 403
rect 1584 369 1600 403
rect 1534 353 1600 369
rect 1634 581 2348 615
rect 1634 530 1722 581
rect 1634 496 1672 530
rect 1706 496 1722 530
rect 1634 426 1722 496
rect 1634 392 1672 426
rect 1706 392 1722 426
rect 1634 376 1722 392
rect 1756 531 2163 547
rect 1756 497 1772 531
rect 1806 513 2163 531
rect 1806 497 1822 513
rect 1756 432 1822 497
rect 1756 424 1772 432
rect 1756 390 1768 424
rect 1806 398 1822 432
rect 1802 390 1822 398
rect 1756 376 1822 390
rect 1856 445 1879 479
rect 1913 445 1962 479
rect 1996 445 2045 479
rect 2079 445 2095 479
rect 1856 424 2095 445
rect 1856 411 1977 424
rect 2011 411 2049 424
rect 1856 377 1879 411
rect 1913 377 1962 411
rect 2011 390 2045 411
rect 2083 390 2095 424
rect 1996 377 2045 390
rect 2079 377 2095 390
rect 1634 242 1668 376
rect 1856 361 2095 377
rect 1702 326 1795 342
rect 1702 292 1718 326
rect 1752 292 1795 326
rect 1702 276 1795 292
rect 1634 226 1727 242
rect 1347 192 1413 226
rect 1347 158 1363 192
rect 1397 158 1413 192
rect 1347 142 1413 158
rect 1447 210 1513 226
rect 1447 176 1463 210
rect 1497 176 1513 210
rect 1634 192 1677 226
rect 1711 192 1727 226
rect 1447 158 1513 176
rect 1761 158 1795 276
rect 1829 294 1895 310
rect 1829 260 1845 294
rect 1879 260 1895 294
rect 1829 236 1895 260
rect 1929 226 1995 361
rect 1929 192 1945 226
rect 1979 192 1995 226
rect 2029 294 2095 310
rect 2029 260 2045 294
rect 2079 260 2095 294
rect 2029 244 2095 260
rect 2029 158 2063 244
rect 2129 210 2163 513
rect 1447 124 2063 158
rect 2097 181 2163 210
rect 2097 147 2113 181
rect 2147 147 2163 181
rect 1447 120 1513 124
rect 519 51 857 85
rect 891 101 941 117
rect 925 85 941 101
rect 1447 86 1463 120
rect 1497 86 1513 120
rect 2097 119 2163 147
rect 2197 528 2231 547
rect 2197 413 2231 494
rect 2197 356 2231 379
rect 2277 528 2348 581
rect 2277 494 2292 528
rect 2326 494 2348 528
rect 2277 415 2348 494
rect 2390 608 2458 649
rect 2390 574 2406 608
rect 2440 574 2458 608
rect 2390 540 2458 574
rect 2390 506 2406 540
rect 2440 506 2458 540
rect 2390 472 2458 506
rect 2390 438 2406 472
rect 2440 466 2458 472
rect 2504 580 2570 596
rect 2504 546 2520 580
rect 2554 546 2570 580
rect 2504 512 2570 546
rect 2504 478 2520 512
rect 2554 478 2570 512
rect 2440 438 2444 466
rect 2390 422 2444 438
rect 2504 444 2570 478
rect 2504 432 2520 444
rect 2478 424 2520 432
rect 2277 381 2292 415
rect 2326 381 2348 415
rect 2478 390 2487 424
rect 2554 410 2570 444
rect 2521 394 2570 410
rect 2610 580 2660 649
rect 2644 546 2660 580
rect 2610 512 2660 546
rect 2644 478 2660 512
rect 2610 444 2660 478
rect 2644 410 2660 444
rect 2610 394 2660 410
rect 2694 580 2766 596
rect 2694 546 2710 580
rect 2744 546 2766 580
rect 2694 512 2766 546
rect 2694 478 2710 512
rect 2744 478 2766 512
rect 2694 444 2766 478
rect 2694 410 2710 444
rect 2744 410 2766 444
rect 2694 394 2766 410
rect 2521 390 2530 394
rect 2478 388 2530 390
rect 2197 350 2243 356
rect 2197 316 2203 350
rect 2237 316 2243 350
rect 2197 310 2243 316
rect 1447 85 1513 86
rect 925 67 1513 85
rect 891 51 1513 67
rect 1549 56 1565 90
rect 1599 56 1615 90
rect 1549 17 1615 56
rect 1779 56 1811 90
rect 1845 85 1877 90
rect 2197 85 2231 310
rect 2277 226 2348 381
rect 1845 56 2231 85
rect 2281 210 2348 226
rect 2281 176 2297 210
rect 2331 176 2348 210
rect 2281 120 2348 176
rect 2382 344 2530 388
rect 2564 344 2698 360
rect 2382 192 2416 344
rect 2564 310 2580 344
rect 2614 310 2648 344
rect 2682 310 2698 344
rect 2450 294 2516 310
rect 2564 294 2698 310
rect 2450 260 2466 294
rect 2500 260 2516 294
rect 2732 260 2766 394
rect 2450 226 2766 260
rect 2382 190 2561 192
rect 2382 158 2511 190
rect 2495 156 2511 158
rect 2545 156 2561 190
rect 2281 86 2297 120
rect 2331 86 2348 120
rect 2281 70 2348 86
rect 2383 108 2449 124
rect 2383 74 2399 108
rect 2433 74 2449 108
rect 1779 51 2231 56
rect 2383 17 2449 74
rect 2495 120 2561 156
rect 2495 86 2511 120
rect 2545 86 2561 120
rect 2495 70 2561 86
rect 2595 190 2661 192
rect 2595 156 2611 190
rect 2645 156 2661 190
rect 2595 120 2661 156
rect 2595 86 2611 120
rect 2645 86 2661 120
rect 2595 17 2661 86
rect 2695 190 2766 226
rect 2695 156 2711 190
rect 2745 156 2766 190
rect 2695 120 2766 156
rect 2695 86 2711 120
rect 2745 86 2766 120
rect 2695 70 2766 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 607 316 641 350
rect 1087 390 1121 424
rect 1279 316 1313 350
rect 1375 316 1409 350
rect 1768 398 1772 424
rect 1772 398 1802 424
rect 1768 390 1802 398
rect 1977 411 2011 424
rect 2049 411 2083 424
rect 1977 390 1996 411
rect 1996 390 2011 411
rect 2049 390 2079 411
rect 2079 390 2083 411
rect 2487 410 2520 424
rect 2520 410 2521 424
rect 2487 390 2521 410
rect 2203 316 2237 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
<< metal1 >>
rect 0 683 2784 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 0 617 2784 649
rect 1075 424 1133 430
rect 1075 390 1087 424
rect 1121 421 1133 424
rect 1756 424 1814 430
rect 1756 421 1768 424
rect 1121 393 1768 421
rect 1121 390 1133 393
rect 1075 384 1133 390
rect 1756 390 1768 393
rect 1802 390 1814 424
rect 1756 384 1814 390
rect 1965 424 2095 430
rect 1965 390 1977 424
rect 2011 390 2049 424
rect 2083 421 2095 424
rect 2475 424 2533 430
rect 2475 421 2487 424
rect 2083 393 2487 421
rect 2083 390 2095 393
rect 1965 384 2095 390
rect 2475 390 2487 393
rect 2521 390 2533 424
rect 2475 384 2533 390
rect 595 350 653 356
rect 595 316 607 350
rect 641 347 653 350
rect 1267 350 1325 356
rect 1267 347 1279 350
rect 641 319 1279 347
rect 641 316 653 319
rect 595 310 653 316
rect 1267 316 1279 319
rect 1313 316 1325 350
rect 1267 310 1325 316
rect 1363 350 1421 356
rect 1363 316 1375 350
rect 1409 347 1421 350
rect 2191 350 2249 356
rect 2191 347 2203 350
rect 1409 319 2203 347
rect 1409 316 1421 319
rect 1363 310 1421 316
rect 2191 316 2203 319
rect 2237 316 2249 350
rect 2191 310 2249 316
rect 0 17 2784 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
rect 0 -49 2784 -17
<< labels >>
rlabel comment s 0 0 0 0 4 fah_1
flabel pwell s 0 0 2784 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 0 617 2784 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 2784 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 2784 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 2623 316 2657 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 CI
port 3 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 SUM
port 9 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 SUM
port 9 nsew
flabel corelocali s 31 390 65 424 0 FreeSans 340 0 0 0 SUM
port 9 nsew
flabel corelocali s 31 464 65 498 0 FreeSans 340 0 0 0 SUM
port 9 nsew
flabel corelocali s 31 538 65 572 0 FreeSans 340 0 0 0 SUM
port 9 nsew
flabel corelocali s 319 94 353 128 0 FreeSans 340 0 0 0 COUT
port 8 nsew
flabel corelocali s 1855 242 1889 276 0 FreeSans 340 0 0 0 B
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 2784 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2253010
string GDS_START 2232684
<< end >>
