magic
tech sky130A
magscale 1 2
timestamp 1604502711
<< locali >>
rect 351 383 443 493
rect 20 265 73 337
rect 20 215 155 265
rect 199 215 267 265
rect 393 109 443 383
rect 331 51 443 109
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 57 393 113 527
rect 147 349 207 459
rect 247 383 313 527
rect 147 315 335 349
rect 301 265 335 315
rect 301 199 359 265
rect 301 181 335 199
rect 57 143 335 181
rect 57 71 123 143
rect 247 17 297 109
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
rlabel locali s 20 265 73 337 6 A
port 1 nsew signal input
rlabel locali s 20 215 155 265 6 A
port 1 nsew signal input
rlabel locali s 199 215 267 265 6 B
port 2 nsew signal input
rlabel locali s 393 109 443 383 6 X
port 3 nsew signal output
rlabel locali s 351 383 443 493 6 X
port 3 nsew signal output
rlabel locali s 331 51 443 109 6 X
port 3 nsew signal output
rlabel metal1 s 0 -48 460 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 460 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 460 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3746536
string GDS_START 3741694
<< end >>
