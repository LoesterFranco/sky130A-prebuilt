magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 1746 409 1812 493
rect 1350 357 1812 409
rect 1746 333 1812 357
rect 1942 333 1992 493
rect 2122 333 2188 493
rect 367 289 1254 323
rect 1746 289 2188 333
rect 367 255 401 289
rect 1220 255 1254 289
rect 98 215 401 255
rect 475 215 1186 255
rect 1220 215 1634 255
rect 2141 181 2188 289
rect 1830 131 2188 181
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 17 323 92 493
rect 136 367 186 527
rect 230 401 280 493
rect 324 435 374 527
rect 418 401 468 493
rect 512 435 562 527
rect 606 401 656 493
rect 700 435 750 527
rect 794 401 844 493
rect 230 357 844 401
rect 885 401 948 493
rect 992 435 1042 527
rect 1086 401 1136 493
rect 1180 435 1230 527
rect 1274 443 1708 493
rect 1274 401 1316 443
rect 885 357 1316 401
rect 1848 367 1898 527
rect 230 323 280 357
rect 2036 367 2086 527
rect 17 289 280 323
rect 1298 289 1712 323
rect 17 181 64 289
rect 1678 255 1712 289
rect 1678 215 2107 255
rect 17 129 382 181
rect 426 145 852 181
rect 426 95 476 145
rect 34 51 476 95
rect 520 17 554 111
rect 588 51 664 145
rect 708 17 742 111
rect 776 51 852 145
rect 886 17 940 181
rect 974 147 1796 181
rect 974 145 1634 147
rect 974 51 1050 145
rect 1094 17 1128 111
rect 1162 51 1238 145
rect 1282 17 1316 111
rect 1350 51 1426 145
rect 1470 17 1504 111
rect 1538 51 1614 145
rect 1658 17 1692 111
rect 1746 95 1796 147
rect 1746 61 2188 95
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
<< metal1 >>
rect 0 561 2208 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 0 496 2208 527
rect 0 17 2208 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
rect 0 -48 2208 -17
<< obsm1 >>
rect 211 320 279 329
rect 1331 320 1401 329
rect 211 292 1401 320
rect 211 283 279 292
rect 1331 283 1401 292
<< labels >>
rlabel locali s 475 215 1186 255 6 A
port 1 nsew signal input
rlabel locali s 1220 255 1254 289 6 B
port 2 nsew signal input
rlabel locali s 1220 215 1634 255 6 B
port 2 nsew signal input
rlabel locali s 367 289 1254 323 6 B
port 2 nsew signal input
rlabel locali s 367 255 401 289 6 B
port 2 nsew signal input
rlabel locali s 98 215 401 255 6 B
port 2 nsew signal input
rlabel locali s 2141 181 2188 289 6 Y
port 3 nsew signal output
rlabel locali s 2122 333 2188 493 6 Y
port 3 nsew signal output
rlabel locali s 1942 333 1992 493 6 Y
port 3 nsew signal output
rlabel locali s 1830 131 2188 181 6 Y
port 3 nsew signal output
rlabel locali s 1746 409 1812 493 6 Y
port 3 nsew signal output
rlabel locali s 1746 333 1812 357 6 Y
port 3 nsew signal output
rlabel locali s 1746 289 2188 333 6 Y
port 3 nsew signal output
rlabel locali s 1350 357 1812 409 6 Y
port 3 nsew signal output
rlabel metal1 s 0 -48 2208 48 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 496 2208 592 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2208 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 710770
string GDS_START 695802
<< end >>
