magic
tech sky130A
magscale 1 2
timestamp 1604502705
<< nwell >>
rect -38 332 1286 704
<< pwell >>
rect 0 0 1248 49
<< scnmos >>
rect 84 74 114 222
rect 180 74 210 222
rect 266 74 296 222
rect 352 74 382 222
rect 564 74 594 222
rect 650 74 680 222
rect 741 74 771 222
rect 850 74 880 222
rect 1048 74 1078 222
rect 1134 74 1164 222
<< pmoshvt >>
rect 87 368 117 592
rect 186 368 216 592
rect 286 368 316 592
rect 386 368 416 592
rect 486 368 516 592
rect 654 368 684 592
rect 744 368 774 592
rect 847 368 877 592
rect 972 368 1002 592
rect 1082 368 1112 592
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 142 180 222
rect 114 108 125 142
rect 159 108 180 142
rect 114 74 180 108
rect 210 210 266 222
rect 210 176 221 210
rect 255 176 266 210
rect 210 120 266 176
rect 210 86 221 120
rect 255 86 266 120
rect 210 74 266 86
rect 296 177 352 222
rect 296 143 307 177
rect 341 143 352 177
rect 296 74 352 143
rect 382 127 453 222
rect 382 93 407 127
rect 441 93 453 127
rect 382 74 453 93
rect 507 127 564 222
rect 507 93 519 127
rect 553 93 564 127
rect 507 74 564 93
rect 594 169 650 222
rect 594 135 605 169
rect 639 135 650 169
rect 594 74 650 135
rect 680 210 741 222
rect 680 176 691 210
rect 725 176 741 210
rect 680 120 741 176
rect 680 86 691 120
rect 725 86 741 120
rect 680 74 741 86
rect 771 169 850 222
rect 771 135 791 169
rect 825 135 850 169
rect 771 74 850 135
rect 880 152 937 222
rect 880 118 891 152
rect 925 118 937 152
rect 880 74 937 118
rect 991 152 1048 222
rect 991 118 1003 152
rect 1037 118 1048 152
rect 991 74 1048 118
rect 1078 210 1134 222
rect 1078 176 1089 210
rect 1123 176 1134 210
rect 1078 120 1134 176
rect 1078 86 1089 120
rect 1123 86 1134 120
rect 1078 74 1134 86
rect 1164 188 1221 222
rect 1164 154 1175 188
rect 1209 154 1221 188
rect 1164 120 1221 154
rect 1164 86 1175 120
rect 1209 86 1221 120
rect 1164 74 1221 86
<< pdiff >>
rect 27 580 87 592
rect 27 546 39 580
rect 73 546 87 580
rect 27 510 87 546
rect 27 476 39 510
rect 73 476 87 510
rect 27 440 87 476
rect 27 406 39 440
rect 73 406 87 440
rect 27 368 87 406
rect 117 546 186 592
rect 117 512 139 546
rect 173 512 186 546
rect 117 478 186 512
rect 117 444 139 478
rect 173 444 186 478
rect 117 410 186 444
rect 117 376 139 410
rect 173 376 186 410
rect 117 368 186 376
rect 216 580 286 592
rect 216 546 239 580
rect 273 546 286 580
rect 216 471 286 546
rect 216 437 239 471
rect 273 437 286 471
rect 216 368 286 437
rect 316 547 386 592
rect 316 513 339 547
rect 373 513 386 547
rect 316 479 386 513
rect 316 445 339 479
rect 373 445 386 479
rect 316 411 386 445
rect 316 377 339 411
rect 373 377 386 411
rect 316 368 386 377
rect 416 584 486 592
rect 416 550 439 584
rect 473 550 486 584
rect 416 516 486 550
rect 416 482 439 516
rect 473 482 486 516
rect 416 446 486 482
rect 416 412 439 446
rect 473 412 486 446
rect 416 368 486 412
rect 516 584 654 592
rect 516 550 530 584
rect 564 550 606 584
rect 640 550 654 584
rect 516 516 654 550
rect 516 482 530 516
rect 564 482 606 516
rect 640 482 654 516
rect 516 368 654 482
rect 684 580 744 592
rect 684 546 697 580
rect 731 546 744 580
rect 684 510 744 546
rect 684 476 697 510
rect 731 476 744 510
rect 684 440 744 476
rect 684 406 697 440
rect 731 406 744 440
rect 684 368 744 406
rect 774 580 847 592
rect 774 546 798 580
rect 832 546 847 580
rect 774 492 847 546
rect 774 458 798 492
rect 832 458 847 492
rect 774 368 847 458
rect 877 580 972 592
rect 877 546 900 580
rect 934 546 972 580
rect 877 497 972 546
rect 877 463 900 497
rect 934 463 972 497
rect 877 414 972 463
rect 877 380 925 414
rect 959 380 972 414
rect 877 368 972 380
rect 1002 584 1082 592
rect 1002 550 1025 584
rect 1059 550 1082 584
rect 1002 516 1082 550
rect 1002 482 1025 516
rect 1059 482 1082 516
rect 1002 448 1082 482
rect 1002 414 1025 448
rect 1059 414 1082 448
rect 1002 368 1082 414
rect 1112 580 1171 592
rect 1112 546 1125 580
rect 1159 546 1171 580
rect 1112 497 1171 546
rect 1112 463 1125 497
rect 1159 463 1171 497
rect 1112 414 1171 463
rect 1112 380 1125 414
rect 1159 380 1171 414
rect 1112 368 1171 380
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 125 108 159 142
rect 221 176 255 210
rect 221 86 255 120
rect 307 143 341 177
rect 407 93 441 127
rect 519 93 553 127
rect 605 135 639 169
rect 691 176 725 210
rect 691 86 725 120
rect 791 135 825 169
rect 891 118 925 152
rect 1003 118 1037 152
rect 1089 176 1123 210
rect 1089 86 1123 120
rect 1175 154 1209 188
rect 1175 86 1209 120
<< pdiffc >>
rect 39 546 73 580
rect 39 476 73 510
rect 39 406 73 440
rect 139 512 173 546
rect 139 444 173 478
rect 139 376 173 410
rect 239 546 273 580
rect 239 437 273 471
rect 339 513 373 547
rect 339 445 373 479
rect 339 377 373 411
rect 439 550 473 584
rect 439 482 473 516
rect 439 412 473 446
rect 530 550 564 584
rect 606 550 640 584
rect 530 482 564 516
rect 606 482 640 516
rect 697 546 731 580
rect 697 476 731 510
rect 697 406 731 440
rect 798 546 832 580
rect 798 458 832 492
rect 900 546 934 580
rect 900 463 934 497
rect 925 380 959 414
rect 1025 550 1059 584
rect 1025 482 1059 516
rect 1025 414 1059 448
rect 1125 546 1159 580
rect 1125 463 1159 497
rect 1125 380 1159 414
<< poly >>
rect 87 592 117 618
rect 186 592 216 618
rect 286 592 316 618
rect 386 592 416 618
rect 486 592 516 618
rect 654 592 684 618
rect 744 592 774 618
rect 847 592 877 618
rect 972 592 1002 618
rect 1082 592 1112 618
rect 87 353 117 368
rect 186 353 216 368
rect 286 353 316 368
rect 386 353 416 368
rect 486 353 516 368
rect 654 353 684 368
rect 744 353 774 368
rect 847 353 877 368
rect 972 353 1002 368
rect 1082 353 1112 368
rect 84 326 120 353
rect 183 326 219 353
rect 84 310 219 326
rect 84 276 100 310
rect 134 276 168 310
rect 202 276 219 310
rect 84 260 219 276
rect 283 310 319 353
rect 383 310 419 353
rect 483 310 519 353
rect 651 310 687 353
rect 283 294 435 310
rect 283 274 317 294
rect 266 260 317 274
rect 351 260 385 294
rect 419 260 435 294
rect 84 222 114 260
rect 180 222 210 260
rect 266 244 435 260
rect 483 294 687 310
rect 483 260 505 294
rect 539 260 687 294
rect 483 244 687 260
rect 741 336 777 353
rect 844 336 880 353
rect 741 320 880 336
rect 741 286 757 320
rect 791 286 825 320
rect 859 286 880 320
rect 741 270 880 286
rect 266 222 296 244
rect 352 222 382 244
rect 564 222 594 244
rect 650 222 680 244
rect 741 222 771 270
rect 850 222 880 270
rect 969 310 1005 353
rect 1079 310 1115 353
rect 969 294 1223 310
rect 969 260 1173 294
rect 1207 260 1223 294
rect 969 244 1223 260
rect 1048 222 1078 244
rect 1134 222 1164 244
rect 84 48 114 74
rect 180 48 210 74
rect 266 48 296 74
rect 352 48 382 74
rect 564 48 594 74
rect 650 48 680 74
rect 741 48 771 74
rect 850 48 880 74
rect 1048 48 1078 74
rect 1134 48 1164 74
<< polycont >>
rect 100 276 134 310
rect 168 276 202 310
rect 317 260 351 294
rect 385 260 419 294
rect 505 260 539 294
rect 757 286 791 320
rect 825 286 859 320
rect 1173 260 1207 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 23 584 480 615
rect 23 581 439 584
rect 23 580 89 581
rect 23 546 39 580
rect 73 546 89 580
rect 223 580 289 581
rect 23 510 89 546
rect 23 476 39 510
rect 73 476 89 510
rect 23 440 89 476
rect 23 406 39 440
rect 73 406 89 440
rect 23 390 89 406
rect 123 546 189 547
rect 123 512 139 546
rect 173 512 189 546
rect 123 478 189 512
rect 123 444 139 478
rect 173 444 189 478
rect 123 410 189 444
rect 223 546 239 580
rect 273 546 289 580
rect 423 550 439 581
rect 473 550 480 584
rect 223 471 289 546
rect 223 437 239 471
rect 273 437 289 471
rect 223 428 289 437
rect 323 513 339 547
rect 373 513 389 547
rect 323 479 389 513
rect 323 445 339 479
rect 373 445 389 479
rect 123 376 139 410
rect 173 394 189 410
rect 323 411 389 445
rect 423 516 480 550
rect 423 482 439 516
rect 473 482 480 516
rect 423 446 480 482
rect 514 584 656 649
rect 514 550 530 584
rect 564 550 606 584
rect 640 550 656 584
rect 514 516 656 550
rect 514 482 530 516
rect 564 482 606 516
rect 640 482 656 516
rect 514 480 656 482
rect 690 580 747 596
rect 690 546 697 580
rect 731 546 747 580
rect 690 510 747 546
rect 690 476 697 510
rect 731 476 747 510
rect 690 446 747 476
rect 781 580 850 649
rect 781 546 798 580
rect 832 546 850 580
rect 781 492 850 546
rect 781 458 798 492
rect 832 458 850 492
rect 884 580 975 596
rect 884 546 900 580
rect 934 546 975 580
rect 884 497 975 546
rect 884 463 900 497
rect 934 463 975 497
rect 423 412 439 446
rect 473 440 747 446
rect 473 412 697 440
rect 323 394 339 411
rect 173 377 339 394
rect 373 378 389 411
rect 681 406 697 412
rect 731 424 747 440
rect 884 424 975 463
rect 731 414 975 424
rect 731 406 925 414
rect 681 390 925 406
rect 909 380 925 390
rect 959 380 975 414
rect 1009 584 1075 649
rect 1009 550 1025 584
rect 1059 550 1075 584
rect 1009 516 1075 550
rect 1009 482 1025 516
rect 1059 482 1075 516
rect 1009 448 1075 482
rect 1009 414 1025 448
rect 1059 414 1075 448
rect 1009 412 1075 414
rect 1109 580 1175 596
rect 1109 546 1125 580
rect 1159 546 1175 580
rect 1109 497 1175 546
rect 1109 463 1125 497
rect 1159 463 1175 497
rect 1109 414 1175 463
rect 909 378 975 380
rect 1109 380 1125 414
rect 1159 380 1175 414
rect 1109 378 1175 380
rect 373 377 647 378
rect 173 376 647 377
rect 123 360 647 376
rect 25 326 71 356
rect 323 344 647 360
rect 25 310 218 326
rect 25 276 100 310
rect 134 276 168 310
rect 202 276 218 310
rect 25 260 218 276
rect 301 294 455 310
rect 301 260 317 294
rect 351 260 385 294
rect 419 260 455 294
rect 301 236 455 260
rect 489 294 555 310
rect 489 260 505 294
rect 539 260 555 294
rect 489 236 555 260
rect 601 247 647 344
rect 697 320 875 356
rect 909 344 1175 378
rect 697 286 757 320
rect 791 286 825 320
rect 859 286 875 320
rect 697 270 875 286
rect 1157 294 1223 310
rect 1157 260 1173 294
rect 1207 260 1223 294
rect 23 210 255 226
rect 23 176 39 210
rect 73 192 221 210
rect 23 120 73 176
rect 601 202 641 247
rect 1157 236 1223 260
rect 23 86 39 120
rect 23 70 73 86
rect 109 142 175 158
rect 109 108 125 142
rect 159 108 175 142
rect 109 17 175 108
rect 221 120 255 176
rect 291 177 641 202
rect 291 143 307 177
rect 341 169 641 177
rect 341 168 605 169
rect 341 143 357 168
rect 291 119 357 143
rect 603 135 605 168
rect 639 135 641 169
rect 391 127 457 134
rect 221 85 255 86
rect 391 93 407 127
rect 441 93 457 127
rect 391 85 457 93
rect 221 51 457 85
rect 503 127 569 134
rect 503 93 519 127
rect 553 93 569 127
rect 603 119 641 135
rect 675 210 741 226
rect 675 176 691 210
rect 725 176 741 210
rect 675 120 741 176
rect 503 85 569 93
rect 675 86 691 120
rect 725 86 741 120
rect 775 210 1123 236
rect 775 202 1089 210
rect 775 169 841 202
rect 775 135 791 169
rect 825 135 841 169
rect 1073 176 1089 202
rect 775 119 841 135
rect 875 152 941 168
rect 675 85 741 86
rect 875 118 891 152
rect 925 118 941 152
rect 875 85 941 118
rect 503 51 941 85
rect 987 152 1037 168
rect 987 118 1003 152
rect 987 17 1037 118
rect 1073 120 1123 176
rect 1073 86 1089 120
rect 1073 70 1123 86
rect 1159 188 1225 202
rect 1159 154 1175 188
rect 1209 154 1225 188
rect 1159 120 1225 154
rect 1159 86 1175 120
rect 1209 86 1225 120
rect 1159 17 1225 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
<< metal1 >>
rect 0 683 1248 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 0 617 1248 649
rect 0 17 1248 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
rect 0 -49 1248 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a32oi_2
flabel pwell s 0 0 1248 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 0 617 1248 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 0 617 1248 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 1248 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 B2
port 5 nsew
flabel corelocali s 319 242 353 276 0 FreeSans 340 0 0 0 B1
port 4 nsew
flabel corelocali s 415 242 449 276 0 FreeSans 340 0 0 0 B1
port 4 nsew
flabel corelocali s 1183 242 1217 276 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 511 242 545 276 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 Y
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 1248 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3751420
string GDS_START 3740926
<< end >>
