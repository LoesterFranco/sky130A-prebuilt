magic
tech sky130A
magscale 1 2
timestamp 1604502729
<< locali >>
rect 121 364 189 547
rect 23 236 89 310
rect 123 70 189 364
rect 361 282 427 321
rect 361 88 455 282
rect 361 51 427 88
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 31 581 261 615
rect 31 364 81 581
rect 23 17 89 202
rect 227 389 261 581
rect 301 423 351 649
rect 391 389 457 596
rect 227 355 457 389
rect 223 17 289 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< metal1 >>
rect 0 683 480 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 0 617 480 649
rect 0 17 480 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
rect 0 -49 480 -17
<< labels >>
rlabel locali s 361 282 427 321 6 A
port 1 nsew signal input
rlabel locali s 361 88 455 282 6 A
port 1 nsew signal input
rlabel locali s 361 51 427 88 6 A
port 1 nsew signal input
rlabel locali s 23 236 89 310 6 B
port 2 nsew signal input
rlabel locali s 123 70 189 364 6 Y
port 3 nsew signal output
rlabel locali s 121 364 189 547 6 Y
port 3 nsew signal output
rlabel metal1 s 0 -49 480 49 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 617 480 715 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 480 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1552180
string GDS_START 1546932
<< end >>
