magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 368 561
rect 18 299 69 527
rect 103 333 169 493
rect 203 367 249 527
rect 283 333 349 493
rect 103 299 349 333
rect 22 149 66 265
rect 103 119 139 299
rect 173 153 248 265
rect 289 199 351 265
rect 283 119 349 165
rect 18 17 69 115
rect 103 51 349 119
rect 0 -17 368 17
<< metal1 >>
rect 0 496 368 592
rect 0 -48 368 48
<< labels >>
rlabel locali s 289 199 351 265 6 A
port 1 nsew signal input
rlabel locali s 173 153 248 265 6 B
port 2 nsew signal input
rlabel locali s 22 149 66 265 6 C
port 3 nsew signal input
rlabel locali s 283 333 349 493 6 Y
port 4 nsew signal output
rlabel locali s 283 119 349 165 6 Y
port 4 nsew signal output
rlabel locali s 103 333 169 493 6 Y
port 4 nsew signal output
rlabel locali s 103 299 349 333 6 Y
port 4 nsew signal output
rlabel locali s 103 119 139 299 6 Y
port 4 nsew signal output
rlabel locali s 103 51 349 119 6 Y
port 4 nsew signal output
rlabel locali s 18 17 69 115 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 368 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 368 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 203 367 249 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 18 299 69 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 368 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 368 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 368 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1793200
string GDS_START 1788858
<< end >>
