magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 2246 704
rect 127 311 1324 332
<< pwell >>
rect 0 0 2208 49
<< scnmos >>
rect 84 74 114 222
rect 302 74 332 222
rect 388 74 418 222
rect 502 74 532 222
rect 610 74 640 222
rect 704 74 734 222
rect 790 74 820 222
rect 908 74 938 222
rect 994 74 1024 222
rect 1130 74 1160 222
rect 1208 74 1238 222
rect 1310 74 1340 222
rect 1428 82 1458 230
rect 1514 82 1544 230
rect 1632 82 1662 230
rect 1718 82 1748 230
rect 1836 82 1866 230
rect 1922 82 1952 230
rect 2008 82 2038 230
rect 2094 82 2124 230
<< pmoshvt >>
rect 86 392 116 592
rect 216 347 246 547
rect 415 347 445 547
rect 505 347 535 547
rect 607 347 637 547
rect 707 347 737 547
rect 797 347 827 547
rect 911 347 941 547
rect 1011 347 1041 547
rect 1111 347 1141 547
rect 1205 347 1235 547
rect 1313 368 1343 568
rect 1422 368 1452 592
rect 1512 368 1542 592
rect 1612 368 1642 592
rect 1702 368 1732 592
rect 1802 368 1832 592
rect 1892 368 1922 592
rect 1992 368 2022 592
rect 2082 368 2112 592
<< ndiff >>
rect 1378 222 1428 230
rect 27 199 84 222
rect 27 165 39 199
rect 73 165 84 199
rect 27 120 84 165
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 82 302 222
rect 114 74 161 82
rect 129 48 161 74
rect 195 74 302 82
rect 332 127 388 222
rect 332 93 343 127
rect 377 93 388 127
rect 332 74 388 93
rect 418 202 502 222
rect 418 168 443 202
rect 477 168 502 202
rect 418 120 502 168
rect 418 86 443 120
rect 477 86 502 120
rect 418 74 502 86
rect 532 74 610 222
rect 640 127 704 222
rect 640 93 651 127
rect 685 93 704 127
rect 640 74 704 93
rect 734 127 790 222
rect 734 93 745 127
rect 779 93 790 127
rect 734 74 790 93
rect 820 82 908 222
rect 820 74 847 82
rect 195 48 227 74
rect 835 48 847 74
rect 881 74 908 82
rect 938 127 994 222
rect 938 93 949 127
rect 983 93 994 127
rect 938 74 994 93
rect 1024 177 1130 222
rect 1024 143 1085 177
rect 1119 143 1130 177
rect 1024 74 1130 143
rect 1160 74 1208 222
rect 1238 74 1310 222
rect 1340 82 1428 222
rect 1458 218 1514 230
rect 1458 184 1469 218
rect 1503 184 1514 218
rect 1458 82 1514 184
rect 1544 82 1632 230
rect 1662 218 1718 230
rect 1662 184 1673 218
rect 1707 184 1718 218
rect 1662 82 1718 184
rect 1748 82 1836 230
rect 1866 214 1922 230
rect 1866 180 1877 214
rect 1911 180 1922 214
rect 1866 128 1922 180
rect 1866 94 1877 128
rect 1911 94 1922 128
rect 1866 82 1922 94
rect 1952 146 2008 230
rect 1952 112 1963 146
rect 1997 112 2008 146
rect 1952 82 2008 112
rect 2038 218 2094 230
rect 2038 184 2049 218
rect 2083 184 2094 218
rect 2038 128 2094 184
rect 2038 94 2049 128
rect 2083 94 2094 128
rect 2038 82 2094 94
rect 2124 218 2181 230
rect 2124 184 2135 218
rect 2169 184 2181 218
rect 2124 128 2181 184
rect 2124 94 2135 128
rect 2169 94 2181 128
rect 2124 82 2181 94
rect 1340 74 1367 82
rect 881 48 893 74
rect 1355 48 1367 74
rect 1401 48 1413 82
rect 129 36 227 48
rect 835 36 893 48
rect 1355 36 1413 48
rect 1559 48 1571 82
rect 1605 48 1617 82
rect 1559 36 1617 48
rect 1763 48 1775 82
rect 1809 48 1821 82
rect 1763 36 1821 48
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 510 86 546
rect 27 476 39 510
rect 73 476 86 510
rect 27 440 86 476
rect 27 406 39 440
rect 73 406 86 440
rect 27 392 86 406
rect 116 547 169 592
rect 264 576 397 588
rect 264 547 276 576
rect 116 535 216 547
rect 116 501 129 535
rect 163 501 216 535
rect 116 392 216 501
rect 163 347 216 392
rect 246 542 276 547
rect 310 542 351 576
rect 385 547 397 576
rect 1363 580 1422 592
rect 1363 568 1375 580
rect 1260 547 1313 568
rect 385 542 415 547
rect 246 347 415 542
rect 445 508 505 547
rect 445 474 458 508
rect 492 474 505 508
rect 445 347 505 474
rect 535 347 607 547
rect 637 535 707 547
rect 637 501 650 535
rect 684 501 707 535
rect 637 451 707 501
rect 637 417 650 451
rect 684 417 707 451
rect 637 347 707 417
rect 737 535 797 547
rect 737 501 750 535
rect 784 501 797 535
rect 737 451 797 501
rect 737 417 750 451
rect 784 417 797 451
rect 737 347 797 417
rect 827 535 911 547
rect 827 501 857 535
rect 891 501 911 535
rect 827 347 911 501
rect 941 535 1011 547
rect 941 501 964 535
rect 998 501 1011 535
rect 941 451 1011 501
rect 941 417 964 451
rect 998 417 1011 451
rect 941 347 1011 417
rect 1041 535 1111 547
rect 1041 501 1064 535
rect 1098 501 1111 535
rect 1041 446 1111 501
rect 1041 412 1064 446
rect 1098 412 1111 446
rect 1041 347 1111 412
rect 1141 347 1205 547
rect 1235 368 1313 547
rect 1343 546 1375 568
rect 1409 546 1422 580
rect 1343 508 1422 546
rect 1343 474 1375 508
rect 1409 474 1422 508
rect 1343 368 1422 474
rect 1452 580 1512 592
rect 1452 546 1465 580
rect 1499 546 1512 580
rect 1452 499 1512 546
rect 1452 465 1465 499
rect 1499 465 1512 499
rect 1452 418 1512 465
rect 1452 384 1465 418
rect 1499 384 1512 418
rect 1452 368 1512 384
rect 1542 580 1612 592
rect 1542 546 1555 580
rect 1589 546 1612 580
rect 1542 486 1612 546
rect 1542 452 1555 486
rect 1589 452 1612 486
rect 1542 368 1612 452
rect 1642 580 1702 592
rect 1642 546 1655 580
rect 1689 546 1702 580
rect 1642 499 1702 546
rect 1642 465 1655 499
rect 1689 465 1702 499
rect 1642 418 1702 465
rect 1642 384 1655 418
rect 1689 384 1702 418
rect 1642 368 1702 384
rect 1732 580 1802 592
rect 1732 546 1745 580
rect 1779 546 1802 580
rect 1732 497 1802 546
rect 1732 463 1745 497
rect 1779 463 1802 497
rect 1732 414 1802 463
rect 1732 380 1745 414
rect 1779 380 1802 414
rect 1732 368 1802 380
rect 1832 580 1892 592
rect 1832 546 1845 580
rect 1879 546 1892 580
rect 1832 497 1892 546
rect 1832 463 1845 497
rect 1879 463 1892 497
rect 1832 414 1892 463
rect 1832 380 1845 414
rect 1879 380 1892 414
rect 1832 368 1892 380
rect 1922 580 1992 592
rect 1922 546 1935 580
rect 1969 546 1992 580
rect 1922 482 1992 546
rect 1922 448 1935 482
rect 1969 448 1992 482
rect 1922 368 1992 448
rect 2022 580 2082 592
rect 2022 546 2035 580
rect 2069 546 2082 580
rect 2022 497 2082 546
rect 2022 463 2035 497
rect 2069 463 2082 497
rect 2022 414 2082 463
rect 2022 380 2035 414
rect 2069 380 2082 414
rect 2022 368 2082 380
rect 2112 580 2171 592
rect 2112 546 2125 580
rect 2159 546 2171 580
rect 2112 497 2171 546
rect 2112 463 2125 497
rect 2159 463 2171 497
rect 2112 414 2171 463
rect 2112 380 2125 414
rect 2159 380 2171 414
rect 2112 368 2171 380
rect 1235 347 1288 368
<< ndiffc >>
rect 39 165 73 199
rect 39 86 73 120
rect 161 48 195 82
rect 343 93 377 127
rect 443 168 477 202
rect 443 86 477 120
rect 651 93 685 127
rect 745 93 779 127
rect 847 48 881 82
rect 949 93 983 127
rect 1085 143 1119 177
rect 1469 184 1503 218
rect 1673 184 1707 218
rect 1877 180 1911 214
rect 1877 94 1911 128
rect 1963 112 1997 146
rect 2049 184 2083 218
rect 2049 94 2083 128
rect 2135 184 2169 218
rect 2135 94 2169 128
rect 1367 48 1401 82
rect 1571 48 1605 82
rect 1775 48 1809 82
<< pdiffc >>
rect 39 546 73 580
rect 39 476 73 510
rect 39 406 73 440
rect 129 501 163 535
rect 276 542 310 576
rect 351 542 385 576
rect 458 474 492 508
rect 650 501 684 535
rect 650 417 684 451
rect 750 501 784 535
rect 750 417 784 451
rect 857 501 891 535
rect 964 501 998 535
rect 964 417 998 451
rect 1064 501 1098 535
rect 1064 412 1098 446
rect 1375 546 1409 580
rect 1375 474 1409 508
rect 1465 546 1499 580
rect 1465 465 1499 499
rect 1465 384 1499 418
rect 1555 546 1589 580
rect 1555 452 1589 486
rect 1655 546 1689 580
rect 1655 465 1689 499
rect 1655 384 1689 418
rect 1745 546 1779 580
rect 1745 463 1779 497
rect 1745 380 1779 414
rect 1845 546 1879 580
rect 1845 463 1879 497
rect 1845 380 1879 414
rect 1935 546 1969 580
rect 1935 448 1969 482
rect 2035 546 2069 580
rect 2035 463 2069 497
rect 2035 380 2069 414
rect 2125 546 2159 580
rect 2125 463 2159 497
rect 2125 380 2159 414
<< poly >>
rect 83 615 1346 645
rect 83 607 119 615
rect 86 592 116 607
rect 216 547 246 573
rect 86 377 116 392
rect 83 315 119 377
rect 415 547 445 573
rect 505 547 535 573
rect 604 562 640 615
rect 607 547 637 562
rect 707 547 737 573
rect 797 547 827 573
rect 908 562 944 615
rect 1310 583 1346 615
rect 1422 592 1452 618
rect 1512 592 1542 618
rect 1612 592 1642 618
rect 1702 592 1732 618
rect 1802 592 1832 618
rect 1892 592 1922 618
rect 1992 592 2022 618
rect 2082 592 2112 618
rect 911 547 941 562
rect 1011 547 1041 573
rect 1111 547 1141 573
rect 1205 547 1235 573
rect 1313 568 1343 583
rect 1313 353 1343 368
rect 1422 353 1452 368
rect 1512 353 1542 368
rect 1612 353 1642 368
rect 1702 353 1732 368
rect 1802 353 1832 368
rect 1892 353 1922 368
rect 1992 353 2022 368
rect 2082 353 2112 368
rect 216 332 246 347
rect 415 332 445 347
rect 505 332 535 347
rect 607 332 637 347
rect 707 332 737 347
rect 797 332 827 347
rect 911 332 941 347
rect 1011 332 1041 347
rect 1111 332 1141 347
rect 1205 332 1235 347
rect 213 315 249 332
rect 25 299 159 315
rect 25 265 41 299
rect 75 265 109 299
rect 143 265 159 299
rect 25 249 159 265
rect 213 299 335 315
rect 412 310 448 332
rect 502 315 538 332
rect 213 265 285 299
rect 319 265 335 299
rect 213 249 335 265
rect 388 294 454 310
rect 388 260 404 294
rect 438 260 454 294
rect 84 222 114 249
rect 302 222 332 249
rect 388 244 454 260
rect 496 299 562 315
rect 496 265 512 299
rect 546 265 562 299
rect 496 249 562 265
rect 388 222 418 244
rect 502 222 532 249
rect 604 237 640 332
rect 704 315 740 332
rect 794 315 830 332
rect 682 299 748 315
rect 682 265 698 299
rect 732 265 748 299
rect 682 249 748 265
rect 790 299 856 315
rect 790 265 806 299
rect 840 265 856 299
rect 790 249 856 265
rect 610 222 640 237
rect 704 222 734 249
rect 790 222 820 249
rect 908 237 944 332
rect 1008 310 1044 332
rect 1108 310 1144 332
rect 1202 315 1238 332
rect 1310 323 1346 353
rect 1419 334 1455 353
rect 1509 334 1545 353
rect 1609 334 1645 353
rect 1699 334 1735 353
rect 986 294 1052 310
rect 986 260 1002 294
rect 1036 260 1052 294
rect 986 244 1052 260
rect 1094 294 1160 310
rect 1094 260 1110 294
rect 1144 260 1160 294
rect 1094 244 1160 260
rect 1202 299 1268 315
rect 1202 265 1218 299
rect 1252 265 1268 299
rect 1202 249 1268 265
rect 908 222 938 237
rect 994 222 1024 244
rect 1130 222 1160 244
rect 1208 222 1238 249
rect 1310 222 1340 323
rect 1419 318 1735 334
rect 1419 284 1435 318
rect 1469 284 1503 318
rect 1537 284 1571 318
rect 1605 298 1735 318
rect 1799 330 1835 353
rect 1889 330 1925 353
rect 1989 330 2025 353
rect 2079 330 2115 353
rect 1799 314 2115 330
rect 1605 284 1748 298
rect 1419 268 1748 284
rect 1428 230 1458 268
rect 1514 230 1544 268
rect 1632 230 1662 268
rect 1718 230 1748 268
rect 1799 280 1815 314
rect 1849 280 1883 314
rect 1917 280 1951 314
rect 1985 294 2115 314
rect 1985 280 2124 294
rect 1799 264 2124 280
rect 1836 230 1866 264
rect 1922 230 1952 264
rect 2008 230 2038 264
rect 2094 230 2124 264
rect 84 48 114 74
rect 302 48 332 74
rect 388 48 418 74
rect 502 48 532 74
rect 610 48 640 74
rect 704 48 734 74
rect 790 48 820 74
rect 908 48 938 74
rect 994 48 1024 74
rect 1130 48 1160 74
rect 1208 48 1238 74
rect 1310 48 1340 74
rect 1428 56 1458 82
rect 1514 56 1544 82
rect 1632 56 1662 82
rect 1718 56 1748 82
rect 1836 56 1866 82
rect 1922 56 1952 82
rect 2008 56 2038 82
rect 2094 56 2124 82
<< polycont >>
rect 41 265 75 299
rect 109 265 143 299
rect 285 265 319 299
rect 404 260 438 294
rect 512 265 546 299
rect 698 265 732 299
rect 806 265 840 299
rect 1002 260 1036 294
rect 1110 260 1144 294
rect 1218 265 1252 299
rect 1435 284 1469 318
rect 1503 284 1537 318
rect 1571 284 1605 318
rect 1815 280 1849 314
rect 1883 280 1917 314
rect 1951 280 1985 314
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 23 580 89 596
rect 23 546 39 580
rect 73 546 89 580
rect 23 510 89 546
rect 23 476 39 510
rect 73 476 89 510
rect 129 535 163 649
rect 129 485 163 501
rect 197 576 401 592
rect 197 542 276 576
rect 310 542 351 576
rect 385 542 401 576
rect 197 526 401 542
rect 23 451 89 476
rect 197 451 231 526
rect 442 508 508 551
rect 442 492 458 508
rect 23 440 231 451
rect 23 406 39 440
rect 73 417 231 440
rect 265 474 458 492
rect 492 474 508 508
rect 265 458 508 474
rect 634 535 700 649
rect 634 501 650 535
rect 684 501 700 535
rect 73 406 89 417
rect 23 390 89 406
rect 265 383 299 458
rect 634 451 700 501
rect 25 299 167 356
rect 25 265 41 299
rect 75 265 109 299
rect 143 265 167 299
rect 25 249 167 265
rect 201 349 299 383
rect 333 390 530 424
rect 634 417 650 451
rect 684 417 700 451
rect 734 535 800 551
rect 734 501 750 535
rect 784 501 800 535
rect 734 451 800 501
rect 834 535 914 649
rect 1359 580 1409 649
rect 834 501 857 535
rect 891 501 914 535
rect 834 485 914 501
rect 948 535 1014 551
rect 948 501 964 535
rect 998 501 1014 535
rect 948 451 1014 501
rect 734 417 750 451
rect 784 417 964 451
rect 998 417 1014 451
rect 1048 535 1114 551
rect 1048 501 1064 535
rect 1098 501 1114 535
rect 1048 446 1114 501
rect 1359 546 1375 580
rect 1359 508 1409 546
rect 1359 474 1375 508
rect 1359 458 1409 474
rect 1449 580 1515 596
rect 1449 546 1465 580
rect 1499 546 1515 580
rect 1449 499 1515 546
rect 1449 465 1465 499
rect 1499 465 1515 499
rect 1048 412 1064 446
rect 1098 424 1285 446
rect 1098 412 1415 424
rect 1251 390 1415 412
rect 201 218 235 349
rect 333 315 367 390
rect 496 383 530 390
rect 496 378 924 383
rect 496 356 1217 378
rect 269 299 367 315
rect 269 265 285 299
rect 319 265 367 299
rect 269 252 367 265
rect 401 294 455 356
rect 401 260 404 294
rect 438 276 455 294
rect 401 242 415 260
rect 449 242 455 276
rect 496 349 1319 356
rect 496 299 562 349
rect 496 265 512 299
rect 546 265 562 299
rect 496 249 562 265
rect 601 299 748 315
rect 601 276 698 299
rect 401 236 455 242
rect 601 242 607 276
rect 641 265 698 276
rect 732 265 748 299
rect 641 252 748 265
rect 790 299 856 349
rect 890 344 1319 349
rect 1183 310 1319 344
rect 1381 334 1415 390
rect 1449 418 1515 465
rect 1555 580 1605 649
rect 1589 546 1605 580
rect 1555 486 1605 546
rect 1589 452 1605 486
rect 1555 436 1605 452
rect 1639 580 1705 596
rect 1639 546 1655 580
rect 1689 546 1705 580
rect 1639 499 1705 546
rect 1639 465 1655 499
rect 1689 465 1705 499
rect 1449 384 1465 418
rect 1499 402 1515 418
rect 1639 418 1705 465
rect 1639 402 1655 418
rect 1499 384 1655 402
rect 1689 384 1705 418
rect 1449 368 1705 384
rect 1381 318 1621 334
rect 790 265 806 299
rect 840 265 856 299
rect 790 252 856 265
rect 986 294 1052 310
rect 986 260 1002 294
rect 1036 260 1052 294
rect 641 242 643 252
rect 601 236 643 242
rect 986 244 1052 260
rect 1086 294 1149 310
rect 1086 276 1110 294
rect 986 218 1051 244
rect 1086 242 1087 276
rect 1144 260 1149 294
rect 1121 242 1149 260
rect 1183 299 1268 310
rect 1183 265 1218 299
rect 1252 265 1268 299
rect 1183 252 1268 265
rect 1381 284 1435 318
rect 1469 284 1503 318
rect 1537 284 1571 318
rect 1605 284 1621 318
rect 1381 268 1621 284
rect 1086 236 1149 242
rect 1381 218 1415 268
rect 1657 234 1705 368
rect 1745 580 1795 649
rect 1779 546 1795 580
rect 1745 497 1795 546
rect 1779 463 1795 497
rect 1745 414 1795 463
rect 1779 380 1795 414
rect 1745 364 1795 380
rect 1829 580 1895 596
rect 1829 546 1845 580
rect 1879 546 1895 580
rect 1829 497 1895 546
rect 1829 463 1845 497
rect 1879 463 1895 497
rect 1829 414 1895 463
rect 1935 580 1985 649
rect 1969 546 1985 580
rect 1935 482 1985 546
rect 1969 448 1985 482
rect 1935 432 1985 448
rect 2019 580 2087 596
rect 2019 546 2035 580
rect 2069 546 2087 580
rect 2019 497 2087 546
rect 2019 463 2035 497
rect 2069 463 2087 497
rect 1829 380 1845 414
rect 1879 398 1895 414
rect 2019 414 2087 463
rect 2019 398 2035 414
rect 1879 380 2035 398
rect 2069 380 2087 414
rect 1829 364 2087 380
rect 2125 580 2175 649
rect 2159 546 2175 580
rect 2125 497 2175 546
rect 2159 463 2175 497
rect 2125 414 2175 463
rect 2159 380 2175 414
rect 2125 364 2175 380
rect 1793 314 1991 330
rect 1793 280 1815 314
rect 1849 280 1883 314
rect 1917 280 1951 314
rect 1985 280 1991 314
rect 1793 264 1991 280
rect 2033 310 2087 364
rect 23 199 89 215
rect 23 165 39 199
rect 73 165 89 199
rect 201 202 367 218
rect 677 202 1051 218
rect 1183 202 1415 218
rect 201 184 443 202
rect 333 168 443 184
rect 477 184 1051 202
rect 477 168 711 184
rect 23 150 89 165
rect 23 134 299 150
rect 23 127 393 134
rect 23 120 343 127
rect 23 86 39 120
rect 73 116 343 120
rect 73 86 89 116
rect 23 70 89 86
rect 265 93 343 116
rect 377 93 393 127
rect 125 48 161 82
rect 195 48 231 82
rect 265 70 393 93
rect 427 120 493 168
rect 427 86 443 120
rect 477 86 493 120
rect 427 70 493 86
rect 635 127 701 134
rect 635 93 651 127
rect 685 93 701 127
rect 125 17 231 48
rect 635 17 701 93
rect 745 127 983 150
rect 779 116 949 127
rect 779 93 795 116
rect 745 70 795 93
rect 933 93 949 116
rect 831 48 847 82
rect 881 48 897 82
rect 933 70 983 93
rect 1017 85 1051 184
rect 1085 184 1415 202
rect 1453 218 1723 234
rect 1453 184 1469 218
rect 1503 184 1673 218
rect 1707 184 1723 218
rect 1085 177 1217 184
rect 1119 168 1217 177
rect 1119 143 1135 168
rect 1793 150 1827 264
rect 2033 230 2085 310
rect 1085 119 1135 143
rect 1251 116 1827 150
rect 1861 218 2085 230
rect 1861 214 2049 218
rect 1861 180 1877 214
rect 1911 196 2049 214
rect 1861 128 1911 180
rect 2033 184 2049 196
rect 2083 184 2085 218
rect 1251 85 1285 116
rect 1017 51 1285 85
rect 1861 94 1877 128
rect 831 17 897 48
rect 1351 48 1367 82
rect 1401 48 1417 82
rect 1351 17 1417 48
rect 1555 48 1571 82
rect 1605 48 1621 82
rect 1555 17 1621 48
rect 1759 48 1775 82
rect 1809 48 1825 82
rect 1861 78 1911 94
rect 1947 146 1997 162
rect 1947 112 1963 146
rect 1759 17 1825 48
rect 1947 17 1997 112
rect 2033 128 2085 184
rect 2033 94 2049 128
rect 2083 94 2085 128
rect 2033 78 2085 94
rect 2119 218 2185 234
rect 2119 184 2135 218
rect 2169 184 2185 218
rect 2119 128 2185 184
rect 2119 94 2135 128
rect 2169 94 2185 128
rect 2119 17 2185 94
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 415 260 438 276
rect 438 260 449 276
rect 415 242 449 260
rect 607 242 641 276
rect 1087 260 1110 276
rect 1110 260 1121 276
rect 1087 242 1121 260
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
<< metal1 >>
rect 0 683 2208 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 0 617 2208 649
rect 403 276 461 282
rect 403 242 415 276
rect 449 273 461 276
rect 595 276 653 282
rect 595 273 607 276
rect 449 245 607 273
rect 449 242 461 245
rect 403 236 461 242
rect 595 242 607 245
rect 641 273 653 276
rect 1075 276 1133 282
rect 1075 273 1087 276
rect 641 245 1087 273
rect 641 242 653 245
rect 595 236 653 242
rect 1075 242 1087 245
rect 1121 242 1133 276
rect 1075 236 1133 242
rect 0 17 2208 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
rect 0 -49 2208 -17
<< labels >>
rlabel comment s 0 0 0 0 4 fa_4
flabel pwell s 0 0 2208 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 0 617 2208 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 415 242 449 276 0 FreeSans 340 0 0 0 CIN
port 3 nsew
flabel metal1 s 0 617 2208 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 2208 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 1183 316 1217 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 1279 316 1313 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 2047 316 2081 350 0 FreeSans 340 0 0 0 COUT
port 8 nsew
flabel corelocali s 2047 390 2081 424 0 FreeSans 340 0 0 0 COUT
port 8 nsew
flabel corelocali s 2047 464 2081 498 0 FreeSans 340 0 0 0 COUT
port 8 nsew
flabel corelocali s 2047 538 2081 572 0 FreeSans 340 0 0 0 COUT
port 8 nsew
flabel corelocali s 1663 390 1697 424 0 FreeSans 340 0 0 0 SUM
port 9 nsew
flabel corelocali s 1663 464 1697 498 0 FreeSans 340 0 0 0 SUM
port 9 nsew
flabel corelocali s 1663 538 1697 572 0 FreeSans 340 0 0 0 SUM
port 9 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 2208 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2232630
string GDS_START 2215556
<< end >>
