magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 129 430 195 547
rect 129 394 359 430
rect 107 360 359 394
rect 107 226 141 360
rect 107 123 175 226
rect 593 236 659 330
rect 697 270 773 356
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 29 581 295 615
rect 336 584 402 649
rect 29 428 95 581
rect 229 550 295 581
rect 443 550 509 596
rect 229 516 509 550
rect 645 522 741 649
rect 229 464 295 516
rect 775 482 841 572
rect 393 448 841 482
rect 393 326 427 448
rect 175 260 427 326
rect 479 364 621 414
rect 775 390 841 448
rect 23 85 73 226
rect 209 192 445 226
rect 209 85 275 192
rect 23 51 275 85
rect 309 17 359 158
rect 395 70 445 192
rect 479 202 545 364
rect 807 206 841 390
rect 479 65 634 202
rect 668 17 734 202
rect 768 70 841 206
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel locali s 697 270 773 356 6 A
port 1 nsew signal input
rlabel locali s 593 236 659 330 6 TE_B
port 2 nsew signal input
rlabel locali s 129 430 195 547 6 Z
port 3 nsew signal output
rlabel locali s 129 394 359 430 6 Z
port 3 nsew signal output
rlabel locali s 107 360 359 394 6 Z
port 3 nsew signal output
rlabel locali s 107 226 141 360 6 Z
port 3 nsew signal output
rlabel locali s 107 123 175 226 6 Z
port 3 nsew signal output
rlabel metal1 s 0 -49 864 49 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 617 864 715 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2050804
string GDS_START 2043612
<< end >>
