magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 87 290 161 356
rect 195 290 261 356
rect 1240 412 1334 596
rect 1085 236 1159 310
rect 1300 236 1334 412
rect 1226 202 1334 236
rect 1543 364 1611 596
rect 1226 70 1292 202
rect 1577 208 1611 364
rect 1542 70 1611 208
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 19 512 89 570
rect 130 546 196 649
rect 470 546 537 649
rect 571 581 803 615
rect 19 478 535 512
rect 19 394 89 478
rect 237 394 329 444
rect 19 256 53 394
rect 295 350 329 394
rect 363 388 443 444
rect 295 284 375 350
rect 295 256 329 284
rect 19 138 89 256
rect 125 17 191 256
rect 237 150 329 256
rect 409 260 443 388
rect 501 360 535 478
rect 571 428 605 581
rect 639 481 703 547
rect 571 394 635 428
rect 501 294 567 360
rect 601 296 635 394
rect 669 364 703 481
rect 737 410 803 581
rect 881 530 1016 649
rect 1050 464 1116 596
rect 845 398 1116 464
rect 1156 412 1206 649
rect 1017 378 1116 398
rect 669 330 983 364
rect 601 260 679 296
rect 409 250 679 260
rect 365 226 679 250
rect 365 184 443 226
rect 716 192 750 330
rect 917 270 983 330
rect 1017 344 1266 378
rect 1017 226 1051 344
rect 1201 270 1266 344
rect 237 116 598 150
rect 638 142 750 192
rect 237 100 329 116
rect 564 102 598 116
rect 464 17 530 82
rect 564 51 781 102
rect 848 17 914 212
rect 960 70 1051 226
rect 1368 330 1402 596
rect 1442 420 1508 649
rect 1368 264 1543 330
rect 1124 17 1190 202
rect 1368 168 1404 264
rect 1338 70 1404 168
rect 1440 17 1506 188
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
rlabel locali s 87 290 161 356 6 D
port 1 nsew signal input
rlabel locali s 1300 236 1334 412 6 Q
port 2 nsew signal output
rlabel locali s 1240 412 1334 596 6 Q
port 2 nsew signal output
rlabel locali s 1226 202 1334 236 6 Q
port 2 nsew signal output
rlabel locali s 1226 70 1292 202 6 Q
port 2 nsew signal output
rlabel locali s 1577 208 1611 364 6 Q_N
port 3 nsew signal output
rlabel locali s 1543 364 1611 596 6 Q_N
port 3 nsew signal output
rlabel locali s 1542 70 1611 208 6 Q_N
port 3 nsew signal output
rlabel locali s 1085 236 1159 310 6 RESET_B
port 4 nsew signal input
rlabel locali s 195 290 261 356 6 GATE
port 5 nsew clock input
rlabel metal1 s 0 -49 1632 49 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1632 715 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2856170
string GDS_START 2843470
<< end >>
