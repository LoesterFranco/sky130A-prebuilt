magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 103 195 157 349
rect 331 370 443 493
rect 191 213 257 265
rect 407 179 443 370
rect 227 145 443 179
rect 227 51 303 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 155 451 221 527
rect 19 383 297 417
rect 19 58 69 383
rect 263 333 297 383
rect 263 299 331 333
rect 297 265 331 299
rect 297 215 373 265
rect 135 17 193 125
rect 347 17 424 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
rlabel locali s 191 213 257 265 6 A
port 1 nsew signal input
rlabel locali s 103 195 157 349 6 B_N
port 2 nsew signal input
rlabel locali s 407 179 443 370 6 Y
port 3 nsew signal output
rlabel locali s 331 370 443 493 6 Y
port 3 nsew signal output
rlabel locali s 227 145 443 179 6 Y
port 3 nsew signal output
rlabel locali s 227 51 303 145 6 Y
port 3 nsew signal output
rlabel metal1 s 0 -48 460 48 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 496 460 592 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 460 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2414358
string GDS_START 2410072
<< end >>
