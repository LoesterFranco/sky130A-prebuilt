magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 828 561
rect 27 391 69 493
rect 103 425 169 527
rect 203 391 237 493
rect 27 357 237 391
rect 543 428 609 527
rect 27 165 69 357
rect 743 383 810 527
rect 469 289 510 323
rect 27 131 169 165
rect 223 149 306 255
rect 469 249 503 289
rect 661 265 709 325
rect 417 215 503 249
rect 537 191 597 265
rect 633 199 709 265
rect 763 199 811 326
rect 18 17 85 93
rect 187 17 328 89
rect 551 122 597 191
rect 551 83 621 122
rect 661 85 709 199
rect 743 17 810 161
rect 0 -17 828 17
<< obsli1 >>
rect 307 459 509 493
rect 307 357 341 459
rect 375 389 441 423
rect 475 393 509 459
rect 675 393 709 493
rect 375 323 425 389
rect 475 359 709 393
rect 107 289 425 323
rect 107 199 141 289
rect 340 157 378 289
rect 340 123 517 157
rect 451 55 517 123
<< metal1 >>
rect 0 496 828 592
rect 0 -48 828 48
<< labels >>
rlabel locali s 551 122 597 191 6 A1
port 1 nsew signal input
rlabel locali s 551 83 621 122 6 A1
port 1 nsew signal input
rlabel locali s 537 191 597 265 6 A1
port 1 nsew signal input
rlabel locali s 661 265 709 325 6 A2
port 2 nsew signal input
rlabel locali s 661 85 709 199 6 A2
port 2 nsew signal input
rlabel locali s 633 199 709 265 6 A2
port 2 nsew signal input
rlabel locali s 763 199 811 326 6 A3
port 3 nsew signal input
rlabel locali s 469 289 510 323 6 B1
port 4 nsew signal input
rlabel locali s 469 249 503 289 6 B1
port 4 nsew signal input
rlabel locali s 417 215 503 249 6 B1
port 4 nsew signal input
rlabel locali s 223 149 306 255 6 B2
port 5 nsew signal input
rlabel locali s 203 391 237 493 6 X
port 6 nsew signal output
rlabel locali s 27 391 69 493 6 X
port 6 nsew signal output
rlabel locali s 27 357 237 391 6 X
port 6 nsew signal output
rlabel locali s 27 165 69 357 6 X
port 6 nsew signal output
rlabel locali s 27 131 169 165 6 X
port 6 nsew signal output
rlabel locali s 743 17 810 161 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 187 17 328 89 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 18 17 85 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 828 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 828 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 743 383 810 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 543 428 609 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 103 425 169 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 828 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 828 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3629138
string GDS_START 3620756
<< end >>
