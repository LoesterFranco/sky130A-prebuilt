magic
tech sky130A
magscale 1 2
timestamp 1601050082
<< locali >>
rect 213 492 279 547
rect 505 492 559 596
rect 213 458 559 492
rect 53 390 455 424
rect 53 270 119 390
rect 169 270 303 356
rect 351 270 455 390
rect 505 364 559 458
rect 505 226 547 364
rect 581 236 647 310
rect 495 143 547 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 23 458 73 649
rect 113 581 379 615
rect 113 458 179 581
rect 313 526 379 581
rect 419 526 469 649
rect 599 364 649 649
rect 23 202 461 236
rect 23 70 89 202
rect 123 17 189 166
rect 225 70 275 202
rect 309 17 375 166
rect 411 104 461 202
rect 583 104 649 202
rect 411 70 649 104
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel locali s 351 270 455 390 6 A1
port 1 nsew signal input
rlabel locali s 53 390 455 424 6 A1
port 1 nsew signal input
rlabel locali s 53 270 119 390 6 A1
port 1 nsew signal input
rlabel locali s 169 270 303 356 6 A2
port 2 nsew signal input
rlabel locali s 581 236 647 310 6 B1
port 3 nsew signal input
rlabel locali s 505 492 559 596 6 Y
port 4 nsew signal output
rlabel locali s 505 364 559 458 6 Y
port 4 nsew signal output
rlabel locali s 505 226 547 364 6 Y
port 4 nsew signal output
rlabel locali s 495 143 547 226 6 Y
port 4 nsew signal output
rlabel locali s 213 492 279 547 6 Y
port 4 nsew signal output
rlabel locali s 213 458 559 492 6 Y
port 4 nsew signal output
rlabel metal1 s 0 -49 672 49 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 617 672 715 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1353620
string GDS_START 1347090
<< end >>
