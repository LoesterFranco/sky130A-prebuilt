magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 1094 704
<< pwell >>
rect 0 0 1056 49
<< scnmos >>
rect 98 74 128 158
rect 184 74 214 158
rect 293 74 323 158
rect 384 74 414 158
rect 498 74 528 158
rect 584 74 614 158
rect 670 74 700 158
rect 756 74 786 158
rect 856 74 886 158
rect 942 74 972 158
<< pmoshvt >>
rect 95 368 125 592
rect 186 368 216 592
rect 296 368 326 592
rect 386 368 416 592
rect 476 368 506 592
rect 566 368 596 592
rect 656 368 686 592
rect 746 368 776 592
rect 846 368 876 592
rect 939 368 969 592
<< ndiff >>
rect 27 133 98 158
rect 27 99 39 133
rect 73 99 98 133
rect 27 74 98 99
rect 128 133 184 158
rect 128 99 139 133
rect 173 99 184 133
rect 128 74 184 99
rect 214 133 293 158
rect 214 99 239 133
rect 273 99 293 133
rect 214 74 293 99
rect 323 133 384 158
rect 323 99 339 133
rect 373 99 384 133
rect 323 74 384 99
rect 414 120 498 158
rect 414 86 439 120
rect 473 86 498 120
rect 414 74 498 86
rect 528 133 584 158
rect 528 99 539 133
rect 573 99 584 133
rect 528 74 584 99
rect 614 120 670 158
rect 614 86 625 120
rect 659 86 670 120
rect 614 74 670 86
rect 700 133 756 158
rect 700 99 711 133
rect 745 99 756 133
rect 700 74 756 99
rect 786 120 856 158
rect 786 86 804 120
rect 838 86 856 120
rect 786 74 856 86
rect 886 133 942 158
rect 886 99 897 133
rect 931 99 942 133
rect 886 74 942 99
rect 972 120 1029 158
rect 972 86 983 120
rect 1017 86 1029 120
rect 972 74 1029 86
<< pdiff >>
rect 27 580 95 592
rect 27 546 39 580
rect 73 546 95 580
rect 27 510 95 546
rect 27 476 39 510
rect 73 476 95 510
rect 27 440 95 476
rect 27 406 39 440
rect 73 406 95 440
rect 27 368 95 406
rect 125 580 186 592
rect 125 546 139 580
rect 173 546 186 580
rect 125 510 186 546
rect 125 476 139 510
rect 173 476 186 510
rect 125 440 186 476
rect 125 406 139 440
rect 173 406 186 440
rect 125 368 186 406
rect 216 580 296 592
rect 216 546 239 580
rect 273 546 296 580
rect 216 508 296 546
rect 216 474 239 508
rect 273 474 296 508
rect 216 368 296 474
rect 326 580 386 592
rect 326 546 339 580
rect 373 546 386 580
rect 326 497 386 546
rect 326 463 339 497
rect 373 463 386 497
rect 326 414 386 463
rect 326 380 339 414
rect 373 380 386 414
rect 326 368 386 380
rect 416 580 476 592
rect 416 546 429 580
rect 463 546 476 580
rect 416 508 476 546
rect 416 474 429 508
rect 463 474 476 508
rect 416 440 476 474
rect 416 406 429 440
rect 463 406 476 440
rect 416 368 476 406
rect 506 580 566 592
rect 506 546 519 580
rect 553 546 566 580
rect 506 497 566 546
rect 506 463 519 497
rect 553 463 566 497
rect 506 414 566 463
rect 506 380 519 414
rect 553 380 566 414
rect 506 368 566 380
rect 596 580 656 592
rect 596 546 609 580
rect 643 546 656 580
rect 596 456 656 546
rect 596 422 609 456
rect 643 422 656 456
rect 596 368 656 422
rect 686 580 746 592
rect 686 546 699 580
rect 733 546 746 580
rect 686 497 746 546
rect 686 463 699 497
rect 733 463 746 497
rect 686 414 746 463
rect 686 380 699 414
rect 733 380 746 414
rect 686 368 746 380
rect 776 580 846 592
rect 776 546 789 580
rect 823 546 846 580
rect 776 508 846 546
rect 776 474 789 508
rect 823 474 846 508
rect 776 440 846 474
rect 776 406 789 440
rect 823 406 846 440
rect 776 368 846 406
rect 876 580 939 592
rect 876 546 890 580
rect 924 546 939 580
rect 876 497 939 546
rect 876 463 890 497
rect 924 463 939 497
rect 876 414 939 463
rect 876 380 890 414
rect 924 380 939 414
rect 876 368 939 380
rect 969 580 1028 592
rect 969 546 982 580
rect 1016 546 1028 580
rect 969 508 1028 546
rect 969 474 982 508
rect 1016 474 1028 508
rect 969 440 1028 474
rect 969 406 982 440
rect 1016 406 1028 440
rect 969 368 1028 406
<< ndiffc >>
rect 39 99 73 133
rect 139 99 173 133
rect 239 99 273 133
rect 339 99 373 133
rect 439 86 473 120
rect 539 99 573 133
rect 625 86 659 120
rect 711 99 745 133
rect 804 86 838 120
rect 897 99 931 133
rect 983 86 1017 120
<< pdiffc >>
rect 39 546 73 580
rect 39 476 73 510
rect 39 406 73 440
rect 139 546 173 580
rect 139 476 173 510
rect 139 406 173 440
rect 239 546 273 580
rect 239 474 273 508
rect 339 546 373 580
rect 339 463 373 497
rect 339 380 373 414
rect 429 546 463 580
rect 429 474 463 508
rect 429 406 463 440
rect 519 546 553 580
rect 519 463 553 497
rect 519 380 553 414
rect 609 546 643 580
rect 609 422 643 456
rect 699 546 733 580
rect 699 463 733 497
rect 699 380 733 414
rect 789 546 823 580
rect 789 474 823 508
rect 789 406 823 440
rect 890 546 924 580
rect 890 463 924 497
rect 890 380 924 414
rect 982 546 1016 580
rect 982 474 1016 508
rect 982 406 1016 440
<< poly >>
rect 95 592 125 618
rect 186 592 216 618
rect 296 592 326 618
rect 386 592 416 618
rect 476 592 506 618
rect 566 592 596 618
rect 656 592 686 618
rect 746 592 776 618
rect 846 592 876 618
rect 939 592 969 618
rect 95 353 125 368
rect 186 353 216 368
rect 296 353 326 368
rect 386 353 416 368
rect 476 353 506 368
rect 566 353 596 368
rect 656 353 686 368
rect 746 353 776 368
rect 846 353 876 368
rect 939 353 969 368
rect 92 336 128 353
rect 183 336 219 353
rect 85 320 219 336
rect 85 286 101 320
rect 135 286 169 320
rect 203 286 219 320
rect 85 270 219 286
rect 293 304 329 353
rect 383 304 419 353
rect 473 304 509 353
rect 563 304 599 353
rect 653 304 689 353
rect 743 304 779 353
rect 843 304 879 353
rect 936 304 972 353
rect 293 288 972 304
rect 98 158 128 270
rect 184 158 214 270
rect 293 254 309 288
rect 343 254 377 288
rect 411 254 445 288
rect 479 254 513 288
rect 547 254 581 288
rect 615 254 649 288
rect 683 254 717 288
rect 751 254 785 288
rect 819 254 853 288
rect 887 254 972 288
rect 293 238 972 254
rect 293 158 323 238
rect 384 158 414 238
rect 498 158 528 238
rect 584 158 614 238
rect 670 158 700 238
rect 756 158 786 238
rect 856 158 886 238
rect 942 158 972 238
rect 98 48 128 74
rect 184 48 214 74
rect 293 48 323 74
rect 384 48 414 74
rect 498 48 528 74
rect 584 48 614 74
rect 670 48 700 74
rect 756 48 786 74
rect 856 48 886 74
rect 942 48 972 74
<< polycont >>
rect 101 286 135 320
rect 169 286 203 320
rect 309 254 343 288
rect 377 254 411 288
rect 445 254 479 288
rect 513 254 547 288
rect 581 254 615 288
rect 649 254 683 288
rect 717 254 751 288
rect 785 254 819 288
rect 853 254 887 288
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 23 580 89 649
rect 23 546 39 580
rect 73 546 89 580
rect 23 510 89 546
rect 23 476 39 510
rect 73 476 89 510
rect 23 440 89 476
rect 23 406 39 440
rect 73 406 89 440
rect 23 390 89 406
rect 123 580 189 596
rect 123 546 139 580
rect 173 546 189 580
rect 123 510 189 546
rect 123 476 139 510
rect 173 476 189 510
rect 123 440 189 476
rect 223 580 289 649
rect 223 546 239 580
rect 273 546 289 580
rect 223 508 289 546
rect 223 474 239 508
rect 273 474 289 508
rect 223 458 289 474
rect 323 580 376 596
rect 323 546 339 580
rect 373 546 376 580
rect 323 497 376 546
rect 323 463 339 497
rect 373 463 376 497
rect 123 406 139 440
rect 173 424 189 440
rect 173 406 289 424
rect 123 390 289 406
rect 25 320 219 356
rect 25 286 101 320
rect 135 286 169 320
rect 203 286 219 320
rect 25 270 219 286
rect 255 304 289 390
rect 323 414 376 463
rect 323 380 339 414
rect 373 380 376 414
rect 413 580 479 649
rect 413 546 429 580
rect 463 546 479 580
rect 413 508 479 546
rect 413 474 429 508
rect 463 474 479 508
rect 413 440 479 474
rect 413 406 429 440
rect 463 406 479 440
rect 517 580 569 596
rect 517 546 519 580
rect 553 546 569 580
rect 517 497 569 546
rect 517 463 519 497
rect 553 463 569 497
rect 517 414 569 463
rect 323 372 376 380
rect 517 380 519 414
rect 553 380 569 414
rect 609 580 643 649
rect 609 456 643 546
rect 609 406 643 422
rect 683 580 736 596
rect 683 546 699 580
rect 733 546 736 580
rect 683 497 736 546
rect 683 463 699 497
rect 733 463 736 497
rect 683 414 736 463
rect 517 372 569 380
rect 683 380 699 414
rect 733 380 736 414
rect 773 580 839 649
rect 773 546 789 580
rect 823 546 839 580
rect 773 508 839 546
rect 773 474 789 508
rect 823 474 839 508
rect 773 440 839 474
rect 773 406 789 440
rect 823 406 839 440
rect 877 580 929 596
rect 877 546 890 580
rect 924 546 929 580
rect 877 497 929 546
rect 877 463 890 497
rect 924 463 929 497
rect 877 414 929 463
rect 683 372 736 380
rect 877 380 890 414
rect 924 380 929 414
rect 966 580 1032 649
rect 966 546 982 580
rect 1016 546 1032 580
rect 966 508 1032 546
rect 966 474 982 508
rect 1016 474 1032 508
rect 966 440 1032 474
rect 966 406 982 440
rect 1016 406 1032 440
rect 877 372 929 380
rect 323 338 1031 372
rect 255 288 903 304
rect 255 254 309 288
rect 343 254 377 288
rect 411 254 445 288
rect 479 254 513 288
rect 547 254 581 288
rect 615 254 649 288
rect 683 254 717 288
rect 751 254 785 288
rect 819 254 853 288
rect 887 254 903 288
rect 255 238 903 254
rect 255 230 289 238
rect 123 196 289 230
rect 942 236 1031 338
rect 942 204 976 236
rect 23 133 89 162
rect 23 99 39 133
rect 73 99 89 133
rect 23 17 89 99
rect 123 133 189 196
rect 323 170 976 204
rect 123 99 139 133
rect 173 99 189 133
rect 123 70 189 99
rect 223 133 289 162
rect 223 99 239 133
rect 273 99 289 133
rect 223 17 289 99
rect 323 133 389 170
rect 323 99 339 133
rect 373 99 389 133
rect 323 70 389 99
rect 423 120 489 136
rect 423 86 439 120
rect 473 86 489 120
rect 423 17 489 86
rect 523 133 573 170
rect 523 99 539 133
rect 523 70 573 99
rect 609 120 675 136
rect 609 86 625 120
rect 659 86 675 120
rect 609 17 675 86
rect 711 133 745 170
rect 711 70 745 99
rect 781 120 861 136
rect 781 86 804 120
rect 838 86 861 120
rect 781 17 861 86
rect 897 133 931 170
rect 897 70 931 99
rect 967 120 1033 136
rect 967 86 983 120
rect 1017 86 1033 120
rect 967 17 1033 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 683 1056 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 0 617 1056 649
rect 0 17 1056 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -49 1056 -17
<< labels >>
rlabel comment s 0 0 0 0 4 clkbuf_8
flabel pwell s 0 0 1056 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew
flabel nwell s 0 617 1056 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew
flabel metal1 s 0 617 1056 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew
flabel metal1 s 0 0 1056 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew
flabel corelocali s 991 242 1025 276 0 FreeSans 340 0 0 0 X
port 6 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 X
port 6 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 1056 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3405152
string GDS_START 3396410
<< end >>
