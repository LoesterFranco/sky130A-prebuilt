magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 89 53 119 137
rect 278 53 308 137
rect 362 53 392 137
rect 480 47 510 177
rect 612 47 642 177
<< pmoshvt >>
rect 81 297 117 381
rect 282 297 318 381
rect 364 297 400 381
rect 472 297 508 497
rect 604 297 640 497
<< ndiff >>
rect 417 137 480 177
rect 27 106 89 137
rect 27 72 35 106
rect 69 72 89 106
rect 27 53 89 72
rect 119 97 278 137
rect 119 63 129 97
rect 163 63 224 97
rect 258 63 278 97
rect 119 53 278 63
rect 308 111 362 137
rect 308 77 318 111
rect 352 77 362 111
rect 308 53 362 77
rect 392 97 480 137
rect 392 63 422 97
rect 456 63 480 97
rect 392 53 480 63
rect 417 47 480 53
rect 510 135 612 177
rect 510 101 558 135
rect 592 101 612 135
rect 510 47 612 101
rect 642 162 699 177
rect 642 128 657 162
rect 691 128 699 162
rect 642 94 699 128
rect 642 60 657 94
rect 691 60 699 94
rect 642 47 699 60
<< pdiff >>
rect 417 485 472 497
rect 417 451 425 485
rect 459 451 472 485
rect 417 417 472 451
rect 417 383 425 417
rect 459 383 472 417
rect 417 381 472 383
rect 27 349 81 381
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 343 171 381
rect 117 309 129 343
rect 163 309 171 343
rect 117 297 171 309
rect 228 354 282 381
rect 228 320 236 354
rect 270 320 282 354
rect 228 297 282 320
rect 318 297 364 381
rect 400 297 472 381
rect 508 454 604 497
rect 508 420 558 454
rect 592 420 604 454
rect 508 386 604 420
rect 508 352 558 386
rect 592 352 604 386
rect 508 297 604 352
rect 640 483 699 497
rect 640 449 657 483
rect 691 449 699 483
rect 640 415 699 449
rect 640 381 657 415
rect 691 381 699 415
rect 640 347 699 381
rect 640 313 657 347
rect 691 313 699 347
rect 640 297 699 313
<< ndiffc >>
rect 35 72 69 106
rect 129 63 163 97
rect 224 63 258 97
rect 318 77 352 111
rect 422 63 456 97
rect 558 101 592 135
rect 657 128 691 162
rect 657 60 691 94
<< pdiffc >>
rect 425 451 459 485
rect 425 383 459 417
rect 35 315 69 349
rect 129 309 163 343
rect 236 320 270 354
rect 558 420 592 454
rect 558 352 592 386
rect 657 449 691 483
rect 657 381 691 415
rect 657 313 691 347
<< poly >>
rect 472 497 508 523
rect 604 497 640 523
rect 178 473 402 483
rect 178 439 194 473
rect 228 453 402 473
rect 228 439 244 453
rect 178 429 244 439
rect 362 407 402 453
rect 81 381 117 407
rect 282 381 318 407
rect 364 381 400 407
rect 81 282 117 297
rect 282 282 318 297
rect 364 282 400 297
rect 472 282 508 297
rect 604 282 640 297
rect 79 265 119 282
rect 280 265 320 282
rect 21 249 119 265
rect 21 215 35 249
rect 69 215 119 249
rect 21 199 119 215
rect 226 249 320 265
rect 226 215 236 249
rect 270 215 320 249
rect 226 199 320 215
rect 89 137 119 199
rect 278 137 308 199
rect 362 192 402 282
rect 470 265 510 282
rect 602 265 642 282
rect 444 249 642 265
rect 444 215 454 249
rect 488 215 642 249
rect 444 199 642 215
rect 362 137 392 192
rect 480 177 510 199
rect 612 177 642 199
rect 89 27 119 53
rect 278 27 308 53
rect 362 27 392 53
rect 480 21 510 47
rect 612 21 642 47
<< polycont >>
rect 194 439 228 473
rect 35 215 69 249
rect 236 215 270 249
rect 454 215 488 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 17 349 69 527
rect 412 485 468 527
rect 108 473 366 483
rect 108 439 194 473
rect 228 439 366 473
rect 108 417 366 439
rect 412 451 425 485
rect 459 451 468 485
rect 412 417 468 451
rect 412 383 425 417
rect 459 383 468 417
rect 17 315 35 349
rect 17 299 69 315
rect 129 343 163 377
rect 129 265 163 309
rect 207 354 291 383
rect 412 367 468 383
rect 558 454 622 493
rect 592 420 622 454
rect 558 386 622 420
rect 207 320 236 354
rect 270 333 291 354
rect 592 352 622 386
rect 270 320 488 333
rect 207 299 488 320
rect 17 249 85 265
rect 17 215 35 249
rect 69 215 85 249
rect 129 249 276 265
rect 129 215 236 249
rect 270 215 276 249
rect 129 199 276 215
rect 454 249 488 299
rect 129 181 178 199
rect 21 147 178 181
rect 454 165 488 215
rect 21 106 84 147
rect 318 131 488 165
rect 558 135 622 352
rect 657 483 704 527
rect 691 449 704 483
rect 657 415 704 449
rect 691 381 704 415
rect 657 347 704 381
rect 691 313 704 347
rect 657 292 704 313
rect 21 72 35 106
rect 69 72 84 106
rect 21 53 84 72
rect 128 97 274 113
rect 128 63 129 97
rect 163 63 224 97
rect 258 63 274 97
rect 128 17 274 63
rect 318 111 352 131
rect 592 101 622 135
rect 318 61 352 77
rect 406 63 422 97
rect 456 63 472 97
rect 558 83 622 101
rect 657 162 704 185
rect 691 128 704 162
rect 657 94 704 128
rect 406 17 472 63
rect 691 60 704 94
rect 657 17 704 60
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel corelocali s 223 425 257 459 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 400 0 0 0 B_N
port 2 nsew
flabel corelocali s 577 357 611 391 0 FreeSans 400 0 0 0 X
port 7 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew
rlabel comment s 0 0 0 0 4 or2b_2
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 654648
string GDS_START 648880
<< end >>
