magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 121 492 171 596
rect 473 492 539 547
rect 873 492 923 547
rect 121 458 923 492
rect 21 260 87 356
rect 121 119 175 458
rect 217 390 681 424
rect 217 270 455 390
rect 504 270 570 356
rect 615 270 681 390
rect 729 390 1127 424
rect 729 270 795 390
rect 869 270 935 356
rect 985 270 1127 390
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 31 390 81 649
rect 211 526 339 649
rect 373 581 639 615
rect 373 526 439 581
rect 573 526 639 581
rect 673 526 739 649
rect 773 581 1029 615
rect 773 526 839 581
rect 963 458 1029 581
rect 1063 458 1129 649
rect 23 85 73 226
rect 211 202 656 236
rect 211 85 261 202
rect 23 51 261 85
rect 307 85 373 164
rect 409 119 443 202
rect 479 85 545 164
rect 579 119 656 202
rect 692 202 1129 236
rect 692 85 742 202
rect 307 51 742 85
rect 776 17 842 164
rect 876 81 942 202
rect 976 17 1042 164
rect 1078 81 1129 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
rlabel locali s 985 270 1127 390 6 A1
port 1 nsew signal input
rlabel locali s 729 390 1127 424 6 A1
port 1 nsew signal input
rlabel locali s 729 270 795 390 6 A1
port 1 nsew signal input
rlabel locali s 869 270 935 356 6 A2
port 2 nsew signal input
rlabel locali s 615 270 681 390 6 B1
port 3 nsew signal input
rlabel locali s 217 390 681 424 6 B1
port 3 nsew signal input
rlabel locali s 217 270 455 390 6 B1
port 3 nsew signal input
rlabel locali s 504 270 570 356 6 B2
port 4 nsew signal input
rlabel locali s 21 260 87 356 6 C1
port 5 nsew signal input
rlabel locali s 873 492 923 547 6 Y
port 6 nsew signal output
rlabel locali s 473 492 539 547 6 Y
port 6 nsew signal output
rlabel locali s 121 492 171 596 6 Y
port 6 nsew signal output
rlabel locali s 121 458 923 492 6 Y
port 6 nsew signal output
rlabel locali s 121 119 175 458 6 Y
port 6 nsew signal output
rlabel metal1 s 0 -49 1152 49 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1152 715 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1484032
string GDS_START 1473870
<< end >>
