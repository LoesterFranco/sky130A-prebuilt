magic
tech sky130A
magscale 1 2
timestamp 1601050047
<< nwell >>
rect -38 332 710 704
<< pwell >>
rect 0 0 672 49
<< scpmos >>
rect 108 368 138 592
rect 192 368 222 592
rect 306 368 336 592
rect 420 368 450 592
rect 534 368 564 592
<< nmoslvt >>
rect 98 74 128 222
rect 189 74 219 222
rect 339 74 369 222
rect 439 74 469 222
rect 531 74 561 222
<< ndiff >>
rect 27 210 98 222
rect 27 176 39 210
rect 73 176 98 210
rect 27 120 98 176
rect 27 86 39 120
rect 73 86 98 120
rect 27 74 98 86
rect 128 210 189 222
rect 128 176 139 210
rect 173 176 189 210
rect 128 120 189 176
rect 128 86 139 120
rect 173 86 189 120
rect 128 74 189 86
rect 219 120 339 222
rect 219 86 264 120
rect 298 86 339 120
rect 219 74 339 86
rect 369 202 439 222
rect 369 168 394 202
rect 428 168 439 202
rect 369 116 439 168
rect 369 82 394 116
rect 428 82 439 116
rect 369 74 439 82
rect 469 74 531 222
rect 561 202 618 222
rect 561 168 572 202
rect 606 168 618 202
rect 561 120 618 168
rect 561 86 572 120
rect 606 86 618 120
rect 561 74 618 86
<< pdiff >>
rect 49 580 108 592
rect 49 546 61 580
rect 95 546 108 580
rect 49 510 108 546
rect 49 476 61 510
rect 95 476 108 510
rect 49 440 108 476
rect 49 406 61 440
rect 95 406 108 440
rect 49 368 108 406
rect 138 368 192 592
rect 222 368 306 592
rect 336 580 420 592
rect 336 546 373 580
rect 407 546 420 580
rect 336 497 420 546
rect 336 463 373 497
rect 407 463 420 497
rect 336 414 420 463
rect 336 380 373 414
rect 407 380 420 414
rect 336 368 420 380
rect 450 582 534 592
rect 450 548 473 582
rect 507 548 534 582
rect 450 514 534 548
rect 450 480 473 514
rect 507 480 534 514
rect 450 446 534 480
rect 450 412 473 446
rect 507 412 534 446
rect 450 368 534 412
rect 564 580 623 592
rect 564 546 577 580
rect 611 546 623 580
rect 564 497 623 546
rect 564 463 577 497
rect 611 463 623 497
rect 564 414 623 463
rect 564 380 577 414
rect 611 380 623 414
rect 564 368 623 380
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 139 176 173 210
rect 139 86 173 120
rect 264 86 298 120
rect 394 168 428 202
rect 394 82 428 116
rect 572 168 606 202
rect 572 86 606 120
<< pdiffc >>
rect 61 546 95 580
rect 61 476 95 510
rect 61 406 95 440
rect 373 546 407 580
rect 373 463 407 497
rect 373 380 407 414
rect 473 548 507 582
rect 473 480 507 514
rect 473 412 507 446
rect 577 546 611 580
rect 577 463 611 497
rect 577 380 611 414
<< poly >>
rect 108 592 138 618
rect 192 592 222 618
rect 306 592 336 618
rect 420 592 450 618
rect 534 592 564 618
rect 108 353 138 368
rect 192 353 222 368
rect 306 353 336 368
rect 420 353 450 368
rect 534 353 564 368
rect 105 336 141 353
rect 75 320 141 336
rect 75 286 91 320
rect 125 286 141 320
rect 75 270 141 286
rect 189 336 225 353
rect 189 320 255 336
rect 189 286 205 320
rect 239 286 255 320
rect 189 270 255 286
rect 303 310 339 353
rect 417 310 453 353
rect 531 310 567 353
rect 303 294 369 310
rect 98 222 128 270
rect 189 222 219 270
rect 303 260 319 294
rect 353 260 369 294
rect 303 244 369 260
rect 417 294 483 310
rect 417 260 433 294
rect 467 260 483 294
rect 417 244 483 260
rect 531 294 651 310
rect 531 260 601 294
rect 635 260 651 294
rect 531 244 651 260
rect 339 222 369 244
rect 439 222 469 244
rect 531 222 561 244
rect 98 48 128 74
rect 189 48 219 74
rect 339 48 369 74
rect 439 48 469 74
rect 531 48 561 74
<< polycont >>
rect 91 286 125 320
rect 205 286 239 320
rect 319 260 353 294
rect 433 260 467 294
rect 601 260 635 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 45 580 111 649
rect 45 546 61 580
rect 95 546 111 580
rect 357 580 423 596
rect 45 510 111 546
rect 45 476 61 510
rect 95 476 111 510
rect 45 440 111 476
rect 45 406 61 440
rect 95 406 111 440
rect 45 390 111 406
rect 25 320 141 356
rect 25 286 91 320
rect 125 286 141 320
rect 25 270 141 286
rect 189 320 263 578
rect 357 546 373 580
rect 407 546 423 580
rect 357 497 423 546
rect 357 463 373 497
rect 407 463 423 497
rect 357 414 423 463
rect 357 380 373 414
rect 407 380 423 414
rect 457 582 523 649
rect 457 548 473 582
rect 507 548 523 582
rect 457 514 523 548
rect 457 480 473 514
rect 507 480 523 514
rect 457 446 523 480
rect 457 412 473 446
rect 507 412 523 446
rect 561 580 647 596
rect 561 546 577 580
rect 611 546 647 580
rect 561 497 647 546
rect 561 463 577 497
rect 611 463 647 497
rect 561 414 647 463
rect 357 378 423 380
rect 561 380 577 414
rect 611 380 647 414
rect 561 378 647 380
rect 357 344 647 378
rect 189 286 205 320
rect 239 286 263 320
rect 189 270 263 286
rect 303 294 369 310
rect 303 260 319 294
rect 353 260 369 294
rect 303 236 369 260
rect 409 294 483 310
rect 409 260 433 294
rect 467 260 483 294
rect 409 236 483 260
rect 23 210 89 226
rect 23 176 39 210
rect 73 176 89 210
rect 23 120 89 176
rect 23 86 39 120
rect 73 86 89 120
rect 23 17 89 86
rect 123 210 189 226
rect 123 176 139 210
rect 173 202 189 210
rect 517 202 551 344
rect 585 294 651 310
rect 585 260 601 294
rect 635 260 651 294
rect 585 236 651 260
rect 173 176 394 202
rect 123 168 394 176
rect 428 168 444 202
rect 123 120 189 168
rect 123 86 139 120
rect 173 86 189 120
rect 123 70 189 86
rect 223 120 335 130
rect 223 86 264 120
rect 298 86 335 120
rect 223 17 335 86
rect 378 116 444 168
rect 378 82 394 116
rect 428 82 444 116
rect 378 66 444 82
rect 517 168 572 202
rect 606 168 622 202
rect 517 120 622 168
rect 517 86 572 120
rect 606 86 622 120
rect 517 70 622 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o311ai_1
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 223 390 257 424 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 223 464 257 498 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 223 538 257 572 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 607 242 641 276 0 FreeSans 340 0 0 0 C1
port 5 nsew
flabel corelocali s 415 242 449 276 0 FreeSans 340 0 0 0 B1
port 4 nsew
flabel corelocali s 607 390 641 424 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 607 464 641 498 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 607 538 641 572 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 319 242 353 276 0 FreeSans 340 0 0 0 A3
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 672 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1352668
string GDS_START 1345892
<< end >>
