magic
tech sky130A
magscale 1 2
timestamp 1604502729
<< locali >>
rect 88 290 163 356
rect 197 339 263 430
rect 1177 360 1318 414
rect 1177 226 1223 360
rect 1645 364 1711 596
rect 1665 226 1699 364
rect 1177 170 1301 226
rect 1249 71 1301 170
rect 1649 70 1699 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 20 420 89 596
rect 130 464 196 649
rect 230 512 297 596
rect 472 546 538 649
rect 230 478 855 512
rect 230 464 331 478
rect 20 250 54 420
rect 297 305 331 464
rect 365 376 431 444
rect 646 410 787 444
rect 365 342 677 376
rect 227 252 377 305
rect 20 150 89 250
rect 227 184 293 252
rect 411 218 445 342
rect 339 184 445 218
rect 503 150 569 308
rect 20 116 569 150
rect 603 294 677 342
rect 603 101 637 294
rect 711 237 745 410
rect 821 350 855 478
rect 934 414 1016 649
rect 1050 482 1131 596
rect 1178 516 1228 649
rect 1342 516 1408 649
rect 1050 448 1391 482
rect 1050 378 1131 448
rect 779 284 855 350
rect 889 344 1131 378
rect 889 271 955 344
rect 997 237 1063 310
rect 711 211 1063 237
rect 671 203 1063 211
rect 671 145 814 203
rect 1097 169 1131 344
rect 1357 326 1391 448
rect 1257 260 1391 326
rect 1443 330 1509 596
rect 1555 364 1605 649
rect 1751 364 1801 649
rect 1443 264 1631 330
rect 1443 226 1503 264
rect 125 17 191 82
rect 457 17 528 82
rect 603 51 853 101
rect 926 17 1003 169
rect 1037 70 1131 169
rect 1165 17 1215 136
rect 1335 17 1401 226
rect 1437 90 1503 226
rect 1549 17 1615 226
rect 1735 17 1801 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
<< metal1 >>
rect 0 683 1824 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 0 617 1824 649
rect 0 17 1824 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
rect 0 -49 1824 -17
<< labels >>
rlabel locali s 88 290 163 356 6 D
port 1 nsew signal input
rlabel locali s 1249 71 1301 170 6 Q
port 2 nsew signal output
rlabel locali s 1177 360 1318 414 6 Q
port 2 nsew signal output
rlabel locali s 1177 226 1223 360 6 Q
port 2 nsew signal output
rlabel locali s 1177 170 1301 226 6 Q
port 2 nsew signal output
rlabel locali s 1665 226 1699 364 6 Q_N
port 3 nsew signal output
rlabel locali s 1649 70 1699 226 6 Q_N
port 3 nsew signal output
rlabel locali s 1645 364 1711 596 6 Q_N
port 3 nsew signal output
rlabel locali s 197 339 263 430 6 GATE_N
port 4 nsew clock input
rlabel metal1 s 0 -49 1824 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 617 1824 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1824 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 2215604
string GDS_START 2201770
<< end >>
