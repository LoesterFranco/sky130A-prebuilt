magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 17 197 66 325
rect 293 191 378 265
rect 1118 83 1175 491
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 35 393 69 493
rect 103 427 179 527
rect 35 359 166 393
rect 132 280 166 359
rect 223 337 268 493
rect 132 214 178 280
rect 132 161 166 214
rect 35 127 166 161
rect 35 69 69 127
rect 103 17 179 93
rect 223 69 257 337
rect 311 333 377 483
rect 421 367 484 527
rect 604 451 770 485
rect 311 299 458 333
rect 424 219 458 299
rect 534 271 591 401
rect 634 283 702 399
rect 424 157 508 219
rect 634 207 668 283
rect 327 153 508 157
rect 327 123 458 153
rect 577 141 668 207
rect 736 265 770 451
rect 810 427 870 527
rect 914 373 958 487
rect 814 307 958 373
rect 924 265 958 307
rect 1004 299 1058 527
rect 736 199 886 265
rect 924 199 1084 265
rect 327 69 361 123
rect 736 107 770 199
rect 924 165 958 199
rect 395 17 471 89
rect 601 73 770 107
rect 804 17 860 165
rect 914 83 958 165
rect 1004 17 1058 165
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< obsm1 >>
rect 222 388 280 397
rect 522 388 580 397
rect 222 360 580 388
rect 222 351 280 360
rect 522 351 580 360
rect 120 320 178 329
rect 623 320 681 329
rect 120 292 681 320
rect 120 283 178 292
rect 623 283 681 292
<< labels >>
rlabel locali s 293 191 378 265 6 D
port 1 nsew signal input
rlabel locali s 17 197 66 325 6 GATE_N
port 2 nsew signal input
rlabel locali s 1118 83 1175 491 6 Q
port 3 nsew signal output
rlabel metal1 s 0 -48 1196 48 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 496 1196 592 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1938136
string GDS_START 1928318
<< end >>
