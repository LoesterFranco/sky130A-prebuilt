magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 17 51 535 493
<< labels >>
rlabel locali s 17 51 535 493 6 DIODE
port 1 nsew signal input
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 552 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3603704
string GDS_START 3598642
<< end >>
