magic
tech sky130A
magscale 1 2
timestamp 1599588244
<< locali >>
rect 25 236 119 370
rect 1446 364 1519 596
rect 1273 270 1343 356
rect 1485 230 1519 364
rect 1447 78 1519 230
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 23 420 89 649
rect 129 420 189 596
rect 155 354 189 420
rect 225 557 291 596
rect 332 591 399 649
rect 433 557 594 597
rect 225 547 594 557
rect 628 569 808 603
rect 968 569 1034 649
rect 225 523 467 547
rect 225 388 291 523
rect 628 513 662 569
rect 1068 535 1305 540
rect 501 489 662 513
rect 416 479 662 489
rect 718 501 1305 535
rect 416 455 535 479
rect 416 388 466 455
rect 569 421 684 445
rect 503 411 684 421
rect 503 387 603 411
rect 155 220 233 354
rect 267 271 469 305
rect 155 202 189 220
rect 23 17 89 202
rect 123 84 189 202
rect 267 186 301 271
rect 235 81 301 186
rect 335 17 401 237
rect 435 185 469 271
rect 503 253 537 387
rect 718 377 752 501
rect 637 353 752 377
rect 571 343 752 353
rect 786 433 1125 467
rect 571 287 671 343
rect 786 309 820 433
rect 854 333 963 399
rect 705 255 820 309
rect 503 221 671 253
rect 503 219 879 221
rect 603 187 879 219
rect 435 153 569 185
rect 813 155 879 187
rect 435 151 779 153
rect 535 119 779 151
rect 913 150 963 333
rect 1075 234 1125 433
rect 1169 390 1305 501
rect 1346 390 1412 649
rect 1169 270 1235 390
rect 1201 234 1235 270
rect 1379 264 1451 330
rect 1075 184 1167 234
rect 1201 184 1282 234
rect 1379 150 1413 264
rect 435 85 501 117
rect 913 116 1413 150
rect 913 85 963 116
rect 435 51 963 85
rect 999 17 1065 82
rect 1318 17 1411 82
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
rlabel locali s 25 236 119 370 6 D
port 1 nsew signal input
rlabel locali s 1485 230 1519 364 6 Q
port 2 nsew signal output
rlabel locali s 1447 78 1519 230 6 Q
port 2 nsew signal output
rlabel locali s 1446 364 1519 596 6 Q
port 2 nsew signal output
rlabel locali s 1273 270 1343 356 6 GATE
port 3 nsew clock input
rlabel metal1 s 0 -49 1536 49 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 5 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 617 1536 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1536 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 2187520
string GDS_START 2176092
<< end >>
