magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 125 265 201 485
rect 313 288 379 493
rect 313 265 372 288
rect 125 199 372 265
rect 125 75 185 199
rect 313 185 372 199
rect 313 70 375 185
rect 649 215 772 265
rect 1631 289 1757 323
rect 1631 199 1675 289
rect 1815 215 1907 265
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 57 298 91 527
rect 245 299 279 527
rect 413 443 490 527
rect 526 447 840 481
rect 991 447 1057 527
rect 1144 455 1803 489
rect 1885 455 1962 527
rect 526 409 570 447
rect 1144 413 1178 455
rect 413 375 570 409
rect 638 379 1178 413
rect 413 265 457 375
rect 503 307 840 341
rect 406 199 457 265
rect 57 17 91 147
rect 245 17 279 147
rect 412 173 457 199
rect 412 139 547 173
rect 409 17 469 105
rect 503 85 547 139
rect 581 119 615 307
rect 806 265 840 307
rect 884 323 961 339
rect 884 305 927 323
rect 905 289 927 305
rect 905 275 961 289
rect 806 199 871 265
rect 675 159 751 181
rect 905 159 939 275
rect 995 241 1029 379
rect 1075 289 1179 343
rect 675 125 939 159
rect 973 207 1029 241
rect 973 91 1007 207
rect 1121 187 1179 289
rect 740 85 837 91
rect 503 51 837 85
rect 881 57 1007 91
rect 1041 17 1075 173
rect 1155 153 1179 187
rect 1121 83 1179 153
rect 1215 119 1249 421
rect 1283 165 1317 455
rect 2006 421 2065 493
rect 1363 323 1446 409
rect 1563 387 2065 421
rect 1363 289 1417 323
rect 1451 289 1529 323
rect 1366 199 1451 254
rect 1409 187 1451 199
rect 1283 131 1375 165
rect 1249 85 1304 97
rect 1215 53 1304 85
rect 1341 64 1375 131
rect 1409 153 1417 187
rect 1409 126 1451 153
rect 1495 85 1529 289
rect 1563 119 1597 387
rect 1958 375 2065 387
rect 1801 299 1975 341
rect 1941 265 1975 299
rect 1709 189 1771 255
rect 1941 199 1997 265
rect 1709 187 1750 189
rect 1709 153 1713 187
rect 1747 153 1750 187
rect 1941 181 1975 199
rect 1709 146 1750 153
rect 1817 150 1975 181
rect 1809 147 1975 150
rect 1809 119 1867 147
rect 1631 85 1734 93
rect 1495 51 1734 85
rect 1809 85 1815 119
rect 1849 85 1867 119
rect 2031 117 2065 375
rect 1809 59 1867 85
rect 1911 17 1945 113
rect 2005 51 2065 117
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 927 289 961 323
rect 1121 153 1155 187
rect 1417 289 1451 323
rect 1215 85 1249 119
rect 1417 153 1451 187
rect 1713 153 1747 187
rect 1815 85 1849 119
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
<< metal1 >>
rect 0 561 2116 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 0 496 2116 527
rect 0 17 2116 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
rect 0 -48 2116 -17
<< obsm1 >>
rect 915 323 973 329
rect 915 289 927 323
rect 961 320 973 323
rect 1405 323 1463 329
rect 1405 320 1417 323
rect 961 292 1417 320
rect 961 289 973 292
rect 915 283 973 289
rect 1405 289 1417 292
rect 1451 289 1463 323
rect 1405 283 1463 289
rect 1109 187 1167 193
rect 1109 153 1121 187
rect 1155 184 1167 187
rect 1405 187 1463 193
rect 1405 184 1417 187
rect 1155 156 1417 184
rect 1155 153 1167 156
rect 1109 147 1167 153
rect 1405 153 1417 156
rect 1451 184 1463 187
rect 1701 187 1759 193
rect 1701 184 1713 187
rect 1451 156 1713 184
rect 1451 153 1463 156
rect 1405 147 1463 153
rect 1701 153 1713 156
rect 1747 153 1759 187
rect 1701 147 1759 153
rect 1203 119 1263 125
rect 1203 85 1215 119
rect 1249 116 1263 119
rect 1803 119 1861 125
rect 1803 116 1815 119
rect 1249 88 1815 116
rect 1249 85 1263 88
rect 1203 79 1263 85
rect 1803 85 1815 88
rect 1849 85 1861 119
rect 1803 79 1861 85
<< labels >>
rlabel locali s 1815 215 1907 265 6 A
port 1 nsew signal input
rlabel locali s 1631 289 1757 323 6 B
port 2 nsew signal input
rlabel locali s 1631 199 1675 289 6 B
port 2 nsew signal input
rlabel locali s 649 215 772 265 6 C
port 3 nsew signal input
rlabel locali s 313 288 379 493 6 X
port 4 nsew signal output
rlabel locali s 313 265 372 288 6 X
port 4 nsew signal output
rlabel locali s 313 185 372 199 6 X
port 4 nsew signal output
rlabel locali s 313 70 375 185 6 X
port 4 nsew signal output
rlabel locali s 125 265 201 485 6 X
port 4 nsew signal output
rlabel locali s 125 199 372 265 6 X
port 4 nsew signal output
rlabel locali s 125 75 185 199 6 X
port 4 nsew signal output
rlabel metal1 s 0 -48 2116 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 2116 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2116 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 749920
string GDS_START 735998
<< end >>
