magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 335 2918 704
rect -38 332 825 335
rect 1117 332 2918 335
rect 1618 311 1956 332
<< pwell >>
rect 0 0 2880 49
<< scnmos >>
rect 84 74 114 158
rect 282 81 312 165
rect 360 81 390 165
rect 515 81 545 165
rect 593 81 623 165
rect 685 81 715 165
rect 904 119 934 267
rect 1014 119 1044 267
rect 1204 119 1234 203
rect 1290 119 1320 203
rect 1367 119 1397 203
rect 1445 119 1475 203
rect 1693 74 1723 222
rect 1794 74 1824 222
rect 2048 74 2078 158
rect 2126 74 2156 158
rect 2212 74 2242 158
rect 2284 74 2314 158
rect 2482 74 2512 202
rect 2680 74 2710 222
rect 2766 74 2796 222
<< pmoshvt >>
rect 86 464 116 592
rect 310 464 340 592
rect 394 464 424 592
rect 482 464 512 592
rect 592 464 622 592
rect 706 464 736 592
rect 914 392 944 592
rect 1004 392 1034 592
rect 1212 457 1242 541
rect 1302 457 1332 541
rect 1374 457 1404 541
rect 1464 457 1494 541
rect 1713 347 1743 547
rect 1837 366 1867 566
rect 2007 508 2037 592
rect 2085 508 2115 592
rect 2255 508 2285 592
rect 2345 508 2375 592
rect 2462 392 2492 592
rect 2664 368 2694 592
rect 2754 368 2784 592
<< ndiff >>
rect 845 180 904 267
rect 27 133 84 158
rect 27 99 39 133
rect 73 99 84 133
rect 27 74 84 99
rect 114 128 171 158
rect 114 94 125 128
rect 159 94 171 128
rect 114 74 171 94
rect 225 127 282 165
rect 225 93 237 127
rect 271 93 282 127
rect 225 81 282 93
rect 312 81 360 165
rect 390 153 515 165
rect 390 119 470 153
rect 504 119 515 153
rect 390 81 515 119
rect 545 81 593 165
rect 623 130 685 165
rect 623 96 638 130
rect 672 96 685 130
rect 623 81 685 96
rect 715 130 781 165
rect 715 96 735 130
rect 769 96 781 130
rect 835 150 904 180
rect 835 116 847 150
rect 881 119 904 150
rect 934 142 1014 267
rect 934 119 957 142
rect 881 116 889 119
rect 835 98 889 116
rect 715 81 781 96
rect 949 108 957 119
rect 991 119 1014 142
rect 1044 241 1097 267
rect 1044 207 1055 241
rect 1089 207 1097 241
rect 1044 173 1097 207
rect 1643 203 1693 222
rect 1044 139 1055 173
rect 1089 139 1097 173
rect 1044 119 1097 139
rect 1151 179 1204 203
rect 1151 145 1159 179
rect 1193 145 1204 179
rect 1151 119 1204 145
rect 1234 179 1290 203
rect 1234 145 1245 179
rect 1279 145 1290 179
rect 1234 119 1290 145
rect 1320 119 1367 203
rect 1397 119 1445 203
rect 1475 119 1693 203
rect 991 108 999 119
rect 949 90 999 108
rect 1491 82 1693 119
rect 1491 48 1502 82
rect 1536 74 1693 82
rect 1723 189 1794 222
rect 1723 155 1734 189
rect 1768 155 1794 189
rect 1723 74 1794 155
rect 1824 158 1874 222
rect 2623 210 2680 222
rect 1824 146 2048 158
rect 1824 112 1902 146
rect 1936 112 2003 146
rect 2037 112 2048 146
rect 1824 74 2048 112
rect 2078 74 2126 158
rect 2156 133 2212 158
rect 2156 99 2167 133
rect 2201 99 2212 133
rect 2156 74 2212 99
rect 2242 74 2284 158
rect 2314 133 2371 158
rect 2314 99 2325 133
rect 2359 99 2371 133
rect 2314 74 2371 99
rect 2425 120 2482 202
rect 2425 86 2437 120
rect 2471 86 2482 120
rect 2425 74 2482 86
rect 2512 190 2569 202
rect 2512 156 2523 190
rect 2557 156 2569 190
rect 2512 120 2569 156
rect 2512 86 2523 120
rect 2557 86 2569 120
rect 2512 74 2569 86
rect 2623 176 2635 210
rect 2669 176 2680 210
rect 2623 120 2680 176
rect 2623 86 2635 120
rect 2669 86 2680 120
rect 2623 74 2680 86
rect 2710 210 2766 222
rect 2710 176 2721 210
rect 2755 176 2766 210
rect 2710 120 2766 176
rect 2710 86 2721 120
rect 2755 86 2766 120
rect 2710 74 2766 86
rect 2796 210 2853 222
rect 2796 176 2807 210
rect 2841 176 2853 210
rect 2796 120 2853 176
rect 2796 86 2807 120
rect 2841 86 2853 120
rect 2796 74 2853 86
rect 1536 48 1549 74
rect 1491 36 1549 48
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 510 86 546
rect 27 476 39 510
rect 73 476 86 510
rect 27 464 86 476
rect 116 580 310 592
rect 116 546 139 580
rect 173 546 263 580
rect 297 546 310 580
rect 116 510 310 546
rect 116 476 139 510
rect 173 476 263 510
rect 297 476 310 510
rect 116 464 310 476
rect 340 464 394 592
rect 424 584 482 592
rect 424 550 435 584
rect 469 550 482 584
rect 424 512 482 550
rect 424 478 435 512
rect 469 478 482 512
rect 424 464 482 478
rect 512 464 592 592
rect 622 580 706 592
rect 622 546 635 580
rect 669 546 706 580
rect 622 464 706 546
rect 736 580 795 592
rect 736 546 749 580
rect 783 546 795 580
rect 736 512 795 546
rect 736 478 749 512
rect 783 478 795 512
rect 736 464 795 478
rect 855 434 914 592
rect 855 400 867 434
rect 901 400 914 434
rect 855 392 914 400
rect 944 584 1004 592
rect 944 550 957 584
rect 991 550 1004 584
rect 944 392 1004 550
rect 1034 443 1093 592
rect 1034 409 1047 443
rect 1081 409 1093 443
rect 1034 392 1093 409
rect 1948 566 2007 592
rect 1761 547 1837 566
rect 1153 516 1212 541
rect 1153 482 1165 516
rect 1199 482 1212 516
rect 1153 457 1212 482
rect 1242 528 1302 541
rect 1242 494 1255 528
rect 1289 494 1302 528
rect 1242 457 1302 494
rect 1332 457 1374 541
rect 1404 533 1464 541
rect 1404 499 1417 533
rect 1451 499 1464 533
rect 1404 457 1464 499
rect 1494 523 1553 541
rect 1494 489 1507 523
rect 1541 489 1553 523
rect 1494 457 1553 489
rect 1654 502 1713 547
rect 1654 468 1666 502
rect 1700 468 1713 502
rect 1654 347 1713 468
rect 1743 535 1837 547
rect 1743 501 1773 535
rect 1807 501 1837 535
rect 1743 464 1837 501
rect 1743 430 1773 464
rect 1807 430 1837 464
rect 1743 393 1837 430
rect 1743 359 1773 393
rect 1807 366 1837 393
rect 1867 554 2007 566
rect 1867 520 1880 554
rect 1914 520 1960 554
rect 1994 520 2007 554
rect 1867 508 2007 520
rect 2037 508 2085 592
rect 2115 580 2255 592
rect 2115 546 2128 580
rect 2162 546 2198 580
rect 2232 546 2255 580
rect 2115 508 2255 546
rect 2285 567 2345 592
rect 2285 533 2298 567
rect 2332 533 2345 567
rect 2285 508 2345 533
rect 2375 580 2462 592
rect 2375 546 2405 580
rect 2439 546 2462 580
rect 2375 509 2462 546
rect 2375 508 2405 509
rect 1867 486 1925 508
rect 1867 452 1880 486
rect 1914 452 1925 486
rect 1867 418 1925 452
rect 1867 384 1880 418
rect 1914 384 1925 418
rect 1867 366 1925 384
rect 1807 359 1819 366
rect 1743 347 1819 359
rect 2393 475 2405 508
rect 2439 475 2462 509
rect 2393 438 2462 475
rect 2393 404 2405 438
rect 2439 404 2462 438
rect 2393 392 2462 404
rect 2492 580 2551 592
rect 2492 546 2505 580
rect 2539 546 2551 580
rect 2492 509 2551 546
rect 2492 475 2505 509
rect 2539 475 2551 509
rect 2492 438 2551 475
rect 2492 404 2505 438
rect 2539 404 2551 438
rect 2492 392 2551 404
rect 2605 580 2664 592
rect 2605 546 2617 580
rect 2651 546 2664 580
rect 2605 497 2664 546
rect 2605 463 2617 497
rect 2651 463 2664 497
rect 2605 414 2664 463
rect 2605 380 2617 414
rect 2651 380 2664 414
rect 2605 368 2664 380
rect 2694 580 2754 592
rect 2694 546 2707 580
rect 2741 546 2754 580
rect 2694 497 2754 546
rect 2694 463 2707 497
rect 2741 463 2754 497
rect 2694 414 2754 463
rect 2694 380 2707 414
rect 2741 380 2754 414
rect 2694 368 2754 380
rect 2784 580 2853 592
rect 2784 546 2807 580
rect 2841 546 2853 580
rect 2784 497 2853 546
rect 2784 463 2807 497
rect 2841 463 2853 497
rect 2784 414 2853 463
rect 2784 380 2807 414
rect 2841 380 2853 414
rect 2784 368 2853 380
<< ndiffc >>
rect 39 99 73 133
rect 125 94 159 128
rect 237 93 271 127
rect 470 119 504 153
rect 638 96 672 130
rect 735 96 769 130
rect 847 116 881 150
rect 957 108 991 142
rect 1055 207 1089 241
rect 1055 139 1089 173
rect 1159 145 1193 179
rect 1245 145 1279 179
rect 1502 48 1536 82
rect 1734 155 1768 189
rect 1902 112 1936 146
rect 2003 112 2037 146
rect 2167 99 2201 133
rect 2325 99 2359 133
rect 2437 86 2471 120
rect 2523 156 2557 190
rect 2523 86 2557 120
rect 2635 176 2669 210
rect 2635 86 2669 120
rect 2721 176 2755 210
rect 2721 86 2755 120
rect 2807 176 2841 210
rect 2807 86 2841 120
<< pdiffc >>
rect 39 546 73 580
rect 39 476 73 510
rect 139 546 173 580
rect 263 546 297 580
rect 139 476 173 510
rect 263 476 297 510
rect 435 550 469 584
rect 435 478 469 512
rect 635 546 669 580
rect 749 546 783 580
rect 749 478 783 512
rect 867 400 901 434
rect 957 550 991 584
rect 1047 409 1081 443
rect 1165 482 1199 516
rect 1255 494 1289 528
rect 1417 499 1451 533
rect 1507 489 1541 523
rect 1666 468 1700 502
rect 1773 501 1807 535
rect 1773 430 1807 464
rect 1773 359 1807 393
rect 1880 520 1914 554
rect 1960 520 1994 554
rect 2128 546 2162 580
rect 2198 546 2232 580
rect 2298 533 2332 567
rect 2405 546 2439 580
rect 1880 452 1914 486
rect 1880 384 1914 418
rect 2405 475 2439 509
rect 2405 404 2439 438
rect 2505 546 2539 580
rect 2505 475 2539 509
rect 2505 404 2539 438
rect 2617 546 2651 580
rect 2617 463 2651 497
rect 2617 380 2651 414
rect 2707 546 2741 580
rect 2707 463 2741 497
rect 2707 380 2741 414
rect 2807 546 2841 580
rect 2807 463 2841 497
rect 2807 380 2841 414
<< poly >>
rect 86 592 116 618
rect 310 592 340 618
rect 394 592 424 618
rect 482 592 512 618
rect 592 592 622 618
rect 706 592 736 618
rect 914 592 944 618
rect 1004 592 1034 618
rect 1108 615 1870 645
rect 86 449 116 464
rect 310 449 340 464
rect 394 449 424 464
rect 482 449 512 464
rect 592 449 622 464
rect 706 449 736 464
rect 83 367 119 449
rect 307 367 343 449
rect 83 351 343 367
rect 83 317 137 351
rect 171 317 205 351
rect 239 317 273 351
rect 307 317 343 351
rect 83 301 343 317
rect 84 158 114 301
rect 391 253 425 449
rect 479 432 515 449
rect 467 416 533 432
rect 467 382 483 416
rect 517 382 533 416
rect 467 366 533 382
rect 577 406 643 449
rect 577 372 593 406
rect 627 372 643 406
rect 577 338 643 372
rect 162 237 228 253
rect 162 203 178 237
rect 212 217 228 237
rect 354 237 425 253
rect 469 302 535 318
rect 469 268 485 302
rect 519 268 535 302
rect 577 304 593 338
rect 627 304 643 338
rect 577 288 643 304
rect 685 432 739 449
rect 685 416 823 432
rect 685 382 773 416
rect 807 382 823 416
rect 685 370 823 382
rect 914 377 944 392
rect 685 366 819 370
rect 469 252 535 268
rect 212 203 312 217
rect 162 187 312 203
rect 354 203 370 237
rect 404 203 425 237
rect 354 187 425 203
rect 505 210 535 252
rect 282 165 312 187
rect 360 165 390 187
rect 505 180 545 210
rect 515 165 545 180
rect 593 165 623 288
rect 685 165 715 366
rect 904 324 944 377
rect 1004 375 1034 392
rect 1108 375 1138 615
rect 1212 541 1242 567
rect 1302 541 1332 615
rect 1834 581 1870 615
rect 2007 592 2037 618
rect 2085 592 2115 618
rect 2255 592 2285 618
rect 2345 592 2375 618
rect 2462 592 2492 618
rect 2664 592 2694 618
rect 2754 592 2784 618
rect 1374 541 1404 567
rect 1464 541 1494 567
rect 1713 547 1743 573
rect 1837 566 1867 581
rect 1212 442 1242 457
rect 1209 375 1245 442
rect 1302 431 1332 457
rect 757 308 944 324
rect 757 274 773 308
rect 807 282 944 308
rect 990 344 1142 375
rect 990 310 1006 344
rect 1040 310 1142 344
rect 990 282 1142 310
rect 1184 359 1250 375
rect 1374 361 1404 457
rect 1464 442 1494 457
rect 1464 429 1542 442
rect 1464 409 1605 429
rect 1464 403 1555 409
rect 1504 375 1555 403
rect 1589 375 1605 409
rect 1184 325 1200 359
rect 1234 345 1250 359
rect 1367 345 1462 361
rect 1234 325 1320 345
rect 1184 309 1320 325
rect 807 274 823 282
rect 757 240 823 274
rect 904 267 934 282
rect 1014 267 1044 282
rect 1112 267 1142 282
rect 757 206 773 240
rect 807 206 823 240
rect 757 190 823 206
rect 904 93 934 119
rect 1112 223 1234 267
rect 1204 203 1234 223
rect 1290 203 1320 309
rect 1367 311 1412 345
rect 1446 311 1462 345
rect 1367 295 1462 311
rect 1504 359 1605 375
rect 1367 203 1397 295
rect 1504 253 1534 359
rect 2007 493 2037 508
rect 2085 493 2115 508
rect 2255 493 2285 508
rect 2345 493 2375 508
rect 2004 466 2040 493
rect 1957 450 2040 466
rect 1957 416 1973 450
rect 2007 416 2040 450
rect 2082 476 2118 493
rect 2082 460 2170 476
rect 2082 446 2120 460
rect 1957 400 2040 416
rect 2088 426 2120 446
rect 2154 426 2170 460
rect 2252 447 2288 493
rect 2088 392 2170 426
rect 2222 431 2288 447
rect 2222 411 2238 431
rect 1837 351 1867 366
rect 2088 358 2120 392
rect 2154 358 2170 392
rect 1713 332 1743 347
rect 1834 345 1870 351
rect 1710 315 1746 332
rect 1834 315 2040 345
rect 1445 223 1534 253
rect 1618 299 1746 315
rect 1618 265 1634 299
rect 1668 285 1746 299
rect 1668 265 1723 285
rect 1618 249 1723 265
rect 1445 203 1475 223
rect 1693 222 1723 249
rect 1794 251 1962 267
rect 1794 237 1912 251
rect 1794 222 1824 237
rect 1014 93 1044 119
rect 1204 93 1234 119
rect 1290 93 1320 119
rect 1367 93 1397 119
rect 84 48 114 74
rect 282 55 312 81
rect 360 55 390 81
rect 515 55 545 81
rect 593 55 623 81
rect 685 51 715 81
rect 1445 51 1475 119
rect 685 21 1475 51
rect 1896 217 1912 237
rect 1946 217 1962 251
rect 1896 201 1962 217
rect 2010 226 2040 315
rect 2088 324 2170 358
rect 2088 290 2120 324
rect 2154 290 2170 324
rect 2088 274 2170 290
rect 2212 397 2238 411
rect 2272 397 2288 431
rect 2212 381 2288 397
rect 2010 196 2078 226
rect 2048 158 2078 196
rect 2126 158 2156 274
rect 2212 158 2242 381
rect 2342 333 2378 493
rect 2462 377 2492 392
rect 2348 285 2378 333
rect 2459 285 2495 377
rect 2664 353 2694 368
rect 2754 353 2784 368
rect 2661 326 2697 353
rect 2751 326 2787 353
rect 2312 269 2495 285
rect 2312 249 2328 269
rect 2284 235 2328 249
rect 2362 249 2495 269
rect 2605 310 2787 326
rect 2605 276 2621 310
rect 2655 290 2787 310
rect 2655 276 2796 290
rect 2605 260 2796 276
rect 2362 235 2512 249
rect 2284 219 2512 235
rect 2680 222 2710 260
rect 2766 222 2796 260
rect 2284 158 2314 219
rect 2482 202 2512 219
rect 1693 48 1723 74
rect 1794 48 1824 74
rect 2048 48 2078 74
rect 2126 48 2156 74
rect 2212 48 2242 74
rect 2284 48 2314 74
rect 2482 48 2512 74
rect 2680 48 2710 74
rect 2766 48 2796 74
<< polycont >>
rect 137 317 171 351
rect 205 317 239 351
rect 273 317 307 351
rect 483 382 517 416
rect 593 372 627 406
rect 178 203 212 237
rect 485 268 519 302
rect 593 304 627 338
rect 773 382 807 416
rect 370 203 404 237
rect 773 274 807 308
rect 1006 310 1040 344
rect 1555 375 1589 409
rect 1200 325 1234 359
rect 773 206 807 240
rect 1412 311 1446 345
rect 1973 416 2007 450
rect 2120 426 2154 460
rect 2120 358 2154 392
rect 1634 265 1668 299
rect 1912 217 1946 251
rect 2120 290 2154 324
rect 2238 397 2272 431
rect 2328 235 2362 269
rect 2621 276 2655 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2880 683
rect 23 580 89 596
rect 23 546 39 580
rect 73 546 89 580
rect 23 510 89 546
rect 23 476 39 510
rect 73 476 89 510
rect 23 435 89 476
rect 123 580 313 649
rect 123 546 139 580
rect 173 546 263 580
rect 297 546 313 580
rect 123 510 313 546
rect 123 476 139 510
rect 173 476 263 510
rect 297 476 313 510
rect 123 469 313 476
rect 419 584 485 596
rect 419 550 435 584
rect 469 550 485 584
rect 419 512 485 550
rect 619 580 685 649
rect 619 546 635 580
rect 669 546 685 580
rect 619 537 685 546
rect 723 580 799 596
rect 723 546 749 580
rect 783 546 799 580
rect 941 584 1007 649
rect 941 550 957 584
rect 991 550 1007 584
rect 419 478 435 512
rect 469 503 485 512
rect 723 524 799 546
rect 723 520 916 524
rect 723 518 922 520
rect 723 517 926 518
rect 723 516 929 517
rect 1165 516 1215 545
rect 723 512 1165 516
rect 723 503 749 512
rect 469 478 749 503
rect 783 484 1165 512
rect 783 480 850 484
rect 911 483 1165 484
rect 914 482 1165 483
rect 1199 482 1215 516
rect 918 480 1215 482
rect 783 478 846 480
rect 419 477 846 478
rect 923 477 1215 480
rect 1250 528 1371 545
rect 1250 494 1255 528
rect 1289 494 1371 528
rect 1250 477 1371 494
rect 419 469 757 477
rect 689 466 757 469
rect 23 416 541 435
rect 23 401 483 416
rect 23 253 57 401
rect 475 382 483 401
rect 517 382 541 416
rect 575 406 655 435
rect 575 400 593 406
rect 91 351 441 367
rect 475 366 541 382
rect 589 372 593 400
rect 627 372 655 406
rect 91 317 137 351
rect 171 317 205 351
rect 239 317 273 351
rect 307 332 441 351
rect 589 338 655 372
rect 307 317 541 332
rect 91 302 541 317
rect 91 298 485 302
rect 475 268 485 298
rect 519 268 541 302
rect 589 304 593 338
rect 627 304 655 338
rect 589 288 655 304
rect 23 237 228 253
rect 23 203 178 237
rect 212 203 228 237
rect 23 187 228 203
rect 313 237 420 253
rect 475 252 541 268
rect 689 254 723 466
rect 867 439 901 450
rect 1165 443 1215 477
rect 784 432 833 438
rect 757 424 833 432
rect 757 416 799 424
rect 757 382 773 416
rect 807 382 833 390
rect 757 366 833 382
rect 867 434 997 439
rect 901 400 997 434
rect 867 364 997 400
rect 1031 409 1047 443
rect 1081 409 1126 443
rect 1165 409 1303 443
rect 1031 391 1126 409
rect 963 355 997 364
rect 1090 375 1126 391
rect 1090 359 1235 375
rect 963 344 1056 355
rect 313 203 370 237
rect 404 203 420 237
rect 23 133 73 187
rect 313 162 420 203
rect 575 187 723 254
rect 571 182 723 187
rect 757 308 929 326
rect 757 274 773 308
rect 807 274 929 308
rect 757 252 929 274
rect 963 310 1006 344
rect 1040 310 1056 344
rect 963 291 1056 310
rect 1090 325 1200 359
rect 1234 325 1235 359
rect 1090 309 1235 325
rect 757 240 839 252
rect 757 206 773 240
rect 807 236 839 240
rect 807 206 812 236
rect 963 216 1009 291
rect 1090 257 1126 309
rect 1269 274 1303 409
rect 757 184 812 206
rect 878 187 1009 216
rect 874 182 1009 187
rect 568 180 723 182
rect 568 178 622 180
rect 871 178 1009 182
rect 566 176 622 178
rect 869 176 1009 178
rect 1043 241 1126 257
rect 1043 207 1055 241
rect 1089 214 1126 241
rect 1160 240 1303 274
rect 1337 433 1371 477
rect 1405 533 1453 649
rect 1405 499 1417 533
rect 1451 499 1453 533
rect 1405 469 1453 499
rect 1487 523 1553 549
rect 1487 489 1507 523
rect 1541 489 1553 523
rect 1487 464 1553 489
rect 1649 502 1716 649
rect 2112 580 2248 649
rect 1864 554 2078 570
rect 1649 468 1666 502
rect 1700 468 1716 502
rect 1649 466 1716 468
rect 1750 535 1823 551
rect 1750 501 1773 535
rect 1807 501 1823 535
rect 1750 464 1823 501
rect 1487 433 1521 464
rect 1337 397 1521 433
rect 1750 430 1773 464
rect 1807 430 1823 464
rect 1089 207 1124 214
rect 562 173 617 176
rect 865 173 925 176
rect 557 171 613 173
rect 860 172 925 173
rect 1043 173 1124 207
rect 1160 199 1195 240
rect 1337 206 1371 397
rect 557 169 611 171
rect 860 169 920 172
rect 23 99 39 133
rect 23 70 73 99
rect 109 128 175 153
rect 109 94 125 128
rect 159 94 175 128
rect 109 17 175 94
rect 221 127 287 128
rect 221 93 237 127
rect 271 93 287 127
rect 321 119 420 162
rect 454 167 611 169
rect 846 167 916 169
rect 454 162 608 167
rect 846 163 914 167
rect 454 153 604 162
rect 454 119 470 153
rect 504 119 604 153
rect 846 158 911 163
rect 846 150 907 158
rect 638 130 686 146
rect 221 85 287 93
rect 672 96 686 130
rect 638 85 686 96
rect 221 51 686 85
rect 722 130 776 146
rect 722 96 735 130
rect 769 96 776 130
rect 827 116 847 150
rect 881 116 907 150
rect 827 100 907 116
rect 941 108 957 142
rect 991 108 1007 142
rect 722 17 776 96
rect 941 17 1007 108
rect 1043 139 1055 173
rect 1089 139 1124 173
rect 1043 85 1124 139
rect 1159 179 1195 199
rect 1193 145 1195 179
rect 1159 119 1195 145
rect 1229 179 1371 206
rect 1405 345 1453 361
rect 1405 311 1412 345
rect 1446 311 1453 345
rect 1405 218 1453 311
rect 1487 309 1521 397
rect 1555 424 1714 430
rect 1555 409 1663 424
rect 1589 390 1663 409
rect 1697 390 1714 424
rect 1589 375 1714 390
rect 1555 359 1714 375
rect 1750 393 1823 430
rect 1750 359 1773 393
rect 1807 359 1823 393
rect 1864 520 1880 554
rect 1914 520 1960 554
rect 1994 520 2078 554
rect 2112 546 2128 580
rect 2162 546 2198 580
rect 2232 546 2248 580
rect 2282 567 2348 596
rect 1864 504 2078 520
rect 2282 533 2298 567
rect 2332 533 2348 567
rect 2282 512 2348 533
rect 1864 486 1920 504
rect 1864 452 1880 486
rect 1914 452 1920 486
rect 1864 418 1920 452
rect 1864 384 1880 418
rect 1914 384 1920 418
rect 1864 368 1920 384
rect 1957 450 2010 466
rect 1957 416 1973 450
rect 2007 416 2010 450
rect 1750 343 1823 359
rect 1487 299 1697 309
rect 1487 265 1634 299
rect 1668 265 1697 299
rect 1487 252 1697 265
rect 1750 218 1784 343
rect 1957 267 2010 416
rect 1405 189 1784 218
rect 1405 184 1734 189
rect 1229 145 1245 179
rect 1279 172 1371 179
rect 1279 145 1294 172
rect 1654 155 1734 184
rect 1768 155 1784 189
rect 1229 119 1294 145
rect 1410 116 1620 150
rect 1654 119 1784 155
rect 1818 251 2010 267
rect 1818 217 1912 251
rect 1946 217 2010 251
rect 1818 201 2010 217
rect 2044 240 2078 504
rect 2112 478 2348 512
rect 2389 580 2455 649
rect 2389 546 2405 580
rect 2439 546 2455 580
rect 2389 509 2455 546
rect 2112 460 2170 478
rect 2112 426 2120 460
rect 2154 426 2170 460
rect 2389 475 2405 509
rect 2439 475 2455 509
rect 2112 392 2170 426
rect 2112 358 2120 392
rect 2154 358 2170 392
rect 2222 431 2288 444
rect 2222 397 2238 431
rect 2272 424 2288 431
rect 2222 390 2239 397
rect 2273 390 2288 424
rect 2222 384 2288 390
rect 2389 438 2455 475
rect 2389 404 2405 438
rect 2439 404 2455 438
rect 2389 388 2455 404
rect 2489 580 2555 596
rect 2489 546 2505 580
rect 2539 546 2555 580
rect 2489 509 2555 546
rect 2489 475 2505 509
rect 2539 475 2555 509
rect 2489 438 2555 475
rect 2489 404 2505 438
rect 2539 404 2555 438
rect 2489 388 2555 404
rect 2112 350 2170 358
rect 2112 324 2446 350
rect 2112 290 2120 324
rect 2154 316 2446 324
rect 2154 290 2170 316
rect 2112 274 2170 290
rect 2204 269 2378 282
rect 2204 240 2328 269
rect 2044 235 2328 240
rect 2362 235 2378 269
rect 2044 222 2378 235
rect 2044 206 2238 222
rect 1410 85 1444 116
rect 1043 51 1444 85
rect 1586 85 1620 116
rect 1818 85 1852 201
rect 2044 162 2078 206
rect 2412 188 2446 316
rect 1886 146 2078 162
rect 1886 112 1902 146
rect 1936 112 2003 146
rect 2037 112 2078 146
rect 1886 96 2078 112
rect 2151 133 2217 162
rect 2151 99 2167 133
rect 2201 99 2217 133
rect 1486 48 1502 82
rect 1536 48 1552 82
rect 1586 51 1852 85
rect 1486 17 1552 48
rect 2151 17 2217 99
rect 2309 154 2446 188
rect 2521 326 2555 388
rect 2601 580 2667 649
rect 2601 546 2617 580
rect 2651 546 2667 580
rect 2601 497 2667 546
rect 2601 463 2617 497
rect 2651 463 2667 497
rect 2601 414 2667 463
rect 2601 380 2617 414
rect 2651 380 2667 414
rect 2601 364 2667 380
rect 2705 580 2757 596
rect 2705 546 2707 580
rect 2741 546 2757 580
rect 2705 497 2757 546
rect 2705 463 2707 497
rect 2741 463 2757 497
rect 2705 414 2757 463
rect 2705 380 2707 414
rect 2741 380 2757 414
rect 2521 310 2671 326
rect 2521 276 2621 310
rect 2655 276 2671 310
rect 2521 260 2671 276
rect 2705 282 2757 380
rect 2791 580 2857 649
rect 2791 546 2807 580
rect 2841 546 2857 580
rect 2791 497 2857 546
rect 2791 463 2807 497
rect 2841 463 2857 497
rect 2791 414 2857 463
rect 2791 380 2807 414
rect 2841 380 2857 414
rect 2791 364 2857 380
rect 2521 190 2573 260
rect 2521 156 2523 190
rect 2557 156 2573 190
rect 2309 133 2375 154
rect 2309 99 2325 133
rect 2359 99 2375 133
rect 2521 120 2573 156
rect 2309 70 2375 99
rect 2421 86 2437 120
rect 2471 86 2487 120
rect 2421 17 2487 86
rect 2521 86 2523 120
rect 2557 86 2573 120
rect 2521 70 2573 86
rect 2619 210 2669 226
rect 2619 176 2635 210
rect 2619 120 2669 176
rect 2619 86 2635 120
rect 2619 17 2669 86
rect 2705 210 2771 282
rect 2705 176 2721 210
rect 2755 176 2771 210
rect 2705 120 2771 176
rect 2705 86 2721 120
rect 2755 86 2771 120
rect 2705 70 2771 86
rect 2807 210 2857 226
rect 2841 176 2857 210
rect 2807 120 2857 176
rect 2841 86 2857 120
rect 2807 17 2857 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2880 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 799 416 833 424
rect 799 390 807 416
rect 807 390 833 416
rect 1663 390 1697 424
rect 2239 397 2272 424
rect 2272 397 2273 424
rect 2239 390 2273 397
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
<< metal1 >>
rect 0 683 2880 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2880 683
rect 0 617 2880 649
rect 787 424 845 430
rect 787 390 799 424
rect 833 421 845 424
rect 1651 424 1709 430
rect 1651 421 1663 424
rect 833 393 1663 421
rect 833 390 845 393
rect 787 384 845 390
rect 1651 390 1663 393
rect 1697 421 1709 424
rect 2227 424 2285 430
rect 2227 421 2239 424
rect 1697 393 2239 421
rect 1697 390 1709 393
rect 1651 384 1709 390
rect 2227 390 2239 393
rect 2273 390 2285 424
rect 2227 384 2285 390
rect 0 17 2880 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2880 17
rect 0 -49 2880 -17
<< labels >>
flabel comment s 1063 36 1063 36 0 FreeSans 300 0 0 0 no_jumper_check
flabel comment s 1503 630 1503 630 0 FreeSans 300 0 0 0 no_jumper_check
rlabel comment s 0 0 0 0 4 sdfrtp_2
flabel pwell s 0 0 2880 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nwell s 0 617 2880 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 2239 390 2273 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew
flabel metal1 s 0 617 2880 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 2880 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 319 168 353 202 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 SCD
port 4 nsew
flabel corelocali s 607 390 641 424 0 FreeSans 340 0 0 0 SCD
port 4 nsew
flabel corelocali s 799 242 833 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 2719 94 2753 128 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2719 168 2753 202 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2719 242 2753 276 0 FreeSans 340 0 0 0 Q
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 2880 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 184708
string GDS_START 162290
<< end >>
