magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 517 333 583 425
rect 695 333 771 493
rect 925 333 993 493
rect 517 299 993 333
rect 18 211 262 265
rect 300 211 484 265
rect 540 211 711 265
rect 815 119 891 299
rect 926 151 994 265
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 18 333 89 493
rect 133 367 167 527
rect 201 333 277 493
rect 321 459 661 493
rect 321 367 355 459
rect 389 333 465 425
rect 18 299 465 333
rect 627 367 661 459
rect 815 367 881 527
rect 18 143 771 177
rect 18 51 89 143
rect 133 17 167 109
rect 201 51 277 143
rect 321 17 433 109
rect 485 51 551 143
rect 585 17 661 109
rect 695 85 771 143
rect 926 85 993 117
rect 695 51 993 85
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
rlabel locali s 18 211 262 265 6 A1
port 1 nsew signal input
rlabel locali s 300 211 484 265 6 A2
port 2 nsew signal input
rlabel locali s 540 211 711 265 6 A3
port 3 nsew signal input
rlabel locali s 926 151 994 265 6 B1
port 4 nsew signal input
rlabel locali s 925 333 993 493 6 Y
port 5 nsew signal output
rlabel locali s 815 119 891 299 6 Y
port 5 nsew signal output
rlabel locali s 695 333 771 493 6 Y
port 5 nsew signal output
rlabel locali s 517 333 583 425 6 Y
port 5 nsew signal output
rlabel locali s 517 299 993 333 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -48 1012 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 1012 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1012 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 559036
string GDS_START 549708
<< end >>
