magic
tech sky130A
magscale 1 2
timestamp 1599588218
<< nwell >>
rect -38 332 1286 704
<< pwell >>
rect 0 0 1248 49
<< scpmos >>
rect 85 368 121 592
rect 183 368 219 592
rect 307 368 343 592
rect 473 368 509 592
rect 705 368 741 592
rect 795 368 831 592
rect 922 368 958 592
rect 1012 368 1048 592
rect 1129 368 1165 568
<< nmoslvt >>
rect 85 74 115 222
rect 189 74 219 222
rect 307 74 337 222
rect 479 74 509 222
rect 705 98 735 246
rect 801 98 831 246
rect 922 98 952 246
rect 1018 98 1048 246
rect 1134 118 1164 246
<< ndiff >>
rect 352 222 410 233
rect 28 202 85 222
rect 28 168 40 202
rect 74 168 85 202
rect 28 120 85 168
rect 28 86 40 120
rect 74 86 85 120
rect 28 74 85 86
rect 115 177 189 222
rect 115 143 144 177
rect 178 143 189 177
rect 115 74 189 143
rect 219 85 307 222
rect 219 74 246 85
rect 234 51 246 74
rect 280 74 307 85
rect 337 221 479 222
rect 337 187 364 221
rect 398 187 479 221
rect 337 74 479 187
rect 509 116 578 222
rect 509 82 532 116
rect 566 82 578 116
rect 509 74 578 82
rect 632 98 705 246
rect 735 234 801 246
rect 735 200 751 234
rect 785 200 801 234
rect 735 98 801 200
rect 831 98 922 246
rect 952 150 1018 246
rect 952 116 968 150
rect 1002 116 1018 150
rect 952 98 1018 116
rect 1048 148 1134 246
rect 1048 114 1073 148
rect 1107 118 1134 148
rect 1164 232 1221 246
rect 1164 198 1175 232
rect 1209 198 1221 232
rect 1164 164 1221 198
rect 1164 130 1175 164
rect 1209 130 1221 164
rect 1164 118 1221 130
rect 1107 114 1119 118
rect 1048 98 1119 114
rect 632 82 690 98
rect 280 51 292 74
rect 234 39 292 51
rect 632 48 644 82
rect 678 48 690 82
rect 846 82 907 98
rect 632 36 690 48
rect 846 48 859 82
rect 893 48 907 82
rect 846 36 907 48
<< pdiff >>
rect 619 627 690 639
rect 619 593 637 627
rect 671 593 690 627
rect 619 592 690 593
rect 846 616 907 632
rect 846 592 859 616
rect 27 580 85 592
rect 27 546 39 580
rect 73 546 85 580
rect 27 497 85 546
rect 27 463 39 497
rect 73 463 85 497
rect 27 414 85 463
rect 27 380 39 414
rect 73 380 85 414
rect 27 368 85 380
rect 121 580 183 592
rect 121 546 139 580
rect 173 546 183 580
rect 121 491 183 546
rect 121 457 139 491
rect 173 457 183 491
rect 121 368 183 457
rect 219 423 307 592
rect 219 389 246 423
rect 280 389 307 423
rect 219 368 307 389
rect 343 575 473 592
rect 343 541 353 575
rect 387 541 429 575
rect 463 541 473 575
rect 343 368 473 541
rect 509 423 565 592
rect 509 389 519 423
rect 553 389 565 423
rect 509 368 565 389
rect 619 368 705 592
rect 741 452 795 592
rect 741 418 751 452
rect 785 418 795 452
rect 741 368 795 418
rect 831 582 859 592
rect 893 592 907 616
rect 893 582 922 592
rect 831 368 922 582
rect 958 580 1012 592
rect 958 546 968 580
rect 1002 546 1012 580
rect 958 470 1012 546
rect 958 436 968 470
rect 1002 436 1012 470
rect 958 368 1012 436
rect 1048 580 1114 592
rect 1048 546 1068 580
rect 1102 568 1114 580
rect 1102 546 1129 568
rect 1048 470 1129 546
rect 1048 436 1068 470
rect 1102 436 1129 470
rect 1048 368 1129 436
rect 1165 556 1221 568
rect 1165 522 1175 556
rect 1209 522 1221 556
rect 1165 470 1221 522
rect 1165 436 1175 470
rect 1209 436 1221 470
rect 1165 368 1221 436
<< ndiffc >>
rect 40 168 74 202
rect 40 86 74 120
rect 144 143 178 177
rect 246 51 280 85
rect 364 187 398 221
rect 532 82 566 116
rect 751 200 785 234
rect 968 116 1002 150
rect 1073 114 1107 148
rect 1175 198 1209 232
rect 1175 130 1209 164
rect 644 48 678 82
rect 859 48 893 82
<< pdiffc >>
rect 637 593 671 627
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 139 546 173 580
rect 139 457 173 491
rect 246 389 280 423
rect 353 541 387 575
rect 429 541 463 575
rect 519 389 553 423
rect 751 418 785 452
rect 859 582 893 616
rect 968 546 1002 580
rect 968 436 1002 470
rect 1068 546 1102 580
rect 1068 436 1102 470
rect 1175 522 1209 556
rect 1175 436 1209 470
<< poly >>
rect 85 592 121 618
rect 183 592 219 618
rect 307 592 343 618
rect 473 592 509 618
rect 705 592 741 618
rect 795 592 831 618
rect 922 592 958 618
rect 1012 592 1048 618
rect 1129 568 1165 594
rect 85 310 121 368
rect 183 310 219 368
rect 85 294 219 310
rect 85 260 101 294
rect 135 260 169 294
rect 203 260 219 294
rect 85 244 219 260
rect 85 222 115 244
rect 189 222 219 244
rect 307 336 343 368
rect 473 336 509 368
rect 307 320 509 336
rect 307 286 323 320
rect 357 286 391 320
rect 425 286 459 320
rect 493 286 509 320
rect 307 270 509 286
rect 307 222 337 270
rect 479 222 509 270
rect 705 336 741 368
rect 795 336 831 368
rect 705 320 839 336
rect 705 286 721 320
rect 755 286 789 320
rect 823 286 839 320
rect 705 270 839 286
rect 922 334 958 368
rect 1012 334 1048 368
rect 1129 336 1165 368
rect 922 318 1048 334
rect 922 284 998 318
rect 1032 284 1048 318
rect 705 246 735 270
rect 801 246 831 270
rect 922 268 1048 284
rect 1096 320 1165 336
rect 1096 286 1112 320
rect 1146 286 1165 320
rect 1096 270 1165 286
rect 922 246 952 268
rect 1018 246 1048 268
rect 1134 246 1164 270
rect 85 48 115 74
rect 189 48 219 74
rect 307 48 337 74
rect 479 48 509 74
rect 705 72 735 98
rect 801 72 831 98
rect 922 72 952 98
rect 1018 72 1048 98
rect 1134 92 1164 118
<< polycont >>
rect 101 260 135 294
rect 169 260 203 294
rect 323 286 357 320
rect 391 286 425 320
rect 459 286 493 320
rect 721 286 755 320
rect 789 286 823 320
rect 998 284 1032 318
rect 1112 286 1146 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 615 627 694 649
rect 17 580 89 596
rect 17 546 39 580
rect 73 546 89 580
rect 17 497 89 546
rect 17 463 39 497
rect 73 463 89 497
rect 17 423 89 463
rect 123 580 189 596
rect 615 593 637 627
rect 671 593 694 627
rect 842 616 911 649
rect 123 546 139 580
rect 173 546 189 580
rect 123 491 189 546
rect 337 575 479 591
rect 337 541 353 575
rect 387 541 429 575
rect 463 559 479 575
rect 842 582 859 616
rect 893 582 911 616
rect 842 570 911 582
rect 952 580 1018 596
rect 463 541 705 559
rect 337 536 705 541
rect 952 546 968 580
rect 1002 546 1018 580
rect 952 536 1018 546
rect 337 525 1018 536
rect 671 502 1018 525
rect 123 457 139 491
rect 173 468 637 491
rect 952 470 1018 502
rect 173 457 801 468
rect 603 452 801 457
rect 17 414 246 423
rect 17 380 39 414
rect 73 389 246 414
rect 280 389 519 423
rect 553 389 569 423
rect 603 418 751 452
rect 785 418 801 452
rect 952 436 968 470
rect 1002 436 1018 470
rect 1052 580 1118 649
rect 1052 546 1068 580
rect 1102 546 1118 580
rect 1052 470 1118 546
rect 1052 436 1068 470
rect 1102 436 1118 470
rect 1159 556 1230 572
rect 1159 522 1175 556
rect 1209 522 1230 556
rect 1159 470 1230 522
rect 1159 436 1175 470
rect 1209 436 1230 470
rect 603 402 801 418
rect 73 380 89 389
rect 17 364 89 380
rect 870 368 1162 402
rect 17 202 51 364
rect 307 320 647 355
rect 85 294 263 310
rect 85 260 101 294
rect 135 260 169 294
rect 203 260 263 294
rect 307 286 323 320
rect 357 286 391 320
rect 425 286 459 320
rect 493 286 647 320
rect 697 320 935 368
rect 697 286 721 320
rect 755 286 789 320
rect 823 286 935 320
rect 982 318 1048 334
rect 85 236 263 260
rect 982 284 998 318
rect 1032 284 1048 318
rect 348 234 806 252
rect 348 221 751 234
rect 17 168 40 202
rect 74 168 90 202
rect 17 120 90 168
rect 17 86 40 120
rect 74 86 90 120
rect 128 177 194 202
rect 348 187 364 221
rect 398 218 751 221
rect 398 187 414 218
rect 730 200 751 218
rect 785 200 806 234
rect 982 236 1048 284
rect 1096 320 1162 368
rect 1096 286 1112 320
rect 1146 286 1162 320
rect 1096 270 1162 286
rect 1196 236 1230 436
rect 982 232 1230 236
rect 982 202 1175 232
rect 1159 198 1175 202
rect 1209 198 1230 232
rect 128 143 144 177
rect 178 153 194 177
rect 448 166 650 184
rect 448 153 1023 166
rect 178 150 1023 153
rect 178 143 482 150
rect 128 119 482 143
rect 616 132 968 150
rect 947 116 968 132
rect 1002 116 1023 150
rect 17 85 90 86
rect 516 85 532 116
rect 17 51 246 85
rect 280 82 532 85
rect 566 82 582 116
rect 947 100 1023 116
rect 1057 148 1123 168
rect 1057 114 1073 148
rect 1107 114 1123 148
rect 1159 164 1230 198
rect 1159 130 1175 164
rect 1209 130 1230 164
rect 1159 114 1230 130
rect 280 51 582 82
rect 628 82 694 98
rect 628 48 644 82
rect 678 48 694 82
rect 628 17 694 48
rect 842 82 911 98
rect 842 48 859 82
rect 893 48 911 82
rect 842 17 911 48
rect 1057 17 1123 114
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
<< metal1 >>
rect 0 683 1248 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 0 617 1248 649
rect 0 17 1248 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
rect 0 -49 1248 -17
<< labels >>
flabel pwell s 0 0 1248 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 0 617 1248 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
rlabel comment s 0 0 0 0 4 mux2i_2
flabel metal1 s 0 617 1248 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 1248 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 127 242 161 276 0 FreeSans 340 0 0 0 A0
port 1 nsew
flabel corelocali s 223 242 257 276 0 FreeSans 340 0 0 0 A0
port 1 nsew
flabel corelocali s 31 390 65 424 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 31 464 65 498 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 31 538 65 572 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 S
port 3 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 S
port 3 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 S
port 3 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A1
port 2 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A1
port 2 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 A1
port 2 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 A1
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 1248 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1961614
string GDS_START 1952024
<< end >>
