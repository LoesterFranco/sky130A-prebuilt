magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1564 561
rect 19 383 85 527
rect 119 333 153 493
rect 187 383 253 527
rect 287 333 321 493
rect 355 383 421 527
rect 523 451 589 527
rect 711 451 777 527
rect 879 451 945 527
rect 24 299 321 333
rect 24 161 68 299
rect 442 215 621 259
rect 667 215 806 265
rect 856 215 1015 265
rect 24 127 321 161
rect 19 17 85 93
rect 119 51 153 127
rect 187 17 253 93
rect 287 51 321 127
rect 1126 215 1356 325
rect 1406 259 1445 327
rect 1406 215 1542 259
rect 355 17 421 93
rect 523 17 589 93
rect 1395 17 1461 93
rect 0 -17 1564 17
<< obsli1 >>
rect 455 417 489 493
rect 643 417 677 493
rect 811 417 845 493
rect 979 451 1545 485
rect 979 417 1013 451
rect 455 383 1013 417
rect 1227 415 1461 417
rect 1056 383 1461 415
rect 1056 381 1240 383
rect 1056 333 1090 381
rect 1495 351 1545 451
rect 360 299 1090 333
rect 360 265 394 299
rect 114 199 394 265
rect 455 131 777 165
rect 1056 161 1090 299
rect 455 51 489 131
rect 879 127 1285 161
rect 1327 129 1529 163
rect 1327 93 1361 129
rect 627 59 1029 93
rect 1134 59 1361 93
rect 1327 51 1361 59
rect 1495 51 1529 129
<< metal1 >>
rect 0 496 1564 592
rect 0 -48 1564 48
<< labels >>
rlabel locali s 856 215 1015 265 6 A1
port 1 nsew signal input
rlabel locali s 667 215 806 265 6 A2
port 2 nsew signal input
rlabel locali s 442 215 621 259 6 A3
port 3 nsew signal input
rlabel locali s 1126 215 1356 325 6 B1
port 4 nsew signal input
rlabel locali s 1406 259 1445 327 6 B2
port 5 nsew signal input
rlabel locali s 1406 215 1542 259 6 B2
port 5 nsew signal input
rlabel locali s 287 333 321 493 6 X
port 6 nsew signal output
rlabel locali s 287 51 321 127 6 X
port 6 nsew signal output
rlabel locali s 119 333 153 493 6 X
port 6 nsew signal output
rlabel locali s 119 51 153 127 6 X
port 6 nsew signal output
rlabel locali s 24 299 321 333 6 X
port 6 nsew signal output
rlabel locali s 24 161 68 299 6 X
port 6 nsew signal output
rlabel locali s 24 127 321 161 6 X
port 6 nsew signal output
rlabel locali s 1395 17 1461 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 523 17 589 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 355 17 421 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 187 17 253 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 19 17 85 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 1564 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1564 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 879 451 945 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 711 451 777 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 523 451 589 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 355 383 421 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 187 383 253 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 19 383 85 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 1564 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 1564 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1564 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3641330
string GDS_START 3629194
<< end >>
