magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 25 236 110 371
rect 505 270 573 356
rect 607 207 645 547
rect 679 236 745 310
rect 499 141 645 207
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 21 420 71 649
rect 111 420 178 596
rect 144 304 178 420
rect 216 424 266 596
rect 306 458 372 649
rect 412 581 747 615
rect 412 458 462 581
rect 501 424 567 547
rect 216 390 567 424
rect 216 364 266 390
rect 360 304 426 336
rect 144 270 426 304
rect 144 181 178 270
rect 23 17 73 181
rect 109 81 178 181
rect 221 202 455 236
rect 681 364 747 581
rect 221 70 287 202
rect 321 17 387 168
rect 421 104 455 202
rect 679 104 736 202
rect 421 70 736 104
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel locali s 505 270 573 356 6 A0
port 1 nsew signal input
rlabel locali s 679 236 745 310 6 A1
port 2 nsew signal input
rlabel locali s 25 236 110 371 6 S
port 3 nsew signal input
rlabel locali s 607 207 645 547 6 Y
port 4 nsew signal output
rlabel locali s 499 141 645 207 6 Y
port 4 nsew signal output
rlabel metal1 s 0 -49 768 49 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 617 768 715 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1606014
string GDS_START 1599034
<< end >>
