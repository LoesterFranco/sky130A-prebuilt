magic
tech sky130A
magscale 1 2
timestamp 1604502711
<< locali >>
rect 1223 325 1273 425
rect 1391 325 1441 425
rect 1223 291 1441 325
rect 79 215 361 257
rect 415 215 750 257
rect 797 215 1137 257
rect 1223 181 1293 291
rect 1562 215 1731 257
rect 103 145 1449 181
rect 103 51 169 145
rect 271 51 337 145
rect 439 51 505 145
rect 607 51 673 145
rect 879 51 945 145
rect 1047 51 1113 145
rect 1215 51 1281 145
rect 1383 51 1449 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 19 325 85 493
rect 119 359 161 527
rect 195 325 245 493
rect 279 359 329 527
rect 363 459 749 493
rect 363 325 413 459
rect 19 291 413 325
rect 447 325 497 425
rect 531 359 581 459
rect 615 325 665 425
rect 699 359 749 459
rect 803 459 1525 493
rect 803 359 853 459
rect 887 325 937 425
rect 971 359 1021 459
rect 1055 325 1105 425
rect 447 291 1105 325
rect 1139 291 1189 459
rect 1307 359 1357 459
rect 1475 359 1525 459
rect 1570 325 1637 493
rect 1494 291 1637 325
rect 1671 291 1717 527
rect 1494 257 1528 291
rect 1327 215 1528 257
rect 1494 181 1528 215
rect 35 17 69 179
rect 1494 147 1637 181
rect 203 17 237 111
rect 371 17 405 111
rect 539 17 573 111
rect 707 17 845 111
rect 979 17 1013 111
rect 1147 17 1181 111
rect 1315 17 1349 111
rect 1483 17 1517 111
rect 1562 51 1637 147
rect 1671 17 1717 181
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
<< metal1 >>
rect 0 561 1748 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 0 496 1748 527
rect 0 17 1748 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
rect 0 -48 1748 -17
<< labels >>
rlabel locali s 79 215 361 257 6 A
port 1 nsew signal input
rlabel locali s 415 215 750 257 6 B
port 2 nsew signal input
rlabel locali s 797 215 1137 257 6 C
port 3 nsew signal input
rlabel locali s 1562 215 1731 257 6 D_N
port 4 nsew signal input
rlabel locali s 1391 325 1441 425 6 Y
port 5 nsew signal output
rlabel locali s 1383 51 1449 145 6 Y
port 5 nsew signal output
rlabel locali s 1223 325 1273 425 6 Y
port 5 nsew signal output
rlabel locali s 1223 291 1441 325 6 Y
port 5 nsew signal output
rlabel locali s 1223 181 1293 291 6 Y
port 5 nsew signal output
rlabel locali s 1215 51 1281 145 6 Y
port 5 nsew signal output
rlabel locali s 1047 51 1113 145 6 Y
port 5 nsew signal output
rlabel locali s 879 51 945 145 6 Y
port 5 nsew signal output
rlabel locali s 607 51 673 145 6 Y
port 5 nsew signal output
rlabel locali s 439 51 505 145 6 Y
port 5 nsew signal output
rlabel locali s 271 51 337 145 6 Y
port 5 nsew signal output
rlabel locali s 103 145 1449 181 6 Y
port 5 nsew signal output
rlabel locali s 103 51 169 145 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -48 1748 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1748 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1748 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1191072
string GDS_START 1177578
<< end >>
