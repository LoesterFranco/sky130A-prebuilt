magic
tech sky130A
magscale 1 2
timestamp 1604502729
<< locali >>
rect 17 368 71 596
rect 17 234 51 368
rect 199 270 265 356
rect 17 88 89 234
rect 741 270 875 356
rect 1369 285 1441 356
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 111 458 161 649
rect 195 581 531 615
rect 195 424 229 581
rect 375 508 425 547
rect 465 542 531 581
rect 679 542 745 649
rect 898 581 1418 615
rect 898 542 964 581
rect 1003 508 1053 515
rect 123 390 229 424
rect 263 390 333 500
rect 375 474 1053 508
rect 375 390 425 474
rect 570 406 637 440
rect 123 334 157 390
rect 85 268 157 334
rect 299 350 333 390
rect 503 350 569 362
rect 299 316 569 350
rect 123 166 157 268
rect 299 234 333 316
rect 503 296 569 316
rect 227 200 333 234
rect 367 262 455 282
rect 603 262 637 406
rect 367 228 637 262
rect 123 132 333 166
rect 125 17 191 98
rect 299 85 333 132
rect 367 119 433 228
rect 671 194 705 474
rect 784 390 943 440
rect 909 337 943 390
rect 1003 371 1053 474
rect 1110 513 1318 547
rect 1110 421 1176 513
rect 1216 387 1250 479
rect 1087 353 1250 387
rect 909 271 1009 337
rect 1087 282 1121 353
rect 1284 319 1318 513
rect 1352 424 1418 581
rect 1452 458 1518 649
rect 1558 438 1615 586
rect 1352 390 1524 424
rect 909 236 943 271
rect 1063 237 1121 282
rect 781 202 943 236
rect 1004 236 1121 237
rect 1155 285 1318 319
rect 1483 351 1524 390
rect 1483 285 1533 351
rect 1004 203 1097 236
rect 467 85 533 194
rect 299 51 533 85
rect 567 168 705 194
rect 1155 187 1217 285
rect 1483 251 1524 285
rect 1567 251 1615 438
rect 567 153 1036 168
rect 1251 153 1307 242
rect 567 134 1307 153
rect 567 70 633 134
rect 1002 119 1307 134
rect 1341 217 1524 251
rect 679 17 745 100
rect 893 85 968 100
rect 1341 85 1407 217
rect 893 51 1407 85
rect 1441 17 1523 183
rect 1559 117 1615 251
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< obsm1 >>
rect 403 273 461 282
rect 1075 273 1133 282
rect 403 245 1133 273
rect 403 236 461 245
rect 1075 236 1133 245
rect 1171 273 1229 282
rect 1555 273 1613 282
rect 1171 245 1613 273
rect 1171 236 1229 245
rect 1555 236 1613 245
<< labels >>
rlabel locali s 1369 285 1441 356 6 A
port 1 nsew signal input
rlabel locali s 741 270 875 356 6 B
port 2 nsew signal input
rlabel locali s 199 270 265 356 6 C
port 3 nsew signal input
rlabel locali s 17 368 71 596 6 X
port 4 nsew signal output
rlabel locali s 17 234 51 368 6 X
port 4 nsew signal output
rlabel locali s 17 88 89 234 6 X
port 4 nsew signal output
rlabel metal1 s 0 -49 1632 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 617 1632 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 515290
string GDS_START 502742
<< end >>
