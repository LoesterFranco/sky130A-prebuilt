magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 920 561
rect 115 359 165 527
rect 283 325 333 425
rect 563 325 613 425
rect 283 289 613 325
rect 731 359 781 527
rect 40 215 197 257
rect 231 215 385 255
rect 419 181 468 289
rect 511 215 645 255
rect 679 215 833 257
rect 107 145 468 181
rect 107 129 173 145
rect 275 129 341 145
rect 571 17 605 111
rect 739 17 773 111
rect 0 -17 920 17
<< obsli1 >>
rect 30 325 81 493
rect 199 459 417 493
rect 199 325 249 459
rect 30 291 249 325
rect 367 359 417 459
rect 479 459 697 493
rect 479 359 529 459
rect 647 325 697 459
rect 815 325 866 493
rect 647 291 866 325
rect 18 95 73 181
rect 502 145 873 181
rect 502 95 536 145
rect 18 61 536 95
rect 639 51 705 145
rect 807 51 873 145
<< metal1 >>
rect 0 496 920 592
rect 0 -48 920 48
<< labels >>
rlabel locali s 679 215 833 257 6 A1
port 1 nsew signal input
rlabel locali s 511 215 645 255 6 A2
port 2 nsew signal input
rlabel locali s 40 215 197 257 6 B1
port 3 nsew signal input
rlabel locali s 231 215 385 255 6 B2
port 4 nsew signal input
rlabel locali s 563 325 613 425 6 Y
port 5 nsew signal output
rlabel locali s 419 181 468 289 6 Y
port 5 nsew signal output
rlabel locali s 283 325 333 425 6 Y
port 5 nsew signal output
rlabel locali s 283 289 613 325 6 Y
port 5 nsew signal output
rlabel locali s 275 129 341 145 6 Y
port 5 nsew signal output
rlabel locali s 107 145 468 181 6 Y
port 5 nsew signal output
rlabel locali s 107 129 173 145 6 Y
port 5 nsew signal output
rlabel locali s 739 17 773 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 571 17 605 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 920 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 920 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 731 359 781 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 115 359 165 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 920 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 920 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 920 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1501952
string GDS_START 1494076
<< end >>
