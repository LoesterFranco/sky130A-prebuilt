magic
tech sky130A
magscale 1 2
timestamp 1599588218
<< nwell >>
rect -38 332 1862 704
<< pwell >>
rect 0 0 1824 49
<< scpmos >>
rect 100 424 136 592
rect 200 424 236 592
rect 425 392 461 560
rect 532 392 568 592
rect 616 392 652 592
rect 781 392 817 476
rect 887 392 923 476
rect 1020 368 1056 592
rect 1222 368 1258 592
rect 1312 368 1348 592
rect 1413 392 1449 592
rect 1615 368 1651 592
rect 1705 368 1741 592
<< nmoslvt >>
rect 84 136 114 246
rect 202 98 232 246
rect 416 74 446 222
rect 539 79 569 207
rect 617 79 647 207
rect 809 123 839 207
rect 901 123 931 207
rect 1012 74 1042 222
rect 1210 74 1240 222
rect 1296 74 1326 222
rect 1412 94 1442 222
rect 1624 74 1654 222
rect 1710 74 1740 222
<< ndiff >>
rect 27 208 84 246
rect 27 174 39 208
rect 73 174 84 208
rect 27 136 84 174
rect 114 136 202 246
rect 129 98 202 136
rect 232 234 289 246
rect 232 200 243 234
rect 277 200 289 234
rect 232 98 289 200
rect 343 222 401 230
rect 343 218 416 222
rect 343 184 355 218
rect 389 184 416 218
rect 129 82 187 98
rect 129 48 141 82
rect 175 48 187 82
rect 343 74 416 184
rect 446 207 496 222
rect 962 207 1012 222
rect 446 82 539 207
rect 446 74 475 82
rect 461 48 475 74
rect 509 79 539 82
rect 569 79 617 207
rect 647 195 809 207
rect 647 161 687 195
rect 721 161 764 195
rect 798 161 809 195
rect 647 123 809 161
rect 839 123 901 207
rect 931 169 1012 207
rect 931 135 947 169
rect 981 135 1012 169
rect 931 123 1012 135
rect 647 79 697 123
rect 509 48 524 79
rect 129 36 187 48
rect 461 36 524 48
rect 962 74 1012 123
rect 1042 136 1099 222
rect 1042 102 1053 136
rect 1087 102 1099 136
rect 1042 74 1099 102
rect 1153 120 1210 222
rect 1153 86 1165 120
rect 1199 86 1210 120
rect 1153 74 1210 86
rect 1240 207 1296 222
rect 1240 173 1251 207
rect 1285 173 1296 207
rect 1240 121 1296 173
rect 1240 87 1251 121
rect 1285 87 1296 121
rect 1240 74 1296 87
rect 1326 210 1412 222
rect 1326 176 1351 210
rect 1385 176 1412 210
rect 1326 120 1412 176
rect 1326 86 1351 120
rect 1385 94 1412 120
rect 1442 210 1499 222
rect 1442 176 1453 210
rect 1487 176 1499 210
rect 1442 140 1499 176
rect 1442 106 1453 140
rect 1487 106 1499 140
rect 1442 94 1499 106
rect 1553 210 1624 222
rect 1553 176 1565 210
rect 1599 176 1624 210
rect 1553 120 1624 176
rect 1385 86 1397 94
rect 1326 74 1397 86
rect 1553 86 1565 120
rect 1599 86 1624 120
rect 1553 74 1624 86
rect 1654 210 1710 222
rect 1654 176 1665 210
rect 1699 176 1710 210
rect 1654 120 1710 176
rect 1654 86 1665 120
rect 1699 86 1710 120
rect 1654 74 1710 86
rect 1740 210 1797 222
rect 1740 176 1751 210
rect 1785 176 1797 210
rect 1740 120 1797 176
rect 1740 86 1751 120
rect 1785 86 1797 120
rect 1740 74 1797 86
<< pdiff >>
rect 27 580 100 592
rect 27 546 39 580
rect 73 546 100 580
rect 27 470 100 546
rect 27 436 39 470
rect 73 436 100 470
rect 27 424 100 436
rect 136 580 200 592
rect 136 546 146 580
rect 180 546 200 580
rect 136 498 200 546
rect 136 464 146 498
rect 180 464 200 498
rect 136 424 200 464
rect 236 580 292 592
rect 236 546 246 580
rect 280 546 292 580
rect 476 580 532 592
rect 476 560 488 580
rect 236 498 292 546
rect 236 464 246 498
rect 280 464 292 498
rect 236 424 292 464
rect 369 441 425 560
rect 369 407 381 441
rect 415 407 425 441
rect 369 392 425 407
rect 461 546 488 560
rect 522 546 532 580
rect 461 392 532 546
rect 568 392 616 592
rect 652 476 702 592
rect 938 584 1020 592
rect 938 550 958 584
rect 992 550 1020 584
rect 938 516 1020 550
rect 938 482 958 516
rect 992 482 1020 516
rect 938 476 1020 482
rect 652 444 781 476
rect 652 410 662 444
rect 696 410 737 444
rect 771 410 781 444
rect 652 392 781 410
rect 817 392 887 476
rect 923 448 1020 476
rect 923 414 958 448
rect 992 414 1020 448
rect 923 392 1020 414
rect 970 368 1020 392
rect 1056 580 1112 592
rect 1056 546 1066 580
rect 1100 546 1112 580
rect 1056 497 1112 546
rect 1056 463 1066 497
rect 1100 463 1112 497
rect 1056 414 1112 463
rect 1056 380 1066 414
rect 1100 380 1112 414
rect 1056 368 1112 380
rect 1166 573 1222 592
rect 1166 539 1178 573
rect 1212 539 1222 573
rect 1166 368 1222 539
rect 1258 414 1312 592
rect 1258 380 1268 414
rect 1302 380 1312 414
rect 1258 368 1312 380
rect 1348 573 1413 592
rect 1348 539 1358 573
rect 1392 539 1413 573
rect 1348 392 1413 539
rect 1449 580 1505 592
rect 1449 546 1459 580
rect 1493 546 1505 580
rect 1449 509 1505 546
rect 1449 475 1459 509
rect 1493 475 1505 509
rect 1449 438 1505 475
rect 1449 404 1459 438
rect 1493 404 1505 438
rect 1449 392 1505 404
rect 1559 580 1615 592
rect 1559 546 1571 580
rect 1605 546 1615 580
rect 1559 497 1615 546
rect 1559 463 1571 497
rect 1605 463 1615 497
rect 1559 414 1615 463
rect 1348 368 1398 392
rect 1559 380 1571 414
rect 1605 380 1615 414
rect 1559 368 1615 380
rect 1651 580 1705 592
rect 1651 546 1661 580
rect 1695 546 1705 580
rect 1651 497 1705 546
rect 1651 463 1661 497
rect 1695 463 1705 497
rect 1651 414 1705 463
rect 1651 380 1661 414
rect 1695 380 1705 414
rect 1651 368 1705 380
rect 1741 580 1797 592
rect 1741 546 1751 580
rect 1785 546 1797 580
rect 1741 497 1797 546
rect 1741 463 1751 497
rect 1785 463 1797 497
rect 1741 414 1797 463
rect 1741 380 1751 414
rect 1785 380 1797 414
rect 1741 368 1797 380
<< ndiffc >>
rect 39 174 73 208
rect 243 200 277 234
rect 355 184 389 218
rect 141 48 175 82
rect 475 48 509 82
rect 687 161 721 195
rect 764 161 798 195
rect 947 135 981 169
rect 1053 102 1087 136
rect 1165 86 1199 120
rect 1251 173 1285 207
rect 1251 87 1285 121
rect 1351 176 1385 210
rect 1351 86 1385 120
rect 1453 176 1487 210
rect 1453 106 1487 140
rect 1565 176 1599 210
rect 1565 86 1599 120
rect 1665 176 1699 210
rect 1665 86 1699 120
rect 1751 176 1785 210
rect 1751 86 1785 120
<< pdiffc >>
rect 39 546 73 580
rect 39 436 73 470
rect 146 546 180 580
rect 146 464 180 498
rect 246 546 280 580
rect 246 464 280 498
rect 381 407 415 441
rect 488 546 522 580
rect 958 550 992 584
rect 958 482 992 516
rect 662 410 696 444
rect 737 410 771 444
rect 958 414 992 448
rect 1066 546 1100 580
rect 1066 463 1100 497
rect 1066 380 1100 414
rect 1178 539 1212 573
rect 1268 380 1302 414
rect 1358 539 1392 573
rect 1459 546 1493 580
rect 1459 475 1493 509
rect 1459 404 1493 438
rect 1571 546 1605 580
rect 1571 463 1605 497
rect 1571 380 1605 414
rect 1661 546 1695 580
rect 1661 463 1695 497
rect 1661 380 1695 414
rect 1751 546 1785 580
rect 1751 463 1785 497
rect 1751 380 1785 414
<< poly >>
rect 100 592 136 618
rect 200 592 236 618
rect 532 592 568 618
rect 616 592 652 618
rect 1020 592 1056 618
rect 1222 592 1258 618
rect 1312 592 1348 618
rect 1413 592 1449 618
rect 1615 592 1651 618
rect 1705 592 1741 618
rect 425 560 461 586
rect 100 356 136 424
rect 200 392 236 424
rect 781 476 817 502
rect 887 476 923 502
rect 197 376 263 392
rect 84 340 154 356
rect 84 306 104 340
rect 138 306 154 340
rect 197 342 213 376
rect 247 342 263 376
rect 197 326 263 342
rect 425 358 461 392
rect 84 290 154 306
rect 84 246 114 290
rect 202 246 232 326
rect 311 302 377 318
rect 311 268 327 302
rect 361 282 377 302
rect 425 282 455 358
rect 532 310 568 392
rect 616 360 652 392
rect 611 344 677 360
rect 781 350 817 392
rect 611 310 627 344
rect 661 310 677 344
rect 361 268 455 282
rect 311 252 455 268
rect 503 294 569 310
rect 611 294 677 310
rect 731 334 845 350
rect 731 300 795 334
rect 829 300 845 334
rect 503 260 519 294
rect 553 260 569 294
rect 84 110 114 136
rect 416 222 446 252
rect 503 244 569 260
rect 731 284 845 300
rect 887 336 923 392
rect 887 320 955 336
rect 887 286 905 320
rect 939 286 955 320
rect 1020 310 1056 368
rect 1222 326 1258 368
rect 1312 326 1348 368
rect 1413 326 1449 392
rect 1615 330 1651 368
rect 1222 310 1449 326
rect 731 252 761 284
rect 887 270 955 286
rect 997 294 1063 310
rect 202 72 232 98
rect 539 207 569 244
rect 617 222 761 252
rect 617 207 647 222
rect 809 207 839 233
rect 901 207 931 270
rect 997 260 1013 294
rect 1047 260 1063 294
rect 1222 290 1273 310
rect 997 244 1063 260
rect 1210 276 1273 290
rect 1307 276 1341 310
rect 1375 276 1449 310
rect 1210 260 1449 276
rect 1497 329 1654 330
rect 1705 329 1741 368
rect 1497 314 1741 329
rect 1497 280 1513 314
rect 1547 280 1581 314
rect 1615 294 1741 314
rect 1615 280 1740 294
rect 1497 264 1740 280
rect 1012 222 1042 244
rect 1210 222 1240 260
rect 1296 222 1326 260
rect 1412 222 1442 260
rect 1624 222 1654 264
rect 1710 222 1740 264
rect 416 48 446 74
rect 809 101 839 123
rect 719 85 853 101
rect 901 97 931 123
rect 539 53 569 79
rect 617 53 647 79
rect 719 51 735 85
rect 769 51 803 85
rect 837 51 853 85
rect 719 35 853 51
rect 1012 48 1042 74
rect 1210 48 1240 74
rect 1296 48 1326 74
rect 1412 68 1442 94
rect 1624 48 1654 74
rect 1710 48 1740 74
<< polycont >>
rect 104 306 138 340
rect 213 342 247 376
rect 327 268 361 302
rect 627 310 661 344
rect 795 300 829 334
rect 519 260 553 294
rect 905 286 939 320
rect 1013 260 1047 294
rect 1273 276 1307 310
rect 1341 276 1375 310
rect 1513 280 1547 314
rect 1581 280 1615 314
rect 735 51 769 85
rect 803 51 837 85
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 20 580 89 596
rect 20 546 39 580
rect 73 546 89 580
rect 20 470 89 546
rect 20 436 39 470
rect 73 436 89 470
rect 130 580 196 649
rect 130 546 146 580
rect 180 546 196 580
rect 130 498 196 546
rect 130 464 146 498
rect 180 464 196 498
rect 230 580 297 596
rect 230 546 246 580
rect 280 546 297 580
rect 472 580 538 649
rect 472 546 488 580
rect 522 546 538 580
rect 934 584 1016 649
rect 934 550 958 584
rect 992 550 1016 584
rect 230 512 297 546
rect 934 516 1016 550
rect 230 498 855 512
rect 230 464 246 498
rect 280 478 855 498
rect 280 464 331 478
rect 20 420 89 436
rect 20 250 54 420
rect 197 376 263 430
rect 88 340 163 356
rect 88 306 104 340
rect 138 306 163 340
rect 197 342 213 376
rect 247 342 263 376
rect 197 339 263 342
rect 88 290 163 306
rect 297 305 331 464
rect 365 441 431 444
rect 365 407 381 441
rect 415 407 431 441
rect 646 410 662 444
rect 696 410 737 444
rect 771 410 787 444
rect 365 376 431 407
rect 365 344 677 376
rect 365 342 627 344
rect 227 302 377 305
rect 227 268 327 302
rect 361 268 377 302
rect 227 252 377 268
rect 20 208 89 250
rect 20 174 39 208
rect 73 174 89 208
rect 227 234 293 252
rect 227 200 243 234
rect 277 200 293 234
rect 411 218 445 342
rect 603 310 627 342
rect 661 310 677 344
rect 227 184 293 200
rect 339 184 355 218
rect 389 184 445 218
rect 503 294 569 308
rect 503 260 519 294
rect 553 260 569 294
rect 20 150 89 174
rect 503 150 569 260
rect 20 116 569 150
rect 603 294 677 310
rect 603 101 637 294
rect 711 237 745 410
rect 821 350 855 478
rect 934 482 958 516
rect 992 482 1016 516
rect 934 448 1016 482
rect 934 414 958 448
rect 992 414 1016 448
rect 1050 580 1131 596
rect 1050 546 1066 580
rect 1100 546 1131 580
rect 1050 497 1131 546
rect 1178 573 1228 649
rect 1212 539 1228 573
rect 1178 516 1228 539
rect 1342 573 1408 649
rect 1342 539 1358 573
rect 1392 539 1408 573
rect 1342 516 1408 539
rect 1443 580 1509 596
rect 1443 546 1459 580
rect 1493 546 1509 580
rect 1050 463 1066 497
rect 1100 482 1131 497
rect 1443 509 1509 546
rect 1100 463 1391 482
rect 1050 448 1391 463
rect 1050 414 1131 448
rect 1050 380 1066 414
rect 1100 380 1131 414
rect 1050 378 1131 380
rect 779 334 855 350
rect 779 300 795 334
rect 829 300 855 334
rect 779 284 855 300
rect 889 344 1131 378
rect 889 320 955 344
rect 889 286 905 320
rect 939 286 955 320
rect 889 271 955 286
rect 997 294 1063 310
rect 997 260 1013 294
rect 1047 260 1063 294
rect 997 237 1063 260
rect 711 211 1063 237
rect 671 203 1063 211
rect 671 195 814 203
rect 671 161 687 195
rect 721 161 764 195
rect 798 161 814 195
rect 1097 169 1131 344
rect 1177 380 1268 414
rect 1302 380 1318 414
rect 1177 360 1318 380
rect 1177 226 1223 360
rect 1357 326 1391 448
rect 1257 310 1391 326
rect 1257 276 1273 310
rect 1307 276 1341 310
rect 1375 276 1391 310
rect 1257 260 1391 276
rect 1443 475 1459 509
rect 1493 475 1509 509
rect 1443 438 1509 475
rect 1443 404 1459 438
rect 1493 404 1509 438
rect 1443 330 1509 404
rect 1555 580 1605 649
rect 1555 546 1571 580
rect 1555 497 1605 546
rect 1555 463 1571 497
rect 1555 414 1605 463
rect 1555 380 1571 414
rect 1555 364 1605 380
rect 1645 580 1711 596
rect 1645 546 1661 580
rect 1695 546 1711 580
rect 1645 497 1711 546
rect 1645 463 1661 497
rect 1695 463 1711 497
rect 1645 414 1711 463
rect 1645 380 1661 414
rect 1695 380 1711 414
rect 1645 364 1711 380
rect 1751 580 1801 649
rect 1785 546 1801 580
rect 1751 497 1801 546
rect 1785 463 1801 497
rect 1751 414 1801 463
rect 1785 380 1801 414
rect 1751 364 1801 380
rect 1443 314 1631 330
rect 1443 280 1513 314
rect 1547 280 1581 314
rect 1615 280 1631 314
rect 1443 264 1631 280
rect 1443 226 1503 264
rect 1665 226 1699 364
rect 1177 207 1301 226
rect 1177 173 1251 207
rect 1285 173 1301 207
rect 1177 170 1301 173
rect 671 145 814 161
rect 926 135 947 169
rect 981 135 1003 169
rect 603 85 853 101
rect 125 48 141 82
rect 175 48 191 82
rect 125 17 191 48
rect 457 48 475 82
rect 509 48 528 82
rect 603 51 735 85
rect 769 51 803 85
rect 837 51 853 85
rect 457 17 528 48
rect 926 17 1003 135
rect 1037 136 1131 169
rect 1037 102 1053 136
rect 1087 102 1131 136
rect 1037 70 1131 102
rect 1165 120 1215 136
rect 1199 86 1215 120
rect 1165 17 1215 86
rect 1249 121 1301 170
rect 1249 87 1251 121
rect 1285 87 1301 121
rect 1249 71 1301 87
rect 1335 210 1401 226
rect 1335 176 1351 210
rect 1385 176 1401 210
rect 1335 120 1401 176
rect 1335 86 1351 120
rect 1385 86 1401 120
rect 1437 210 1503 226
rect 1437 176 1453 210
rect 1487 176 1503 210
rect 1437 140 1503 176
rect 1437 106 1453 140
rect 1487 106 1503 140
rect 1437 90 1503 106
rect 1549 210 1615 226
rect 1549 176 1565 210
rect 1599 176 1615 210
rect 1549 120 1615 176
rect 1335 17 1401 86
rect 1549 86 1565 120
rect 1599 86 1615 120
rect 1549 17 1615 86
rect 1649 210 1699 226
rect 1649 176 1665 210
rect 1649 120 1699 176
rect 1649 86 1665 120
rect 1649 70 1699 86
rect 1735 210 1801 226
rect 1735 176 1751 210
rect 1785 176 1801 210
rect 1735 120 1801 176
rect 1735 86 1751 120
rect 1785 86 1801 120
rect 1735 17 1801 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
<< metal1 >>
rect 0 683 1824 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 0 617 1824 649
rect 0 17 1824 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
rect 0 -49 1824 -17
<< labels >>
flabel pwell s 0 0 1824 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nwell s 0 617 1824 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
rlabel comment s 0 0 0 0 4 dlxbn_2
flabel metal1 s 0 617 1824 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 1824 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 1 nsew
flabel corelocali s 223 390 257 424 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew
flabel corelocali s 1183 242 1217 276 0 FreeSans 340 0 0 0 Q
port 7 nsew
flabel corelocali s 1183 316 1217 350 0 FreeSans 340 0 0 0 Q
port 7 nsew
flabel corelocali s 1663 390 1697 424 0 FreeSans 340 0 0 0 Q_N
port 8 nsew
flabel corelocali s 1663 464 1697 498 0 FreeSans 340 0 0 0 Q_N
port 8 nsew
flabel corelocali s 1663 538 1697 572 0 FreeSans 340 0 0 0 Q_N
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 1824 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 2156788
string GDS_START 2143354
<< end >>
