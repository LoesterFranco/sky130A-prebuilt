magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1840 561
rect 103 451 169 527
rect 30 195 66 349
rect 202 289 279 323
rect 245 257 279 289
rect 168 153 248 219
rect 520 411 566 527
rect 103 17 169 93
rect 205 79 248 153
rect 483 203 524 264
rect 449 143 524 203
rect 558 143 616 264
rect 491 17 557 109
rect 952 401 1021 527
rect 950 143 1024 279
rect 960 17 1026 109
rect 1404 367 1438 527
rect 1472 367 1554 491
rect 1226 249 1294 329
rect 1492 299 1554 367
rect 1588 299 1638 527
rect 1328 215 1390 265
rect 1308 199 1390 215
rect 1520 261 1554 299
rect 1672 261 1737 491
rect 1771 299 1821 527
rect 1520 213 1737 261
rect 1308 75 1370 199
rect 1404 17 1454 163
rect 1520 145 1554 213
rect 1488 53 1554 145
rect 1588 17 1638 177
rect 1672 53 1737 213
rect 1771 17 1821 177
rect 0 -17 1840 17
<< obsli1 >>
rect 27 417 69 475
rect 283 425 398 459
rect 432 425 449 459
rect 27 391 134 417
rect 27 383 306 391
rect 100 357 306 383
rect 340 357 381 391
rect 100 161 134 357
rect 313 315 381 357
rect 27 127 134 161
rect 313 207 347 315
rect 415 281 449 425
rect 662 425 674 459
rect 708 425 765 459
rect 595 357 664 391
rect 715 362 765 425
rect 630 332 664 357
rect 630 298 684 332
rect 27 69 69 127
rect 282 141 347 207
rect 381 247 449 281
rect 650 278 684 298
rect 381 107 415 247
rect 650 212 697 278
rect 295 73 415 107
rect 650 93 684 212
rect 731 135 765 362
rect 598 59 684 93
rect 718 69 765 135
rect 799 425 858 459
rect 892 425 904 459
rect 799 69 837 425
rect 1066 431 1256 465
rect 880 347 918 379
rect 1066 347 1100 431
rect 1306 425 1318 459
rect 1352 425 1370 459
rect 880 313 1100 347
rect 880 117 914 313
rect 880 51 921 117
rect 1066 93 1100 313
rect 1134 391 1192 397
rect 1168 357 1192 391
rect 1134 207 1192 357
rect 1336 333 1370 425
rect 1336 299 1458 333
rect 1424 265 1458 299
rect 1134 141 1258 207
rect 1424 199 1486 265
rect 1066 59 1245 93
<< obsli1c >>
rect 398 425 432 459
rect 306 357 340 391
rect 674 425 708 459
rect 858 425 892 459
rect 1318 425 1352 459
rect 1134 357 1168 391
<< metal1 >>
rect 0 496 1840 592
rect 17 320 76 329
rect 202 320 260 329
rect 1214 320 1272 329
rect 17 292 1272 320
rect 17 283 76 292
rect 202 283 260 292
rect 1214 283 1272 292
rect 0 -48 1840 48
<< obsm1 >>
rect 386 459 444 465
rect 386 425 398 459
rect 432 456 444 459
rect 662 459 720 465
rect 662 456 674 459
rect 432 428 674 456
rect 432 425 444 428
rect 386 419 444 425
rect 662 425 674 428
rect 708 425 720 459
rect 662 419 720 425
rect 846 459 904 465
rect 846 425 858 459
rect 892 456 904 459
rect 1306 459 1364 465
rect 1306 456 1318 459
rect 892 428 1318 456
rect 892 425 904 428
rect 846 419 904 425
rect 1306 425 1318 428
rect 1352 425 1364 459
rect 1306 419 1364 425
rect 294 391 352 397
rect 294 357 306 391
rect 340 388 352 391
rect 1122 391 1180 397
rect 1122 388 1134 391
rect 340 360 1134 388
rect 340 357 352 360
rect 294 351 352 357
rect 1122 357 1134 360
rect 1168 357 1180 391
rect 1122 351 1180 357
<< labels >>
rlabel locali s 1328 215 1390 265 6 A0
port 1 nsew signal input
rlabel locali s 1308 199 1390 215 6 A0
port 1 nsew signal input
rlabel locali s 1308 75 1370 199 6 A0
port 1 nsew signal input
rlabel locali s 950 143 1024 279 6 A1
port 2 nsew signal input
rlabel locali s 205 79 248 153 6 A2
port 3 nsew signal input
rlabel locali s 168 153 248 219 6 A2
port 3 nsew signal input
rlabel locali s 483 203 524 264 6 A3
port 4 nsew signal input
rlabel locali s 449 143 524 203 6 A3
port 4 nsew signal input
rlabel locali s 30 195 66 349 6 S0
port 5 nsew signal input
rlabel locali s 245 257 279 289 6 S0
port 5 nsew signal input
rlabel locali s 202 289 279 323 6 S0
port 5 nsew signal input
rlabel locali s 1226 249 1294 329 6 S0
port 5 nsew signal input
rlabel metal1 s 1214 320 1272 329 6 S0
port 5 nsew signal input
rlabel metal1 s 1214 283 1272 292 6 S0
port 5 nsew signal input
rlabel metal1 s 202 320 260 329 6 S0
port 5 nsew signal input
rlabel metal1 s 202 283 260 292 6 S0
port 5 nsew signal input
rlabel metal1 s 17 320 76 329 6 S0
port 5 nsew signal input
rlabel metal1 s 17 292 1272 320 6 S0
port 5 nsew signal input
rlabel metal1 s 17 283 76 292 6 S0
port 5 nsew signal input
rlabel locali s 558 143 616 264 6 S1
port 6 nsew signal input
rlabel locali s 1672 261 1737 491 6 X
port 7 nsew signal output
rlabel locali s 1672 53 1737 213 6 X
port 7 nsew signal output
rlabel locali s 1520 261 1554 299 6 X
port 7 nsew signal output
rlabel locali s 1520 213 1737 261 6 X
port 7 nsew signal output
rlabel locali s 1520 145 1554 213 6 X
port 7 nsew signal output
rlabel locali s 1492 299 1554 367 6 X
port 7 nsew signal output
rlabel locali s 1488 53 1554 145 6 X
port 7 nsew signal output
rlabel locali s 1472 367 1554 491 6 X
port 7 nsew signal output
rlabel locali s 1771 17 1821 177 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 1588 17 1638 177 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 1404 17 1454 163 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 960 17 1026 109 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 491 17 557 109 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 103 17 169 93 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 0 -17 1840 17 8 VGND
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1840 48 8 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 1771 299 1821 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 1588 299 1638 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 1404 367 1438 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 952 401 1021 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 520 411 566 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 103 451 169 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 0 527 1840 561 6 VPWR
port 9 nsew power bidirectional abutment
rlabel metal1 s 0 496 1840 592 6 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1840 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1779688
string GDS_START 1764080
<< end >>
