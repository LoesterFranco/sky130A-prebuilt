magic
tech sky130A
magscale 1 2
timestamp 1601050047
<< nwell >>
rect -38 332 614 704
<< pwell >>
rect 0 0 576 49
<< scpmos >>
rect 112 368 142 592
rect 196 368 226 592
rect 310 368 340 592
rect 424 368 454 592
<< nmoslvt >>
rect 84 74 114 222
rect 229 74 259 222
rect 329 74 359 222
rect 443 74 473 222
<< ndiff >>
rect 27 202 84 222
rect 27 168 39 202
rect 73 168 84 202
rect 27 120 84 168
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 185 229 222
rect 114 151 154 185
rect 188 151 229 185
rect 114 74 229 151
rect 259 210 329 222
rect 259 176 284 210
rect 318 176 329 210
rect 259 120 329 176
rect 259 86 284 120
rect 318 86 329 120
rect 259 74 329 86
rect 359 142 443 222
rect 359 108 384 142
rect 418 108 443 142
rect 359 74 443 108
rect 473 210 530 222
rect 473 176 484 210
rect 518 176 530 210
rect 473 120 530 176
rect 473 86 484 120
rect 518 86 530 120
rect 473 74 530 86
<< pdiff >>
rect 29 580 112 592
rect 29 546 41 580
rect 75 546 112 580
rect 29 497 112 546
rect 29 463 41 497
rect 75 463 112 497
rect 29 414 112 463
rect 29 380 41 414
rect 75 380 112 414
rect 29 368 112 380
rect 142 368 196 592
rect 226 580 310 592
rect 226 546 250 580
rect 284 546 310 580
rect 226 510 310 546
rect 226 476 250 510
rect 284 476 310 510
rect 226 440 310 476
rect 226 406 250 440
rect 284 406 310 440
rect 226 368 310 406
rect 340 368 424 592
rect 454 580 513 592
rect 454 546 467 580
rect 501 546 513 580
rect 454 510 513 546
rect 454 476 467 510
rect 501 476 513 510
rect 454 440 513 476
rect 454 406 467 440
rect 501 406 513 440
rect 454 368 513 406
<< ndiffc >>
rect 39 168 73 202
rect 39 86 73 120
rect 154 151 188 185
rect 284 176 318 210
rect 284 86 318 120
rect 384 108 418 142
rect 484 176 518 210
rect 484 86 518 120
<< pdiffc >>
rect 41 546 75 580
rect 41 463 75 497
rect 41 380 75 414
rect 250 546 284 580
rect 250 476 284 510
rect 250 406 284 440
rect 467 546 501 580
rect 467 476 501 510
rect 467 406 501 440
<< poly >>
rect 112 592 142 618
rect 196 592 226 618
rect 310 592 340 618
rect 424 592 454 618
rect 112 353 142 368
rect 196 353 226 368
rect 310 353 340 368
rect 424 353 454 368
rect 109 310 145 353
rect 23 294 145 310
rect 23 260 39 294
rect 73 280 145 294
rect 193 336 229 353
rect 307 336 343 353
rect 193 320 259 336
rect 193 286 209 320
rect 243 286 259 320
rect 73 260 114 280
rect 193 270 259 286
rect 307 320 373 336
rect 307 286 323 320
rect 357 286 373 320
rect 307 270 373 286
rect 421 326 457 353
rect 421 310 555 326
rect 421 276 437 310
rect 471 276 505 310
rect 539 276 555 310
rect 23 244 114 260
rect 84 222 114 244
rect 229 222 259 270
rect 329 222 359 270
rect 421 260 555 276
rect 443 222 473 260
rect 84 48 114 74
rect 229 48 259 74
rect 329 48 359 74
rect 443 48 473 74
<< polycont >>
rect 39 260 73 294
rect 209 286 243 320
rect 323 286 357 320
rect 437 276 471 310
rect 505 276 539 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 25 580 91 649
rect 25 546 41 580
rect 75 546 91 580
rect 25 497 91 546
rect 25 463 41 497
rect 75 463 91 497
rect 25 414 91 463
rect 25 380 41 414
rect 75 380 91 414
rect 25 364 91 380
rect 125 580 310 596
rect 125 546 250 580
rect 284 546 310 580
rect 125 510 310 546
rect 125 476 250 510
rect 284 476 310 510
rect 125 440 310 476
rect 125 406 250 440
rect 284 406 310 440
rect 125 390 310 406
rect 451 580 517 649
rect 451 546 467 580
rect 501 546 517 580
rect 451 510 517 546
rect 451 476 467 510
rect 501 476 517 510
rect 451 440 517 476
rect 451 406 467 440
rect 501 406 517 440
rect 451 390 517 406
rect 23 294 89 310
rect 23 260 39 294
rect 73 260 89 294
rect 23 236 89 260
rect 125 226 159 390
rect 193 320 263 356
rect 193 286 209 320
rect 243 286 263 320
rect 193 270 263 286
rect 307 320 373 356
rect 307 286 323 320
rect 357 286 373 320
rect 307 270 373 286
rect 409 310 555 356
rect 409 276 437 310
rect 471 276 505 310
rect 539 276 555 310
rect 409 260 555 276
rect 23 168 39 202
rect 73 168 89 202
rect 23 120 89 168
rect 123 185 213 226
rect 123 151 154 185
rect 188 151 213 185
rect 123 131 213 151
rect 268 210 534 226
rect 268 176 284 210
rect 318 192 484 210
rect 318 176 334 192
rect 23 86 39 120
rect 73 97 89 120
rect 268 120 334 176
rect 468 176 484 192
rect 518 176 534 210
rect 268 97 284 120
rect 73 86 284 97
rect 318 86 334 120
rect 23 63 334 86
rect 368 142 434 158
rect 368 108 384 142
rect 418 108 434 142
rect 368 17 434 108
rect 468 120 534 176
rect 468 86 484 120
rect 518 86 534 120
rect 468 70 534 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o22ai_1
flabel pwell s 0 0 576 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 576 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 576 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 576 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 223 464 257 498 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 223 538 257 572 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 576 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1297950
string GDS_START 1292270
<< end >>
