magic
tech sky130A
magscale 1 2
timestamp 1601050088
<< locali >>
rect 121 394 187 596
rect 311 424 377 596
rect 491 424 557 596
rect 783 424 849 547
rect 311 394 849 424
rect 121 390 849 394
rect 121 360 377 390
rect 21 236 87 310
rect 121 236 187 360
rect 269 260 403 326
rect 505 270 743 356
rect 793 270 935 356
rect 985 270 1127 356
rect 313 236 359 260
rect 138 226 187 236
rect 138 119 188 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 31 364 81 649
rect 221 428 271 649
rect 417 458 451 649
rect 597 458 647 649
rect 693 581 923 615
rect 693 458 743 581
rect 889 424 923 581
rect 963 458 1029 649
rect 1063 424 1129 596
rect 889 390 1129 424
rect 36 85 102 202
rect 224 202 258 226
rect 394 202 460 226
rect 224 168 460 202
rect 224 85 258 168
rect 36 51 258 85
rect 294 85 360 134
rect 394 119 460 168
rect 506 202 1120 236
rect 506 119 572 202
rect 606 85 672 168
rect 294 51 672 85
rect 708 70 742 202
rect 778 17 844 168
rect 884 70 934 202
rect 968 17 1034 168
rect 1070 70 1120 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
rlabel locali s 985 270 1127 356 6 A1
port 1 nsew signal input
rlabel locali s 793 270 935 356 6 A2
port 2 nsew signal input
rlabel locali s 505 270 743 356 6 B1
port 3 nsew signal input
rlabel locali s 313 236 359 260 6 C1
port 4 nsew signal input
rlabel locali s 269 260 403 326 6 C1
port 4 nsew signal input
rlabel locali s 21 236 87 310 6 D1
port 5 nsew signal input
rlabel locali s 783 424 849 547 6 Y
port 6 nsew signal output
rlabel locali s 491 424 557 596 6 Y
port 6 nsew signal output
rlabel locali s 311 424 377 596 6 Y
port 6 nsew signal output
rlabel locali s 311 394 849 424 6 Y
port 6 nsew signal output
rlabel locali s 138 226 187 236 6 Y
port 6 nsew signal output
rlabel locali s 138 119 188 226 6 Y
port 6 nsew signal output
rlabel locali s 121 394 187 596 6 Y
port 6 nsew signal output
rlabel locali s 121 390 849 394 6 Y
port 6 nsew signal output
rlabel locali s 121 360 377 390 6 Y
port 6 nsew signal output
rlabel locali s 121 236 187 360 6 Y
port 6 nsew signal output
rlabel metal1 s 0 -49 1152 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 617 1152 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1705216
string GDS_START 1694620
<< end >>
