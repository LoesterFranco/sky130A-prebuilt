magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 19 195 89 325
rect 359 153 431 344
rect 465 237 505 274
rect 465 153 553 237
rect 1121 221 1177 323
rect 1289 221 1390 333
rect 2587 260 2663 493
rect 2587 213 2686 260
rect 2620 51 2686 213
rect 3064 51 3140 484
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3157 561
rect 3191 527 3249 561
rect 3283 527 3312 561
rect 35 393 69 493
rect 103 427 179 527
rect 35 391 179 393
rect 35 359 137 391
rect 133 357 137 359
rect 171 357 179 391
rect 133 161 179 357
rect 35 127 179 161
rect 223 323 257 493
rect 35 69 69 127
rect 103 17 179 93
rect 223 69 257 289
rect 291 378 377 493
rect 477 378 553 527
rect 291 119 325 378
rect 591 344 657 485
rect 703 365 742 527
rect 885 404 961 493
rect 1007 442 1073 493
rect 885 364 973 404
rect 539 271 657 344
rect 596 235 657 271
rect 821 264 905 330
rect 596 169 777 235
rect 821 187 855 264
rect 939 230 973 364
rect 325 85 377 103
rect 291 51 377 85
rect 477 17 553 103
rect 596 51 641 169
rect 821 137 855 153
rect 889 196 973 230
rect 1017 357 1073 442
rect 1158 401 1226 493
rect 1270 435 1339 527
rect 1492 430 1558 493
rect 1600 435 1838 475
rect 1158 367 1474 401
rect 677 17 753 122
rect 889 119 953 196
rect 1017 165 1051 357
rect 1211 187 1245 367
rect 1424 271 1474 367
rect 1508 373 1558 430
rect 1657 391 1760 401
rect 1508 237 1542 373
rect 1657 357 1669 391
rect 1703 357 1760 391
rect 889 85 907 119
rect 941 85 953 119
rect 889 51 953 85
rect 999 129 1051 165
rect 999 119 1039 129
rect 999 85 1003 119
rect 1037 85 1039 119
rect 1179 103 1245 187
rect 999 51 1039 85
rect 1073 51 1245 103
rect 1289 17 1339 181
rect 1460 119 1542 237
rect 1576 323 1623 344
rect 1576 289 1582 323
rect 1616 289 1623 323
rect 1576 225 1623 289
rect 1657 331 1760 357
rect 1657 191 1691 331
rect 1794 315 1838 435
rect 1872 367 1919 527
rect 1794 297 1919 315
rect 1580 147 1691 191
rect 1739 263 1919 297
rect 1460 85 1463 119
rect 1497 113 1542 119
rect 1739 113 1773 263
rect 1885 249 1919 263
rect 1953 275 2029 493
rect 2071 421 2129 527
rect 2252 433 2475 471
rect 2225 391 2273 393
rect 2225 357 2232 391
rect 2266 357 2273 391
rect 1811 213 1861 219
rect 1953 213 2146 275
rect 2225 249 2273 357
rect 2307 323 2381 399
rect 2307 289 2326 323
rect 2360 289 2381 323
rect 1811 209 2146 213
rect 1811 153 2044 209
rect 2307 207 2381 289
rect 1497 85 1584 113
rect 1460 51 1584 85
rect 1628 51 1773 113
rect 1836 17 1915 112
rect 1953 51 2044 153
rect 2278 141 2381 207
rect 2425 391 2475 433
rect 2425 357 2433 391
rect 2467 357 2475 391
rect 2090 17 2145 123
rect 2425 107 2475 357
rect 2519 299 2553 527
rect 2707 293 2757 527
rect 2791 391 2837 402
rect 2791 357 2797 391
rect 2831 357 2837 391
rect 2791 315 2837 357
rect 2871 244 2939 493
rect 2983 293 3030 527
rect 2282 66 2475 107
rect 2526 17 2576 180
rect 2814 187 2939 244
rect 2730 17 2780 180
rect 2814 178 2889 187
rect 2871 153 2889 178
rect 2923 153 2939 187
rect 2871 51 2939 153
rect 2983 17 3030 180
rect 3184 293 3236 527
rect 3184 17 3236 180
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3312 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 2881 527 2915 561
rect 2973 527 3007 561
rect 3065 527 3099 561
rect 3157 527 3191 561
rect 3249 527 3283 561
rect 137 357 171 391
rect 223 289 257 323
rect 291 85 325 119
rect 821 153 855 187
rect 1669 357 1703 391
rect 907 85 941 119
rect 1003 85 1037 119
rect 1582 289 1616 323
rect 1463 85 1497 119
rect 2232 357 2266 391
rect 2326 289 2360 323
rect 2433 357 2467 391
rect 2797 357 2831 391
rect 2889 153 2923 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
rect 2881 -17 2915 17
rect 2973 -17 3007 17
rect 3065 -17 3099 17
rect 3157 -17 3191 17
rect 3249 -17 3283 17
<< metal1 >>
rect 0 561 3312 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3157 561
rect 3191 527 3249 561
rect 3283 527 3312 561
rect 0 496 3312 527
rect 0 17 3312 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3312 17
rect 0 -48 3312 -17
<< obsm1 >>
rect 125 391 183 397
rect 125 357 137 391
rect 171 388 183 391
rect 1657 391 1725 397
rect 1657 388 1669 391
rect 171 360 1669 388
rect 171 357 183 360
rect 125 351 183 357
rect 1657 357 1669 360
rect 1703 388 1725 391
rect 2215 391 2283 397
rect 2215 388 2232 391
rect 1703 360 2232 388
rect 1703 357 1725 360
rect 1657 351 1725 357
rect 2215 357 2232 360
rect 2266 357 2283 391
rect 2215 351 2283 357
rect 2421 391 2479 397
rect 2421 357 2433 391
rect 2467 388 2479 391
rect 2785 391 2843 397
rect 2785 388 2797 391
rect 2467 360 2797 388
rect 2467 357 2479 360
rect 2421 351 2479 357
rect 2785 357 2797 360
rect 2831 357 2843 391
rect 2785 351 2843 357
rect 201 323 269 329
rect 201 289 223 323
rect 257 320 269 323
rect 1565 323 1633 329
rect 1565 320 1582 323
rect 257 292 1582 320
rect 257 289 269 292
rect 201 283 269 289
rect 1565 289 1582 292
rect 1616 320 1633 323
rect 2309 323 2377 329
rect 2309 320 2326 323
rect 1616 292 2326 320
rect 1616 289 1633 292
rect 1565 283 1633 289
rect 2309 289 2326 292
rect 2360 289 2377 323
rect 2309 283 2377 289
rect 809 187 867 193
rect 809 153 821 187
rect 855 184 867 187
rect 2877 187 2935 193
rect 2877 184 2889 187
rect 855 156 2889 184
rect 855 153 867 156
rect 809 147 867 153
rect 2877 153 2889 156
rect 2923 153 2935 187
rect 2877 147 2935 153
rect 279 119 337 125
rect 279 85 291 119
rect 325 116 337 119
rect 885 119 953 125
rect 885 116 907 119
rect 325 85 907 116
rect 941 85 953 119
rect 279 79 953 85
rect 981 119 1049 125
rect 981 85 1003 119
rect 1037 116 1049 119
rect 1441 119 1509 125
rect 1441 116 1463 119
rect 1037 85 1463 116
rect 1497 85 1509 119
rect 981 79 1509 85
<< labels >>
rlabel locali s 19 195 89 325 6 CLK
port 1 nsew signal input
rlabel locali s 359 153 431 344 6 D
port 2 nsew signal input
rlabel locali s 465 237 505 274 6 DE
port 3 nsew signal input
rlabel locali s 465 153 553 237 6 DE
port 3 nsew signal input
rlabel locali s 3064 51 3140 484 6 Q
port 4 nsew signal output
rlabel locali s 2620 51 2686 213 6 Q_N
port 5 nsew signal output
rlabel locali s 2587 260 2663 493 6 Q_N
port 5 nsew signal output
rlabel locali s 2587 213 2686 260 6 Q_N
port 5 nsew signal output
rlabel locali s 1289 221 1390 333 6 SCD
port 6 nsew signal input
rlabel locali s 1121 221 1177 323 6 SCE
port 7 nsew signal input
rlabel metal1 s 0 -48 3312 48 8 VGND
port 8 nsew ground bidirectional
rlabel metal1 s 0 496 3312 592 6 VPWR
port 9 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 3312 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 453582
string GDS_START 429700
<< end >>
