magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 23 215 134 323
rect 90 199 134 215
rect 336 341 589 407
rect 336 317 626 341
rect 564 179 626 317
rect 660 296 1424 341
rect 660 213 739 296
rect 773 213 1088 262
rect 1145 215 1424 296
rect 564 173 1077 179
rect 275 139 1077 173
rect 275 123 505 139
rect 711 135 1077 139
rect 275 74 313 123
rect 467 51 505 123
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 19 401 85 493
rect 129 435 181 527
rect 236 443 673 493
rect 707 455 783 527
rect 899 455 975 527
rect 19 357 202 401
rect 236 359 285 443
rect 411 441 673 443
rect 633 421 673 441
rect 1019 421 1057 493
rect 1091 455 1167 527
rect 1210 421 1247 493
rect 1283 455 1359 527
rect 1398 421 1448 493
rect 168 269 202 357
rect 633 375 1448 421
rect 168 207 524 269
rect 168 159 231 207
rect 18 123 231 159
rect 1121 147 1365 181
rect 18 51 89 123
rect 154 17 231 89
rect 357 17 433 89
rect 549 17 677 105
rect 1121 101 1173 147
rect 713 51 1173 101
rect 1217 17 1255 113
rect 1289 51 1365 147
rect 1400 17 1448 177
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< labels >>
rlabel locali s 773 213 1088 262 6 A1
port 1 nsew signal input
rlabel locali s 1145 215 1424 296 6 A2
port 2 nsew signal input
rlabel locali s 660 296 1424 341 6 A2
port 2 nsew signal input
rlabel locali s 660 213 739 296 6 A2
port 2 nsew signal input
rlabel locali s 90 199 134 215 6 B1_N
port 3 nsew signal input
rlabel locali s 23 215 134 323 6 B1_N
port 3 nsew signal input
rlabel locali s 711 135 1077 139 6 Y
port 4 nsew signal output
rlabel locali s 564 179 626 317 6 Y
port 4 nsew signal output
rlabel locali s 564 173 1077 179 6 Y
port 4 nsew signal output
rlabel locali s 467 51 505 123 6 Y
port 4 nsew signal output
rlabel locali s 336 341 589 407 6 Y
port 4 nsew signal output
rlabel locali s 336 317 626 341 6 Y
port 4 nsew signal output
rlabel locali s 275 139 1077 173 6 Y
port 4 nsew signal output
rlabel locali s 275 123 505 139 6 Y
port 4 nsew signal output
rlabel locali s 275 74 313 123 6 Y
port 4 nsew signal output
rlabel metal1 s 0 -48 1472 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 1472 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1472 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1173848
string GDS_START 1163978
<< end >>
