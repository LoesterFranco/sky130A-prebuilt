magic
tech sky130A
magscale 1 2
timestamp 1601050088
<< locali >>
rect 25 284 130 356
rect 184 284 259 356
rect 298 284 364 356
rect 409 270 478 356
rect 580 364 655 596
rect 621 226 655 364
rect 592 70 655 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 40 424 106 596
rect 430 458 513 649
rect 40 390 546 424
rect 512 326 546 390
rect 512 260 587 326
rect 512 236 546 260
rect 23 17 89 226
rect 123 202 546 236
rect 123 108 189 202
rect 225 17 320 168
rect 372 108 438 202
rect 490 17 556 168
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel locali s 409 270 478 356 6 A
port 1 nsew signal input
rlabel locali s 298 284 364 356 6 B
port 2 nsew signal input
rlabel locali s 184 284 259 356 6 C
port 3 nsew signal input
rlabel locali s 25 284 130 356 6 D
port 4 nsew signal input
rlabel locali s 621 226 655 364 6 X
port 5 nsew signal output
rlabel locali s 592 70 655 226 6 X
port 5 nsew signal output
rlabel locali s 580 364 655 596 6 X
port 5 nsew signal output
rlabel metal1 s 0 -49 672 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 672 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 813974
string GDS_START 808088
<< end >>
