magic
tech sky130A
magscale 1 2
timestamp 1604502710
<< nwell >>
rect -38 332 710 704
<< pwell >>
rect 0 0 672 49
<< scpmos >>
rect 93 424 129 592
rect 193 424 229 592
rect 335 424 371 592
rect 435 424 471 592
rect 552 368 588 592
<< nmoslvt >>
rect 149 74 179 202
rect 227 74 257 202
rect 305 74 335 202
rect 419 74 449 202
rect 521 74 551 222
<< ndiff >>
rect 471 202 521 222
rect 96 190 149 202
rect 96 156 104 190
rect 138 156 149 190
rect 96 120 149 156
rect 96 86 104 120
rect 138 86 149 120
rect 96 74 149 86
rect 179 74 227 202
rect 257 74 305 202
rect 335 74 419 202
rect 449 190 521 202
rect 449 156 460 190
rect 494 156 521 190
rect 449 120 521 156
rect 449 86 460 120
rect 494 86 521 120
rect 449 74 521 86
rect 551 210 608 222
rect 551 176 562 210
rect 596 176 608 210
rect 551 120 608 176
rect 551 86 562 120
rect 596 86 608 120
rect 551 74 608 86
<< pdiff >>
rect 27 580 93 592
rect 27 546 39 580
rect 73 546 93 580
rect 27 504 93 546
rect 27 470 39 504
rect 73 470 93 504
rect 27 424 93 470
rect 129 580 193 592
rect 129 546 139 580
rect 173 546 193 580
rect 129 473 193 546
rect 129 439 139 473
rect 173 439 193 473
rect 129 424 193 439
rect 229 580 335 592
rect 229 546 265 580
rect 299 546 335 580
rect 229 504 335 546
rect 229 470 265 504
rect 299 470 335 504
rect 229 424 335 470
rect 371 580 435 592
rect 371 546 391 580
rect 425 546 435 580
rect 371 473 435 546
rect 371 439 391 473
rect 425 439 435 473
rect 371 424 435 439
rect 471 580 552 592
rect 471 546 498 580
rect 532 546 552 580
rect 471 510 552 546
rect 471 476 498 510
rect 532 476 552 510
rect 471 424 552 476
rect 502 368 552 424
rect 588 580 644 592
rect 588 546 598 580
rect 632 546 644 580
rect 588 497 644 546
rect 588 463 598 497
rect 632 463 644 497
rect 588 414 644 463
rect 588 380 598 414
rect 632 380 644 414
rect 588 368 644 380
<< ndiffc >>
rect 104 156 138 190
rect 104 86 138 120
rect 460 156 494 190
rect 460 86 494 120
rect 562 176 596 210
rect 562 86 596 120
<< pdiffc >>
rect 39 546 73 580
rect 39 470 73 504
rect 139 546 173 580
rect 139 439 173 473
rect 265 546 299 580
rect 265 470 299 504
rect 391 546 425 580
rect 391 439 425 473
rect 498 546 532 580
rect 498 476 532 510
rect 598 546 632 580
rect 598 463 632 497
rect 598 380 632 414
<< poly >>
rect 93 592 129 618
rect 193 592 229 618
rect 335 592 371 618
rect 435 592 471 618
rect 552 592 588 618
rect 93 358 129 424
rect 193 361 229 424
rect 85 342 151 358
rect 85 308 101 342
rect 135 308 151 342
rect 85 274 151 308
rect 193 345 263 361
rect 335 358 371 424
rect 193 311 213 345
rect 247 311 263 345
rect 193 295 263 311
rect 305 342 371 358
rect 305 308 321 342
rect 355 308 371 342
rect 435 336 471 424
rect 85 240 101 274
rect 135 247 151 274
rect 135 240 179 247
rect 85 217 179 240
rect 149 202 179 217
rect 227 202 257 295
rect 305 274 371 308
rect 305 240 321 274
rect 355 240 371 274
rect 413 320 479 336
rect 552 330 588 368
rect 413 286 429 320
rect 463 286 479 320
rect 413 270 479 286
rect 521 314 588 330
rect 521 280 537 314
rect 571 280 588 314
rect 305 224 371 240
rect 305 202 335 224
rect 419 202 449 270
rect 521 264 588 280
rect 521 222 551 264
rect 149 48 179 74
rect 227 48 257 74
rect 305 48 335 74
rect 419 48 449 74
rect 521 48 551 74
<< polycont >>
rect 101 308 135 342
rect 213 311 247 345
rect 321 308 355 342
rect 101 240 135 274
rect 321 240 355 274
rect 429 286 463 320
rect 537 280 571 314
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 23 580 89 649
rect 23 546 39 580
rect 73 546 89 580
rect 23 504 89 546
rect 23 470 39 504
rect 73 470 89 504
rect 23 463 89 470
rect 123 580 189 596
rect 123 546 139 580
rect 173 546 189 580
rect 123 473 189 546
rect 123 439 139 473
rect 173 439 189 473
rect 223 580 341 649
rect 223 546 265 580
rect 299 546 341 580
rect 223 504 341 546
rect 223 470 265 504
rect 299 470 341 504
rect 223 463 341 470
rect 375 580 441 596
rect 375 546 391 580
rect 425 546 441 580
rect 375 473 441 546
rect 123 429 189 439
rect 375 439 391 473
rect 425 439 441 473
rect 482 580 548 649
rect 482 546 498 580
rect 532 546 548 580
rect 482 510 548 546
rect 482 476 498 510
rect 532 476 548 510
rect 482 460 548 476
rect 582 580 655 596
rect 582 546 598 580
rect 632 546 655 580
rect 582 497 655 546
rect 582 463 598 497
rect 632 463 655 497
rect 375 429 441 439
rect 17 426 441 429
rect 17 395 548 426
rect 17 190 51 395
rect 375 392 548 395
rect 85 342 163 358
rect 85 308 101 342
rect 135 308 163 342
rect 85 274 163 308
rect 85 240 101 274
rect 135 240 163 274
rect 85 224 163 240
rect 197 345 263 361
rect 197 311 213 345
rect 247 311 263 345
rect 17 156 104 190
rect 138 156 154 190
rect 17 120 154 156
rect 17 86 104 120
rect 138 86 154 120
rect 197 88 263 311
rect 305 342 371 358
rect 305 308 321 342
rect 355 308 371 342
rect 305 274 371 308
rect 305 240 321 274
rect 355 240 371 274
rect 409 320 479 356
rect 409 286 429 320
rect 463 286 479 320
rect 409 270 479 286
rect 514 330 548 392
rect 582 414 655 463
rect 582 380 598 414
rect 632 380 655 414
rect 582 364 655 380
rect 514 314 587 330
rect 514 280 537 314
rect 571 280 587 314
rect 514 264 587 280
rect 305 88 371 240
rect 621 226 655 364
rect 546 210 655 226
rect 444 190 510 206
rect 444 156 460 190
rect 494 156 510 190
rect 444 120 510 156
rect 17 71 154 86
rect 444 86 460 120
rect 494 86 510 120
rect 444 17 510 86
rect 546 176 562 210
rect 596 176 655 210
rect 546 120 655 176
rect 546 86 562 120
rect 596 86 655 120
rect 546 70 655 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
rlabel comment s 0 0 0 0 4 and4_1
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 127 242 161 276 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 223 94 257 128 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 223 168 257 202 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 223 242 257 276 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 319 94 353 128 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 319 168 353 202 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 319 242 353 276 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 D
port 4 nsew
flabel corelocali s 607 94 641 128 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 607 168 641 202 0 FreeSans 340 0 0 0 X
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 672 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3166682
string GDS_START 3159544
<< end >>
