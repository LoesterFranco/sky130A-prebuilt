magic
tech sky130A
magscale 1 2
timestamp 1599588244
<< locali >>
rect 114 424 164 596
rect 312 424 346 596
rect 114 390 455 424
rect 121 270 263 356
rect 297 270 363 356
rect 409 236 455 390
rect 291 202 455 236
rect 291 119 357 202
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 24 364 74 649
rect 204 458 270 649
rect 386 458 452 649
rect 23 202 255 236
rect 23 70 73 202
rect 109 17 175 168
rect 221 85 255 202
rect 391 85 457 168
rect 221 51 457 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< metal1 >>
rect 0 683 480 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 0 617 480 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 480 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
rect 0 -49 480 -17
<< labels >>
rlabel locali s 297 270 363 356 6 A
port 1 nsew signal input
rlabel locali s 121 270 263 356 6 B
port 2 nsew signal input
rlabel locali s 409 236 455 390 6 Y
port 3 nsew signal output
rlabel locali s 312 424 346 596 6 Y
port 3 nsew signal output
rlabel locali s 291 202 455 236 6 Y
port 3 nsew signal output
rlabel locali s 291 119 357 202 6 Y
port 3 nsew signal output
rlabel locali s 114 424 164 596 6 Y
port 3 nsew signal output
rlabel locali s 114 390 455 424 6 Y
port 3 nsew signal output
rlabel metal1 s 0 -49 480 49 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 5 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 617 480 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 480 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1880436
string GDS_START 1875472
<< end >>
