magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 25 270 110 430
rect 554 364 651 596
rect 409 270 475 356
rect 617 230 651 364
rect 583 74 651 230
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 23 464 233 530
rect 162 236 228 464
rect 273 364 307 649
rect 341 390 413 540
rect 454 390 520 649
rect 23 202 228 236
rect 341 230 375 390
rect 515 264 583 330
rect 515 230 549 264
rect 23 70 89 202
rect 262 196 549 230
rect 123 17 189 168
rect 262 94 328 196
rect 426 17 549 162
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel locali s 25 270 110 430 6 A_N
port 1 nsew signal input
rlabel locali s 409 270 475 356 6 B
port 2 nsew signal input
rlabel locali s 617 230 651 364 6 X
port 3 nsew signal output
rlabel locali s 583 74 651 230 6 X
port 3 nsew signal output
rlabel locali s 554 364 651 596 6 X
port 3 nsew signal output
rlabel metal1 s 0 -49 672 49 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 617 672 715 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3855920
string GDS_START 3849834
<< end >>
