magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 808 325 858 425
rect 808 291 990 325
rect 40 215 203 257
rect 247 215 428 257
rect 482 215 671 257
rect 728 215 855 257
rect 923 181 990 291
rect 114 145 990 181
rect 114 51 190 145
rect 302 51 378 145
rect 602 51 678 145
rect 790 51 866 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 30 325 81 493
rect 125 359 175 527
rect 219 325 269 493
rect 313 459 663 493
rect 313 359 363 459
rect 407 325 457 425
rect 30 291 457 325
rect 519 325 569 425
rect 613 359 663 459
rect 707 459 945 493
rect 707 325 757 459
rect 519 291 757 325
rect 895 359 945 459
rect 18 17 73 181
rect 227 17 261 111
rect 415 17 561 111
rect 715 17 749 111
rect 903 17 961 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
rlabel locali s 40 215 203 257 6 A
port 1 nsew signal input
rlabel locali s 247 215 428 257 6 B
port 2 nsew signal input
rlabel locali s 482 215 671 257 6 C
port 3 nsew signal input
rlabel locali s 728 215 855 257 6 D
port 4 nsew signal input
rlabel locali s 923 181 990 291 6 Y
port 5 nsew signal output
rlabel locali s 808 325 858 425 6 Y
port 5 nsew signal output
rlabel locali s 808 291 990 325 6 Y
port 5 nsew signal output
rlabel locali s 790 51 866 145 6 Y
port 5 nsew signal output
rlabel locali s 602 51 678 145 6 Y
port 5 nsew signal output
rlabel locali s 302 51 378 145 6 Y
port 5 nsew signal output
rlabel locali s 114 145 990 181 6 Y
port 5 nsew signal output
rlabel locali s 114 51 190 145 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -48 1012 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 1012 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1012 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2487712
string GDS_START 2479646
<< end >>
