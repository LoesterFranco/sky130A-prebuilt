magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 644 561
rect 18 327 69 527
rect 21 17 69 177
rect 106 51 155 493
rect 189 437 359 527
rect 289 202 371 323
rect 481 280 522 397
rect 559 330 624 527
rect 405 205 522 280
rect 573 199 625 290
rect 189 17 255 93
rect 469 17 535 93
rect 0 -17 644 17
<< obsli1 >>
rect 393 401 445 493
rect 221 357 445 401
rect 221 266 255 357
rect 189 168 255 266
rect 189 127 359 168
rect 293 51 359 127
rect 393 127 624 165
rect 393 93 435 127
rect 569 99 624 127
<< metal1 >>
rect 0 496 644 592
rect 0 -48 644 48
<< labels >>
rlabel locali s 573 199 625 290 6 A1
port 1 nsew signal input
rlabel locali s 481 280 522 397 6 A2
port 2 nsew signal input
rlabel locali s 405 205 522 280 6 A2
port 2 nsew signal input
rlabel locali s 289 202 371 323 6 B1
port 3 nsew signal input
rlabel locali s 106 51 155 493 6 X
port 4 nsew signal output
rlabel locali s 469 17 535 93 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 189 17 255 93 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 21 17 69 177 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 644 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 644 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 559 330 624 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 189 437 359 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 18 327 69 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 644 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 644 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1352670
string GDS_START 1347162
<< end >>
