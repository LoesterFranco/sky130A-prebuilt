magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 17 211 121 323
rect 556 299 622 493
rect 572 165 622 299
rect 556 51 622 165
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 17 401 76 493
rect 120 435 163 527
rect 197 435 284 493
rect 17 357 189 401
rect 155 265 189 357
rect 155 199 216 265
rect 250 255 284 435
rect 323 349 368 416
rect 429 383 503 527
rect 323 315 522 349
rect 480 265 522 315
rect 250 215 419 255
rect 155 177 189 199
rect 19 143 189 177
rect 19 51 76 143
rect 250 109 284 215
rect 480 199 538 265
rect 480 181 522 199
rect 120 17 163 109
rect 197 51 284 109
rect 323 147 522 181
rect 323 102 368 147
rect 429 17 511 113
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 17 211 121 323 6 A
port 1 nsew signal input
rlabel locali s 572 165 622 299 6 X
port 2 nsew signal output
rlabel locali s 556 299 622 493 6 X
port 2 nsew signal output
rlabel locali s 556 51 622 165 6 X
port 2 nsew signal output
rlabel metal1 s 0 -48 644 48 8 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 4 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3299132
string GDS_START 3293176
<< end >>
