magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 89 47 119 131
rect 186 47 216 177
rect 321 47 351 177
rect 432 53 462 137
rect 518 53 548 137
rect 608 53 638 137
<< pmoshvt >>
rect 81 360 117 444
rect 188 297 224 497
rect 304 297 340 497
rect 412 297 448 381
rect 510 297 546 381
rect 600 297 636 381
<< ndiff >>
rect 134 131 186 177
rect 27 108 89 131
rect 27 74 35 108
rect 69 74 89 108
rect 27 47 89 74
rect 119 97 186 131
rect 119 63 129 97
rect 163 63 186 97
rect 119 47 186 63
rect 216 103 321 177
rect 216 69 236 103
rect 270 69 321 103
rect 216 47 321 69
rect 351 137 401 177
rect 351 97 432 137
rect 351 63 373 97
rect 407 63 432 97
rect 351 53 432 63
rect 462 111 518 137
rect 462 77 473 111
rect 507 77 518 111
rect 462 53 518 77
rect 548 97 608 137
rect 548 63 564 97
rect 598 63 608 97
rect 548 53 608 63
rect 638 111 690 137
rect 638 77 648 111
rect 682 77 690 111
rect 638 53 690 77
rect 351 47 412 53
<< pdiff >>
rect 134 476 188 497
rect 134 444 142 476
rect 27 412 81 444
rect 27 378 35 412
rect 69 378 81 412
rect 27 360 81 378
rect 117 442 142 444
rect 176 442 188 476
rect 117 360 188 442
rect 134 297 188 360
rect 224 340 304 497
rect 224 306 236 340
rect 270 306 304 340
rect 224 297 304 306
rect 340 476 395 497
rect 340 442 353 476
rect 387 442 395 476
rect 340 381 395 442
rect 340 297 412 381
rect 448 297 510 381
rect 546 297 600 381
rect 636 354 690 381
rect 636 320 648 354
rect 682 320 690 354
rect 636 297 690 320
<< ndiffc >>
rect 35 74 69 108
rect 129 63 163 97
rect 236 69 270 103
rect 373 63 407 97
rect 473 77 507 111
rect 564 63 598 97
rect 648 77 682 111
<< pdiffc >>
rect 35 378 69 412
rect 142 442 176 476
rect 236 306 270 340
rect 353 442 387 476
rect 648 320 682 354
<< poly >>
rect 188 497 224 523
rect 304 497 340 523
rect 81 444 117 470
rect 81 345 117 360
rect 79 265 119 345
rect 486 473 562 483
rect 486 439 502 473
rect 536 439 562 473
rect 486 429 562 439
rect 508 407 548 429
rect 412 381 448 407
rect 510 381 546 407
rect 600 381 636 407
rect 188 282 224 297
rect 304 282 340 297
rect 412 282 448 297
rect 510 282 546 297
rect 600 282 636 297
rect 22 249 119 265
rect 22 215 35 249
rect 69 215 119 249
rect 22 199 119 215
rect 89 131 119 199
rect 186 265 226 282
rect 302 265 342 282
rect 410 265 450 282
rect 186 249 351 265
rect 186 215 297 249
rect 331 215 351 249
rect 186 199 351 215
rect 398 249 462 265
rect 398 215 408 249
rect 442 215 462 249
rect 508 222 548 282
rect 598 265 638 282
rect 398 199 462 215
rect 186 177 216 199
rect 321 177 351 199
rect 432 137 462 199
rect 518 137 548 222
rect 590 249 650 265
rect 590 215 600 249
rect 634 215 650 249
rect 590 199 650 215
rect 608 137 638 199
rect 89 21 119 47
rect 186 21 216 47
rect 321 21 351 47
rect 432 27 462 53
rect 518 27 548 53
rect 608 27 638 53
<< polycont >>
rect 502 439 536 473
rect 35 215 69 249
rect 297 215 331 249
rect 408 215 442 249
rect 600 215 634 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 120 476 192 527
rect 17 412 69 444
rect 120 442 142 476
rect 176 442 192 476
rect 337 476 403 527
rect 337 442 353 476
rect 387 442 403 476
rect 439 439 502 473
rect 536 439 709 473
rect 439 425 709 439
rect 17 378 35 412
rect 69 391 396 408
rect 69 378 604 391
rect 17 374 604 378
rect 17 362 163 374
rect 17 249 85 328
rect 17 215 35 249
rect 69 215 85 249
rect 129 181 163 362
rect 362 357 604 374
rect 17 147 163 181
rect 197 306 236 340
rect 270 306 286 340
rect 197 299 286 306
rect 17 108 69 147
rect 197 119 247 299
rect 297 249 331 265
rect 391 249 508 323
rect 391 215 408 249
rect 442 215 508 249
rect 570 265 604 357
rect 648 354 709 385
rect 682 320 709 354
rect 648 299 709 320
rect 570 249 640 265
rect 570 215 600 249
rect 634 215 640 249
rect 297 181 331 215
rect 570 199 640 215
rect 297 165 507 181
rect 675 165 709 299
rect 297 147 709 165
rect 473 131 709 147
rect 17 74 35 108
rect 17 58 69 74
rect 129 97 163 113
rect 129 17 163 63
rect 197 103 277 119
rect 197 69 236 103
rect 270 69 277 103
rect 197 53 277 69
rect 373 97 407 113
rect 373 17 407 63
rect 473 111 507 131
rect 648 111 709 131
rect 473 61 507 77
rect 548 63 564 97
rect 598 63 614 97
rect 548 17 614 63
rect 682 77 709 111
rect 648 61 709 77
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel corelocali s 437 238 437 238 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 575 442 575 442 0 FreeSans 400 180 0 0 B
port 2 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 400 0 0 0 C_N
port 3 nsew
flabel corelocali s 231 102 231 102 0 FreeSans 200 180 0 0 X
port 8 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
rlabel comment s 0 0 0 0 4 or3b_2
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 485170
string GDS_START 479060
<< end >>
