magic
tech sky130A
magscale 1 2
timestamp 1604502705
<< nwell >>
rect -38 332 1766 704
<< pwell >>
rect 0 0 1728 49
<< scnmos >>
rect 79 47 1649 202
<< scpmos >>
rect 79 368 1649 619
<< ndiff >>
rect 27 190 79 202
rect 27 156 35 190
rect 69 156 79 190
rect 27 93 79 156
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 1649 190 1701 202
rect 1649 156 1659 190
rect 1693 156 1701 190
rect 1649 93 1701 156
rect 1649 59 1659 93
rect 1693 59 1701 93
rect 1649 47 1701 59
<< pdiff >>
rect 27 607 79 619
rect 27 573 35 607
rect 69 573 79 607
rect 27 510 79 573
rect 27 476 35 510
rect 69 476 79 510
rect 27 414 79 476
rect 27 380 35 414
rect 69 380 79 414
rect 27 368 79 380
rect 1649 607 1701 619
rect 1649 573 1659 607
rect 1693 573 1701 607
rect 1649 511 1701 573
rect 1649 477 1659 511
rect 1693 477 1701 511
rect 1649 414 1701 477
rect 1649 380 1659 414
rect 1693 380 1701 414
rect 1649 368 1701 380
<< ndiffc >>
rect 35 156 69 190
rect 35 59 69 93
rect 1659 156 1693 190
rect 1659 59 1693 93
<< pdiffc >>
rect 35 573 69 607
rect 35 476 69 510
rect 35 380 69 414
rect 1659 573 1693 607
rect 1659 477 1693 511
rect 1659 380 1693 414
<< poly >>
rect 79 619 1649 645
rect 79 342 1649 368
rect 79 320 225 342
rect 79 286 107 320
rect 141 286 175 320
rect 209 286 225 320
rect 443 320 577 342
rect 79 270 225 286
rect 267 284 401 300
rect 267 250 283 284
rect 317 250 351 284
rect 385 250 401 284
rect 443 286 459 320
rect 493 286 527 320
rect 561 286 577 320
rect 795 320 929 342
rect 443 270 577 286
rect 619 284 753 300
rect 267 228 401 250
rect 619 250 635 284
rect 669 250 703 284
rect 737 250 753 284
rect 795 286 811 320
rect 845 286 879 320
rect 913 286 929 320
rect 1147 320 1281 342
rect 795 270 929 286
rect 971 284 1105 300
rect 619 228 753 250
rect 971 250 987 284
rect 1021 250 1055 284
rect 1089 250 1105 284
rect 1147 286 1163 320
rect 1197 286 1231 320
rect 1265 286 1281 320
rect 1499 320 1649 342
rect 1147 270 1281 286
rect 1323 284 1457 300
rect 971 228 1105 250
rect 1323 250 1339 284
rect 1373 250 1407 284
rect 1441 250 1457 284
rect 1499 286 1515 320
rect 1549 286 1583 320
rect 1617 286 1649 320
rect 1499 270 1649 286
rect 1323 228 1457 250
rect 79 202 1649 228
rect 79 21 1649 47
<< polycont >>
rect 107 286 141 320
rect 175 286 209 320
rect 283 250 317 284
rect 351 250 385 284
rect 459 286 493 320
rect 527 286 561 320
rect 635 250 669 284
rect 703 250 737 284
rect 811 286 845 320
rect 879 286 913 320
rect 987 250 1021 284
rect 1055 250 1089 284
rect 1163 286 1197 320
rect 1231 286 1265 320
rect 1339 250 1373 284
rect 1407 250 1441 284
rect 1515 286 1549 320
rect 1583 286 1617 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 17 607 1711 649
rect 17 573 35 607
rect 69 573 1659 607
rect 1693 573 1711 607
rect 17 511 1711 573
rect 17 510 1659 511
rect 17 476 35 510
rect 69 477 1659 510
rect 1693 477 1711 511
rect 69 476 1711 477
rect 17 414 1711 476
rect 17 380 35 414
rect 69 380 1659 414
rect 1693 380 1711 414
rect 17 354 1711 380
rect 17 286 107 320
rect 141 286 175 320
rect 209 286 231 320
rect 17 216 231 286
rect 265 284 403 354
rect 265 250 283 284
rect 317 250 351 284
rect 385 250 403 284
rect 441 286 459 320
rect 493 286 527 320
rect 561 286 579 320
rect 441 216 579 286
rect 617 284 755 354
rect 617 250 635 284
rect 669 250 703 284
rect 737 250 755 284
rect 793 286 811 320
rect 845 286 879 320
rect 913 286 931 320
rect 793 216 931 286
rect 969 284 1107 354
rect 969 250 987 284
rect 1021 250 1055 284
rect 1089 250 1107 284
rect 1145 286 1163 320
rect 1197 286 1231 320
rect 1265 286 1283 320
rect 1145 216 1283 286
rect 1321 284 1459 354
rect 1321 250 1339 284
rect 1373 250 1407 284
rect 1441 250 1459 284
rect 1497 286 1515 320
rect 1549 286 1583 320
rect 1617 286 1711 320
rect 1497 216 1711 286
rect 17 190 1711 216
rect 17 156 35 190
rect 69 156 1659 190
rect 1693 156 1711 190
rect 17 93 1711 156
rect 17 59 35 93
rect 69 59 1659 93
rect 1693 59 1711 93
rect 17 17 1711 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
<< metal1 >>
rect 0 683 1728 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 0 617 1728 649
rect 0 17 1728 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
rect 0 -49 1728 -17
<< labels >>
flabel pwell s 0 0 1728 49 0 FreeSans 200 0 0 0 VNB
port 2 nsew
flabel nbase s 0 617 1728 666 0 FreeSans 200 0 0 0 VPB
port 3 nsew
rlabel comment s 0 0 0 0 4 decaphe_18
flabel metal1 s 0 0 1728 49 0 FreeSans 340 0 0 0 VGND
port 1 nsew
flabel metal1 s 0 617 1728 666 0 FreeSans 340 0 0 0 VPWR
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 1728 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3443966
string GDS_START 3437870
<< end >>
