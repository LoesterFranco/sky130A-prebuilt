magic
tech sky130A
magscale 1 2
timestamp 1604502710
<< nwell >>
rect -38 332 3398 704
rect 1223 325 1436 332
<< pwell >>
rect 0 0 3360 49
<< scpmos >>
rect 93 464 129 592
rect 177 464 213 592
rect 403 463 439 591
rect 539 463 575 591
rect 617 463 653 591
rect 707 463 743 591
rect 902 455 938 583
rect 1038 455 1074 583
rect 1116 455 1152 583
rect 1312 361 1348 585
rect 1582 368 1618 592
rect 1776 508 1812 592
rect 1866 508 1902 592
rect 1962 508 1998 592
rect 2065 398 2101 566
rect 2259 392 2295 592
rect 2451 392 2487 592
rect 2553 508 2589 592
rect 2637 508 2673 592
rect 2779 464 2815 592
rect 2973 368 3009 592
rect 3063 368 3099 592
rect 3153 368 3189 592
rect 3243 368 3279 592
<< nmoslvt >>
rect 105 74 135 158
rect 183 74 213 158
rect 381 113 411 197
rect 467 113 497 197
rect 545 113 575 197
rect 631 113 661 197
rect 928 125 958 209
rect 1014 125 1044 209
rect 1086 125 1116 209
rect 1283 74 1313 222
rect 1480 74 1510 222
rect 1726 97 1756 181
rect 1828 79 1858 163
rect 1943 79 1973 163
rect 2079 79 2109 207
rect 2301 74 2331 202
rect 2373 74 2403 202
rect 2468 74 2498 158
rect 2546 74 2576 158
rect 2776 74 2806 158
rect 2974 116 3004 264
rect 3060 116 3090 264
rect 3160 116 3190 264
rect 3249 116 3279 264
<< ndiff >>
rect 324 172 381 197
rect 48 132 105 158
rect 48 98 60 132
rect 94 98 105 132
rect 48 74 105 98
rect 135 74 183 158
rect 213 133 270 158
rect 213 99 224 133
rect 258 99 270 133
rect 324 138 336 172
rect 370 138 381 172
rect 324 113 381 138
rect 411 172 467 197
rect 411 138 422 172
rect 456 138 467 172
rect 411 113 467 138
rect 497 113 545 197
rect 575 172 631 197
rect 575 138 586 172
rect 620 138 631 172
rect 575 113 631 138
rect 661 185 761 197
rect 661 151 700 185
rect 734 151 761 185
rect 661 113 761 151
rect 213 74 270 99
rect 871 178 928 209
rect 871 144 883 178
rect 917 144 928 178
rect 871 125 928 144
rect 958 178 1014 209
rect 958 144 969 178
rect 1003 144 1014 178
rect 958 125 1014 144
rect 1044 125 1086 209
rect 1116 184 1172 209
rect 1116 150 1127 184
rect 1161 150 1172 184
rect 1116 125 1172 150
rect 1226 141 1283 222
rect 1226 107 1238 141
rect 1272 107 1283 141
rect 1226 74 1283 107
rect 1313 202 1369 222
rect 1313 168 1324 202
rect 1358 168 1369 202
rect 1313 120 1369 168
rect 1313 86 1324 120
rect 1358 86 1369 120
rect 1313 74 1369 86
rect 1423 127 1480 222
rect 1423 93 1435 127
rect 1469 93 1480 127
rect 1423 74 1480 93
rect 1510 210 1566 222
rect 1510 176 1521 210
rect 1555 176 1566 210
rect 1510 120 1566 176
rect 1510 86 1521 120
rect 1555 86 1566 120
rect 1620 169 1726 181
rect 1620 135 1631 169
rect 1665 135 1726 169
rect 1620 97 1726 135
rect 1756 169 1813 181
rect 1756 135 1767 169
rect 1801 163 1813 169
rect 2029 163 2079 207
rect 1801 135 1828 163
rect 1756 97 1828 135
rect 1510 74 1566 86
rect 1778 79 1828 97
rect 1858 79 1943 163
rect 1973 122 2079 163
rect 1973 88 1984 122
rect 2018 88 2079 122
rect 1973 79 2079 88
rect 2109 182 2166 207
rect 2109 148 2120 182
rect 2154 148 2166 182
rect 2109 79 2166 148
rect 2244 121 2301 202
rect 2244 87 2256 121
rect 2290 87 2301 121
rect 2244 74 2301 87
rect 2331 74 2373 202
rect 2403 158 2453 202
rect 2917 252 2974 264
rect 2917 218 2929 252
rect 2963 218 2974 252
rect 2917 162 2974 218
rect 2403 133 2468 158
rect 2403 99 2423 133
rect 2457 99 2468 133
rect 2403 74 2468 99
rect 2498 74 2546 158
rect 2576 120 2776 158
rect 2576 86 2587 120
rect 2621 86 2717 120
rect 2751 86 2776 120
rect 2576 74 2776 86
rect 2806 133 2863 158
rect 2806 99 2817 133
rect 2851 99 2863 133
rect 2917 128 2929 162
rect 2963 128 2974 162
rect 2917 116 2974 128
rect 3004 252 3060 264
rect 3004 218 3015 252
rect 3049 218 3060 252
rect 3004 162 3060 218
rect 3004 128 3015 162
rect 3049 128 3060 162
rect 3004 116 3060 128
rect 3090 165 3160 264
rect 3090 131 3115 165
rect 3149 131 3160 165
rect 3090 116 3160 131
rect 3190 252 3249 264
rect 3190 218 3202 252
rect 3236 218 3249 252
rect 3190 165 3249 218
rect 3190 131 3202 165
rect 3236 131 3249 165
rect 3190 116 3249 131
rect 3279 165 3333 264
rect 3279 131 3290 165
rect 3324 131 3333 165
rect 3279 116 3333 131
rect 2806 74 2863 99
<< pdiff >>
rect 37 580 93 592
rect 37 546 49 580
rect 83 546 93 580
rect 37 510 93 546
rect 37 476 49 510
rect 83 476 93 510
rect 37 464 93 476
rect 129 464 177 592
rect 213 578 269 592
rect 213 544 223 578
rect 257 544 269 578
rect 213 464 269 544
rect 347 520 403 591
rect 347 486 359 520
rect 393 486 403 520
rect 347 463 403 486
rect 439 577 539 591
rect 439 543 495 577
rect 529 543 539 577
rect 439 463 539 543
rect 575 463 617 591
rect 653 579 707 591
rect 653 545 663 579
rect 697 545 707 579
rect 653 509 707 545
rect 653 475 663 509
rect 697 475 707 509
rect 653 463 707 475
rect 743 579 795 591
rect 743 545 753 579
rect 787 545 795 579
rect 743 509 795 545
rect 743 475 753 509
rect 787 475 795 509
rect 743 463 795 475
rect 849 516 902 583
rect 849 482 858 516
rect 892 482 902 516
rect 849 455 902 482
rect 938 570 1038 583
rect 938 536 994 570
rect 1028 536 1038 570
rect 938 455 1038 536
rect 1074 455 1116 583
rect 1152 571 1205 583
rect 1152 537 1162 571
rect 1196 537 1205 571
rect 1152 501 1205 537
rect 1152 467 1162 501
rect 1196 467 1205 501
rect 1152 455 1205 467
rect 1259 571 1312 585
rect 1259 537 1268 571
rect 1302 537 1312 571
rect 1259 361 1312 537
rect 1348 412 1400 585
rect 1530 574 1582 592
rect 1530 540 1538 574
rect 1572 540 1582 574
rect 1348 378 1358 412
rect 1392 378 1400 412
rect 1348 361 1400 378
rect 1530 368 1582 540
rect 1618 415 1670 592
rect 1724 567 1776 592
rect 1724 533 1732 567
rect 1766 533 1776 567
rect 1724 508 1776 533
rect 1812 567 1866 592
rect 1812 533 1822 567
rect 1856 533 1866 567
rect 1812 508 1866 533
rect 1902 508 1962 592
rect 1998 580 2050 592
rect 1998 546 2008 580
rect 2042 566 2050 580
rect 2207 580 2259 592
rect 2042 546 2065 566
rect 1998 508 2065 546
rect 1618 381 1628 415
rect 1662 381 1670 415
rect 1618 368 1670 381
rect 2015 398 2065 508
rect 2101 444 2153 566
rect 2101 410 2111 444
rect 2145 410 2153 444
rect 2101 398 2153 410
rect 2207 546 2215 580
rect 2249 546 2259 580
rect 2207 392 2259 546
rect 2295 392 2451 592
rect 2487 567 2553 592
rect 2487 533 2509 567
rect 2543 533 2553 567
rect 2487 508 2553 533
rect 2589 508 2637 592
rect 2673 580 2779 592
rect 2673 546 2704 580
rect 2738 546 2779 580
rect 2673 508 2779 546
rect 2487 392 2537 508
rect 2729 464 2779 508
rect 2815 580 2867 592
rect 2815 546 2825 580
rect 2859 546 2867 580
rect 2815 510 2867 546
rect 2815 476 2825 510
rect 2859 476 2867 510
rect 2815 464 2867 476
rect 2921 580 2973 592
rect 2921 546 2929 580
rect 2963 546 2973 580
rect 2921 506 2973 546
rect 2921 472 2929 506
rect 2963 472 2973 506
rect 2921 424 2973 472
rect 2921 390 2929 424
rect 2963 390 2973 424
rect 2921 368 2973 390
rect 3009 580 3063 592
rect 3009 546 3019 580
rect 3053 546 3063 580
rect 3009 506 3063 546
rect 3009 472 3019 506
rect 3053 472 3063 506
rect 3009 414 3063 472
rect 3009 380 3019 414
rect 3053 380 3063 414
rect 3009 368 3063 380
rect 3099 580 3153 592
rect 3099 546 3109 580
rect 3143 546 3153 580
rect 3099 498 3153 546
rect 3099 464 3109 498
rect 3143 464 3153 498
rect 3099 368 3153 464
rect 3189 580 3243 592
rect 3189 546 3199 580
rect 3233 546 3243 580
rect 3189 506 3243 546
rect 3189 472 3199 506
rect 3233 472 3243 506
rect 3189 414 3243 472
rect 3189 380 3199 414
rect 3233 380 3243 414
rect 3189 368 3243 380
rect 3279 580 3333 592
rect 3279 546 3289 580
rect 3323 546 3333 580
rect 3279 498 3333 546
rect 3279 464 3289 498
rect 3323 464 3333 498
rect 3279 368 3333 464
<< ndiffc >>
rect 60 98 94 132
rect 224 99 258 133
rect 336 138 370 172
rect 422 138 456 172
rect 586 138 620 172
rect 700 151 734 185
rect 883 144 917 178
rect 969 144 1003 178
rect 1127 150 1161 184
rect 1238 107 1272 141
rect 1324 168 1358 202
rect 1324 86 1358 120
rect 1435 93 1469 127
rect 1521 176 1555 210
rect 1521 86 1555 120
rect 1631 135 1665 169
rect 1767 135 1801 169
rect 1984 88 2018 122
rect 2120 148 2154 182
rect 2256 87 2290 121
rect 2929 218 2963 252
rect 2423 99 2457 133
rect 2587 86 2621 120
rect 2717 86 2751 120
rect 2817 99 2851 133
rect 2929 128 2963 162
rect 3015 218 3049 252
rect 3015 128 3049 162
rect 3115 131 3149 165
rect 3202 218 3236 252
rect 3202 131 3236 165
rect 3290 131 3324 165
<< pdiffc >>
rect 49 546 83 580
rect 49 476 83 510
rect 223 544 257 578
rect 359 486 393 520
rect 495 543 529 577
rect 663 545 697 579
rect 663 475 697 509
rect 753 545 787 579
rect 753 475 787 509
rect 858 482 892 516
rect 994 536 1028 570
rect 1162 537 1196 571
rect 1162 467 1196 501
rect 1268 537 1302 571
rect 1538 540 1572 574
rect 1358 378 1392 412
rect 1732 533 1766 567
rect 1822 533 1856 567
rect 2008 546 2042 580
rect 1628 381 1662 415
rect 2111 410 2145 444
rect 2215 546 2249 580
rect 2509 533 2543 567
rect 2704 546 2738 580
rect 2825 546 2859 580
rect 2825 476 2859 510
rect 2929 546 2963 580
rect 2929 472 2963 506
rect 2929 390 2963 424
rect 3019 546 3053 580
rect 3019 472 3053 506
rect 3019 380 3053 414
rect 3109 546 3143 580
rect 3109 464 3143 498
rect 3199 546 3233 580
rect 3199 472 3233 506
rect 3199 380 3233 414
rect 3289 546 3323 580
rect 3289 464 3323 498
<< poly >>
rect 93 592 129 618
rect 177 592 213 618
rect 403 591 439 617
rect 539 591 575 617
rect 617 591 653 617
rect 707 606 938 636
rect 707 591 743 606
rect 93 398 129 464
rect 177 424 213 464
rect 902 583 938 606
rect 1038 583 1074 609
rect 1116 583 1152 609
rect 1312 585 1348 611
rect 1582 592 1618 618
rect 1776 592 1812 618
rect 1866 592 1902 618
rect 1962 592 1998 618
rect 2259 592 2295 618
rect 2451 592 2487 618
rect 2553 592 2589 618
rect 2637 592 2673 618
rect 2779 592 2815 618
rect 2973 592 3009 618
rect 3063 592 3099 618
rect 3153 592 3189 618
rect 3243 592 3279 618
rect 403 448 439 463
rect 539 448 575 463
rect 177 408 265 424
rect 69 382 135 398
rect 69 348 85 382
rect 119 348 135 382
rect 69 314 135 348
rect 69 280 85 314
rect 119 280 135 314
rect 177 374 215 408
rect 249 374 265 408
rect 177 340 265 374
rect 177 306 215 340
rect 249 306 265 340
rect 337 418 575 448
rect 337 330 367 418
rect 617 370 653 463
rect 707 437 743 463
rect 415 354 497 370
rect 177 290 265 306
rect 307 314 373 330
rect 69 246 135 280
rect 69 212 85 246
rect 119 212 135 246
rect 307 280 323 314
rect 357 280 373 314
rect 415 320 431 354
rect 465 320 497 354
rect 415 304 497 320
rect 307 242 373 280
rect 69 196 135 212
rect 105 158 135 196
rect 183 212 411 242
rect 183 158 213 212
rect 381 197 411 212
rect 467 197 497 304
rect 545 354 653 370
rect 545 320 561 354
rect 595 320 653 354
rect 545 304 653 320
rect 783 373 849 389
rect 783 339 799 373
rect 833 339 849 373
rect 783 305 849 339
rect 545 197 575 304
rect 783 271 799 305
rect 833 271 849 305
rect 902 302 938 455
rect 1038 349 1074 455
rect 1008 333 1074 349
rect 783 242 849 271
rect 631 237 849 242
rect 631 212 799 237
rect 631 197 661 212
rect 783 203 799 212
rect 833 203 849 237
rect 891 286 958 302
rect 891 252 907 286
rect 941 252 958 286
rect 1008 299 1024 333
rect 1058 299 1074 333
rect 1008 283 1074 299
rect 1116 417 1152 455
rect 1116 401 1182 417
rect 1116 367 1132 401
rect 1166 367 1182 401
rect 1116 333 1182 367
rect 1432 407 1510 423
rect 1432 373 1448 407
rect 1482 373 1510 407
rect 1116 299 1132 333
rect 1166 299 1182 333
rect 1312 310 1348 361
rect 1432 353 1510 373
rect 2065 566 2101 592
rect 1776 467 1812 508
rect 1702 451 1812 467
rect 1866 466 1902 508
rect 1702 417 1718 451
rect 1752 437 1812 451
rect 1854 450 1920 466
rect 1752 417 1768 437
rect 1702 401 1768 417
rect 1854 416 1870 450
rect 1904 416 1920 450
rect 1854 400 1920 416
rect 1582 353 1618 368
rect 1854 353 1884 400
rect 1432 323 1884 353
rect 1116 283 1182 299
rect 1283 294 1349 310
rect 891 236 958 252
rect 928 209 958 236
rect 1014 209 1044 283
rect 1283 260 1299 294
rect 1333 260 1349 294
rect 1283 244 1349 260
rect 1086 209 1116 235
rect 1283 222 1313 244
rect 1480 222 1510 323
rect 783 169 849 203
rect 783 135 799 169
rect 833 135 849 169
rect 381 87 411 113
rect 467 87 497 113
rect 545 87 575 113
rect 631 87 661 113
rect 783 101 849 135
rect 105 48 135 74
rect 183 48 213 74
rect 783 67 799 101
rect 833 67 849 101
rect 783 51 849 67
rect 928 51 958 125
rect 1014 99 1044 125
rect 1086 51 1116 125
rect 1726 181 1756 323
rect 1962 296 1998 508
rect 2065 364 2101 398
rect 2051 348 2117 364
rect 2051 314 2067 348
rect 2101 314 2117 348
rect 2051 298 2117 314
rect 2259 306 2295 392
rect 2451 360 2487 392
rect 1943 280 2009 296
rect 1828 235 1901 251
rect 1828 201 1851 235
rect 1885 201 1901 235
rect 1828 185 1901 201
rect 1943 246 1959 280
rect 1993 246 2009 280
rect 1943 230 2009 246
rect 1828 163 1858 185
rect 1943 163 1973 230
rect 2079 207 2109 298
rect 2229 290 2295 306
rect 2337 344 2403 360
rect 2337 310 2353 344
rect 2387 310 2403 344
rect 2337 294 2403 310
rect 2445 344 2511 360
rect 2445 310 2461 344
rect 2495 310 2511 344
rect 2445 294 2511 310
rect 2553 317 2589 508
rect 2637 476 2673 508
rect 2631 460 2697 476
rect 2631 426 2647 460
rect 2681 426 2697 460
rect 2631 410 2697 426
rect 2553 301 2619 317
rect 2229 256 2245 290
rect 2279 256 2295 290
rect 2229 252 2295 256
rect 2229 222 2331 252
rect 928 21 1116 51
rect 1283 48 1313 74
rect 1480 48 1510 74
rect 1726 71 1756 97
rect 2301 202 2331 222
rect 2373 202 2403 294
rect 1828 53 1858 79
rect 1943 53 1973 79
rect 2079 53 2109 79
rect 2468 158 2498 294
rect 2553 267 2569 301
rect 2603 267 2619 301
rect 2553 251 2619 267
rect 2667 203 2697 410
rect 2779 398 2815 464
rect 2546 173 2697 203
rect 2745 382 2815 398
rect 2745 348 2761 382
rect 2795 348 2815 382
rect 2745 336 2815 348
rect 2973 336 3009 368
rect 3063 336 3099 368
rect 3153 336 3189 368
rect 3243 336 3279 368
rect 2745 314 3279 336
rect 2745 280 2761 314
rect 2795 280 3279 314
rect 2745 279 3279 280
rect 2745 246 2815 279
rect 2974 264 3004 279
rect 3060 264 3090 279
rect 3160 264 3190 279
rect 3249 264 3279 279
rect 2745 212 2761 246
rect 2795 212 2815 246
rect 2745 196 2815 212
rect 2546 158 2576 173
rect 2776 158 2806 196
rect 2974 90 3004 116
rect 3060 90 3090 116
rect 3160 90 3190 116
rect 3249 90 3279 116
rect 2301 48 2331 74
rect 2373 48 2403 74
rect 2468 48 2498 74
rect 2546 48 2576 74
rect 2776 48 2806 74
<< polycont >>
rect 85 348 119 382
rect 85 280 119 314
rect 215 374 249 408
rect 215 306 249 340
rect 85 212 119 246
rect 323 280 357 314
rect 431 320 465 354
rect 561 320 595 354
rect 799 339 833 373
rect 799 271 833 305
rect 799 203 833 237
rect 907 252 941 286
rect 1024 299 1058 333
rect 1132 367 1166 401
rect 1448 373 1482 407
rect 1132 299 1166 333
rect 1718 417 1752 451
rect 1870 416 1904 450
rect 1299 260 1333 294
rect 799 135 833 169
rect 799 67 833 101
rect 2067 314 2101 348
rect 1851 201 1885 235
rect 1959 246 1993 280
rect 2353 310 2387 344
rect 2461 310 2495 344
rect 2647 426 2681 460
rect 2245 256 2279 290
rect 2569 267 2603 301
rect 2761 348 2795 382
rect 2761 280 2795 314
rect 2761 212 2795 246
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3360 683
rect 17 580 99 596
rect 17 546 49 580
rect 83 546 99 580
rect 17 510 99 546
rect 207 578 257 649
rect 207 544 223 578
rect 207 526 257 544
rect 291 581 461 615
rect 17 476 49 510
rect 83 492 99 510
rect 291 492 325 581
rect 83 476 325 492
rect 17 458 325 476
rect 359 520 393 547
rect 17 162 51 458
rect 359 424 393 486
rect 427 492 461 581
rect 495 577 545 649
rect 529 543 545 577
rect 495 526 545 543
rect 647 579 697 595
rect 647 545 663 579
rect 647 509 697 545
rect 647 492 663 509
rect 427 475 663 492
rect 427 458 697 475
rect 199 408 473 424
rect 85 382 165 398
rect 119 348 165 382
rect 85 314 165 348
rect 119 280 165 314
rect 85 246 165 280
rect 119 212 165 246
rect 85 196 165 212
rect 199 374 215 408
rect 249 390 473 408
rect 249 374 265 390
rect 199 340 265 374
rect 199 306 215 340
rect 249 306 265 340
rect 199 230 265 306
rect 307 314 373 356
rect 307 280 323 314
rect 357 280 373 314
rect 423 354 473 390
rect 423 320 431 354
rect 465 320 473 354
rect 423 304 473 320
rect 507 354 611 370
rect 507 350 561 354
rect 507 316 511 350
rect 545 320 561 350
rect 595 320 611 354
rect 545 316 611 320
rect 507 304 611 316
rect 307 264 373 280
rect 663 269 697 458
rect 570 235 697 269
rect 731 581 960 615
rect 731 579 787 581
rect 731 545 753 579
rect 731 509 787 545
rect 731 475 753 509
rect 731 459 787 475
rect 821 516 892 547
rect 821 482 858 516
rect 199 196 370 230
rect 320 172 370 196
rect 17 132 110 162
rect 17 98 60 132
rect 94 98 110 132
rect 17 68 110 98
rect 208 133 274 162
rect 208 99 224 133
rect 258 99 274 133
rect 320 138 336 172
rect 320 109 370 138
rect 406 172 472 201
rect 406 138 422 172
rect 456 138 472 172
rect 208 17 274 99
rect 406 17 472 138
rect 570 172 636 235
rect 731 201 765 459
rect 821 451 892 482
rect 926 485 960 581
rect 994 570 1044 649
rect 1028 536 1044 570
rect 994 519 1044 536
rect 1146 571 1212 587
rect 1146 537 1162 571
rect 1196 537 1212 571
rect 1146 501 1212 537
rect 1252 571 1318 649
rect 1252 537 1268 571
rect 1302 537 1318 571
rect 1252 535 1318 537
rect 1522 574 1588 649
rect 1522 540 1538 574
rect 1572 540 1588 574
rect 1522 535 1588 540
rect 1631 567 1766 596
rect 1631 533 1732 567
rect 1631 501 1766 533
rect 1800 567 1872 596
rect 1800 533 1822 567
rect 1856 533 1872 567
rect 1992 580 2058 649
rect 1992 546 2008 580
rect 2042 546 2058 580
rect 2199 580 2265 649
rect 2199 546 2215 580
rect 2249 546 2265 580
rect 2493 567 2579 596
rect 1800 504 1872 533
rect 2493 533 2509 567
rect 2543 533 2579 567
rect 1146 485 1162 501
rect 926 467 1162 485
rect 1196 467 1665 501
rect 926 451 1240 467
rect 821 417 855 451
rect 570 138 586 172
rect 620 138 636 172
rect 570 109 636 138
rect 670 185 765 201
rect 670 151 700 185
rect 734 151 765 185
rect 670 135 765 151
rect 799 401 1172 417
rect 799 383 1132 401
rect 799 373 855 383
rect 833 339 855 373
rect 1116 367 1132 383
rect 1166 367 1172 401
rect 799 305 855 339
rect 833 271 855 305
rect 991 333 1074 349
rect 799 237 855 271
rect 833 203 855 237
rect 889 286 957 302
rect 889 252 907 286
rect 941 252 957 286
rect 889 236 957 252
rect 991 299 1024 333
rect 1058 299 1074 333
rect 991 236 1074 299
rect 1116 333 1172 367
rect 1116 299 1132 333
rect 1166 299 1172 333
rect 1116 283 1172 299
rect 1206 249 1240 451
rect 1342 412 1498 433
rect 1342 378 1358 412
rect 1392 407 1498 412
rect 1392 378 1448 407
rect 1342 373 1448 378
rect 1482 373 1498 407
rect 1342 357 1498 373
rect 799 202 855 203
rect 1111 215 1240 249
rect 1291 294 1415 310
rect 1291 260 1299 294
rect 1333 260 1415 294
rect 1291 236 1415 260
rect 799 178 917 202
rect 799 169 883 178
rect 833 144 883 169
rect 833 135 917 144
rect 799 121 917 135
rect 953 178 1019 202
rect 953 144 969 178
rect 1003 144 1019 178
rect 799 101 855 121
rect 833 67 855 101
rect 799 51 855 67
rect 953 17 1019 144
rect 1111 184 1177 215
rect 1449 202 1483 357
rect 1544 330 1578 467
rect 1699 451 1766 467
rect 1699 433 1718 451
rect 1612 417 1718 433
rect 1752 417 1766 451
rect 1612 415 1766 417
rect 1612 381 1628 415
rect 1662 399 1766 415
rect 1662 381 1733 399
rect 1612 364 1733 381
rect 1544 296 1665 330
rect 1111 150 1127 184
rect 1161 150 1177 184
rect 1111 121 1177 150
rect 1222 141 1272 181
rect 1222 107 1238 141
rect 1222 17 1272 107
rect 1308 168 1324 202
rect 1358 168 1483 202
rect 1521 210 1571 226
rect 1555 176 1571 210
rect 1308 120 1374 168
rect 1308 86 1324 120
rect 1358 86 1374 120
rect 1308 70 1374 86
rect 1419 127 1485 134
rect 1419 93 1435 127
rect 1469 93 1485 127
rect 1419 17 1485 93
rect 1521 120 1571 176
rect 1555 86 1571 120
rect 1615 169 1665 296
rect 1615 135 1631 169
rect 1615 119 1665 135
rect 1521 85 1571 86
rect 1699 85 1733 364
rect 1800 360 1834 504
rect 1906 478 2459 512
rect 1906 466 1940 478
rect 1868 450 1940 466
rect 1868 416 1870 450
rect 1904 416 1940 450
rect 1868 400 1940 416
rect 2095 410 2111 444
rect 2145 410 2185 444
rect 2095 394 2185 410
rect 1767 348 2117 360
rect 1767 326 2067 348
rect 1767 169 1801 326
rect 2051 314 2067 326
rect 2101 314 2117 348
rect 2051 308 2117 314
rect 2151 306 2185 394
rect 2337 344 2391 360
rect 2337 310 2353 344
rect 2387 310 2391 344
rect 2151 290 2295 306
rect 1943 280 2009 281
rect 1767 119 1801 135
rect 1835 235 1901 251
rect 1943 246 1959 280
rect 1993 274 2009 280
rect 2151 274 2245 290
rect 1993 256 2245 274
rect 2279 256 2295 290
rect 1993 246 2295 256
rect 1943 240 2295 246
rect 2337 272 2391 310
rect 2425 351 2459 478
rect 2493 385 2579 533
rect 2667 580 2775 649
rect 2667 546 2704 580
rect 2738 546 2775 580
rect 2667 530 2775 546
rect 2809 580 2879 596
rect 2809 546 2825 580
rect 2859 546 2879 580
rect 2809 510 2879 546
rect 2809 476 2825 510
rect 2859 476 2879 510
rect 2809 470 2879 476
rect 2631 460 2879 470
rect 2631 426 2647 460
rect 2681 436 2879 460
rect 2681 426 2697 436
rect 2631 419 2697 426
rect 2745 385 2811 398
rect 2545 382 2811 385
rect 2545 351 2761 382
rect 2425 344 2511 351
rect 2425 310 2461 344
rect 2495 310 2511 344
rect 2653 348 2761 351
rect 2795 348 2811 382
rect 2425 306 2511 310
rect 2553 301 2619 317
rect 2553 272 2569 301
rect 2337 267 2569 272
rect 2603 267 2619 301
rect 1835 201 1851 235
rect 1885 206 1901 235
rect 1885 201 2086 206
rect 1835 172 2086 201
rect 1835 85 1901 172
rect 1521 51 1901 85
rect 1968 122 2018 138
rect 1968 88 1984 122
rect 1968 17 2018 88
rect 2052 85 2086 172
rect 2120 182 2154 240
rect 2337 238 2619 267
rect 2653 314 2811 348
rect 2653 280 2761 314
rect 2795 280 2811 314
rect 2653 246 2811 280
rect 2337 206 2371 238
rect 2120 119 2154 148
rect 2188 172 2371 206
rect 2653 212 2761 246
rect 2795 212 2811 246
rect 2653 204 2811 212
rect 2407 198 2811 204
rect 2188 85 2222 172
rect 2407 170 2687 198
rect 2745 196 2811 198
rect 2845 356 2879 436
rect 2913 580 2979 649
rect 2913 546 2929 580
rect 2963 546 2979 580
rect 2913 506 2979 546
rect 2913 472 2929 506
rect 2963 472 2979 506
rect 2913 424 2979 472
rect 2913 390 2929 424
rect 2963 390 2979 424
rect 3013 580 3057 596
rect 3013 546 3019 580
rect 3053 546 3057 580
rect 3013 506 3057 546
rect 3013 472 3019 506
rect 3053 472 3057 506
rect 3013 430 3057 472
rect 3093 580 3159 649
rect 3093 546 3109 580
rect 3143 546 3159 580
rect 3093 498 3159 546
rect 3093 464 3109 498
rect 3143 464 3159 498
rect 3194 580 3237 596
rect 3194 546 3199 580
rect 3233 546 3237 580
rect 3194 506 3237 546
rect 3194 472 3199 506
rect 3233 472 3237 506
rect 3194 430 3237 472
rect 3273 580 3339 649
rect 3273 546 3289 580
rect 3323 546 3339 580
rect 3273 498 3339 546
rect 3273 464 3289 498
rect 3323 464 3339 498
rect 3013 414 3335 430
rect 3013 380 3019 414
rect 3053 380 3199 414
rect 3233 380 3335 414
rect 3013 364 3335 380
rect 2845 350 2951 356
rect 2845 316 2911 350
rect 2945 316 2951 350
rect 2845 310 2951 316
rect 2052 51 2222 85
rect 2256 121 2306 138
rect 2290 87 2306 121
rect 2256 17 2306 87
rect 2407 133 2473 170
rect 2845 162 2879 310
rect 3033 268 3335 364
rect 2407 99 2423 133
rect 2457 99 2473 133
rect 2407 70 2473 99
rect 2571 120 2767 136
rect 2571 86 2587 120
rect 2621 86 2717 120
rect 2751 86 2767 120
rect 2571 17 2767 86
rect 2801 133 2879 162
rect 2801 99 2817 133
rect 2851 99 2879 133
rect 2801 70 2879 99
rect 2913 252 2979 268
rect 2913 218 2929 252
rect 2963 218 2979 252
rect 2913 162 2979 218
rect 2913 128 2929 162
rect 2963 128 2979 162
rect 2913 17 2979 128
rect 3015 252 3335 268
rect 3049 218 3202 252
rect 3236 218 3335 252
rect 3015 162 3065 218
rect 3049 128 3065 162
rect 3015 112 3065 128
rect 3099 165 3165 184
rect 3099 131 3115 165
rect 3149 131 3165 165
rect 3099 17 3165 131
rect 3199 165 3240 218
rect 3199 131 3202 165
rect 3236 131 3240 165
rect 3199 115 3240 131
rect 3274 165 3340 184
rect 3274 131 3290 165
rect 3324 131 3340 165
rect 3274 17 3340 131
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3360 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 3199 649 3233 683
rect 3295 649 3329 683
rect 511 316 545 350
rect 2911 316 2945 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
<< metal1 >>
rect 0 683 3360 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3360 683
rect 0 617 3360 649
rect 499 350 557 356
rect 499 316 511 350
rect 545 347 557 350
rect 2899 350 2957 356
rect 2899 347 2911 350
rect 545 319 2911 347
rect 545 316 557 319
rect 499 310 557 316
rect 2899 316 2911 319
rect 2945 316 2957 350
rect 2899 310 2957 316
rect 0 17 3360 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3360 17
rect 0 -49 3360 -17
<< labels >>
flabel pwell s 0 0 3360 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 0 617 3360 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
rlabel comment s 0 0 0 0 4 sedfxtp_4
flabel comment s 1663 341 1663 341 0 FreeSans 200 0 0 0 no_jumper_check
flabel metal1 s 0 617 3360 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 3360 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 895 242 929 276 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 1375 242 1409 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 127 242 161 276 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 DE
port 3 nsew
flabel corelocali s 991 242 1025 276 0 FreeSans 340 0 0 0 SCD
port 4 nsew
flabel corelocali s 3295 242 3329 276 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 3295 316 3329 350 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 3295 390 3329 424 0 FreeSans 340 0 0 0 Q
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 3360 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 492310
string GDS_START 469782
<< end >>
