magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 123 378 189 547
rect 318 378 455 430
rect 123 344 455 378
rect 23 236 89 310
rect 123 202 157 344
rect 191 236 263 310
rect 305 236 371 310
rect 123 70 366 202
rect 409 88 505 310
rect 553 236 647 310
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 23 581 289 615
rect 23 364 89 581
rect 223 498 289 581
rect 335 532 469 649
rect 503 498 559 596
rect 223 464 559 498
rect 223 412 284 464
rect 493 364 559 464
rect 599 364 649 649
rect 23 17 89 202
rect 578 17 644 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel locali s 305 236 371 310 6 A1
port 1 nsew signal input
rlabel locali s 409 88 505 310 6 A2
port 2 nsew signal input
rlabel locali s 553 236 647 310 6 A3
port 3 nsew signal input
rlabel locali s 191 236 263 310 6 B1
port 4 nsew signal input
rlabel locali s 23 236 89 310 6 B2
port 5 nsew signal input
rlabel locali s 318 378 455 430 6 Y
port 6 nsew signal output
rlabel locali s 123 378 189 547 6 Y
port 6 nsew signal output
rlabel locali s 123 344 455 378 6 Y
port 6 nsew signal output
rlabel locali s 123 202 157 344 6 Y
port 6 nsew signal output
rlabel locali s 123 70 366 202 6 Y
port 6 nsew signal output
rlabel metal1 s 0 -49 672 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 617 672 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3823500
string GDS_START 3816974
<< end >>
