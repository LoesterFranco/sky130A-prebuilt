magic
tech sky130A
magscale 1 2
timestamp 1604502693
<< nwell >>
rect -38 261 3350 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 157 47 187 177
rect 241 47 271 177
rect 325 47 355 177
rect 409 47 439 177
rect 561 47 591 177
rect 645 47 675 177
rect 729 47 759 177
rect 813 47 843 177
rect 897 47 927 177
rect 981 47 1011 177
rect 1065 47 1095 177
rect 1149 47 1179 177
rect 1233 47 1263 177
rect 1317 47 1347 177
rect 1401 47 1431 177
rect 1485 47 1515 177
rect 1569 47 1599 177
rect 1653 47 1683 177
rect 1737 47 1767 177
rect 1821 47 1851 177
rect 1905 47 1935 177
rect 1989 47 2019 177
rect 2073 47 2103 177
rect 2157 47 2187 177
rect 2241 47 2271 177
rect 2325 47 2355 177
rect 2409 47 2439 177
rect 2493 47 2523 177
rect 2577 47 2607 177
rect 2661 47 2691 177
rect 2745 47 2775 177
rect 2829 47 2859 177
rect 2913 47 2943 177
rect 2997 47 3027 177
rect 3081 47 3111 177
rect 3165 47 3195 177
<< pmoshvt >>
rect 113 297 143 497
rect 197 297 227 497
rect 281 297 311 497
rect 365 297 395 497
rect 561 297 591 497
rect 645 297 675 497
rect 729 297 759 497
rect 813 297 843 497
rect 897 297 927 497
rect 981 297 1011 497
rect 1065 297 1095 497
rect 1149 297 1179 497
rect 1233 297 1263 497
rect 1317 297 1347 497
rect 1401 297 1431 497
rect 1485 297 1515 497
rect 1569 297 1599 497
rect 1653 297 1683 497
rect 1737 297 1767 497
rect 1821 297 1851 497
rect 1905 297 1935 497
rect 1989 297 2019 497
rect 2073 297 2103 497
rect 2157 297 2187 497
rect 2241 297 2271 497
rect 2325 297 2355 497
rect 2409 297 2439 497
rect 2493 297 2523 497
rect 2577 297 2607 497
rect 2661 297 2691 497
rect 2745 297 2775 497
rect 2829 297 2859 497
rect 2913 297 2943 497
rect 2997 297 3027 497
rect 3081 297 3111 497
rect 3165 297 3195 497
<< ndiff >>
rect 105 163 157 177
rect 105 129 113 163
rect 147 129 157 163
rect 105 95 157 129
rect 105 61 113 95
rect 147 61 157 95
rect 105 47 157 61
rect 187 169 241 177
rect 187 135 197 169
rect 231 135 241 169
rect 187 101 241 135
rect 187 67 197 101
rect 231 67 241 101
rect 187 47 241 67
rect 271 163 325 177
rect 271 129 281 163
rect 315 129 325 163
rect 271 95 325 129
rect 271 61 281 95
rect 315 61 325 95
rect 271 47 325 61
rect 355 169 409 177
rect 355 135 365 169
rect 399 135 409 169
rect 355 101 409 135
rect 355 67 365 101
rect 399 67 409 101
rect 355 47 409 67
rect 439 163 561 177
rect 439 61 449 163
rect 551 61 561 163
rect 439 47 561 61
rect 591 163 645 177
rect 591 129 601 163
rect 635 129 645 163
rect 591 95 645 129
rect 591 61 601 95
rect 635 61 645 95
rect 591 47 645 61
rect 675 95 729 177
rect 675 61 685 95
rect 719 61 729 95
rect 675 47 729 61
rect 759 163 813 177
rect 759 129 769 163
rect 803 129 813 163
rect 759 95 813 129
rect 759 61 769 95
rect 803 61 813 95
rect 759 47 813 61
rect 843 95 897 177
rect 843 61 853 95
rect 887 61 897 95
rect 843 47 897 61
rect 927 163 981 177
rect 927 129 937 163
rect 971 129 981 163
rect 927 95 981 129
rect 927 61 937 95
rect 971 61 981 95
rect 927 47 981 61
rect 1011 95 1065 177
rect 1011 61 1021 95
rect 1055 61 1065 95
rect 1011 47 1065 61
rect 1095 163 1149 177
rect 1095 129 1105 163
rect 1139 129 1149 163
rect 1095 95 1149 129
rect 1095 61 1105 95
rect 1139 61 1149 95
rect 1095 47 1149 61
rect 1179 95 1233 177
rect 1179 61 1189 95
rect 1223 61 1233 95
rect 1179 47 1233 61
rect 1263 163 1317 177
rect 1263 129 1273 163
rect 1307 129 1317 163
rect 1263 95 1317 129
rect 1263 61 1273 95
rect 1307 61 1317 95
rect 1263 47 1317 61
rect 1347 95 1401 177
rect 1347 61 1357 95
rect 1391 61 1401 95
rect 1347 47 1401 61
rect 1431 163 1485 177
rect 1431 129 1441 163
rect 1475 129 1485 163
rect 1431 95 1485 129
rect 1431 61 1441 95
rect 1475 61 1485 95
rect 1431 47 1485 61
rect 1515 95 1569 177
rect 1515 61 1525 95
rect 1559 61 1569 95
rect 1515 47 1569 61
rect 1599 163 1653 177
rect 1599 129 1609 163
rect 1643 129 1653 163
rect 1599 95 1653 129
rect 1599 61 1609 95
rect 1643 61 1653 95
rect 1599 47 1653 61
rect 1683 95 1737 177
rect 1683 61 1693 95
rect 1727 61 1737 95
rect 1683 47 1737 61
rect 1767 163 1821 177
rect 1767 129 1777 163
rect 1811 129 1821 163
rect 1767 95 1821 129
rect 1767 61 1777 95
rect 1811 61 1821 95
rect 1767 47 1821 61
rect 1851 95 1905 177
rect 1851 61 1861 95
rect 1895 61 1905 95
rect 1851 47 1905 61
rect 1935 163 1989 177
rect 1935 129 1945 163
rect 1979 129 1989 163
rect 1935 95 1989 129
rect 1935 61 1945 95
rect 1979 61 1989 95
rect 1935 47 1989 61
rect 2019 95 2073 177
rect 2019 61 2029 95
rect 2063 61 2073 95
rect 2019 47 2073 61
rect 2103 163 2157 177
rect 2103 129 2113 163
rect 2147 129 2157 163
rect 2103 95 2157 129
rect 2103 61 2113 95
rect 2147 61 2157 95
rect 2103 47 2157 61
rect 2187 95 2241 177
rect 2187 61 2197 95
rect 2231 61 2241 95
rect 2187 47 2241 61
rect 2271 163 2325 177
rect 2271 129 2281 163
rect 2315 129 2325 163
rect 2271 95 2325 129
rect 2271 61 2281 95
rect 2315 61 2325 95
rect 2271 47 2325 61
rect 2355 95 2409 177
rect 2355 61 2365 95
rect 2399 61 2409 95
rect 2355 47 2409 61
rect 2439 163 2493 177
rect 2439 129 2449 163
rect 2483 129 2493 163
rect 2439 95 2493 129
rect 2439 61 2449 95
rect 2483 61 2493 95
rect 2439 47 2493 61
rect 2523 95 2577 177
rect 2523 61 2533 95
rect 2567 61 2577 95
rect 2523 47 2577 61
rect 2607 163 2661 177
rect 2607 129 2617 163
rect 2651 129 2661 163
rect 2607 95 2661 129
rect 2607 61 2617 95
rect 2651 61 2661 95
rect 2607 47 2661 61
rect 2691 95 2745 177
rect 2691 61 2701 95
rect 2735 61 2745 95
rect 2691 47 2745 61
rect 2775 163 2829 177
rect 2775 129 2785 163
rect 2819 129 2829 163
rect 2775 95 2829 129
rect 2775 61 2785 95
rect 2819 61 2829 95
rect 2775 47 2829 61
rect 2859 95 2913 177
rect 2859 61 2869 95
rect 2903 61 2913 95
rect 2859 47 2913 61
rect 2943 163 2997 177
rect 2943 129 2953 163
rect 2987 129 2997 163
rect 2943 95 2997 129
rect 2943 61 2953 95
rect 2987 61 2997 95
rect 2943 47 2997 61
rect 3027 95 3081 177
rect 3027 61 3037 95
rect 3071 61 3081 95
rect 3027 47 3081 61
rect 3111 163 3165 177
rect 3111 129 3121 163
rect 3155 129 3165 163
rect 3111 95 3165 129
rect 3111 61 3121 95
rect 3155 61 3165 95
rect 3111 47 3165 61
rect 3195 95 3247 177
rect 3195 61 3205 95
rect 3239 61 3247 95
rect 3195 47 3247 61
<< pdiff >>
rect 61 485 113 497
rect 61 451 69 485
rect 103 451 113 485
rect 61 417 113 451
rect 61 383 69 417
rect 103 383 113 417
rect 61 349 113 383
rect 61 315 69 349
rect 103 315 113 349
rect 61 297 113 315
rect 143 477 197 497
rect 143 443 153 477
rect 187 443 197 477
rect 143 409 197 443
rect 143 375 153 409
rect 187 375 197 409
rect 143 341 197 375
rect 143 307 153 341
rect 187 307 197 341
rect 143 297 197 307
rect 227 485 281 497
rect 227 451 237 485
rect 271 451 281 485
rect 227 415 281 451
rect 227 381 237 415
rect 271 381 281 415
rect 227 345 281 381
rect 227 311 237 345
rect 271 311 281 345
rect 227 297 281 311
rect 311 477 365 497
rect 311 443 321 477
rect 355 443 365 477
rect 311 409 365 443
rect 311 375 321 409
rect 355 375 365 409
rect 311 341 365 375
rect 311 307 321 341
rect 355 307 365 341
rect 311 297 365 307
rect 395 485 451 497
rect 395 451 405 485
rect 439 451 451 485
rect 395 415 451 451
rect 395 381 405 415
rect 439 381 451 415
rect 395 345 451 381
rect 395 311 405 345
rect 439 311 451 345
rect 395 297 451 311
rect 505 477 561 497
rect 505 443 517 477
rect 551 443 561 477
rect 505 409 561 443
rect 505 375 517 409
rect 551 375 561 409
rect 505 341 561 375
rect 505 307 517 341
rect 551 307 561 341
rect 505 297 561 307
rect 591 485 645 497
rect 591 451 601 485
rect 635 451 645 485
rect 591 417 645 451
rect 591 383 601 417
rect 635 383 645 417
rect 591 297 645 383
rect 675 477 729 497
rect 675 443 685 477
rect 719 443 729 477
rect 675 409 729 443
rect 675 375 685 409
rect 719 375 729 409
rect 675 341 729 375
rect 675 307 685 341
rect 719 307 729 341
rect 675 297 729 307
rect 759 485 813 497
rect 759 451 769 485
rect 803 451 813 485
rect 759 417 813 451
rect 759 383 769 417
rect 803 383 813 417
rect 759 297 813 383
rect 843 477 897 497
rect 843 443 853 477
rect 887 443 897 477
rect 843 409 897 443
rect 843 375 853 409
rect 887 375 897 409
rect 843 341 897 375
rect 843 307 853 341
rect 887 307 897 341
rect 843 297 897 307
rect 927 485 981 497
rect 927 451 937 485
rect 971 451 981 485
rect 927 417 981 451
rect 927 383 937 417
rect 971 383 981 417
rect 927 297 981 383
rect 1011 477 1065 497
rect 1011 443 1021 477
rect 1055 443 1065 477
rect 1011 409 1065 443
rect 1011 375 1021 409
rect 1055 375 1065 409
rect 1011 341 1065 375
rect 1011 307 1021 341
rect 1055 307 1065 341
rect 1011 297 1065 307
rect 1095 485 1149 497
rect 1095 451 1105 485
rect 1139 451 1149 485
rect 1095 417 1149 451
rect 1095 383 1105 417
rect 1139 383 1149 417
rect 1095 297 1149 383
rect 1179 477 1233 497
rect 1179 443 1189 477
rect 1223 443 1233 477
rect 1179 409 1233 443
rect 1179 375 1189 409
rect 1223 375 1233 409
rect 1179 341 1233 375
rect 1179 307 1189 341
rect 1223 307 1233 341
rect 1179 297 1233 307
rect 1263 485 1317 497
rect 1263 451 1273 485
rect 1307 451 1317 485
rect 1263 417 1317 451
rect 1263 383 1273 417
rect 1307 383 1317 417
rect 1263 297 1317 383
rect 1347 477 1401 497
rect 1347 443 1357 477
rect 1391 443 1401 477
rect 1347 409 1401 443
rect 1347 375 1357 409
rect 1391 375 1401 409
rect 1347 341 1401 375
rect 1347 307 1357 341
rect 1391 307 1401 341
rect 1347 297 1401 307
rect 1431 485 1485 497
rect 1431 451 1441 485
rect 1475 451 1485 485
rect 1431 417 1485 451
rect 1431 383 1441 417
rect 1475 383 1485 417
rect 1431 297 1485 383
rect 1515 477 1569 497
rect 1515 443 1525 477
rect 1559 443 1569 477
rect 1515 409 1569 443
rect 1515 375 1525 409
rect 1559 375 1569 409
rect 1515 341 1569 375
rect 1515 307 1525 341
rect 1559 307 1569 341
rect 1515 297 1569 307
rect 1599 485 1653 497
rect 1599 451 1609 485
rect 1643 451 1653 485
rect 1599 417 1653 451
rect 1599 383 1609 417
rect 1643 383 1653 417
rect 1599 297 1653 383
rect 1683 477 1737 497
rect 1683 443 1693 477
rect 1727 443 1737 477
rect 1683 409 1737 443
rect 1683 375 1693 409
rect 1727 375 1737 409
rect 1683 341 1737 375
rect 1683 307 1693 341
rect 1727 307 1737 341
rect 1683 297 1737 307
rect 1767 485 1821 497
rect 1767 451 1777 485
rect 1811 451 1821 485
rect 1767 417 1821 451
rect 1767 383 1777 417
rect 1811 383 1821 417
rect 1767 297 1821 383
rect 1851 477 1905 497
rect 1851 443 1861 477
rect 1895 443 1905 477
rect 1851 409 1905 443
rect 1851 375 1861 409
rect 1895 375 1905 409
rect 1851 341 1905 375
rect 1851 307 1861 341
rect 1895 307 1905 341
rect 1851 297 1905 307
rect 1935 409 1989 497
rect 1935 375 1945 409
rect 1979 375 1989 409
rect 1935 341 1989 375
rect 1935 307 1945 341
rect 1979 307 1989 341
rect 1935 297 1989 307
rect 2019 477 2073 497
rect 2019 443 2029 477
rect 2063 443 2073 477
rect 2019 409 2073 443
rect 2019 375 2029 409
rect 2063 375 2073 409
rect 2019 297 2073 375
rect 2103 409 2157 497
rect 2103 375 2113 409
rect 2147 375 2157 409
rect 2103 341 2157 375
rect 2103 307 2113 341
rect 2147 307 2157 341
rect 2103 297 2157 307
rect 2187 477 2241 497
rect 2187 443 2197 477
rect 2231 443 2241 477
rect 2187 409 2241 443
rect 2187 375 2197 409
rect 2231 375 2241 409
rect 2187 297 2241 375
rect 2271 409 2325 497
rect 2271 375 2281 409
rect 2315 375 2325 409
rect 2271 341 2325 375
rect 2271 307 2281 341
rect 2315 307 2325 341
rect 2271 297 2325 307
rect 2355 477 2409 497
rect 2355 443 2365 477
rect 2399 443 2409 477
rect 2355 409 2409 443
rect 2355 375 2365 409
rect 2399 375 2409 409
rect 2355 297 2409 375
rect 2439 409 2493 497
rect 2439 375 2449 409
rect 2483 375 2493 409
rect 2439 341 2493 375
rect 2439 307 2449 341
rect 2483 307 2493 341
rect 2439 297 2493 307
rect 2523 477 2577 497
rect 2523 443 2533 477
rect 2567 443 2577 477
rect 2523 409 2577 443
rect 2523 375 2533 409
rect 2567 375 2577 409
rect 2523 297 2577 375
rect 2607 409 2661 497
rect 2607 375 2617 409
rect 2651 375 2661 409
rect 2607 341 2661 375
rect 2607 307 2617 341
rect 2651 307 2661 341
rect 2607 297 2661 307
rect 2691 477 2745 497
rect 2691 443 2701 477
rect 2735 443 2745 477
rect 2691 409 2745 443
rect 2691 375 2701 409
rect 2735 375 2745 409
rect 2691 297 2745 375
rect 2775 409 2829 497
rect 2775 375 2785 409
rect 2819 375 2829 409
rect 2775 341 2829 375
rect 2775 307 2785 341
rect 2819 307 2829 341
rect 2775 297 2829 307
rect 2859 477 2913 497
rect 2859 443 2869 477
rect 2903 443 2913 477
rect 2859 409 2913 443
rect 2859 375 2869 409
rect 2903 375 2913 409
rect 2859 297 2913 375
rect 2943 409 2997 497
rect 2943 375 2953 409
rect 2987 375 2997 409
rect 2943 341 2997 375
rect 2943 307 2953 341
rect 2987 307 2997 341
rect 2943 297 2997 307
rect 3027 477 3081 497
rect 3027 443 3037 477
rect 3071 443 3081 477
rect 3027 409 3081 443
rect 3027 375 3037 409
rect 3071 375 3081 409
rect 3027 297 3081 375
rect 3111 409 3165 497
rect 3111 375 3121 409
rect 3155 375 3165 409
rect 3111 341 3165 375
rect 3111 307 3121 341
rect 3155 307 3165 341
rect 3111 297 3165 307
rect 3195 477 3249 497
rect 3195 443 3205 477
rect 3239 443 3249 477
rect 3195 409 3249 443
rect 3195 375 3205 409
rect 3239 375 3249 409
rect 3195 297 3249 375
<< ndiffc >>
rect 113 129 147 163
rect 113 61 147 95
rect 197 135 231 169
rect 197 67 231 101
rect 281 129 315 163
rect 281 61 315 95
rect 365 135 399 169
rect 365 67 399 101
rect 449 61 551 163
rect 601 129 635 163
rect 601 61 635 95
rect 685 61 719 95
rect 769 129 803 163
rect 769 61 803 95
rect 853 61 887 95
rect 937 129 971 163
rect 937 61 971 95
rect 1021 61 1055 95
rect 1105 129 1139 163
rect 1105 61 1139 95
rect 1189 61 1223 95
rect 1273 129 1307 163
rect 1273 61 1307 95
rect 1357 61 1391 95
rect 1441 129 1475 163
rect 1441 61 1475 95
rect 1525 61 1559 95
rect 1609 129 1643 163
rect 1609 61 1643 95
rect 1693 61 1727 95
rect 1777 129 1811 163
rect 1777 61 1811 95
rect 1861 61 1895 95
rect 1945 129 1979 163
rect 1945 61 1979 95
rect 2029 61 2063 95
rect 2113 129 2147 163
rect 2113 61 2147 95
rect 2197 61 2231 95
rect 2281 129 2315 163
rect 2281 61 2315 95
rect 2365 61 2399 95
rect 2449 129 2483 163
rect 2449 61 2483 95
rect 2533 61 2567 95
rect 2617 129 2651 163
rect 2617 61 2651 95
rect 2701 61 2735 95
rect 2785 129 2819 163
rect 2785 61 2819 95
rect 2869 61 2903 95
rect 2953 129 2987 163
rect 2953 61 2987 95
rect 3037 61 3071 95
rect 3121 129 3155 163
rect 3121 61 3155 95
rect 3205 61 3239 95
<< pdiffc >>
rect 69 451 103 485
rect 69 383 103 417
rect 69 315 103 349
rect 153 443 187 477
rect 153 375 187 409
rect 153 307 187 341
rect 237 451 271 485
rect 237 381 271 415
rect 237 311 271 345
rect 321 443 355 477
rect 321 375 355 409
rect 321 307 355 341
rect 405 451 439 485
rect 405 381 439 415
rect 405 311 439 345
rect 517 443 551 477
rect 517 375 551 409
rect 517 307 551 341
rect 601 451 635 485
rect 601 383 635 417
rect 685 443 719 477
rect 685 375 719 409
rect 685 307 719 341
rect 769 451 803 485
rect 769 383 803 417
rect 853 443 887 477
rect 853 375 887 409
rect 853 307 887 341
rect 937 451 971 485
rect 937 383 971 417
rect 1021 443 1055 477
rect 1021 375 1055 409
rect 1021 307 1055 341
rect 1105 451 1139 485
rect 1105 383 1139 417
rect 1189 443 1223 477
rect 1189 375 1223 409
rect 1189 307 1223 341
rect 1273 451 1307 485
rect 1273 383 1307 417
rect 1357 443 1391 477
rect 1357 375 1391 409
rect 1357 307 1391 341
rect 1441 451 1475 485
rect 1441 383 1475 417
rect 1525 443 1559 477
rect 1525 375 1559 409
rect 1525 307 1559 341
rect 1609 451 1643 485
rect 1609 383 1643 417
rect 1693 443 1727 477
rect 1693 375 1727 409
rect 1693 307 1727 341
rect 1777 451 1811 485
rect 1777 383 1811 417
rect 1861 443 1895 477
rect 1861 375 1895 409
rect 1861 307 1895 341
rect 1945 375 1979 409
rect 1945 307 1979 341
rect 2029 443 2063 477
rect 2029 375 2063 409
rect 2113 375 2147 409
rect 2113 307 2147 341
rect 2197 443 2231 477
rect 2197 375 2231 409
rect 2281 375 2315 409
rect 2281 307 2315 341
rect 2365 443 2399 477
rect 2365 375 2399 409
rect 2449 375 2483 409
rect 2449 307 2483 341
rect 2533 443 2567 477
rect 2533 375 2567 409
rect 2617 375 2651 409
rect 2617 307 2651 341
rect 2701 443 2735 477
rect 2701 375 2735 409
rect 2785 375 2819 409
rect 2785 307 2819 341
rect 2869 443 2903 477
rect 2869 375 2903 409
rect 2953 375 2987 409
rect 2953 307 2987 341
rect 3037 443 3071 477
rect 3037 375 3071 409
rect 3121 375 3155 409
rect 3121 307 3155 341
rect 3205 443 3239 477
rect 3205 375 3239 409
<< poly >>
rect 113 497 143 523
rect 197 497 227 523
rect 281 497 311 523
rect 365 497 395 523
rect 561 497 591 523
rect 645 497 675 523
rect 729 497 759 523
rect 813 497 843 523
rect 897 497 927 523
rect 981 497 1011 523
rect 1065 497 1095 523
rect 1149 497 1179 523
rect 1233 497 1263 523
rect 1317 497 1347 523
rect 1401 497 1431 523
rect 1485 497 1515 523
rect 1569 497 1599 523
rect 1653 497 1683 523
rect 1737 497 1767 523
rect 1821 497 1851 523
rect 1905 497 1935 523
rect 1989 497 2019 523
rect 2073 497 2103 523
rect 2157 497 2187 523
rect 2241 497 2271 523
rect 2325 497 2355 523
rect 2409 497 2439 523
rect 2493 497 2523 523
rect 2577 497 2607 523
rect 2661 497 2691 523
rect 2745 497 2775 523
rect 2829 497 2859 523
rect 2913 497 2943 523
rect 2997 497 3027 523
rect 3081 497 3111 523
rect 3165 497 3195 523
rect 113 265 143 297
rect 197 265 227 297
rect 281 265 311 297
rect 365 265 395 297
rect 561 265 591 297
rect 645 265 675 297
rect 729 265 759 297
rect 813 265 843 297
rect 897 265 927 297
rect 981 265 1011 297
rect 1065 265 1095 297
rect 1149 265 1179 297
rect 1233 265 1263 297
rect 1317 265 1347 297
rect 1401 265 1431 297
rect 1485 265 1515 297
rect 1569 265 1599 297
rect 1653 265 1683 297
rect 1737 265 1767 297
rect 1821 265 1851 297
rect 21 249 439 265
rect 21 215 31 249
rect 65 215 99 249
rect 133 215 439 249
rect 21 199 439 215
rect 157 177 187 199
rect 241 177 271 199
rect 325 177 355 199
rect 409 177 439 199
rect 561 249 1851 265
rect 561 215 577 249
rect 611 215 645 249
rect 679 215 713 249
rect 747 215 781 249
rect 815 215 849 249
rect 883 215 917 249
rect 951 215 985 249
rect 1019 215 1053 249
rect 1087 215 1121 249
rect 1155 215 1189 249
rect 1223 215 1257 249
rect 1291 215 1325 249
rect 1359 215 1393 249
rect 1427 215 1461 249
rect 1495 215 1529 249
rect 1563 215 1597 249
rect 1631 215 1665 249
rect 1699 215 1733 249
rect 1767 215 1801 249
rect 1835 215 1851 249
rect 561 199 1851 215
rect 561 177 591 199
rect 645 177 675 199
rect 729 177 759 199
rect 813 177 843 199
rect 897 177 927 199
rect 981 177 1011 199
rect 1065 177 1095 199
rect 1149 177 1179 199
rect 1233 177 1263 199
rect 1317 177 1347 199
rect 1401 177 1431 199
rect 1485 177 1515 199
rect 1569 177 1599 199
rect 1653 177 1683 199
rect 1737 177 1767 199
rect 1821 177 1851 199
rect 1905 265 1935 297
rect 1989 265 2019 297
rect 2073 265 2103 297
rect 2157 265 2187 297
rect 2241 265 2271 297
rect 2325 265 2355 297
rect 2409 265 2439 297
rect 2493 265 2523 297
rect 2577 265 2607 297
rect 2661 265 2691 297
rect 2745 265 2775 297
rect 2829 265 2859 297
rect 2913 265 2943 297
rect 2997 265 3027 297
rect 3081 265 3111 297
rect 3165 265 3195 297
rect 1905 249 3195 265
rect 1905 215 1921 249
rect 1955 215 1989 249
rect 2023 215 2057 249
rect 2091 215 2125 249
rect 2159 215 2193 249
rect 2227 215 2261 249
rect 2295 215 2329 249
rect 2363 215 2397 249
rect 2431 215 2465 249
rect 2499 215 2533 249
rect 2567 215 2601 249
rect 2635 215 2669 249
rect 2703 215 2737 249
rect 2771 215 2805 249
rect 2839 215 2873 249
rect 2907 215 2941 249
rect 2975 215 3009 249
rect 3043 215 3077 249
rect 3111 215 3195 249
rect 1905 199 3195 215
rect 1905 177 1935 199
rect 1989 177 2019 199
rect 2073 177 2103 199
rect 2157 177 2187 199
rect 2241 177 2271 199
rect 2325 177 2355 199
rect 2409 177 2439 199
rect 2493 177 2523 199
rect 2577 177 2607 199
rect 2661 177 2691 199
rect 2745 177 2775 199
rect 2829 177 2859 199
rect 2913 177 2943 199
rect 2997 177 3027 199
rect 3081 177 3111 199
rect 3165 177 3195 199
rect 157 21 187 47
rect 241 21 271 47
rect 325 21 355 47
rect 409 21 439 47
rect 561 21 591 47
rect 645 21 675 47
rect 729 21 759 47
rect 813 21 843 47
rect 897 21 927 47
rect 981 21 1011 47
rect 1065 21 1095 47
rect 1149 21 1179 47
rect 1233 21 1263 47
rect 1317 21 1347 47
rect 1401 21 1431 47
rect 1485 21 1515 47
rect 1569 21 1599 47
rect 1653 21 1683 47
rect 1737 21 1767 47
rect 1821 21 1851 47
rect 1905 21 1935 47
rect 1989 21 2019 47
rect 2073 21 2103 47
rect 2157 21 2187 47
rect 2241 21 2271 47
rect 2325 21 2355 47
rect 2409 21 2439 47
rect 2493 21 2523 47
rect 2577 21 2607 47
rect 2661 21 2691 47
rect 2745 21 2775 47
rect 2829 21 2859 47
rect 2913 21 2943 47
rect 2997 21 3027 47
rect 3081 21 3111 47
rect 3165 21 3195 47
<< polycont >>
rect 31 215 65 249
rect 99 215 133 249
rect 577 215 611 249
rect 645 215 679 249
rect 713 215 747 249
rect 781 215 815 249
rect 849 215 883 249
rect 917 215 951 249
rect 985 215 1019 249
rect 1053 215 1087 249
rect 1121 215 1155 249
rect 1189 215 1223 249
rect 1257 215 1291 249
rect 1325 215 1359 249
rect 1393 215 1427 249
rect 1461 215 1495 249
rect 1529 215 1563 249
rect 1597 215 1631 249
rect 1665 215 1699 249
rect 1733 215 1767 249
rect 1801 215 1835 249
rect 1921 215 1955 249
rect 1989 215 2023 249
rect 2057 215 2091 249
rect 2125 215 2159 249
rect 2193 215 2227 249
rect 2261 215 2295 249
rect 2329 215 2363 249
rect 2397 215 2431 249
rect 2465 215 2499 249
rect 2533 215 2567 249
rect 2601 215 2635 249
rect 2669 215 2703 249
rect 2737 215 2771 249
rect 2805 215 2839 249
rect 2873 215 2907 249
rect 2941 215 2975 249
rect 3009 215 3043 249
rect 3077 215 3111 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3157 561
rect 3191 527 3249 561
rect 3283 527 3312 561
rect 60 485 103 527
rect 60 451 69 485
rect 60 417 103 451
rect 60 383 69 417
rect 60 349 103 383
rect 60 315 69 349
rect 60 299 103 315
rect 137 477 203 493
rect 137 443 153 477
rect 187 443 203 477
rect 137 409 203 443
rect 137 375 153 409
rect 187 375 203 409
rect 137 341 203 375
rect 137 307 153 341
rect 187 307 203 341
rect 137 299 203 307
rect 17 249 133 265
rect 17 215 31 249
rect 65 215 99 249
rect 17 199 133 215
rect 167 257 203 299
rect 237 485 271 527
rect 237 415 271 451
rect 237 345 271 381
rect 237 291 271 311
rect 305 477 371 493
rect 305 443 321 477
rect 355 443 371 477
rect 305 409 371 443
rect 305 375 321 409
rect 355 375 371 409
rect 305 341 371 375
rect 305 307 321 341
rect 355 307 371 341
rect 305 257 371 307
rect 405 485 454 527
rect 439 451 454 485
rect 405 415 454 451
rect 439 381 454 415
rect 405 345 454 381
rect 439 311 454 345
rect 405 291 454 311
rect 495 477 559 493
rect 495 443 517 477
rect 551 443 559 477
rect 495 409 559 443
rect 495 375 517 409
rect 551 375 559 409
rect 495 341 559 375
rect 593 485 643 527
rect 593 451 601 485
rect 635 451 643 485
rect 593 417 643 451
rect 593 383 601 417
rect 635 383 643 417
rect 593 367 643 383
rect 677 477 727 493
rect 677 443 685 477
rect 719 443 727 477
rect 677 409 727 443
rect 677 375 685 409
rect 719 375 727 409
rect 495 307 517 341
rect 551 333 559 341
rect 677 341 727 375
rect 761 485 811 527
rect 761 451 769 485
rect 803 451 811 485
rect 761 417 811 451
rect 761 383 769 417
rect 803 383 811 417
rect 761 367 811 383
rect 845 477 895 493
rect 845 443 853 477
rect 887 443 895 477
rect 845 409 895 443
rect 845 375 853 409
rect 887 375 895 409
rect 677 333 685 341
rect 551 307 685 333
rect 719 333 727 341
rect 845 341 895 375
rect 929 485 979 527
rect 929 451 937 485
rect 971 451 979 485
rect 929 417 979 451
rect 929 383 937 417
rect 971 383 979 417
rect 929 367 979 383
rect 1013 477 1063 493
rect 1013 443 1021 477
rect 1055 443 1063 477
rect 1013 409 1063 443
rect 1013 375 1021 409
rect 1055 375 1063 409
rect 845 333 853 341
rect 719 307 853 333
rect 887 333 895 341
rect 1013 341 1063 375
rect 1097 485 1147 527
rect 1097 451 1105 485
rect 1139 451 1147 485
rect 1097 417 1147 451
rect 1097 383 1105 417
rect 1139 383 1147 417
rect 1097 367 1147 383
rect 1181 477 1231 493
rect 1181 443 1189 477
rect 1223 443 1231 477
rect 1181 409 1231 443
rect 1181 375 1189 409
rect 1223 375 1231 409
rect 1013 333 1021 341
rect 887 307 1021 333
rect 1055 333 1063 341
rect 1181 341 1231 375
rect 1265 485 1315 527
rect 1265 451 1273 485
rect 1307 451 1315 485
rect 1265 417 1315 451
rect 1265 383 1273 417
rect 1307 383 1315 417
rect 1265 367 1315 383
rect 1349 477 1399 493
rect 1349 443 1357 477
rect 1391 443 1399 477
rect 1349 409 1399 443
rect 1349 375 1357 409
rect 1391 375 1399 409
rect 1181 333 1189 341
rect 1055 307 1189 333
rect 1223 333 1231 341
rect 1349 341 1399 375
rect 1433 485 1483 527
rect 1433 451 1441 485
rect 1475 451 1483 485
rect 1433 417 1483 451
rect 1433 383 1441 417
rect 1475 383 1483 417
rect 1433 367 1483 383
rect 1517 477 1567 493
rect 1517 443 1525 477
rect 1559 443 1567 477
rect 1517 409 1567 443
rect 1517 375 1525 409
rect 1559 375 1567 409
rect 1349 333 1357 341
rect 1223 307 1357 333
rect 1391 333 1399 341
rect 1517 341 1567 375
rect 1601 485 1651 527
rect 1601 451 1609 485
rect 1643 451 1651 485
rect 1601 417 1651 451
rect 1601 383 1609 417
rect 1643 383 1651 417
rect 1601 367 1651 383
rect 1685 477 1735 493
rect 1685 443 1693 477
rect 1727 443 1735 477
rect 1685 409 1735 443
rect 1685 375 1693 409
rect 1727 375 1735 409
rect 1517 333 1525 341
rect 1391 307 1525 333
rect 1559 333 1567 341
rect 1685 341 1735 375
rect 1769 485 1819 527
rect 1769 451 1777 485
rect 1811 451 1819 485
rect 1769 417 1819 451
rect 1769 383 1777 417
rect 1811 383 1819 417
rect 1769 367 1819 383
rect 1853 477 3247 493
rect 1853 443 1861 477
rect 1895 459 2029 477
rect 1895 443 1903 459
rect 1853 409 1903 443
rect 2021 443 2029 459
rect 2063 459 2197 477
rect 2063 443 2071 459
rect 1853 375 1861 409
rect 1895 375 1903 409
rect 1685 333 1693 341
rect 1559 307 1693 333
rect 1727 333 1735 341
rect 1853 341 1903 375
rect 1853 333 1861 341
rect 1727 307 1861 333
rect 1895 307 1903 341
rect 495 291 1903 307
rect 1937 409 1987 425
rect 1937 375 1945 409
rect 1979 375 1987 409
rect 1937 341 1987 375
rect 2021 409 2071 443
rect 2189 443 2197 459
rect 2231 459 2365 477
rect 2231 443 2239 459
rect 2021 375 2029 409
rect 2063 375 2071 409
rect 2021 359 2071 375
rect 2105 409 2155 425
rect 2105 375 2113 409
rect 2147 375 2155 409
rect 1937 307 1945 341
rect 1979 325 1987 341
rect 2105 341 2155 375
rect 2189 409 2239 443
rect 2357 443 2365 459
rect 2399 459 2533 477
rect 2399 443 2407 459
rect 2189 375 2197 409
rect 2231 375 2239 409
rect 2189 359 2239 375
rect 2273 409 2323 425
rect 2273 375 2281 409
rect 2315 375 2323 409
rect 2105 325 2113 341
rect 1979 307 2113 325
rect 2147 325 2155 341
rect 2273 341 2323 375
rect 2357 409 2407 443
rect 2525 443 2533 459
rect 2567 459 2701 477
rect 2567 443 2575 459
rect 2357 375 2365 409
rect 2399 375 2407 409
rect 2357 359 2407 375
rect 2441 409 2491 425
rect 2441 375 2449 409
rect 2483 375 2491 409
rect 2273 325 2281 341
rect 2147 307 2281 325
rect 2315 325 2323 341
rect 2441 341 2491 375
rect 2525 409 2575 443
rect 2693 443 2701 459
rect 2735 459 2869 477
rect 2735 443 2743 459
rect 2525 375 2533 409
rect 2567 375 2575 409
rect 2525 359 2575 375
rect 2609 409 2659 425
rect 2609 375 2617 409
rect 2651 375 2659 409
rect 2441 325 2449 341
rect 2315 307 2449 325
rect 2483 325 2491 341
rect 2609 341 2659 375
rect 2693 409 2743 443
rect 2861 443 2869 459
rect 2903 459 3037 477
rect 2903 443 2911 459
rect 2693 375 2701 409
rect 2735 375 2743 409
rect 2693 359 2743 375
rect 2777 409 2827 425
rect 2777 375 2785 409
rect 2819 375 2827 409
rect 2609 325 2617 341
rect 2483 307 2617 325
rect 2651 325 2659 341
rect 2777 341 2827 375
rect 2861 409 2911 443
rect 3029 443 3037 459
rect 3071 459 3205 477
rect 3071 443 3079 459
rect 2861 375 2869 409
rect 2903 375 2911 409
rect 2861 359 2911 375
rect 2945 409 2995 425
rect 2945 375 2953 409
rect 2987 375 2995 409
rect 2777 325 2785 341
rect 2651 307 2785 325
rect 2819 325 2827 341
rect 2945 341 2995 375
rect 3029 409 3079 443
rect 3197 443 3205 459
rect 3239 443 3247 477
rect 3029 375 3037 409
rect 3071 375 3079 409
rect 3029 359 3079 375
rect 3113 409 3163 425
rect 3113 375 3121 409
rect 3155 375 3163 409
rect 2945 325 2953 341
rect 2819 307 2953 325
rect 2987 325 2995 341
rect 3113 341 3163 375
rect 3197 409 3247 443
rect 3197 375 3205 409
rect 3239 375 3247 409
rect 3197 359 3247 375
rect 3113 325 3121 341
rect 2987 307 3121 325
rect 3155 325 3163 341
rect 3155 307 3295 325
rect 1937 291 3295 307
rect 167 249 1856 257
rect 167 215 577 249
rect 611 215 645 249
rect 679 215 713 249
rect 747 215 781 249
rect 815 215 849 249
rect 883 215 917 249
rect 951 215 985 249
rect 1019 215 1053 249
rect 1087 215 1121 249
rect 1155 215 1189 249
rect 1223 215 1257 249
rect 1291 215 1325 249
rect 1359 215 1393 249
rect 1427 215 1461 249
rect 1495 215 1529 249
rect 1563 215 1597 249
rect 1631 215 1665 249
rect 1699 215 1733 249
rect 1767 215 1801 249
rect 1835 215 1856 249
rect 1890 249 3130 257
rect 1890 215 1921 249
rect 1955 215 1989 249
rect 2023 215 2057 249
rect 2091 215 2125 249
rect 2159 215 2193 249
rect 2227 215 2261 249
rect 2295 215 2329 249
rect 2363 215 2397 249
rect 2431 215 2465 249
rect 2499 215 2533 249
rect 2567 215 2601 249
rect 2635 215 2669 249
rect 2703 215 2737 249
rect 2771 215 2805 249
rect 2839 215 2873 249
rect 2907 215 2941 249
rect 2975 215 3009 249
rect 3043 215 3077 249
rect 3111 215 3130 249
rect 167 213 407 215
rect 17 51 63 199
rect 197 169 239 213
rect 97 163 163 165
rect 97 129 113 163
rect 147 129 163 163
rect 97 95 163 129
rect 97 61 113 95
rect 147 61 163 95
rect 97 17 163 61
rect 231 135 239 169
rect 197 101 239 135
rect 231 67 239 101
rect 197 51 239 67
rect 273 163 323 179
rect 273 129 281 163
rect 315 129 323 163
rect 273 95 323 129
rect 273 61 281 95
rect 315 61 323 95
rect 273 17 323 61
rect 357 169 407 213
rect 3164 181 3295 291
rect 357 135 365 169
rect 399 135 407 169
rect 357 101 407 135
rect 357 67 365 101
rect 399 67 407 101
rect 357 51 407 67
rect 441 163 551 181
rect 441 61 449 163
rect 441 17 551 61
rect 585 163 3295 181
rect 585 129 601 163
rect 635 145 769 163
rect 635 129 651 145
rect 585 95 651 129
rect 753 129 769 145
rect 803 145 937 163
rect 803 129 819 145
rect 585 61 601 95
rect 635 61 651 95
rect 585 51 651 61
rect 685 95 719 111
rect 685 17 719 61
rect 753 95 819 129
rect 921 129 937 145
rect 971 145 1105 163
rect 971 129 987 145
rect 753 61 769 95
rect 803 61 819 95
rect 753 51 819 61
rect 853 95 887 111
rect 853 17 887 61
rect 921 95 987 129
rect 1089 129 1105 145
rect 1139 145 1273 163
rect 1139 129 1155 145
rect 921 61 937 95
rect 971 61 987 95
rect 921 51 987 61
rect 1021 95 1055 111
rect 1021 17 1055 61
rect 1089 95 1155 129
rect 1257 129 1273 145
rect 1307 145 1441 163
rect 1307 129 1323 145
rect 1089 61 1105 95
rect 1139 61 1155 95
rect 1089 51 1155 61
rect 1189 95 1223 111
rect 1189 17 1223 61
rect 1257 95 1323 129
rect 1425 129 1441 145
rect 1475 145 1609 163
rect 1475 129 1491 145
rect 1257 61 1273 95
rect 1307 61 1323 95
rect 1257 51 1323 61
rect 1357 95 1391 111
rect 1357 17 1391 61
rect 1425 95 1491 129
rect 1593 129 1609 145
rect 1643 145 1777 163
rect 1643 129 1659 145
rect 1425 61 1441 95
rect 1475 61 1491 95
rect 1425 51 1491 61
rect 1525 95 1559 111
rect 1525 17 1559 61
rect 1593 95 1659 129
rect 1761 129 1777 145
rect 1811 145 1945 163
rect 1811 129 1827 145
rect 1593 61 1609 95
rect 1643 61 1659 95
rect 1593 51 1659 61
rect 1693 95 1727 111
rect 1693 17 1727 61
rect 1761 95 1827 129
rect 1929 129 1945 145
rect 1979 145 2113 163
rect 1979 129 1995 145
rect 1761 61 1777 95
rect 1811 61 1827 95
rect 1761 51 1827 61
rect 1861 95 1895 111
rect 1861 17 1895 61
rect 1929 95 1995 129
rect 2097 129 2113 145
rect 2147 145 2281 163
rect 2147 129 2163 145
rect 1929 61 1945 95
rect 1979 61 1995 95
rect 1929 51 1995 61
rect 2029 95 2063 111
rect 2029 17 2063 61
rect 2097 95 2163 129
rect 2265 129 2281 145
rect 2315 145 2449 163
rect 2315 129 2331 145
rect 2097 61 2113 95
rect 2147 61 2163 95
rect 2097 51 2163 61
rect 2197 95 2231 111
rect 2197 17 2231 61
rect 2265 95 2331 129
rect 2433 129 2449 145
rect 2483 145 2617 163
rect 2483 129 2499 145
rect 2265 61 2281 95
rect 2315 61 2331 95
rect 2265 51 2331 61
rect 2365 95 2399 111
rect 2365 17 2399 61
rect 2433 95 2499 129
rect 2601 129 2617 145
rect 2651 145 2785 163
rect 2651 129 2667 145
rect 2433 61 2449 95
rect 2483 61 2499 95
rect 2433 51 2499 61
rect 2533 95 2567 111
rect 2533 17 2567 61
rect 2601 95 2667 129
rect 2769 129 2785 145
rect 2819 145 2953 163
rect 2819 129 2835 145
rect 2601 61 2617 95
rect 2651 61 2667 95
rect 2601 51 2667 61
rect 2701 95 2735 111
rect 2701 17 2735 61
rect 2769 95 2835 129
rect 2937 129 2953 145
rect 2987 145 3121 163
rect 2987 129 3003 145
rect 2769 61 2785 95
rect 2819 61 2835 95
rect 2769 51 2835 61
rect 2869 95 2903 111
rect 2869 17 2903 61
rect 2937 95 3003 129
rect 3105 129 3121 145
rect 3155 145 3295 163
rect 3155 129 3171 145
rect 2937 61 2953 95
rect 2987 61 3003 95
rect 2937 51 3003 61
rect 3037 95 3071 111
rect 3037 17 3071 61
rect 3105 95 3171 129
rect 3105 61 3121 95
rect 3155 61 3171 95
rect 3105 51 3171 61
rect 3205 95 3259 111
rect 3239 61 3259 95
rect 3205 17 3259 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3312 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 2881 527 2915 561
rect 2973 527 3007 561
rect 3065 527 3099 561
rect 3157 527 3191 561
rect 3249 527 3283 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
rect 2881 -17 2915 17
rect 2973 -17 3007 17
rect 3065 -17 3099 17
rect 3157 -17 3191 17
rect 3249 -17 3283 17
<< metal1 >>
rect 0 561 3312 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3157 561
rect 3191 527 3249 561
rect 3283 527 3312 561
rect 0 496 3312 527
rect 0 17 3312 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3312 17
rect 0 -48 3312 -17
<< labels >>
flabel corelocali s 59 221 93 255 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 3194 289 3228 323 0 FreeSans 400 0 0 0 X
port 7 nsew
flabel corelocali s 2499 221 2533 255 0 FreeSans 400 0 0 0 SLEEP
port 2 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew
rlabel comment s 0 0 0 0 4 lpflow_isobufsrc_16
<< properties >>
string FIXED_BBOX 0 0 3312 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2363660
string GDS_START 2340052
string path 0.000 0.000 82.800 0.000 
<< end >>
