magic
tech sky130A
magscale 1 2
timestamp 1599588218
<< nwell >>
rect -38 332 806 704
<< pwell >>
rect 0 0 768 49
<< scpmos >>
rect 84 424 120 592
rect 322 368 358 536
rect 431 368 467 536
rect 522 368 558 536
rect 639 368 675 592
<< nmoslvt >>
rect 84 74 114 184
rect 323 94 353 222
rect 401 94 431 222
rect 509 94 539 222
rect 652 74 682 222
<< ndiff >>
rect 266 210 323 222
rect 27 146 84 184
rect 27 112 39 146
rect 73 112 84 146
rect 27 74 84 112
rect 114 146 185 184
rect 114 112 139 146
rect 173 112 185 146
rect 114 74 185 112
rect 266 176 278 210
rect 312 176 323 210
rect 266 140 323 176
rect 266 106 278 140
rect 312 106 323 140
rect 266 94 323 106
rect 353 94 401 222
rect 431 94 509 222
rect 539 176 652 222
rect 539 142 550 176
rect 584 142 652 176
rect 539 116 652 142
rect 539 94 607 116
rect 581 82 607 94
rect 641 82 652 116
rect 581 74 652 82
rect 682 210 739 222
rect 682 176 693 210
rect 727 176 739 210
rect 682 120 739 176
rect 682 86 693 120
rect 727 86 739 120
rect 682 74 739 86
<< pdiff >>
rect 27 580 84 592
rect 27 546 39 580
rect 73 546 84 580
rect 27 470 84 546
rect 27 436 39 470
rect 73 436 84 470
rect 27 424 84 436
rect 120 580 185 592
rect 120 546 139 580
rect 173 546 185 580
rect 120 470 185 546
rect 573 536 639 592
rect 120 436 139 470
rect 173 436 185 470
rect 120 424 185 436
rect 266 524 322 536
rect 266 490 278 524
rect 312 490 322 524
rect 266 414 322 490
rect 266 380 278 414
rect 312 380 322 414
rect 266 368 322 380
rect 358 508 431 536
rect 358 474 378 508
rect 412 474 431 508
rect 358 368 431 474
rect 467 524 522 536
rect 467 490 478 524
rect 512 490 522 524
rect 467 440 522 490
rect 467 406 478 440
rect 512 406 522 440
rect 467 368 522 406
rect 558 524 639 536
rect 558 490 585 524
rect 619 490 639 524
rect 558 440 639 490
rect 558 406 585 440
rect 619 406 639 440
rect 558 368 639 406
rect 675 580 731 592
rect 675 546 685 580
rect 719 546 731 580
rect 675 497 731 546
rect 675 463 685 497
rect 719 463 731 497
rect 675 414 731 463
rect 675 380 685 414
rect 719 380 731 414
rect 675 368 731 380
<< ndiffc >>
rect 39 112 73 146
rect 139 112 173 146
rect 278 176 312 210
rect 278 106 312 140
rect 550 142 584 176
rect 607 82 641 116
rect 693 176 727 210
rect 693 86 727 120
<< pdiffc >>
rect 39 546 73 580
rect 39 436 73 470
rect 139 546 173 580
rect 139 436 173 470
rect 278 490 312 524
rect 278 380 312 414
rect 378 474 412 508
rect 478 490 512 524
rect 478 406 512 440
rect 585 490 619 524
rect 585 406 619 440
rect 685 546 719 580
rect 685 463 719 497
rect 685 380 719 414
<< poly >>
rect 84 592 120 618
rect 639 592 675 618
rect 322 536 358 562
rect 431 536 467 562
rect 522 536 558 562
rect 84 388 120 424
rect 84 356 114 388
rect 48 340 114 356
rect 48 306 64 340
rect 98 306 114 340
rect 48 272 114 306
rect 48 238 64 272
rect 98 238 114 272
rect 48 222 114 238
rect 84 184 114 222
rect 162 324 228 340
rect 162 290 178 324
rect 212 290 228 324
rect 162 267 228 290
rect 322 267 358 368
rect 431 336 467 368
rect 522 336 558 368
rect 401 320 467 336
rect 401 286 417 320
rect 451 286 467 320
rect 401 270 467 286
rect 509 320 575 336
rect 639 326 675 368
rect 509 286 525 320
rect 559 286 575 320
rect 509 270 575 286
rect 617 310 683 326
rect 617 276 633 310
rect 667 276 683 310
rect 162 256 353 267
rect 162 222 178 256
rect 212 237 353 256
rect 212 222 228 237
rect 323 222 353 237
rect 401 222 431 270
rect 509 222 539 270
rect 617 260 683 276
rect 652 222 682 260
rect 162 206 228 222
rect 84 48 114 74
rect 323 68 353 94
rect 401 68 431 94
rect 509 68 539 94
rect 652 48 682 74
<< polycont >>
rect 64 306 98 340
rect 64 238 98 272
rect 178 290 212 324
rect 417 286 451 320
rect 525 286 559 320
rect 633 276 667 310
rect 178 222 212 256
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 23 580 89 649
rect 23 546 39 580
rect 73 546 89 580
rect 23 470 89 546
rect 23 436 39 470
rect 73 436 89 470
rect 23 420 89 436
rect 123 580 189 596
rect 123 546 139 580
rect 173 546 189 580
rect 123 470 189 546
rect 123 436 139 470
rect 173 436 189 470
rect 123 420 189 436
rect 25 340 114 356
rect 25 306 64 340
rect 98 306 114 340
rect 25 272 114 306
rect 25 238 64 272
rect 98 238 114 272
rect 25 222 114 238
rect 155 340 189 420
rect 262 524 328 540
rect 262 490 278 524
rect 312 490 328 524
rect 262 424 328 490
rect 362 508 428 649
rect 362 474 378 508
rect 412 474 428 508
rect 362 458 428 474
rect 462 524 528 540
rect 462 490 478 524
rect 512 490 528 524
rect 462 440 528 490
rect 462 424 478 440
rect 262 414 478 424
rect 262 380 278 414
rect 312 406 478 414
rect 512 406 528 440
rect 312 390 528 406
rect 569 524 635 649
rect 569 490 585 524
rect 619 490 635 524
rect 569 440 635 490
rect 569 406 585 440
rect 619 406 635 440
rect 569 390 635 406
rect 669 580 751 596
rect 669 546 685 580
rect 719 546 751 580
rect 669 497 751 546
rect 669 463 685 497
rect 719 463 751 497
rect 669 414 751 463
rect 312 380 328 390
rect 155 324 228 340
rect 155 290 178 324
rect 212 290 228 324
rect 155 256 228 290
rect 155 222 178 256
rect 212 222 228 256
rect 155 206 228 222
rect 262 244 328 380
rect 669 380 685 414
rect 719 380 751 414
rect 669 364 751 380
rect 401 320 467 356
rect 401 286 417 320
rect 451 286 467 320
rect 401 278 467 286
rect 505 320 575 356
rect 505 286 525 320
rect 559 286 575 320
rect 505 278 575 286
rect 609 310 683 326
rect 609 276 633 310
rect 667 276 683 310
rect 609 260 683 276
rect 609 244 643 260
rect 262 210 643 244
rect 717 226 751 364
rect 677 210 751 226
rect 155 188 189 206
rect 23 146 89 188
rect 23 112 39 146
rect 73 112 89 146
rect 23 17 89 112
rect 123 146 189 188
rect 123 112 139 146
rect 173 112 189 146
rect 123 70 189 112
rect 262 176 278 210
rect 312 176 328 210
rect 677 176 693 210
rect 727 176 751 210
rect 262 140 328 176
rect 262 106 278 140
rect 312 106 328 140
rect 262 90 328 106
rect 525 142 550 176
rect 584 142 643 176
rect 525 116 643 142
rect 525 82 607 116
rect 641 82 643 116
rect 525 17 643 82
rect 677 120 751 176
rect 677 86 693 120
rect 727 86 751 120
rect 677 70 751 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
rlabel comment s 0 0 0 0 4 and3b_1
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 703 390 737 424 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 703 464 737 498 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 703 538 737 572 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 A_N
port 1 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 B
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 768 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3137048
string GDS_START 3130228
<< end >>
