magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 644 561
rect 103 379 179 527
rect 282 451 455 527
rect 17 199 65 277
rect 557 339 627 493
rect 389 289 627 339
rect 473 169 523 289
rect 557 215 627 255
rect 103 17 169 97
rect 290 17 356 97
rect 473 119 539 169
rect 0 -17 644 17
<< obsli1 >>
rect 17 345 69 493
rect 214 417 248 493
rect 489 417 523 493
rect 214 373 523 417
rect 17 311 179 345
rect 99 255 179 311
rect 214 289 355 373
rect 99 199 407 255
rect 99 165 168 199
rect 17 131 168 165
rect 203 131 439 165
rect 17 51 69 131
rect 203 51 256 131
rect 390 85 439 131
rect 573 85 627 155
rect 390 51 627 85
<< metal1 >>
rect 0 496 644 592
rect 0 -48 644 48
<< labels >>
rlabel locali s 557 215 627 255 6 A
port 1 nsew signal input
rlabel locali s 17 199 65 277 6 TE_B
port 2 nsew signal input
rlabel locali s 557 339 627 493 6 Z
port 3 nsew signal output
rlabel locali s 473 169 523 289 6 Z
port 3 nsew signal output
rlabel locali s 473 119 539 169 6 Z
port 3 nsew signal output
rlabel locali s 389 289 627 339 6 Z
port 3 nsew signal output
rlabel locali s 290 17 356 97 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 103 17 169 97 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 644 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 644 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 282 451 455 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 103 379 179 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 644 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 644 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2900138
string GDS_START 2893852
<< end >>
