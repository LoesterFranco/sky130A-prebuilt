magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 644 561
rect 17 165 69 490
rect 419 437 485 527
rect 197 199 257 323
rect 291 199 357 323
rect 391 199 455 323
rect 489 199 559 323
rect 17 131 385 165
rect 71 17 137 96
rect 171 60 211 131
rect 245 17 311 97
rect 345 62 385 131
rect 419 17 485 165
rect 0 -17 644 17
<< obsli1 >>
rect 105 359 627 401
rect 105 199 149 359
rect 593 165 627 359
rect 532 131 627 165
rect 532 81 566 131
<< metal1 >>
rect 0 496 644 592
rect 0 -48 644 48
<< labels >>
rlabel locali s 391 199 455 323 6 A
port 1 nsew signal input
rlabel locali s 291 199 357 323 6 B
port 2 nsew signal input
rlabel locali s 197 199 257 323 6 C
port 3 nsew signal input
rlabel locali s 489 199 559 323 6 D_N
port 4 nsew signal input
rlabel locali s 345 62 385 131 6 Y
port 5 nsew signal output
rlabel locali s 171 60 211 131 6 Y
port 5 nsew signal output
rlabel locali s 17 165 69 490 6 Y
port 5 nsew signal output
rlabel locali s 17 131 385 165 6 Y
port 5 nsew signal output
rlabel locali s 419 17 485 165 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 245 17 311 97 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 71 17 137 96 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 644 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 644 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 419 437 485 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 644 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 644 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1168196
string GDS_START 1162990
<< end >>
