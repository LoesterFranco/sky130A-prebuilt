magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1656 561
rect 103 451 169 527
rect 29 195 65 349
rect 201 289 278 323
rect 244 257 278 289
rect 167 153 247 219
rect 519 411 565 527
rect 103 17 169 93
rect 204 79 247 153
rect 482 203 523 264
rect 448 143 523 203
rect 557 143 615 264
rect 490 17 556 109
rect 951 401 1020 527
rect 949 143 1023 279
rect 959 17 1025 109
rect 1403 367 1437 527
rect 1471 367 1553 491
rect 1225 249 1293 329
rect 1491 299 1553 367
rect 1587 299 1637 527
rect 1327 215 1389 265
rect 1307 199 1389 215
rect 1307 75 1369 199
rect 1403 17 1453 163
rect 1519 145 1553 299
rect 1487 53 1553 145
rect 1587 17 1638 177
rect 0 -17 1656 17
<< obsli1 >>
rect 35 417 69 475
rect 282 425 397 459
rect 431 425 448 459
rect 35 391 133 417
rect 35 383 305 391
rect 99 357 305 383
rect 339 357 380 391
rect 99 161 133 357
rect 312 315 380 357
rect 34 127 133 161
rect 312 207 346 315
rect 414 281 448 425
rect 661 425 673 459
rect 707 425 764 459
rect 594 357 663 391
rect 713 362 764 425
rect 629 332 663 357
rect 629 298 683 332
rect 34 69 69 127
rect 281 141 346 207
rect 380 247 448 281
rect 649 278 683 298
rect 380 107 414 247
rect 649 212 696 278
rect 294 73 414 107
rect 649 93 683 212
rect 730 135 764 362
rect 597 59 683 93
rect 717 69 764 135
rect 798 425 857 459
rect 891 425 903 459
rect 798 69 836 425
rect 1065 431 1255 465
rect 879 347 917 379
rect 1065 347 1099 431
rect 1305 425 1317 459
rect 1351 425 1369 459
rect 879 313 1099 347
rect 879 117 913 313
rect 879 51 920 117
rect 1065 93 1099 313
rect 1133 391 1191 397
rect 1167 357 1191 391
rect 1133 207 1191 357
rect 1335 333 1369 425
rect 1335 299 1457 333
rect 1423 265 1457 299
rect 1133 141 1257 207
rect 1423 199 1485 265
rect 1065 59 1244 93
<< obsli1c >>
rect 397 425 431 459
rect 305 357 339 391
rect 673 425 707 459
rect 857 425 891 459
rect 1317 425 1351 459
rect 1133 357 1167 391
<< metal1 >>
rect 0 496 1656 592
rect 17 320 75 329
rect 201 320 259 329
rect 1213 320 1271 329
rect 17 292 1271 320
rect 17 283 75 292
rect 201 283 259 292
rect 1213 283 1271 292
rect 0 -48 1656 48
<< obsm1 >>
rect 385 459 443 465
rect 385 425 397 459
rect 431 456 443 459
rect 661 459 719 465
rect 661 456 673 459
rect 431 428 673 456
rect 431 425 443 428
rect 385 419 443 425
rect 661 425 673 428
rect 707 425 719 459
rect 661 419 719 425
rect 845 459 903 465
rect 845 425 857 459
rect 891 456 903 459
rect 1305 459 1363 465
rect 1305 456 1317 459
rect 891 428 1317 456
rect 891 425 903 428
rect 845 419 903 425
rect 1305 425 1317 428
rect 1351 425 1363 459
rect 1305 419 1363 425
rect 293 391 351 397
rect 293 357 305 391
rect 339 388 351 391
rect 1121 391 1179 397
rect 1121 388 1133 391
rect 339 360 1133 388
rect 339 357 351 360
rect 293 351 351 357
rect 1121 357 1133 360
rect 1167 357 1179 391
rect 1121 351 1179 357
<< labels >>
rlabel locali s 1327 215 1389 265 6 A0
port 1 nsew signal input
rlabel locali s 1307 199 1389 215 6 A0
port 1 nsew signal input
rlabel locali s 1307 75 1369 199 6 A0
port 1 nsew signal input
rlabel locali s 949 143 1023 279 6 A1
port 2 nsew signal input
rlabel locali s 204 79 247 153 6 A2
port 3 nsew signal input
rlabel locali s 167 153 247 219 6 A2
port 3 nsew signal input
rlabel locali s 482 203 523 264 6 A3
port 4 nsew signal input
rlabel locali s 448 143 523 203 6 A3
port 4 nsew signal input
rlabel locali s 29 195 65 349 6 S0
port 5 nsew signal input
rlabel locali s 244 257 278 289 6 S0
port 5 nsew signal input
rlabel locali s 201 289 278 323 6 S0
port 5 nsew signal input
rlabel locali s 1225 249 1293 329 6 S0
port 5 nsew signal input
rlabel metal1 s 1213 320 1271 329 6 S0
port 5 nsew signal input
rlabel metal1 s 1213 283 1271 292 6 S0
port 5 nsew signal input
rlabel metal1 s 201 320 259 329 6 S0
port 5 nsew signal input
rlabel metal1 s 201 283 259 292 6 S0
port 5 nsew signal input
rlabel metal1 s 17 320 75 329 6 S0
port 5 nsew signal input
rlabel metal1 s 17 292 1271 320 6 S0
port 5 nsew signal input
rlabel metal1 s 17 283 75 292 6 S0
port 5 nsew signal input
rlabel locali s 557 143 615 264 6 S1
port 6 nsew signal input
rlabel locali s 1519 145 1553 299 6 X
port 7 nsew signal output
rlabel locali s 1491 299 1553 367 6 X
port 7 nsew signal output
rlabel locali s 1487 53 1553 145 6 X
port 7 nsew signal output
rlabel locali s 1471 367 1553 491 6 X
port 7 nsew signal output
rlabel locali s 1587 17 1638 177 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 1403 17 1453 163 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 959 17 1025 109 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 490 17 556 109 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 103 17 169 93 6 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 0 -17 1656 17 8 VGND
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1656 48 8 VGND
port 8 nsew ground bidirectional abutment
rlabel locali s 1587 299 1637 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 1403 367 1437 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 951 401 1020 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 519 411 565 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 103 451 169 527 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 0 527 1656 561 6 VPWR
port 9 nsew power bidirectional abutment
rlabel metal1 s 0 496 1656 592 6 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1656 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1764024
string GDS_START 1749786
<< end >>
