magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 131 409 181 493
rect 66 288 181 409
rect 66 185 139 288
rect 66 132 186 185
rect 136 70 186 132
rect 451 199 588 265
rect 1476 289 1602 333
rect 1476 199 1520 289
rect 1660 215 1752 265
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 21 443 87 527
rect 225 443 292 527
rect 329 447 668 481
rect 721 447 802 481
rect 836 447 902 527
rect 989 455 1648 489
rect 1730 455 1807 527
rect 329 409 373 447
rect 768 413 802 447
rect 989 413 1023 455
rect 225 375 373 409
rect 453 379 734 413
rect 768 379 1023 413
rect 225 265 259 375
rect 306 307 656 341
rect 219 199 259 265
rect 225 173 259 199
rect 225 139 349 173
rect 21 17 87 93
rect 221 17 271 105
rect 305 85 349 139
rect 383 119 417 307
rect 622 265 656 307
rect 700 339 734 379
rect 700 305 806 339
rect 749 275 806 305
rect 622 199 687 265
rect 473 131 715 165
rect 557 85 638 91
rect 305 51 638 85
rect 672 85 715 131
rect 749 119 783 275
rect 840 241 874 379
rect 920 289 1023 343
rect 817 207 874 241
rect 817 85 851 207
rect 672 51 851 85
rect 885 17 919 173
rect 965 83 1023 289
rect 1058 119 1092 421
rect 1126 178 1160 455
rect 1851 421 1910 493
rect 1208 323 1291 409
rect 1408 387 1910 421
rect 1208 289 1374 323
rect 1211 199 1296 254
rect 1126 165 1180 178
rect 1126 144 1219 165
rect 1136 131 1219 144
rect 1058 97 1102 119
rect 1058 53 1141 97
rect 1185 64 1219 131
rect 1253 126 1296 199
rect 1340 85 1374 289
rect 1408 119 1442 387
rect 1803 375 1910 387
rect 1646 299 1820 341
rect 1786 265 1820 299
rect 1554 189 1618 255
rect 1786 199 1842 265
rect 1554 146 1595 189
rect 1786 181 1820 199
rect 1662 150 1820 181
rect 1654 147 1820 150
rect 1476 85 1579 93
rect 1340 51 1579 85
rect 1654 59 1712 147
rect 1876 117 1910 375
rect 1756 17 1790 113
rect 1850 51 1910 117
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< obsm1 >>
rect 760 320 818 329
rect 1250 320 1308 329
rect 760 292 1308 320
rect 760 283 818 292
rect 1250 283 1308 292
rect 954 184 1012 193
rect 1250 184 1308 193
rect 1546 184 1604 193
rect 954 156 1604 184
rect 954 147 1012 156
rect 1250 147 1308 156
rect 1546 147 1604 156
rect 1056 116 1114 125
rect 1648 116 1706 125
rect 1056 88 1706 116
rect 1056 79 1114 88
rect 1648 79 1706 88
<< labels >>
rlabel locali s 1660 215 1752 265 6 A
port 1 nsew signal input
rlabel locali s 1476 289 1602 333 6 B
port 2 nsew signal input
rlabel locali s 1476 199 1520 289 6 B
port 2 nsew signal input
rlabel locali s 451 199 588 265 6 C
port 3 nsew signal input
rlabel locali s 136 70 186 132 6 X
port 4 nsew signal output
rlabel locali s 131 409 181 493 6 X
port 4 nsew signal output
rlabel locali s 66 288 181 409 6 X
port 4 nsew signal output
rlabel locali s 66 185 139 288 6 X
port 4 nsew signal output
rlabel locali s 66 132 186 185 6 X
port 4 nsew signal output
rlabel metal1 s 0 -48 1932 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 1932 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1932 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 805980
string GDS_START 793160
<< end >>
