magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 368 561
rect 18 456 234 490
rect 18 299 85 456
rect 119 265 166 401
rect 200 333 234 456
rect 287 367 350 527
rect 200 299 263 333
rect 18 199 85 265
rect 119 199 195 265
rect 229 165 263 299
rect 18 131 263 165
rect 297 131 351 333
rect 18 77 69 131
rect 103 17 169 97
rect 203 77 237 131
rect 271 17 337 97
rect 0 -17 368 17
<< metal1 >>
rect 0 496 368 592
rect 0 -48 368 48
<< labels >>
rlabel locali s 297 131 351 333 6 A
port 1 nsew signal input
rlabel locali s 119 265 166 401 6 B
port 2 nsew signal input
rlabel locali s 119 199 195 265 6 B
port 2 nsew signal input
rlabel locali s 18 199 85 265 6 C
port 3 nsew signal input
rlabel locali s 229 165 263 299 6 Y
port 4 nsew signal output
rlabel locali s 203 77 237 131 6 Y
port 4 nsew signal output
rlabel locali s 200 333 234 456 6 Y
port 4 nsew signal output
rlabel locali s 200 299 263 333 6 Y
port 4 nsew signal output
rlabel locali s 18 456 234 490 6 Y
port 4 nsew signal output
rlabel locali s 18 299 85 456 6 Y
port 4 nsew signal output
rlabel locali s 18 131 263 165 6 Y
port 4 nsew signal output
rlabel locali s 18 77 69 131 6 Y
port 4 nsew signal output
rlabel locali s 271 17 337 97 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 103 17 169 97 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 368 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 368 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 287 367 350 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 368 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 368 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 368 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1972612
string GDS_START 1968432
<< end >>
