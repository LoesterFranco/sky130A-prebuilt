magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 2062 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 89 47 119 131
rect 183 47 213 131
rect 408 47 438 131
rect 504 47 534 119
rect 612 47 642 119
rect 775 47 805 131
rect 847 47 877 131
rect 999 47 1029 175
rect 1098 47 1128 119
rect 1207 47 1237 119
rect 1323 47 1353 131
rect 1512 47 1542 131
rect 1618 47 1648 131
rect 1806 47 1836 177
rect 1910 47 1940 177
<< pmoshvt >>
rect 81 363 117 491
rect 175 363 211 491
rect 400 413 436 497
rect 504 413 540 497
rect 613 413 649 497
rect 753 413 789 497
rect 860 413 896 497
rect 1077 329 1113 497
rect 1186 413 1222 497
rect 1294 413 1330 497
rect 1376 413 1412 497
rect 1514 413 1550 497
rect 1610 413 1646 497
rect 1808 297 1844 497
rect 1902 297 1938 497
<< ndiff >>
rect 27 119 89 131
rect 27 85 35 119
rect 69 85 89 119
rect 27 47 89 85
rect 119 93 183 131
rect 119 59 129 93
rect 163 59 183 93
rect 119 47 183 59
rect 213 119 265 131
rect 213 85 223 119
rect 257 85 265 119
rect 213 47 265 85
rect 319 89 408 131
rect 319 55 331 89
rect 365 55 408 89
rect 319 47 408 55
rect 438 119 488 131
rect 939 131 999 175
rect 657 119 775 131
rect 438 95 504 119
rect 438 61 449 95
rect 483 61 504 95
rect 438 47 504 61
rect 534 95 612 119
rect 534 61 555 95
rect 589 61 612 95
rect 534 47 612 61
rect 642 47 775 119
rect 805 47 847 131
rect 877 93 999 131
rect 877 59 921 93
rect 955 59 999 93
rect 877 47 999 59
rect 1029 119 1083 175
rect 1754 163 1806 177
rect 1273 119 1323 131
rect 1029 89 1098 119
rect 1029 55 1043 89
rect 1077 55 1098 89
rect 1029 47 1098 55
rect 1128 93 1207 119
rect 1128 59 1163 93
rect 1197 59 1207 93
rect 1128 47 1207 59
rect 1237 47 1323 119
rect 1353 89 1512 131
rect 1353 55 1365 89
rect 1399 55 1512 89
rect 1353 47 1512 55
rect 1542 47 1618 131
rect 1648 109 1700 131
rect 1648 75 1658 109
rect 1692 75 1700 109
rect 1648 47 1700 75
rect 1754 129 1762 163
rect 1796 129 1806 163
rect 1754 95 1806 129
rect 1754 61 1762 95
rect 1796 61 1806 95
rect 1754 47 1806 61
rect 1836 163 1910 177
rect 1836 129 1856 163
rect 1890 129 1910 163
rect 1836 95 1910 129
rect 1836 61 1856 95
rect 1890 61 1910 95
rect 1836 47 1910 61
rect 1940 95 1992 177
rect 1940 61 1950 95
rect 1984 61 1992 95
rect 1940 47 1992 61
<< pdiff >>
rect 27 477 81 491
rect 27 443 35 477
rect 69 443 81 477
rect 27 409 81 443
rect 27 375 35 409
rect 69 375 81 409
rect 27 363 81 375
rect 117 461 175 491
rect 117 427 129 461
rect 163 427 175 461
rect 117 363 175 427
rect 211 477 265 491
rect 211 443 223 477
rect 257 443 265 477
rect 211 409 265 443
rect 346 485 400 497
rect 346 451 354 485
rect 388 451 400 485
rect 346 413 400 451
rect 436 477 504 497
rect 436 443 450 477
rect 484 443 504 477
rect 436 413 504 443
rect 540 483 613 497
rect 540 449 553 483
rect 587 449 613 483
rect 540 413 613 449
rect 649 459 753 497
rect 649 425 707 459
rect 741 425 753 459
rect 649 413 753 425
rect 789 475 860 497
rect 789 441 814 475
rect 848 441 860 475
rect 789 413 860 441
rect 896 459 950 497
rect 896 425 908 459
rect 942 425 950 459
rect 896 413 950 425
rect 1013 485 1077 497
rect 1013 451 1031 485
rect 1065 451 1077 485
rect 211 375 223 409
rect 257 375 265 409
rect 211 363 265 375
rect 1013 329 1077 451
rect 1113 477 1186 497
rect 1113 443 1129 477
rect 1163 443 1186 477
rect 1113 413 1186 443
rect 1222 484 1294 497
rect 1222 450 1236 484
rect 1270 450 1294 484
rect 1222 413 1294 450
rect 1330 413 1376 497
rect 1412 485 1514 497
rect 1412 451 1468 485
rect 1502 451 1514 485
rect 1412 413 1514 451
rect 1550 459 1610 497
rect 1550 425 1562 459
rect 1596 425 1610 459
rect 1550 413 1610 425
rect 1646 485 1700 497
rect 1646 451 1658 485
rect 1692 451 1700 485
rect 1646 413 1700 451
rect 1754 485 1808 497
rect 1754 451 1762 485
rect 1796 451 1808 485
rect 1754 417 1808 451
rect 1113 329 1169 413
rect 1754 383 1762 417
rect 1796 383 1808 417
rect 1754 297 1808 383
rect 1844 477 1902 497
rect 1844 443 1856 477
rect 1890 443 1902 477
rect 1844 409 1902 443
rect 1844 375 1856 409
rect 1890 375 1902 409
rect 1844 341 1902 375
rect 1844 307 1856 341
rect 1890 307 1902 341
rect 1844 297 1902 307
rect 1938 477 1992 497
rect 1938 443 1950 477
rect 1984 443 1992 477
rect 1938 409 1992 443
rect 1938 375 1950 409
rect 1984 375 1992 409
rect 1938 297 1992 375
<< ndiffc >>
rect 35 85 69 119
rect 129 59 163 93
rect 223 85 257 119
rect 331 55 365 89
rect 449 61 483 95
rect 555 61 589 95
rect 921 59 955 93
rect 1043 55 1077 89
rect 1163 59 1197 93
rect 1365 55 1399 89
rect 1658 75 1692 109
rect 1762 129 1796 163
rect 1762 61 1796 95
rect 1856 129 1890 163
rect 1856 61 1890 95
rect 1950 61 1984 95
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 129 427 163 461
rect 223 443 257 477
rect 354 451 388 485
rect 450 443 484 477
rect 553 449 587 483
rect 707 425 741 459
rect 814 441 848 475
rect 908 425 942 459
rect 1031 451 1065 485
rect 223 375 257 409
rect 1129 443 1163 477
rect 1236 450 1270 484
rect 1468 451 1502 485
rect 1562 425 1596 459
rect 1658 451 1692 485
rect 1762 451 1796 485
rect 1762 383 1796 417
rect 1856 443 1890 477
rect 1856 375 1890 409
rect 1856 307 1890 341
rect 1950 443 1984 477
rect 1950 375 1984 409
<< poly >>
rect 81 491 117 517
rect 175 491 211 517
rect 400 497 436 523
rect 504 497 540 523
rect 613 497 649 523
rect 753 497 789 523
rect 860 497 896 523
rect 1077 497 1113 523
rect 1186 497 1222 523
rect 1294 497 1330 523
rect 1376 497 1412 523
rect 1514 497 1550 523
rect 1610 497 1646 523
rect 1808 497 1844 523
rect 1902 497 1938 523
rect 400 398 436 413
rect 504 398 540 413
rect 613 398 649 413
rect 753 398 789 413
rect 860 398 896 413
rect 81 348 117 363
rect 175 348 211 363
rect 46 318 119 348
rect 46 265 76 318
rect 173 274 213 348
rect 398 326 438 398
rect 502 375 542 398
rect 22 249 76 265
rect 22 215 32 249
rect 66 215 76 249
rect 128 264 213 274
rect 128 230 144 264
rect 178 230 213 264
rect 337 310 438 326
rect 486 365 562 375
rect 486 331 502 365
rect 536 331 562 365
rect 486 321 562 331
rect 337 276 347 310
rect 381 276 438 310
rect 611 279 651 398
rect 751 355 791 398
rect 751 339 816 355
rect 751 305 761 339
rect 795 305 816 339
rect 751 289 816 305
rect 337 260 438 276
rect 128 220 213 230
rect 22 199 76 215
rect 46 176 76 199
rect 46 146 119 176
rect 89 131 119 146
rect 183 131 213 220
rect 408 131 438 260
rect 493 249 651 279
rect 493 219 534 249
rect 480 203 534 219
rect 480 169 490 203
rect 524 169 534 203
rect 480 153 534 169
rect 576 197 642 207
rect 576 163 592 197
rect 626 163 642 197
rect 576 153 642 163
rect 504 119 534 153
rect 612 119 642 153
rect 775 131 805 289
rect 858 219 898 398
rect 1186 398 1222 413
rect 1294 398 1330 413
rect 1376 398 1412 413
rect 1514 398 1550 413
rect 1610 398 1646 413
rect 1077 314 1113 329
rect 989 284 1115 314
rect 989 267 1029 284
rect 953 251 1029 267
rect 847 203 911 219
rect 847 169 857 203
rect 891 169 911 203
rect 953 217 963 251
rect 997 217 1029 251
rect 1184 279 1224 398
rect 1292 381 1332 398
rect 1266 365 1332 381
rect 1266 331 1282 365
rect 1316 331 1332 365
rect 1266 321 1332 331
rect 1184 249 1261 279
rect 953 201 1029 217
rect 1207 239 1261 249
rect 999 175 1029 201
rect 1098 191 1165 207
rect 847 153 911 169
rect 847 131 877 153
rect 1098 157 1121 191
rect 1155 157 1165 191
rect 1098 141 1165 157
rect 1207 205 1217 239
rect 1251 205 1261 239
rect 1207 189 1261 205
rect 1374 229 1414 398
rect 1512 257 1552 398
rect 1608 365 1648 398
rect 1594 349 1648 365
rect 1594 315 1604 349
rect 1638 315 1648 349
rect 1594 299 1648 315
rect 1512 241 1568 257
rect 1374 213 1445 229
rect 1374 193 1391 213
rect 1098 119 1128 141
rect 1207 119 1237 189
rect 1323 179 1391 193
rect 1425 179 1445 213
rect 1323 163 1445 179
rect 1512 207 1522 241
rect 1556 207 1568 241
rect 1512 191 1568 207
rect 1323 131 1353 163
rect 1512 131 1542 191
rect 1618 131 1648 299
rect 1808 282 1844 297
rect 1902 282 1938 297
rect 1806 265 1846 282
rect 1900 265 1940 282
rect 1806 249 1940 265
rect 1806 215 1817 249
rect 1851 215 1940 249
rect 1806 199 1940 215
rect 1806 177 1836 199
rect 1910 177 1940 199
rect 89 21 119 47
rect 183 21 213 47
rect 408 21 438 47
rect 504 21 534 47
rect 612 21 642 47
rect 775 21 805 47
rect 847 21 877 47
rect 999 21 1029 47
rect 1098 21 1128 47
rect 1207 21 1237 47
rect 1323 21 1353 47
rect 1512 21 1542 47
rect 1618 21 1648 47
rect 1806 21 1836 47
rect 1910 21 1940 47
<< polycont >>
rect 32 215 66 249
rect 144 230 178 264
rect 502 331 536 365
rect 347 276 381 310
rect 761 305 795 339
rect 490 169 524 203
rect 592 163 626 197
rect 857 169 891 203
rect 963 217 997 251
rect 1282 331 1316 365
rect 1121 157 1155 191
rect 1217 205 1251 239
rect 1604 315 1638 349
rect 1391 179 1425 213
rect 1522 207 1556 241
rect 1817 215 1851 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 18 477 69 493
rect 18 443 35 477
rect 18 409 69 443
rect 103 461 179 527
rect 103 427 129 461
rect 163 427 179 461
rect 223 477 257 493
rect 18 375 35 409
rect 223 409 257 443
rect 354 485 388 527
rect 354 435 388 451
rect 434 477 484 493
rect 434 443 450 477
rect 69 375 178 393
rect 18 359 178 375
rect 18 249 88 325
rect 18 215 32 249
rect 66 215 88 249
rect 18 195 88 215
rect 132 264 178 359
rect 132 255 144 264
rect 166 221 178 230
rect 132 161 178 221
rect 18 127 178 161
rect 434 427 484 443
rect 537 483 673 493
rect 537 449 553 483
rect 587 449 673 483
rect 798 475 864 527
rect 1001 485 1085 527
rect 537 427 673 449
rect 434 401 468 427
rect 18 119 69 127
rect 18 85 35 119
rect 223 119 257 357
rect 291 333 354 401
rect 415 367 468 401
rect 502 391 605 393
rect 291 310 381 333
rect 291 276 347 310
rect 291 123 381 276
rect 18 69 69 85
rect 103 59 129 93
rect 163 59 179 93
rect 223 69 257 85
rect 103 17 179 59
rect 315 55 331 89
rect 365 55 381 89
rect 415 61 449 367
rect 502 365 545 391
rect 536 357 545 365
rect 579 357 605 391
rect 536 331 605 357
rect 502 315 605 331
rect 485 255 537 277
rect 485 221 496 255
rect 530 221 537 255
rect 485 203 537 221
rect 485 169 490 203
rect 524 169 537 203
rect 485 153 537 169
rect 571 197 605 315
rect 639 271 673 427
rect 707 459 741 475
rect 798 441 814 475
rect 848 441 864 475
rect 908 459 942 475
rect 707 407 741 425
rect 1001 451 1031 485
rect 1065 451 1085 485
rect 1001 435 1085 451
rect 1129 477 1163 493
rect 908 407 942 425
rect 707 373 942 407
rect 1129 401 1163 443
rect 1210 484 1401 493
rect 1210 450 1236 484
rect 1270 450 1401 484
rect 1210 425 1401 450
rect 1468 485 1518 527
rect 1502 451 1518 485
rect 1632 485 1708 527
rect 1468 435 1518 451
rect 1562 459 1596 475
rect 1031 367 1163 401
rect 1031 339 1065 367
rect 745 305 761 339
rect 795 305 1065 339
rect 1229 365 1294 391
rect 1229 333 1282 365
rect 1328 357 1332 391
rect 639 251 997 271
rect 639 237 963 251
rect 571 163 592 197
rect 626 163 642 197
rect 571 153 642 163
rect 686 95 720 237
rect 761 187 857 203
rect 761 153 821 187
rect 855 169 857 187
rect 891 187 929 203
rect 963 201 997 217
rect 891 169 893 187
rect 855 153 893 169
rect 927 153 929 187
rect 1031 167 1065 305
rect 483 61 499 95
rect 539 61 555 95
rect 589 61 720 95
rect 905 93 971 109
rect 315 17 381 55
rect 905 59 921 93
rect 955 59 971 93
rect 905 17 971 59
rect 1013 89 1065 167
rect 1121 331 1282 333
rect 1316 331 1332 357
rect 1367 349 1401 425
rect 1632 451 1658 485
rect 1692 451 1708 485
rect 1762 485 1796 527
rect 1562 417 1596 425
rect 1762 417 1796 451
rect 1562 383 1722 417
rect 1121 299 1263 331
rect 1367 315 1604 349
rect 1638 315 1654 349
rect 1121 191 1155 299
rect 1367 297 1411 315
rect 1121 141 1155 157
rect 1189 255 1263 265
rect 1189 221 1204 255
rect 1238 239 1263 255
rect 1189 205 1217 221
rect 1251 205 1263 239
rect 1189 141 1263 205
rect 1297 263 1411 297
rect 1297 107 1331 263
rect 1501 241 1581 281
rect 1688 259 1722 383
rect 1762 315 1796 383
rect 1848 477 1906 493
rect 1848 443 1856 477
rect 1890 443 1906 477
rect 1848 409 1906 443
rect 1848 375 1856 409
rect 1890 375 1906 409
rect 1848 341 1906 375
rect 1950 477 1984 527
rect 1950 409 1984 443
rect 1950 359 1984 375
rect 1848 307 1856 341
rect 1890 325 1906 341
rect 1890 307 2002 325
rect 1848 291 2002 307
rect 1391 213 1445 229
rect 1425 179 1445 213
rect 1391 173 1445 179
rect 1501 207 1522 241
rect 1556 207 1581 241
rect 1501 187 1581 207
rect 1391 139 1467 173
rect 1147 93 1331 107
rect 1013 55 1043 89
rect 1077 55 1093 89
rect 1147 59 1163 93
rect 1197 59 1331 93
rect 1147 51 1331 59
rect 1365 89 1399 105
rect 1433 93 1467 139
rect 1501 153 1527 187
rect 1561 153 1581 187
rect 1501 127 1581 153
rect 1658 257 1722 259
rect 1658 249 1867 257
rect 1658 215 1817 249
rect 1851 215 1867 249
rect 1658 109 1727 215
rect 1925 181 2002 291
rect 1433 75 1658 93
rect 1692 75 1727 109
rect 1433 59 1727 75
rect 1762 163 1796 179
rect 1762 95 1796 129
rect 1365 17 1399 55
rect 1762 17 1796 61
rect 1830 163 2002 181
rect 1830 129 1856 163
rect 1890 147 2002 163
rect 1890 129 1906 147
rect 1830 95 1906 129
rect 1830 61 1856 95
rect 1890 61 1906 95
rect 1830 51 1906 61
rect 1950 95 1984 111
rect 1950 17 1984 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 132 230 144 255
rect 144 230 166 255
rect 132 221 166 230
rect 223 375 257 391
rect 223 357 257 375
rect 545 357 579 391
rect 496 221 530 255
rect 1294 365 1328 391
rect 1294 357 1316 365
rect 1316 357 1328 365
rect 821 153 855 187
rect 893 153 927 187
rect 1204 239 1238 255
rect 1204 221 1217 239
rect 1217 221 1238 239
rect 1527 153 1561 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
<< metal1 >>
rect 0 561 2024 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 0 496 2024 527
rect 201 391 269 397
rect 201 357 223 391
rect 257 388 269 391
rect 533 391 591 397
rect 533 388 545 391
rect 257 360 545 388
rect 257 357 269 360
rect 201 351 269 357
rect 533 357 545 360
rect 579 388 591 391
rect 1282 391 1340 397
rect 1282 388 1294 391
rect 579 360 1294 388
rect 579 357 591 360
rect 533 351 591 357
rect 1282 357 1294 360
rect 1328 357 1340 391
rect 1282 351 1340 357
rect 120 255 178 261
rect 120 221 132 255
rect 166 252 178 255
rect 484 255 542 261
rect 484 252 496 255
rect 166 224 496 252
rect 166 221 178 224
rect 120 215 178 221
rect 484 221 496 224
rect 530 252 542 255
rect 1192 255 1250 261
rect 1192 252 1204 255
rect 530 224 1204 252
rect 530 221 542 224
rect 484 215 542 221
rect 1192 221 1204 224
rect 1238 221 1250 255
rect 1192 215 1250 221
rect 799 187 949 193
rect 799 153 821 187
rect 855 153 893 187
rect 927 184 949 187
rect 1515 187 1573 193
rect 1515 184 1527 187
rect 927 156 1527 184
rect 927 153 949 156
rect 799 147 949 153
rect 1515 153 1527 156
rect 1561 153 1573 187
rect 1515 147 1573 153
rect 0 17 2024 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
rect 0 -48 2024 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dfrtp_4
flabel metal1 s 1527 153 1561 187 0 FreeSans 400 0 0 0 RESET_B
port 3 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel corelocali s 1958 221 1992 255 0 FreeSans 400 0 0 0 Q
port 8 nsew
flabel corelocali s 1958 153 1992 187 0 FreeSans 400 0 0 0 Q
port 8 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 400 0 0 0 CLK
port 1 nsew
flabel corelocali s 30 289 64 323 0 FreeSans 400 0 0 0 CLK
port 1 nsew
flabel corelocali s 305 289 339 323 0 FreeSans 400 0 0 0 D
port 2 nsew
flabel corelocali s 1958 289 1992 323 0 FreeSans 400 0 0 0 Q
port 8 nsew
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 2024 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1860434
string GDS_START 1845400
<< end >>
