magic
tech sky130A
magscale 1 2
timestamp 1604502705
<< nwell >>
rect -38 332 1670 704
<< pwell >>
rect 0 0 1632 49
<< scnmos >>
rect 84 136 114 246
rect 202 98 232 246
rect 435 82 465 230
rect 667 74 697 202
rect 745 74 775 202
rect 840 74 870 158
rect 925 74 955 158
rect 1123 74 1153 222
rect 1201 74 1231 222
rect 1416 74 1446 222
rect 1502 74 1532 222
<< pmoshvt >>
rect 120 394 150 562
rect 230 394 260 562
rect 432 392 462 560
rect 556 392 586 592
rect 640 392 670 592
rect 748 504 778 588
rect 916 504 946 588
rect 1114 368 1144 592
rect 1206 368 1236 592
rect 1414 368 1444 592
rect 1504 368 1534 592
<< ndiff >>
rect 27 208 84 246
rect 27 174 39 208
rect 73 174 84 208
rect 27 136 84 174
rect 114 136 202 246
rect 129 98 202 136
rect 232 225 293 246
rect 232 191 243 225
rect 277 191 293 225
rect 232 98 293 191
rect 373 218 435 230
rect 373 184 387 218
rect 421 184 435 218
rect 129 82 187 98
rect 129 48 141 82
rect 175 48 187 82
rect 373 82 435 184
rect 465 202 515 230
rect 465 82 667 202
rect 129 36 187 48
rect 480 48 492 82
rect 526 48 606 82
rect 640 74 667 82
rect 697 74 745 202
rect 775 158 825 202
rect 1066 210 1123 222
rect 1066 176 1078 210
rect 1112 176 1123 210
rect 775 133 840 158
rect 775 99 795 133
rect 829 99 840 133
rect 775 74 840 99
rect 870 74 925 158
rect 955 120 1012 158
rect 955 86 966 120
rect 1000 86 1012 120
rect 955 74 1012 86
rect 1066 120 1123 176
rect 1066 86 1078 120
rect 1112 86 1123 120
rect 1066 74 1123 86
rect 1153 74 1201 222
rect 1231 188 1416 222
rect 1231 154 1242 188
rect 1276 154 1357 188
rect 1391 154 1416 188
rect 1231 120 1416 154
rect 1231 86 1242 120
rect 1276 86 1357 120
rect 1391 86 1416 120
rect 1231 74 1416 86
rect 1446 210 1502 222
rect 1446 176 1457 210
rect 1491 176 1502 210
rect 1446 120 1502 176
rect 1446 86 1457 120
rect 1491 86 1502 120
rect 1446 74 1502 86
rect 1532 210 1603 222
rect 1532 176 1557 210
rect 1591 176 1603 210
rect 1532 120 1603 176
rect 1532 86 1557 120
rect 1591 86 1603 120
rect 1532 74 1603 86
rect 640 48 652 74
rect 480 36 652 48
<< pdiff >>
rect 480 622 538 634
rect 480 588 492 622
rect 526 592 538 622
rect 526 588 556 592
rect 61 550 120 562
rect 61 516 73 550
rect 107 516 120 550
rect 61 440 120 516
rect 61 406 73 440
rect 107 406 120 440
rect 61 394 120 406
rect 150 550 230 562
rect 150 516 173 550
rect 207 516 230 550
rect 150 440 230 516
rect 150 406 173 440
rect 207 406 230 440
rect 150 394 230 406
rect 260 550 319 562
rect 480 560 556 588
rect 260 516 273 550
rect 307 516 319 550
rect 260 440 319 516
rect 260 406 273 440
rect 307 406 319 440
rect 260 394 319 406
rect 373 446 432 560
rect 373 412 385 446
rect 419 412 432 446
rect 373 392 432 412
rect 462 392 556 560
rect 586 392 640 592
rect 670 588 723 592
rect 1061 588 1114 592
rect 670 504 748 588
rect 778 504 916 588
rect 946 576 1114 588
rect 946 542 959 576
rect 993 542 1059 576
rect 1093 542 1114 576
rect 946 504 1114 542
rect 670 470 730 504
rect 670 436 683 470
rect 717 436 730 470
rect 670 392 730 436
rect 1061 368 1114 504
rect 1144 580 1206 592
rect 1144 546 1159 580
rect 1193 546 1206 580
rect 1144 497 1206 546
rect 1144 463 1159 497
rect 1193 463 1206 497
rect 1144 414 1206 463
rect 1144 380 1159 414
rect 1193 380 1206 414
rect 1144 368 1206 380
rect 1236 580 1414 592
rect 1236 546 1280 580
rect 1314 546 1414 580
rect 1236 462 1414 546
rect 1236 428 1280 462
rect 1314 428 1414 462
rect 1236 368 1414 428
rect 1444 580 1504 592
rect 1444 546 1457 580
rect 1491 546 1504 580
rect 1444 497 1504 546
rect 1444 463 1457 497
rect 1491 463 1504 497
rect 1444 414 1504 463
rect 1444 380 1457 414
rect 1491 380 1504 414
rect 1444 368 1504 380
rect 1534 580 1605 592
rect 1534 546 1558 580
rect 1592 546 1605 580
rect 1534 497 1605 546
rect 1534 463 1558 497
rect 1592 463 1605 497
rect 1534 414 1605 463
rect 1534 380 1558 414
rect 1592 380 1605 414
rect 1534 368 1605 380
<< ndiffc >>
rect 39 174 73 208
rect 243 191 277 225
rect 387 184 421 218
rect 141 48 175 82
rect 492 48 526 82
rect 606 48 640 82
rect 1078 176 1112 210
rect 795 99 829 133
rect 966 86 1000 120
rect 1078 86 1112 120
rect 1242 154 1276 188
rect 1357 154 1391 188
rect 1242 86 1276 120
rect 1357 86 1391 120
rect 1457 176 1491 210
rect 1457 86 1491 120
rect 1557 176 1591 210
rect 1557 86 1591 120
<< pdiffc >>
rect 492 588 526 622
rect 73 516 107 550
rect 73 406 107 440
rect 173 516 207 550
rect 173 406 207 440
rect 273 516 307 550
rect 273 406 307 440
rect 385 412 419 446
rect 959 542 993 576
rect 1059 542 1093 576
rect 683 436 717 470
rect 1159 546 1193 580
rect 1159 463 1193 497
rect 1159 380 1193 414
rect 1280 546 1314 580
rect 1280 428 1314 462
rect 1457 546 1491 580
rect 1457 463 1491 497
rect 1457 380 1491 414
rect 1558 546 1592 580
rect 1558 463 1592 497
rect 1558 380 1592 414
<< poly >>
rect 556 592 586 618
rect 640 592 670 618
rect 120 562 150 588
rect 230 562 260 588
rect 432 560 462 586
rect 120 379 150 394
rect 230 379 260 394
rect 748 588 778 614
rect 916 588 946 614
rect 1114 592 1144 618
rect 1206 592 1236 618
rect 1414 592 1444 618
rect 1504 592 1534 618
rect 748 489 778 504
rect 916 489 946 504
rect 745 472 781 489
rect 913 472 949 489
rect 745 456 865 472
rect 745 422 815 456
rect 849 422 865 456
rect 745 406 865 422
rect 913 456 979 472
rect 913 422 929 456
rect 963 422 979 456
rect 913 406 979 422
rect 117 356 153 379
rect 227 356 263 379
rect 432 377 462 392
rect 556 377 586 392
rect 640 377 670 392
rect 84 340 153 356
rect 84 306 103 340
rect 137 306 153 340
rect 84 290 153 306
rect 201 340 267 356
rect 201 306 217 340
rect 251 306 267 340
rect 201 290 267 306
rect 315 318 381 334
rect 84 246 114 290
rect 202 246 232 290
rect 315 284 331 318
rect 365 298 381 318
rect 429 298 465 377
rect 553 318 589 377
rect 637 360 673 377
rect 365 284 465 298
rect 315 268 465 284
rect 84 110 114 136
rect 435 230 465 268
rect 523 302 589 318
rect 523 268 539 302
rect 573 268 589 302
rect 631 344 697 360
rect 631 310 647 344
rect 681 310 697 344
rect 631 294 697 310
rect 523 252 589 268
rect 202 72 232 98
rect 559 222 697 252
rect 667 202 697 222
rect 745 202 775 406
rect 925 336 961 406
rect 1114 353 1144 368
rect 1206 353 1236 368
rect 1414 353 1444 368
rect 1504 353 1534 368
rect 1111 336 1147 353
rect 817 288 883 304
rect 817 254 833 288
rect 867 254 883 288
rect 817 238 883 254
rect 435 56 465 82
rect 840 158 870 238
rect 925 158 955 336
rect 1009 320 1147 336
rect 1009 286 1025 320
rect 1059 300 1147 320
rect 1203 310 1239 353
rect 1303 314 1369 330
rect 1059 286 1153 300
rect 1009 270 1153 286
rect 1123 222 1153 270
rect 1195 294 1261 310
rect 1195 260 1211 294
rect 1245 260 1261 294
rect 1303 280 1319 314
rect 1353 294 1369 314
rect 1411 294 1447 353
rect 1501 294 1537 353
rect 1353 280 1537 294
rect 1303 264 1537 280
rect 1195 244 1261 260
rect 1201 222 1231 244
rect 1416 222 1446 264
rect 1502 222 1532 264
rect 667 48 697 74
rect 745 48 775 74
rect 840 48 870 74
rect 925 48 955 74
rect 1123 48 1153 74
rect 1201 48 1231 74
rect 1416 48 1446 74
rect 1502 48 1532 74
<< polycont >>
rect 815 422 849 456
rect 929 422 963 456
rect 103 306 137 340
rect 217 306 251 340
rect 331 284 365 318
rect 539 268 573 302
rect 647 310 681 344
rect 833 254 867 288
rect 1025 286 1059 320
rect 1211 260 1245 294
rect 1319 280 1353 314
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 19 550 123 566
rect 19 516 73 550
rect 107 516 123 550
rect 19 440 123 516
rect 19 406 73 440
rect 107 406 123 440
rect 19 390 123 406
rect 157 550 223 649
rect 476 622 542 649
rect 476 588 492 622
rect 526 588 542 622
rect 476 572 542 588
rect 943 576 1109 649
rect 157 516 173 550
rect 207 516 223 550
rect 157 440 223 516
rect 157 406 173 440
rect 207 406 223 440
rect 157 390 223 406
rect 257 550 335 566
rect 257 516 273 550
rect 307 538 335 550
rect 943 542 959 576
rect 993 542 1059 576
rect 1093 542 1109 576
rect 307 516 865 538
rect 943 526 1109 542
rect 1143 580 1209 596
rect 1143 546 1159 580
rect 1193 546 1209 580
rect 257 504 865 516
rect 257 440 335 504
rect 257 406 273 440
rect 307 406 335 440
rect 257 390 335 406
rect 19 250 53 390
rect 87 340 167 356
rect 87 306 103 340
rect 137 306 167 340
rect 87 290 167 306
rect 201 340 267 356
rect 201 306 217 340
rect 251 306 267 340
rect 201 290 267 306
rect 301 334 335 390
rect 369 446 449 470
rect 369 412 385 446
rect 419 412 449 446
rect 667 436 683 470
rect 717 436 765 470
rect 369 402 449 412
rect 369 368 697 402
rect 301 318 381 334
rect 301 284 331 318
rect 365 284 381 318
rect 301 268 381 284
rect 301 250 335 268
rect 19 208 89 250
rect 19 174 39 208
rect 73 174 89 208
rect 227 225 335 250
rect 415 234 449 368
rect 631 344 697 368
rect 227 191 243 225
rect 277 191 335 225
rect 227 184 335 191
rect 369 218 449 234
rect 369 184 387 218
rect 421 184 449 218
rect 523 302 589 318
rect 523 268 539 302
rect 573 268 589 302
rect 19 150 89 174
rect 523 150 589 268
rect 631 310 647 344
rect 681 310 697 344
rect 731 372 765 436
rect 799 456 865 504
rect 1143 497 1209 546
rect 1143 472 1159 497
rect 799 422 815 456
rect 849 422 865 456
rect 799 406 865 422
rect 913 463 1159 472
rect 1193 463 1209 497
rect 913 456 1209 463
rect 913 422 929 456
rect 963 422 1209 456
rect 913 414 1209 422
rect 913 406 1159 414
rect 1109 380 1159 406
rect 1193 380 1209 414
rect 1264 580 1330 649
rect 1264 546 1280 580
rect 1314 546 1330 580
rect 1264 462 1330 546
rect 1264 428 1280 462
rect 1314 428 1330 462
rect 1264 412 1330 428
rect 1369 580 1507 596
rect 1369 546 1457 580
rect 1491 546 1507 580
rect 1369 497 1507 546
rect 1369 463 1457 497
rect 1491 463 1507 497
rect 1369 414 1507 463
rect 1109 378 1209 380
rect 1369 380 1457 414
rect 1491 380 1507 414
rect 731 338 1075 372
rect 631 304 697 310
rect 994 320 1075 338
rect 631 288 883 304
rect 631 254 833 288
rect 867 254 883 288
rect 631 238 883 254
rect 994 286 1025 320
rect 1059 286 1075 320
rect 994 270 1075 286
rect 1109 344 1335 378
rect 1369 364 1507 380
rect 1541 580 1609 649
rect 1541 546 1558 580
rect 1592 546 1609 580
rect 1541 497 1609 546
rect 1541 463 1558 497
rect 1592 463 1609 497
rect 1541 414 1609 463
rect 1541 380 1558 414
rect 1592 380 1609 414
rect 1541 364 1609 380
rect 994 204 1028 270
rect 1109 226 1143 344
rect 1301 330 1335 344
rect 1301 314 1369 330
rect 1177 294 1261 310
rect 1177 260 1211 294
rect 1245 260 1261 294
rect 1301 280 1319 314
rect 1353 280 1369 314
rect 1473 294 1507 364
rect 1301 264 1369 280
rect 1177 236 1261 260
rect 19 116 589 150
rect 779 170 1028 204
rect 1062 210 1143 226
rect 1062 176 1078 210
rect 1112 176 1143 210
rect 1441 210 1507 294
rect 779 133 845 170
rect 779 99 795 133
rect 829 99 845 133
rect 125 48 141 82
rect 175 48 191 82
rect 125 17 191 48
rect 476 48 492 82
rect 526 48 606 82
rect 640 48 656 82
rect 779 70 845 99
rect 950 120 1016 136
rect 950 86 966 120
rect 1000 86 1016 120
rect 476 17 656 48
rect 950 17 1016 86
rect 1062 120 1143 176
rect 1062 86 1078 120
rect 1112 86 1143 120
rect 1062 70 1143 86
rect 1226 188 1407 202
rect 1226 154 1242 188
rect 1276 154 1357 188
rect 1391 154 1407 188
rect 1226 120 1407 154
rect 1226 86 1242 120
rect 1276 86 1357 120
rect 1391 86 1407 120
rect 1226 17 1407 86
rect 1441 176 1457 210
rect 1491 176 1507 210
rect 1441 120 1507 176
rect 1441 86 1457 120
rect 1491 86 1507 120
rect 1441 70 1507 86
rect 1541 210 1607 226
rect 1541 176 1557 210
rect 1591 176 1607 210
rect 1541 120 1607 176
rect 1541 86 1557 120
rect 1591 86 1607 120
rect 1541 17 1607 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dlrtn_2
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 1 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew
flabel corelocali s 1183 242 1217 276 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew
flabel corelocali s 1375 390 1409 424 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 1375 464 1409 498 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 1375 538 1409 572 0 FreeSans 340 0 0 0 Q
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 1632 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2818636
string GDS_START 2807072
<< end >>
