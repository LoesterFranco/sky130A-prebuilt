magic
tech sky130A
magscale 1 2
timestamp 1599588244
<< locali >>
rect 25 260 91 356
rect 202 364 288 414
rect 202 226 236 364
rect 544 236 647 310
rect 681 236 747 310
rect 202 70 268 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 23 482 89 540
rect 130 516 196 649
rect 313 516 447 649
rect 489 482 555 572
rect 23 448 442 482
rect 23 390 159 448
rect 125 226 159 390
rect 21 192 159 226
rect 270 260 336 326
rect 378 270 442 448
rect 476 364 555 482
rect 681 364 747 649
rect 302 236 336 260
rect 476 236 510 364
rect 21 91 71 192
rect 107 17 157 158
rect 302 202 510 236
rect 304 17 354 164
rect 396 70 446 202
rect 682 168 748 202
rect 482 134 748 168
rect 482 70 548 134
rect 582 17 648 100
rect 682 70 748 134
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel locali s 681 236 747 310 6 A1
port 1 nsew signal input
rlabel locali s 544 236 647 310 6 A2
port 2 nsew signal input
rlabel locali s 25 260 91 356 6 B1_N
port 3 nsew signal input
rlabel locali s 202 364 288 414 6 X
port 4 nsew signal output
rlabel locali s 202 226 236 364 6 X
port 4 nsew signal output
rlabel locali s 202 70 268 226 6 X
port 4 nsew signal output
rlabel metal1 s 0 -49 768 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 6 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 617 768 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1017820
string GDS_START 1011190
<< end >>
