magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 828 561
rect 18 299 69 527
rect 103 333 169 493
rect 203 367 237 527
rect 271 333 337 493
rect 371 367 405 527
rect 439 333 505 493
rect 539 367 573 527
rect 607 333 673 493
rect 707 367 757 527
rect 103 299 673 333
rect 22 215 346 265
rect 382 215 489 299
rect 523 215 811 265
rect 119 17 153 109
rect 287 17 321 109
rect 439 161 489 215
rect 439 127 673 161
rect 0 -17 828 17
<< obsli1 >>
rect 18 143 405 181
rect 18 51 85 143
rect 187 51 253 143
rect 355 93 405 143
rect 707 93 757 177
rect 355 51 757 93
<< metal1 >>
rect 0 496 828 592
rect 0 -48 828 48
<< labels >>
rlabel locali s 523 215 811 265 6 A
port 1 nsew signal input
rlabel locali s 22 215 346 265 6 B
port 2 nsew signal input
rlabel locali s 607 333 673 493 6 Y
port 3 nsew signal output
rlabel locali s 439 333 505 493 6 Y
port 3 nsew signal output
rlabel locali s 439 161 489 215 6 Y
port 3 nsew signal output
rlabel locali s 439 127 673 161 6 Y
port 3 nsew signal output
rlabel locali s 382 215 489 299 6 Y
port 3 nsew signal output
rlabel locali s 271 333 337 493 6 Y
port 3 nsew signal output
rlabel locali s 103 333 169 493 6 Y
port 3 nsew signal output
rlabel locali s 103 299 673 333 6 Y
port 3 nsew signal output
rlabel locali s 287 17 321 109 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 119 17 153 109 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 828 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 828 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 707 367 757 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 539 367 573 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 371 367 405 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 203 367 237 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 18 299 69 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 828 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 828 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1698444
string GDS_START 1690862
<< end >>
