magic
tech sky130A
magscale 1 2
timestamp 1601050047
<< nwell >>
rect -38 332 710 704
<< pwell >>
rect 0 0 672 49
<< scpmos >>
rect 84 368 114 592
rect 334 392 364 592
rect 424 392 454 592
rect 520 392 550 592
<< nmoslvt >>
rect 226 116 256 264
rect 336 136 366 264
rect 422 136 452 264
rect 517 136 547 264
<< ndiff >>
rect 173 194 226 264
rect 173 160 181 194
rect 215 160 226 194
rect 173 116 226 160
rect 256 172 336 264
rect 256 138 267 172
rect 301 138 336 172
rect 256 136 336 138
rect 366 246 422 264
rect 366 212 377 246
rect 411 212 422 246
rect 366 178 422 212
rect 366 144 377 178
rect 411 144 422 178
rect 366 136 422 144
rect 452 136 517 264
rect 547 235 600 264
rect 547 201 558 235
rect 592 201 600 235
rect 547 136 600 201
rect 256 116 313 136
<< pdiff >>
rect 29 580 84 592
rect 29 546 37 580
rect 71 546 84 580
rect 29 497 84 546
rect 29 463 37 497
rect 71 463 84 497
rect 29 414 84 463
rect 29 380 37 414
rect 71 380 84 414
rect 29 368 84 380
rect 114 580 169 592
rect 114 546 127 580
rect 161 546 169 580
rect 114 497 169 546
rect 114 463 127 497
rect 161 463 169 497
rect 114 414 169 463
rect 114 380 127 414
rect 161 380 169 414
rect 279 580 334 592
rect 279 546 287 580
rect 321 546 334 580
rect 279 510 334 546
rect 279 476 287 510
rect 321 476 334 510
rect 279 440 334 476
rect 279 406 287 440
rect 321 406 334 440
rect 279 392 334 406
rect 364 580 424 592
rect 364 546 377 580
rect 411 546 424 580
rect 364 510 424 546
rect 364 476 377 510
rect 411 476 424 510
rect 364 440 424 476
rect 364 406 377 440
rect 411 406 424 440
rect 364 392 424 406
rect 454 580 520 592
rect 454 546 470 580
rect 504 546 520 580
rect 454 508 520 546
rect 454 474 470 508
rect 504 474 520 508
rect 454 392 520 474
rect 550 580 605 592
rect 550 546 563 580
rect 597 546 605 580
rect 550 509 605 546
rect 550 475 563 509
rect 597 475 605 509
rect 550 438 605 475
rect 550 404 563 438
rect 597 404 605 438
rect 550 392 605 404
rect 114 368 169 380
<< ndiffc >>
rect 181 160 215 194
rect 267 138 301 172
rect 377 212 411 246
rect 377 144 411 178
rect 558 201 592 235
<< pdiffc >>
rect 37 546 71 580
rect 37 463 71 497
rect 37 380 71 414
rect 127 546 161 580
rect 127 463 161 497
rect 127 380 161 414
rect 287 546 321 580
rect 287 476 321 510
rect 287 406 321 440
rect 377 546 411 580
rect 377 476 411 510
rect 377 406 411 440
rect 470 546 504 580
rect 470 474 504 508
rect 563 546 597 580
rect 563 475 597 509
rect 563 404 597 438
<< poly >>
rect 84 592 114 618
rect 334 592 364 618
rect 424 592 454 618
rect 520 592 550 618
rect 334 377 364 392
rect 424 377 454 392
rect 520 377 550 392
rect 84 353 114 368
rect 331 356 367 377
rect 421 356 457 377
rect 81 330 117 353
rect 301 340 367 356
rect 81 314 151 330
rect 81 280 101 314
rect 135 309 151 314
rect 135 280 256 309
rect 301 306 317 340
rect 351 306 367 340
rect 301 290 367 306
rect 409 340 475 356
rect 409 306 425 340
rect 459 306 475 340
rect 409 290 475 306
rect 81 279 256 280
rect 81 264 151 279
rect 226 264 256 279
rect 336 264 366 290
rect 422 264 452 290
rect 517 279 553 377
rect 517 264 547 279
rect 226 90 256 116
rect 336 110 366 136
rect 422 110 452 136
rect 517 114 547 136
rect 517 98 595 114
rect 517 64 545 98
rect 579 64 595 98
rect 517 48 595 64
<< polycont >>
rect 101 280 135 314
rect 317 306 351 340
rect 425 306 459 340
rect 545 64 579 98
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 17 580 87 596
rect 17 546 37 580
rect 71 546 87 580
rect 17 497 87 546
rect 17 463 37 497
rect 71 463 87 497
rect 17 414 87 463
rect 17 380 37 414
rect 71 380 87 414
rect 17 364 87 380
rect 127 580 177 649
rect 161 546 177 580
rect 127 497 177 546
rect 161 463 177 497
rect 127 414 177 463
rect 161 380 177 414
rect 127 364 177 380
rect 249 580 321 596
rect 249 546 287 580
rect 249 510 321 546
rect 249 476 287 510
rect 249 440 321 476
rect 249 406 287 440
rect 249 390 321 406
rect 361 580 427 596
rect 361 546 377 580
rect 411 546 427 580
rect 361 510 427 546
rect 361 476 377 510
rect 411 476 427 510
rect 361 440 427 476
rect 467 580 507 649
rect 467 546 470 580
rect 504 546 507 580
rect 467 508 507 546
rect 467 474 470 508
rect 504 474 507 508
rect 467 458 507 474
rect 547 580 613 596
rect 547 546 563 580
rect 597 546 613 580
rect 547 509 613 546
rect 547 475 563 509
rect 597 475 613 509
rect 361 406 377 440
rect 411 424 427 440
rect 547 438 613 475
rect 547 424 563 438
rect 411 406 563 424
rect 361 404 563 406
rect 597 404 613 438
rect 361 390 613 404
rect 17 230 51 364
rect 249 330 283 390
rect 547 388 613 390
rect 85 314 283 330
rect 85 280 101 314
rect 135 280 283 314
rect 317 340 367 356
rect 351 306 367 340
rect 317 290 367 306
rect 409 340 475 356
rect 409 306 425 340
rect 459 306 475 340
rect 409 290 475 306
rect 85 264 283 280
rect 249 256 283 264
rect 249 246 427 256
rect 17 196 215 230
rect 249 222 377 246
rect 165 194 215 196
rect 165 160 181 194
rect 361 212 377 222
rect 411 212 427 246
rect 165 134 215 160
rect 251 172 317 188
rect 251 138 267 172
rect 301 138 317 172
rect 251 17 317 138
rect 361 178 427 212
rect 542 235 608 268
rect 542 202 558 235
rect 361 144 377 178
rect 411 144 427 178
rect 361 132 427 144
rect 461 201 558 202
rect 592 201 608 235
rect 461 168 608 201
rect 461 17 495 168
rect 601 114 647 134
rect 529 98 647 114
rect 529 64 545 98
rect 579 64 647 98
rect 529 51 647 64
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a21o_1
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 607 94 641 128 0 FreeSans 340 0 0 0 A2
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 672 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 4084908
string GDS_START 4078508
<< end >>
