magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 25 258 109 392
rect 161 326 257 430
rect 1066 271 1132 356
rect 1447 364 1517 596
rect 1483 226 1517 364
rect 1448 70 1517 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 23 426 89 649
rect 191 498 257 596
rect 303 532 369 649
rect 522 498 572 551
rect 191 464 572 498
rect 612 485 678 551
rect 797 488 863 649
rect 898 533 964 580
rect 1117 567 1198 649
rect 898 499 1200 533
rect 291 292 325 464
rect 143 258 325 292
rect 359 343 476 430
rect 522 377 572 464
rect 359 309 580 343
rect 143 224 177 258
rect 359 224 393 309
rect 525 277 580 309
rect 614 310 678 485
rect 898 424 964 499
rect 720 348 964 424
rect 998 399 1076 465
rect 23 17 73 224
rect 109 142 177 224
rect 313 190 393 224
rect 427 240 483 272
rect 614 244 864 310
rect 427 206 543 240
rect 313 176 379 190
rect 425 142 475 156
rect 109 108 475 142
rect 211 17 277 74
rect 425 70 475 108
rect 509 85 543 206
rect 614 185 648 244
rect 898 210 936 348
rect 998 226 1032 399
rect 1166 310 1200 499
rect 1239 378 1305 575
rect 1339 412 1405 649
rect 1239 344 1329 378
rect 1295 326 1329 344
rect 1166 244 1261 310
rect 1295 260 1449 326
rect 577 119 648 185
rect 682 176 852 210
rect 682 85 716 176
rect 509 51 716 85
rect 750 17 784 142
rect 818 85 852 176
rect 886 119 936 210
rect 980 85 1046 226
rect 818 51 1046 85
rect 1082 17 1132 226
rect 1295 210 1329 260
rect 1233 90 1329 210
rect 1363 17 1413 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
rlabel locali s 161 326 257 430 6 GATE
port 1 nsew signal input
rlabel locali s 1483 226 1517 364 6 GCLK
port 2 nsew signal output
rlabel locali s 1448 70 1517 226 6 GCLK
port 2 nsew signal output
rlabel locali s 1447 364 1517 596 6 GCLK
port 2 nsew signal output
rlabel locali s 25 258 109 392 6 SCE
port 3 nsew signal input
rlabel locali s 1066 271 1132 356 6 CLK
port 4 nsew clock input
rlabel metal1 s 0 -49 1536 49 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1536 715 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1536 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 420810
string GDS_START 409002
<< end >>
