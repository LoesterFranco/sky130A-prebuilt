magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 103 333 179 419
rect 605 333 681 417
rect 103 299 681 333
rect 18 215 179 265
rect 213 215 363 265
rect 397 221 474 299
rect 397 181 449 221
rect 531 215 673 265
rect 744 215 986 265
rect 1040 215 1259 265
rect 103 131 449 181
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 18 459 273 493
rect 18 299 69 459
rect 223 401 273 459
rect 317 435 351 527
rect 385 401 461 491
rect 223 367 461 401
rect 517 451 967 489
rect 517 367 567 451
rect 725 299 759 451
rect 803 333 869 417
rect 917 367 967 451
rect 1014 367 1055 527
rect 1099 333 1165 492
rect 803 299 1165 333
rect 1209 299 1253 527
rect 18 97 69 181
rect 497 143 1261 181
rect 497 97 531 143
rect 18 51 531 97
rect 574 17 650 109
rect 687 51 763 143
rect 807 17 841 109
rect 901 51 1035 143
rect 1071 17 1147 109
rect 1195 51 1261 143
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
rlabel locali s 1040 215 1259 265 6 A1
port 1 nsew signal input
rlabel locali s 744 215 986 265 6 A2
port 2 nsew signal input
rlabel locali s 531 215 673 265 6 A3
port 3 nsew signal input
rlabel locali s 213 215 363 265 6 B1
port 4 nsew signal input
rlabel locali s 18 215 179 265 6 B2
port 5 nsew signal input
rlabel locali s 605 333 681 417 6 Y
port 6 nsew signal output
rlabel locali s 397 221 474 299 6 Y
port 6 nsew signal output
rlabel locali s 397 181 449 221 6 Y
port 6 nsew signal output
rlabel locali s 103 333 179 419 6 Y
port 6 nsew signal output
rlabel locali s 103 299 681 333 6 Y
port 6 nsew signal output
rlabel locali s 103 131 449 181 6 Y
port 6 nsew signal output
rlabel metal1 s 0 -48 1288 48 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 496 1288 592 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1288 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 591166
string GDS_START 580822
<< end >>
