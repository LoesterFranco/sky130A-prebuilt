magic
tech sky130A
magscale 1 2
timestamp 1599588238
<< locali >>
rect 105 316 171 430
rect 221 364 315 430
rect 105 282 409 316
rect 343 250 409 282
rect 511 220 567 430
rect 669 236 743 310
rect 2809 430 2865 596
rect 3005 430 3039 596
rect 2809 364 3039 430
rect 3005 356 3039 364
rect 3005 322 3143 356
rect 3097 288 3143 322
rect 2979 254 3143 288
rect 2979 230 3045 254
rect 2779 196 3045 230
rect 2779 70 2845 196
rect 2979 70 3045 196
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3168 683
rect 21 498 71 596
rect 111 532 177 649
rect 285 532 477 582
rect 512 566 578 649
rect 443 498 635 532
rect 714 516 780 649
rect 814 579 1166 613
rect 814 516 880 579
rect 21 464 409 498
rect 21 248 71 464
rect 357 366 409 464
rect 21 182 228 248
rect 443 216 477 498
rect 601 482 635 498
rect 940 482 1006 545
rect 601 448 1006 482
rect 601 364 843 414
rect 358 182 477 216
rect 601 202 635 364
rect 777 270 843 364
rect 882 380 1006 448
rect 1040 455 1096 545
rect 1132 492 1166 579
rect 1255 526 1305 649
rect 1339 579 1509 613
rect 1339 492 1373 579
rect 1132 458 1373 492
rect 21 70 89 182
rect 358 148 392 182
rect 123 17 189 148
rect 295 82 392 148
rect 490 17 556 148
rect 601 70 678 202
rect 712 17 778 202
rect 814 85 848 226
rect 882 185 916 380
rect 950 253 1006 346
rect 1040 321 1074 455
rect 1132 421 1166 458
rect 1407 424 1441 545
rect 1108 355 1166 421
rect 1208 390 1441 424
rect 1475 424 1509 579
rect 1543 458 1577 649
rect 1617 458 1673 543
rect 1707 492 1773 649
rect 1819 572 2075 615
rect 1819 520 1875 572
rect 1909 458 1975 538
rect 2009 496 2075 572
rect 2109 530 2191 596
rect 2225 530 2275 649
rect 2315 496 2381 596
rect 2427 530 2510 596
rect 2009 462 2442 496
rect 1617 424 1975 458
rect 1475 390 1579 424
rect 1909 420 1975 424
rect 1208 356 1274 390
rect 1545 386 1875 390
rect 2087 386 2153 427
rect 1545 356 2153 386
rect 1325 321 1391 356
rect 1040 287 1391 321
rect 1439 350 1511 356
rect 1439 316 1471 350
rect 1505 316 1511 350
rect 1439 290 1511 316
rect 1809 352 2153 356
rect 1809 290 1875 352
rect 2187 314 2221 462
rect 950 219 1028 253
rect 882 119 960 185
rect 994 85 1028 219
rect 814 51 1028 85
rect 1062 77 1128 287
rect 1325 256 1391 287
rect 1587 256 1653 290
rect 2042 280 2221 314
rect 2294 350 2374 428
rect 2294 316 2335 350
rect 2369 316 2374 350
rect 2294 294 2374 316
rect 2408 402 2442 462
rect 2476 470 2510 530
rect 2544 504 2594 649
rect 2476 436 2542 470
rect 1201 188 1267 253
rect 1325 222 1653 256
rect 1688 222 2006 256
rect 1201 154 1420 188
rect 1242 17 1308 120
rect 1354 70 1420 154
rect 1518 17 1652 186
rect 1688 70 1722 222
rect 1758 17 1824 188
rect 1870 85 1936 188
rect 1972 119 2006 222
rect 2042 85 2108 280
rect 2408 268 2474 402
rect 2191 214 2257 246
rect 2508 214 2542 436
rect 2634 330 2668 596
rect 2708 420 2774 649
rect 2899 464 2965 649
rect 3079 390 3145 649
rect 2634 298 2939 330
rect 2191 180 2542 214
rect 1870 51 2108 85
rect 2330 17 2430 136
rect 2464 70 2542 180
rect 2576 264 2939 298
rect 2576 70 2642 264
rect 2676 17 2742 226
rect 2879 17 2945 162
rect 3079 17 3145 220
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3168 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 1471 316 1505 350
rect 2335 316 2369 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
<< metal1 >>
rect 0 683 3168 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3168 683
rect 0 617 3168 649
rect 1459 350 1517 356
rect 1459 316 1471 350
rect 1505 347 1517 350
rect 2323 350 2381 356
rect 2323 347 2335 350
rect 1505 319 2335 347
rect 1505 316 1517 319
rect 1459 310 1517 316
rect 2323 316 2335 319
rect 2369 316 2381 350
rect 2323 310 2381 316
rect 0 17 3168 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3168 17
rect 0 -49 3168 -17
<< labels >>
rlabel locali s 221 364 315 430 6 D
port 1 nsew signal input
rlabel locali s 3097 288 3143 322 6 Q
port 2 nsew signal output
rlabel locali s 3005 430 3039 596 6 Q
port 2 nsew signal output
rlabel locali s 3005 356 3039 364 6 Q
port 2 nsew signal output
rlabel locali s 3005 322 3143 356 6 Q
port 2 nsew signal output
rlabel locali s 2979 254 3143 288 6 Q
port 2 nsew signal output
rlabel locali s 2979 230 3045 254 6 Q
port 2 nsew signal output
rlabel locali s 2979 70 3045 196 6 Q
port 2 nsew signal output
rlabel locali s 2809 430 2865 596 6 Q
port 2 nsew signal output
rlabel locali s 2809 364 3039 430 6 Q
port 2 nsew signal output
rlabel locali s 2779 196 3045 230 6 Q
port 2 nsew signal output
rlabel locali s 2779 70 2845 196 6 Q
port 2 nsew signal output
rlabel locali s 511 220 567 430 6 SCD
port 3 nsew signal input
rlabel locali s 343 250 409 282 6 SCE
port 4 nsew signal input
rlabel locali s 105 316 171 430 6 SCE
port 4 nsew signal input
rlabel locali s 105 282 409 316 6 SCE
port 4 nsew signal input
rlabel metal1 s 2323 347 2381 356 6 SET_B
port 5 nsew signal input
rlabel metal1 s 2323 310 2381 319 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1459 347 1517 356 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1459 319 2381 347 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1459 310 1517 319 6 SET_B
port 5 nsew signal input
rlabel locali s 669 236 743 310 6 CLK
port 6 nsew clock input
rlabel metal1 s 0 -49 3168 49 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 617 3168 715 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 3168 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 319886
string GDS_START 296922
<< end >>
