magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 736 561
rect 104 441 182 527
rect 283 441 446 527
rect 119 265 155 339
rect 85 199 155 265
rect 189 299 270 339
rect 119 17 155 165
rect 189 119 223 299
rect 640 375 706 527
rect 489 215 586 257
rect 620 215 719 325
rect 189 51 248 119
rect 282 17 354 97
rect 583 17 617 111
rect 0 -17 736 17
<< obsli1 >>
rect 480 407 545 493
rect 17 373 387 407
rect 17 299 79 373
rect 17 165 51 299
rect 17 86 69 165
rect 257 212 291 265
rect 257 178 319 212
rect 353 199 387 373
rect 421 291 545 407
rect 285 165 319 178
rect 421 165 455 291
rect 285 131 455 165
rect 388 51 455 131
rect 489 147 718 181
rect 489 73 549 147
rect 651 54 718 147
<< metal1 >>
rect 0 496 736 592
rect 0 -48 736 48
<< labels >>
rlabel locali s 620 215 719 325 6 A1
port 1 nsew signal input
rlabel locali s 489 215 586 257 6 A2
port 2 nsew signal input
rlabel locali s 119 265 155 339 6 B1_N
port 3 nsew signal input
rlabel locali s 85 199 155 265 6 B1_N
port 3 nsew signal input
rlabel locali s 189 299 270 339 6 X
port 4 nsew signal output
rlabel locali s 189 119 223 299 6 X
port 4 nsew signal output
rlabel locali s 189 51 248 119 6 X
port 4 nsew signal output
rlabel locali s 583 17 617 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 282 17 354 97 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 119 17 155 165 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 736 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 736 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 640 375 706 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 283 441 446 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 104 441 182 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 736 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 736 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1379784
string GDS_START 1373496
<< end >>
