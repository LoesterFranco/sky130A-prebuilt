magic
tech sky130A
magscale 1 2
timestamp 1604502729
<< locali >>
rect 313 378 363 596
rect 21 236 87 310
rect 121 270 210 356
rect 244 344 363 378
rect 244 236 278 344
rect 312 238 363 310
rect 184 202 278 236
rect 184 70 258 202
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 384 683
rect 21 446 80 596
rect 114 480 180 649
rect 214 446 273 596
rect 21 412 273 446
rect 21 397 191 412
rect 21 364 87 397
rect 26 17 92 202
rect 312 17 358 204
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 384 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
<< metal1 >>
rect 0 683 384 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 384 683
rect 0 617 384 649
rect 0 17 384 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 384 17
rect 0 -49 384 -17
<< labels >>
rlabel locali s 121 270 210 356 6 A1
port 1 nsew signal input
rlabel locali s 21 236 87 310 6 A2
port 2 nsew signal input
rlabel locali s 312 238 363 310 6 B1
port 3 nsew signal input
rlabel locali s 313 378 363 596 6 Y
port 4 nsew signal output
rlabel locali s 244 344 363 378 6 Y
port 4 nsew signal output
rlabel locali s 244 236 278 344 6 Y
port 4 nsew signal output
rlabel locali s 184 202 278 236 6 Y
port 4 nsew signal output
rlabel locali s 184 70 258 202 6 Y
port 4 nsew signal output
rlabel metal1 s 0 -49 384 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 617 384 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 384 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 4110954
string GDS_START 4106040
<< end >>
