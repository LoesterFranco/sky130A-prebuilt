magic
tech sky130A
magscale 1 2
timestamp 1604502729
<< locali >>
rect 87 256 161 310
rect 195 290 263 356
rect 297 256 369 318
rect 87 252 369 256
rect 87 236 331 252
rect 127 222 331 236
rect 297 118 331 222
rect 567 256 621 356
rect 663 290 737 356
rect 771 290 839 356
rect 879 256 945 310
rect 1095 256 1149 350
rect 567 222 1149 256
rect 1183 236 1269 356
rect 1380 290 1511 356
rect 567 118 621 222
rect 297 84 621 118
rect 1930 364 2000 596
rect 1930 88 1996 364
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 51 430 117 596
rect 19 384 117 430
rect 151 390 217 649
rect 19 202 53 384
rect 409 290 465 430
rect 499 424 689 596
rect 723 458 789 649
rect 1011 532 1189 582
rect 1233 542 1299 649
rect 1440 581 1826 615
rect 1440 542 1506 581
rect 1155 508 1189 532
rect 1562 513 1758 547
rect 1562 508 1596 513
rect 823 464 1121 498
rect 1155 474 1596 508
rect 823 424 857 464
rect 1087 440 1121 464
rect 499 390 857 424
rect 19 100 93 202
rect 164 17 230 188
rect 499 218 533 390
rect 370 152 533 218
rect 985 292 1053 430
rect 1087 392 1416 440
rect 1312 390 1416 392
rect 1530 390 1596 474
rect 1312 256 1346 390
rect 1640 356 1690 479
rect 1545 290 1690 356
rect 1312 222 1591 256
rect 689 17 785 188
rect 906 154 1603 188
rect 1637 187 1690 290
rect 906 70 1021 154
rect 1228 17 1294 120
rect 1338 70 1388 154
rect 1569 153 1603 154
rect 1724 153 1758 513
rect 1424 85 1490 120
rect 1569 119 1758 153
rect 1792 336 1826 581
rect 1860 370 1894 649
rect 2040 364 2090 649
rect 1792 270 1877 336
rect 1792 85 1826 270
rect 1424 51 1826 85
rect 1860 17 1894 236
rect 2032 17 2082 252
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
<< metal1 >>
rect 0 683 2112 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 0 617 2112 649
rect 0 17 2112 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
rect 0 -49 2112 -17
<< obsm1 >>
rect 19 421 77 430
rect 403 421 461 430
rect 979 421 1037 430
rect 19 393 1037 421
rect 19 384 77 393
rect 403 384 461 393
rect 979 384 1037 393
<< labels >>
rlabel locali s 663 290 737 356 6 A0
port 1 nsew signal input
rlabel locali s 195 290 263 356 6 A1
port 2 nsew signal input
rlabel locali s 1183 236 1269 356 6 A2
port 3 nsew signal input
rlabel locali s 771 290 839 356 6 A3
port 4 nsew signal input
rlabel locali s 1095 256 1149 350 6 S0
port 5 nsew signal input
rlabel locali s 879 256 945 310 6 S0
port 5 nsew signal input
rlabel locali s 567 256 621 356 6 S0
port 5 nsew signal input
rlabel locali s 567 222 1149 256 6 S0
port 5 nsew signal input
rlabel locali s 567 118 621 222 6 S0
port 5 nsew signal input
rlabel locali s 297 256 369 318 6 S0
port 5 nsew signal input
rlabel locali s 297 118 331 222 6 S0
port 5 nsew signal input
rlabel locali s 297 84 621 118 6 S0
port 5 nsew signal input
rlabel locali s 127 222 331 236 6 S0
port 5 nsew signal input
rlabel locali s 87 256 161 310 6 S0
port 5 nsew signal input
rlabel locali s 87 252 369 256 6 S0
port 5 nsew signal input
rlabel locali s 87 236 331 252 6 S0
port 5 nsew signal input
rlabel locali s 1380 290 1511 356 6 S1
port 6 nsew signal input
rlabel locali s 1930 364 2000 596 6 X
port 7 nsew signal output
rlabel locali s 1930 88 1996 364 6 X
port 7 nsew signal output
rlabel metal1 s 0 -49 2112 49 8 VGND
port 8 nsew ground bidirectional
rlabel metal1 s 0 617 2112 715 6 VPWR
port 9 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2112 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1976282
string GDS_START 1960810
<< end >>
