magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1196 561
rect 127 379 193 527
rect 483 345 533 425
rect 667 345 701 493
rect 735 379 869 527
rect 903 345 965 493
rect 999 379 1065 527
rect 1099 345 1179 493
rect 483 297 1179 345
rect 17 211 221 263
rect 255 211 431 263
rect 465 211 615 263
rect 673 211 877 263
rect 911 177 983 297
rect 1017 211 1179 263
rect 911 131 1179 177
rect 131 17 197 97
rect 299 17 365 97
rect 467 17 621 97
rect 1103 51 1179 131
rect 0 -17 1196 17
<< obsli1 >>
rect 17 345 93 493
rect 227 345 261 493
rect 295 459 633 493
rect 295 379 361 459
rect 395 345 445 425
rect 17 297 445 345
rect 567 379 633 459
rect 17 131 877 177
rect 17 51 97 131
rect 231 51 265 131
rect 399 51 433 131
rect 655 51 689 131
rect 723 51 1069 97
<< metal1 >>
rect 0 496 1196 592
rect 0 -48 1196 48
<< labels >>
rlabel locali s 17 211 221 263 6 A1
port 1 nsew signal input
rlabel locali s 255 211 431 263 6 A2
port 2 nsew signal input
rlabel locali s 465 211 615 263 6 A3
port 3 nsew signal input
rlabel locali s 673 211 877 263 6 B1
port 4 nsew signal input
rlabel locali s 1017 211 1179 263 6 C1
port 5 nsew signal input
rlabel locali s 1103 51 1179 131 6 Y
port 6 nsew signal output
rlabel locali s 1099 345 1179 493 6 Y
port 6 nsew signal output
rlabel locali s 911 177 983 297 6 Y
port 6 nsew signal output
rlabel locali s 911 131 1179 177 6 Y
port 6 nsew signal output
rlabel locali s 903 345 965 493 6 Y
port 6 nsew signal output
rlabel locali s 667 345 701 493 6 Y
port 6 nsew signal output
rlabel locali s 483 345 533 425 6 Y
port 6 nsew signal output
rlabel locali s 483 297 1179 345 6 Y
port 6 nsew signal output
rlabel locali s 467 17 621 97 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 299 17 365 97 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 131 17 197 97 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 1196 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1196 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 999 379 1065 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 735 379 869 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 127 379 193 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 1196 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 1196 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 793012
string GDS_START 782616
<< end >>
