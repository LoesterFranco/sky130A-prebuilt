magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 2024 561
rect 501 451 635 527
rect 21 261 65 393
rect 103 349 169 417
rect 270 349 337 417
rect 737 383 803 527
rect 103 337 337 349
rect 924 383 990 527
rect 1099 383 1233 527
rect 1345 383 1411 527
rect 1513 383 1579 527
rect 1681 383 1747 527
rect 1849 383 1915 527
rect 103 315 431 337
rect 270 299 431 315
rect 21 215 349 261
rect 387 161 431 299
rect 477 199 841 265
rect 881 215 1263 257
rect 1312 215 1591 260
rect 1657 215 1995 256
rect 119 127 803 161
rect 18 17 85 93
rect 119 51 153 127
rect 187 17 253 93
rect 287 51 321 127
rect 355 17 421 93
rect 1681 17 1747 93
rect 1849 17 1915 93
rect 0 -17 2024 17
<< obsli1 >>
rect 433 485 467 493
rect 18 451 467 485
rect 433 415 467 451
rect 669 415 703 493
rect 433 381 703 415
rect 669 349 703 381
rect 837 349 871 485
rect 1024 349 1058 493
rect 1277 349 1311 493
rect 1445 349 1479 493
rect 1613 349 1647 493
rect 1781 349 1815 493
rect 1955 349 1989 493
rect 669 315 1989 349
rect 905 127 1579 161
rect 1613 127 1983 161
rect 1613 93 1647 127
rect 485 59 1223 93
rect 1261 59 1647 93
rect 1613 51 1647 59
rect 1781 51 1815 127
rect 1949 51 1983 127
<< metal1 >>
rect 0 496 2024 592
rect 0 -48 2024 48
<< labels >>
rlabel locali s 477 199 841 265 6 A1
port 1 nsew signal input
rlabel locali s 881 215 1263 257 6 A2
port 2 nsew signal input
rlabel locali s 1312 215 1591 260 6 A3
port 3 nsew signal input
rlabel locali s 1657 215 1995 256 6 A4
port 4 nsew signal input
rlabel locali s 21 261 65 393 6 B1
port 5 nsew signal input
rlabel locali s 21 215 349 261 6 B1
port 5 nsew signal input
rlabel locali s 387 161 431 299 6 Y
port 6 nsew signal output
rlabel locali s 287 51 321 127 6 Y
port 6 nsew signal output
rlabel locali s 270 349 337 417 6 Y
port 6 nsew signal output
rlabel locali s 270 299 431 315 6 Y
port 6 nsew signal output
rlabel locali s 119 127 803 161 6 Y
port 6 nsew signal output
rlabel locali s 119 51 153 127 6 Y
port 6 nsew signal output
rlabel locali s 103 349 169 417 6 Y
port 6 nsew signal output
rlabel locali s 103 337 337 349 6 Y
port 6 nsew signal output
rlabel locali s 103 315 431 337 6 Y
port 6 nsew signal output
rlabel locali s 1849 17 1915 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1681 17 1747 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 355 17 421 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 187 17 253 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 18 17 85 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 2024 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 2024 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1849 383 1915 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1681 383 1747 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1513 383 1579 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1345 383 1411 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1099 383 1233 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 924 383 990 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 737 383 803 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 501 451 635 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 2024 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 2024 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2024 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3737160
string GDS_START 3720602
<< end >>
