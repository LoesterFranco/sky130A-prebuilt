magic
tech sky130A
magscale 1 2
timestamp 1601050047
<< nwell >>
rect -38 332 710 704
<< pwell >>
rect 0 0 672 49
<< scpmos >>
rect 87 392 117 592
rect 165 392 195 592
rect 369 368 399 592
rect 459 368 489 592
rect 555 368 585 592
<< nmoslvt >>
rect 96 112 126 222
rect 182 112 212 222
rect 372 74 402 222
rect 458 74 488 222
rect 552 74 582 222
<< ndiff >>
rect 43 180 96 222
rect 43 146 51 180
rect 85 146 96 180
rect 43 112 96 146
rect 126 184 182 222
rect 126 150 137 184
rect 171 150 182 184
rect 126 112 182 150
rect 212 158 372 222
rect 212 124 237 158
rect 271 142 372 158
rect 271 124 327 142
rect 212 112 327 124
rect 319 108 327 112
rect 361 108 372 142
rect 319 74 372 108
rect 402 194 458 222
rect 402 160 413 194
rect 447 160 458 194
rect 402 120 458 160
rect 402 86 413 120
rect 447 86 458 120
rect 402 74 458 86
rect 488 74 552 222
rect 582 196 635 222
rect 582 162 593 196
rect 627 162 635 196
rect 582 120 635 162
rect 582 86 593 120
rect 627 86 635 120
rect 582 74 635 86
<< pdiff >>
rect 32 580 87 592
rect 32 546 40 580
rect 74 546 87 580
rect 32 510 87 546
rect 32 476 40 510
rect 74 476 87 510
rect 32 440 87 476
rect 32 406 40 440
rect 74 406 87 440
rect 32 392 87 406
rect 117 392 165 592
rect 195 580 250 592
rect 195 546 208 580
rect 242 546 250 580
rect 195 510 250 546
rect 195 476 208 510
rect 242 476 250 510
rect 195 440 250 476
rect 195 406 208 440
rect 242 406 250 440
rect 195 392 250 406
rect 314 580 369 592
rect 314 546 322 580
rect 356 546 369 580
rect 314 497 369 546
rect 314 463 322 497
rect 356 463 369 497
rect 314 414 369 463
rect 314 380 322 414
rect 356 380 369 414
rect 314 368 369 380
rect 399 554 459 592
rect 399 520 412 554
rect 446 520 459 554
rect 399 368 459 520
rect 489 580 555 592
rect 489 546 505 580
rect 539 546 555 580
rect 489 368 555 546
rect 585 580 640 592
rect 585 546 598 580
rect 632 546 640 580
rect 585 497 640 546
rect 585 463 598 497
rect 632 463 640 497
rect 585 414 640 463
rect 585 380 598 414
rect 632 380 640 414
rect 585 368 640 380
<< ndiffc >>
rect 51 146 85 180
rect 137 150 171 184
rect 237 124 271 158
rect 327 108 361 142
rect 413 160 447 194
rect 413 86 447 120
rect 593 162 627 196
rect 593 86 627 120
<< pdiffc >>
rect 40 546 74 580
rect 40 476 74 510
rect 40 406 74 440
rect 208 546 242 580
rect 208 476 242 510
rect 208 406 242 440
rect 322 546 356 580
rect 322 463 356 497
rect 322 380 356 414
rect 412 520 446 554
rect 505 546 539 580
rect 598 546 632 580
rect 598 463 632 497
rect 598 380 632 414
<< poly >>
rect 87 592 117 618
rect 165 592 195 618
rect 369 592 399 618
rect 459 592 489 618
rect 555 592 585 618
rect 87 377 117 392
rect 165 377 195 392
rect 84 318 120 377
rect 21 302 120 318
rect 162 366 198 377
rect 162 340 234 366
rect 369 353 399 368
rect 459 353 489 368
rect 555 353 585 368
rect 162 306 184 340
rect 218 306 234 340
rect 366 310 402 353
rect 456 310 492 353
rect 552 310 588 353
rect 162 305 234 306
rect 21 268 37 302
rect 71 282 120 302
rect 168 290 234 305
rect 276 294 402 310
rect 71 268 126 282
rect 21 252 126 268
rect 96 222 126 252
rect 182 222 212 290
rect 276 260 292 294
rect 326 260 402 294
rect 276 244 402 260
rect 444 294 510 310
rect 444 260 460 294
rect 494 260 510 294
rect 444 244 510 260
rect 552 294 651 310
rect 552 260 601 294
rect 635 260 651 294
rect 552 244 651 260
rect 372 222 402 244
rect 458 222 488 244
rect 552 222 582 244
rect 96 86 126 112
rect 182 86 212 112
rect 372 48 402 74
rect 458 48 488 74
rect 552 48 582 74
<< polycont >>
rect 184 306 218 340
rect 37 268 71 302
rect 292 260 326 294
rect 460 260 494 294
rect 601 260 635 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 24 580 90 649
rect 486 596 520 649
rect 24 546 40 580
rect 74 546 90 580
rect 24 510 90 546
rect 24 476 40 510
rect 74 476 90 510
rect 24 440 90 476
rect 24 406 40 440
rect 74 406 90 440
rect 24 390 90 406
rect 192 580 258 596
rect 192 546 208 580
rect 242 546 258 580
rect 192 510 258 546
rect 192 476 208 510
rect 242 476 258 510
rect 192 440 258 476
rect 306 580 356 596
rect 306 546 322 580
rect 306 497 356 546
rect 306 463 322 497
rect 396 554 446 596
rect 396 520 412 554
rect 486 580 558 596
rect 486 546 505 580
rect 539 546 558 580
rect 598 580 648 596
rect 632 546 648 580
rect 396 512 446 520
rect 598 512 648 546
rect 396 497 648 512
rect 396 478 598 497
rect 306 458 356 463
rect 192 406 208 440
rect 242 424 258 440
rect 322 444 356 458
rect 632 463 648 497
rect 242 406 288 424
rect 192 390 288 406
rect 21 302 87 356
rect 21 268 37 302
rect 71 268 87 302
rect 121 340 220 356
rect 121 306 184 340
rect 218 306 220 340
rect 121 290 220 306
rect 254 310 288 390
rect 322 414 455 444
rect 356 384 455 414
rect 356 380 410 384
rect 322 350 410 380
rect 254 294 342 310
rect 21 252 87 268
rect 254 260 292 294
rect 326 260 342 294
rect 254 244 342 260
rect 254 226 288 244
rect 35 180 85 218
rect 35 146 51 180
rect 35 17 85 146
rect 121 192 288 226
rect 376 210 410 350
rect 505 308 551 430
rect 598 414 648 463
rect 632 380 648 414
rect 598 364 648 380
rect 444 294 551 308
rect 444 260 460 294
rect 494 260 551 294
rect 444 244 551 260
rect 585 294 651 310
rect 585 260 601 294
rect 635 260 651 294
rect 585 236 651 260
rect 376 194 463 210
rect 121 184 187 192
rect 121 150 137 184
rect 171 150 187 184
rect 376 176 413 194
rect 411 160 413 176
rect 447 160 463 194
rect 121 108 187 150
rect 221 124 237 158
rect 271 142 342 158
rect 271 124 327 142
rect 221 108 327 124
rect 361 108 377 142
rect 221 17 377 108
rect 411 120 463 160
rect 411 86 413 120
rect 447 86 463 120
rect 411 70 463 86
rect 577 196 643 202
rect 577 162 593 196
rect 627 162 643 196
rect 577 120 643 162
rect 577 86 593 120
rect 627 86 643 120
rect 577 17 643 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a2bb2oi_1
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 415 390 449 424 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 A2_N
port 2 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 A1_N
port 1 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 511 390 545 424 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 607 242 641 276 0 FreeSans 340 0 0 0 B1
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 672 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3763852
string GDS_START 3757220
<< end >>
