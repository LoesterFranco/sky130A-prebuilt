magic
tech sky130A
magscale 1 2
timestamp 1604502705
<< nwell >>
rect -38 332 1766 704
<< pwell >>
rect 0 0 1728 49
<< scnmos >>
rect 93 74 123 222
rect 357 74 387 222
rect 457 74 487 222
rect 727 74 757 222
rect 827 74 857 222
rect 913 74 943 222
rect 1409 74 1439 222
rect 1581 74 1611 222
<< pmoshvt >>
rect 96 368 126 592
rect 186 368 216 592
rect 276 368 306 592
rect 376 368 406 592
rect 466 368 496 592
rect 556 368 586 592
rect 646 368 676 592
rect 736 368 766 592
rect 938 368 968 592
rect 1028 368 1058 592
rect 1122 368 1152 592
rect 1212 368 1242 592
rect 1302 368 1332 592
rect 1412 368 1442 592
rect 1502 368 1532 592
rect 1612 368 1642 592
<< ndiff >>
rect 27 152 93 222
rect 27 118 39 152
rect 73 118 93 152
rect 27 74 93 118
rect 123 210 357 222
rect 123 176 134 210
rect 168 176 218 210
rect 252 176 312 210
rect 346 176 357 210
rect 123 120 357 176
rect 123 86 134 120
rect 168 86 218 120
rect 252 86 312 120
rect 346 86 357 120
rect 123 74 357 86
rect 387 152 457 222
rect 387 118 398 152
rect 432 118 457 152
rect 387 74 457 118
rect 487 210 727 222
rect 487 176 498 210
rect 532 176 583 210
rect 617 176 682 210
rect 716 176 727 210
rect 487 120 727 176
rect 487 86 498 120
rect 532 86 583 120
rect 617 86 682 120
rect 716 86 727 120
rect 487 74 727 86
rect 757 152 827 222
rect 757 118 768 152
rect 802 118 827 152
rect 757 74 827 118
rect 857 210 913 222
rect 857 176 868 210
rect 902 176 913 210
rect 857 120 913 176
rect 857 86 868 120
rect 902 86 913 120
rect 857 74 913 86
rect 943 142 1409 222
rect 943 108 954 142
rect 988 108 1039 142
rect 1073 108 1118 142
rect 1152 108 1198 142
rect 1232 108 1277 142
rect 1311 108 1364 142
rect 1398 108 1409 142
rect 943 74 1409 108
rect 1439 210 1581 222
rect 1439 176 1450 210
rect 1484 186 1581 210
rect 1484 176 1536 186
rect 1439 152 1536 176
rect 1570 152 1581 186
rect 1439 120 1581 152
rect 1439 86 1450 120
rect 1484 118 1581 120
rect 1484 86 1536 118
rect 1439 84 1536 86
rect 1570 84 1581 118
rect 1439 74 1581 84
rect 1611 202 1668 222
rect 1611 168 1622 202
rect 1656 168 1668 202
rect 1611 120 1668 168
rect 1611 86 1622 120
rect 1656 86 1668 120
rect 1611 74 1668 86
<< pdiff >>
rect 27 580 96 592
rect 27 546 39 580
rect 73 546 96 580
rect 27 508 96 546
rect 27 474 39 508
rect 73 474 96 508
rect 27 368 96 474
rect 126 531 186 592
rect 126 497 139 531
rect 173 497 186 531
rect 126 440 186 497
rect 126 406 139 440
rect 173 406 186 440
rect 126 368 186 406
rect 216 580 276 592
rect 216 546 229 580
rect 263 546 276 580
rect 216 508 276 546
rect 216 474 229 508
rect 263 474 276 508
rect 216 368 276 474
rect 306 531 376 592
rect 306 497 329 531
rect 363 497 376 531
rect 306 440 376 497
rect 306 406 329 440
rect 363 406 376 440
rect 306 368 376 406
rect 406 580 466 592
rect 406 546 419 580
rect 453 546 466 580
rect 406 497 466 546
rect 406 463 419 497
rect 453 463 466 497
rect 406 414 466 463
rect 406 380 419 414
rect 453 380 466 414
rect 406 368 466 380
rect 496 580 556 592
rect 496 546 509 580
rect 543 546 556 580
rect 496 492 556 546
rect 496 458 509 492
rect 543 458 556 492
rect 496 368 556 458
rect 586 531 646 592
rect 586 497 599 531
rect 633 497 646 531
rect 586 424 646 497
rect 586 390 599 424
rect 633 390 646 424
rect 586 368 646 390
rect 676 580 736 592
rect 676 546 689 580
rect 723 546 736 580
rect 676 492 736 546
rect 676 458 689 492
rect 723 458 736 492
rect 676 368 736 458
rect 766 531 825 592
rect 766 497 779 531
rect 813 497 825 531
rect 766 440 825 497
rect 766 406 779 440
rect 813 406 825 440
rect 766 368 825 406
rect 879 531 938 592
rect 879 497 891 531
rect 925 497 938 531
rect 879 424 938 497
rect 879 390 891 424
rect 925 390 938 424
rect 879 368 938 390
rect 968 580 1028 592
rect 968 546 981 580
rect 1015 546 1028 580
rect 968 494 1028 546
rect 968 460 981 494
rect 1015 460 1028 494
rect 968 368 1028 460
rect 1058 531 1122 592
rect 1058 497 1073 531
rect 1107 497 1122 531
rect 1058 424 1122 497
rect 1058 390 1073 424
rect 1107 390 1122 424
rect 1058 368 1122 390
rect 1152 580 1212 592
rect 1152 546 1165 580
rect 1199 546 1212 580
rect 1152 494 1212 546
rect 1152 460 1165 494
rect 1199 460 1212 494
rect 1152 368 1212 460
rect 1242 580 1302 592
rect 1242 546 1255 580
rect 1289 546 1302 580
rect 1242 506 1302 546
rect 1242 472 1255 506
rect 1289 472 1302 506
rect 1242 424 1302 472
rect 1242 390 1255 424
rect 1289 390 1302 424
rect 1242 368 1302 390
rect 1332 580 1412 592
rect 1332 546 1355 580
rect 1389 546 1412 580
rect 1332 492 1412 546
rect 1332 458 1355 492
rect 1389 458 1412 492
rect 1332 368 1412 458
rect 1442 580 1502 592
rect 1442 546 1455 580
rect 1489 546 1502 580
rect 1442 506 1502 546
rect 1442 472 1455 506
rect 1489 472 1502 506
rect 1442 424 1502 472
rect 1442 390 1455 424
rect 1489 390 1502 424
rect 1442 368 1502 390
rect 1532 580 1612 592
rect 1532 546 1555 580
rect 1589 546 1612 580
rect 1532 492 1612 546
rect 1532 458 1555 492
rect 1589 458 1612 492
rect 1532 368 1612 458
rect 1642 580 1701 592
rect 1642 546 1655 580
rect 1689 546 1701 580
rect 1642 497 1701 546
rect 1642 463 1655 497
rect 1689 463 1701 497
rect 1642 414 1701 463
rect 1642 380 1655 414
rect 1689 380 1701 414
rect 1642 368 1701 380
<< ndiffc >>
rect 39 118 73 152
rect 134 176 168 210
rect 218 176 252 210
rect 312 176 346 210
rect 134 86 168 120
rect 218 86 252 120
rect 312 86 346 120
rect 398 118 432 152
rect 498 176 532 210
rect 583 176 617 210
rect 682 176 716 210
rect 498 86 532 120
rect 583 86 617 120
rect 682 86 716 120
rect 768 118 802 152
rect 868 176 902 210
rect 868 86 902 120
rect 954 108 988 142
rect 1039 108 1073 142
rect 1118 108 1152 142
rect 1198 108 1232 142
rect 1277 108 1311 142
rect 1364 108 1398 142
rect 1450 176 1484 210
rect 1536 152 1570 186
rect 1450 86 1484 120
rect 1536 84 1570 118
rect 1622 168 1656 202
rect 1622 86 1656 120
<< pdiffc >>
rect 39 546 73 580
rect 39 474 73 508
rect 139 497 173 531
rect 139 406 173 440
rect 229 546 263 580
rect 229 474 263 508
rect 329 497 363 531
rect 329 406 363 440
rect 419 546 453 580
rect 419 463 453 497
rect 419 380 453 414
rect 509 546 543 580
rect 509 458 543 492
rect 599 497 633 531
rect 599 390 633 424
rect 689 546 723 580
rect 689 458 723 492
rect 779 497 813 531
rect 779 406 813 440
rect 891 497 925 531
rect 891 390 925 424
rect 981 546 1015 580
rect 981 460 1015 494
rect 1073 497 1107 531
rect 1073 390 1107 424
rect 1165 546 1199 580
rect 1165 460 1199 494
rect 1255 546 1289 580
rect 1255 472 1289 506
rect 1255 390 1289 424
rect 1355 546 1389 580
rect 1355 458 1389 492
rect 1455 546 1489 580
rect 1455 472 1489 506
rect 1455 390 1489 424
rect 1555 546 1589 580
rect 1555 458 1589 492
rect 1655 546 1689 580
rect 1655 463 1689 497
rect 1655 380 1689 414
<< poly >>
rect 96 592 126 618
rect 186 592 216 618
rect 276 592 306 618
rect 376 592 406 618
rect 466 592 496 618
rect 556 592 586 618
rect 646 592 676 618
rect 736 592 766 618
rect 938 592 968 618
rect 1028 592 1058 618
rect 1122 592 1152 618
rect 1212 592 1242 618
rect 1302 592 1332 618
rect 1412 592 1442 618
rect 1502 592 1532 618
rect 1612 592 1642 618
rect 96 353 126 368
rect 186 353 216 368
rect 276 353 306 368
rect 376 353 406 368
rect 466 353 496 368
rect 556 353 586 368
rect 646 353 676 368
rect 736 353 766 368
rect 938 353 968 368
rect 1028 353 1058 368
rect 1122 353 1152 368
rect 1212 353 1242 368
rect 1302 353 1332 368
rect 1412 353 1442 368
rect 1502 353 1532 368
rect 1612 353 1642 368
rect 93 336 129 353
rect 183 336 219 353
rect 273 336 309 353
rect 373 336 409 353
rect 463 336 499 353
rect 553 336 589 353
rect 643 336 679 353
rect 733 336 769 353
rect 935 336 971 353
rect 1025 336 1061 353
rect 1119 336 1155 353
rect 1209 336 1245 353
rect 93 320 409 336
rect 93 286 121 320
rect 155 286 189 320
rect 223 286 257 320
rect 291 286 325 320
rect 359 306 409 320
rect 457 320 769 336
rect 359 286 387 306
rect 93 270 387 286
rect 93 222 123 270
rect 357 222 387 270
rect 457 286 503 320
rect 537 286 571 320
rect 605 286 639 320
rect 673 286 707 320
rect 741 306 769 320
rect 827 320 1245 336
rect 741 286 757 306
rect 457 270 757 286
rect 457 222 487 270
rect 727 222 757 270
rect 827 286 843 320
rect 877 286 911 320
rect 945 286 979 320
rect 1013 286 1047 320
rect 1081 286 1115 320
rect 1149 286 1183 320
rect 1217 286 1245 320
rect 1299 326 1335 353
rect 1409 326 1445 353
rect 1499 326 1535 353
rect 1609 326 1645 353
rect 1299 310 1645 326
rect 1299 296 1425 310
rect 827 270 1245 286
rect 1409 276 1425 296
rect 1459 276 1493 310
rect 1527 276 1561 310
rect 1595 296 1645 310
rect 1595 276 1611 296
rect 827 222 857 270
rect 913 222 943 270
rect 1409 260 1611 276
rect 1409 222 1439 260
rect 1581 222 1611 260
rect 93 48 123 74
rect 357 48 387 74
rect 457 48 487 74
rect 727 48 757 74
rect 827 48 857 74
rect 913 48 943 74
rect 1409 48 1439 74
rect 1581 48 1611 74
<< polycont >>
rect 121 286 155 320
rect 189 286 223 320
rect 257 286 291 320
rect 325 286 359 320
rect 503 286 537 320
rect 571 286 605 320
rect 639 286 673 320
rect 707 286 741 320
rect 843 286 877 320
rect 911 286 945 320
rect 979 286 1013 320
rect 1047 286 1081 320
rect 1115 286 1149 320
rect 1183 286 1217 320
rect 1425 276 1459 310
rect 1493 276 1527 310
rect 1561 276 1595 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 23 581 453 615
rect 23 580 89 581
rect 23 546 39 580
rect 73 546 89 580
rect 229 580 279 581
rect 23 508 89 546
rect 23 474 39 508
rect 73 474 89 508
rect 23 458 89 474
rect 123 531 189 547
rect 123 497 139 531
rect 173 497 189 531
rect 123 440 189 497
rect 263 546 279 580
rect 419 580 453 581
rect 229 508 279 546
rect 263 474 279 508
rect 229 458 279 474
rect 313 531 379 547
rect 313 497 329 531
rect 363 497 379 531
rect 123 424 139 440
rect 25 406 139 424
rect 173 424 189 440
rect 313 440 379 497
rect 313 424 329 440
rect 173 406 329 424
rect 363 406 379 440
rect 25 390 379 406
rect 419 497 453 546
rect 419 424 453 463
rect 493 581 1215 615
rect 493 580 559 581
rect 493 546 509 580
rect 543 546 559 580
rect 673 580 739 581
rect 493 492 559 546
rect 493 458 509 492
rect 543 458 559 492
rect 594 531 638 547
rect 594 497 599 531
rect 633 497 638 531
rect 594 424 638 497
rect 673 546 689 580
rect 723 546 739 580
rect 965 580 1031 581
rect 673 492 739 546
rect 673 458 689 492
rect 723 458 739 492
rect 779 531 829 547
rect 813 497 829 531
rect 779 440 829 497
rect 419 414 599 424
rect 25 236 71 390
rect 453 390 599 414
rect 633 406 779 424
rect 813 406 829 440
rect 633 390 829 406
rect 875 531 925 547
rect 875 497 891 531
rect 875 424 925 497
rect 965 546 981 580
rect 1015 546 1031 580
rect 1149 580 1215 581
rect 965 494 1031 546
rect 965 460 981 494
rect 1015 460 1031 494
rect 1068 531 1112 547
rect 1068 497 1073 531
rect 1107 497 1112 531
rect 1068 424 1112 497
rect 1149 546 1165 580
rect 1199 546 1215 580
rect 1149 494 1215 546
rect 1149 460 1165 494
rect 1199 460 1215 494
rect 1251 580 1305 596
rect 1251 546 1255 580
rect 1289 546 1305 580
rect 1251 506 1305 546
rect 1251 472 1255 506
rect 1289 472 1305 506
rect 1251 424 1305 472
rect 1339 580 1405 649
rect 1339 546 1355 580
rect 1389 546 1405 580
rect 1339 492 1405 546
rect 1339 458 1355 492
rect 1389 458 1405 492
rect 1439 580 1505 596
rect 1439 546 1455 580
rect 1489 546 1505 580
rect 1439 506 1505 546
rect 1439 472 1455 506
rect 1489 472 1505 506
rect 1439 424 1505 472
rect 1539 580 1605 649
rect 1539 546 1555 580
rect 1589 546 1605 580
rect 1539 492 1605 546
rect 1539 458 1555 492
rect 1589 458 1605 492
rect 1639 580 1705 596
rect 1639 546 1655 580
rect 1689 546 1705 580
rect 1639 497 1705 546
rect 1639 463 1655 497
rect 1689 463 1705 497
rect 1639 424 1705 463
rect 875 390 891 424
rect 925 390 1073 424
rect 1107 390 1255 424
rect 1289 390 1455 424
rect 1489 414 1705 424
rect 1489 390 1655 414
rect 419 364 453 380
rect 1639 380 1655 390
rect 1689 380 1705 414
rect 1639 364 1705 380
rect 105 320 375 356
rect 105 286 121 320
rect 155 286 189 320
rect 223 286 257 320
rect 291 286 325 320
rect 359 286 375 320
rect 105 270 375 286
rect 487 320 757 356
rect 487 286 503 320
rect 537 286 571 320
rect 605 286 639 320
rect 673 286 707 320
rect 741 286 757 320
rect 487 270 757 286
rect 793 320 1319 356
rect 793 286 843 320
rect 877 286 911 320
rect 945 286 979 320
rect 1013 286 1047 320
rect 1081 286 1115 320
rect 1149 286 1183 320
rect 1217 286 1319 320
rect 793 270 1319 286
rect 1409 310 1703 326
rect 1409 276 1425 310
rect 1459 276 1493 310
rect 1527 276 1561 310
rect 1595 276 1703 310
rect 1409 260 1703 276
rect 1561 236 1703 260
rect 25 226 918 236
rect 25 210 1514 226
rect 25 202 134 210
rect 123 176 134 202
rect 168 176 218 210
rect 252 176 312 210
rect 346 202 498 210
rect 346 176 348 202
rect 23 152 89 168
rect 23 118 39 152
rect 73 118 89 152
rect 23 17 89 118
rect 123 120 348 176
rect 482 176 498 202
rect 532 176 583 210
rect 617 176 682 210
rect 716 202 868 210
rect 716 176 718 202
rect 123 86 134 120
rect 168 86 218 120
rect 252 86 312 120
rect 346 86 348 120
rect 123 70 348 86
rect 382 152 448 168
rect 382 118 398 152
rect 432 118 448 152
rect 382 17 448 118
rect 482 120 718 176
rect 852 176 868 202
rect 902 192 1450 210
rect 902 176 918 192
rect 482 86 498 120
rect 532 86 583 120
rect 617 86 682 120
rect 716 86 718 120
rect 482 70 718 86
rect 752 152 818 168
rect 752 118 768 152
rect 802 118 818 152
rect 752 17 818 118
rect 852 120 918 176
rect 1448 176 1450 192
rect 1484 202 1514 210
rect 1484 186 1572 202
rect 1484 176 1536 186
rect 852 86 868 120
rect 902 86 918 120
rect 852 70 918 86
rect 952 142 1414 158
rect 952 108 954 142
rect 988 108 1039 142
rect 1073 108 1118 142
rect 1152 108 1198 142
rect 1232 108 1277 142
rect 1311 108 1364 142
rect 1398 108 1414 142
rect 952 17 1414 108
rect 1448 152 1536 176
rect 1570 152 1572 186
rect 1448 120 1572 152
rect 1448 86 1450 120
rect 1484 118 1572 120
rect 1484 86 1536 118
rect 1448 84 1536 86
rect 1570 84 1572 118
rect 1448 68 1572 84
rect 1606 168 1622 202
rect 1656 168 1672 202
rect 1606 120 1672 168
rect 1606 86 1622 120
rect 1656 86 1672 120
rect 1606 17 1672 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
<< metal1 >>
rect 0 683 1728 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 0 617 1728 649
rect 0 17 1728 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
rect 0 -49 1728 -17
<< labels >>
rlabel comment s 0 0 0 0 4 nor4_4
flabel pwell s 0 0 1728 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 1728 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 1728 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 1728 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 1567 242 1601 276 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 1663 242 1697 276 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 1087 316 1121 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 1183 316 1217 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 1279 316 1313 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 4 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 D
port 4 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 D
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 1728 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2000124
string GDS_START 1986126
<< end >>
