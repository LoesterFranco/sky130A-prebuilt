magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 2116 561
rect 103 427 169 527
rect 18 195 88 325
rect 291 427 357 527
rect 686 451 762 527
rect 103 17 169 93
rect 354 201 436 325
rect 866 451 932 527
rect 1186 451 1268 527
rect 291 17 357 93
rect 722 147 804 213
rect 1402 389 1468 527
rect 722 17 804 105
rect 948 17 1016 109
rect 1332 201 1398 213
rect 1332 147 1464 201
rect 1604 296 1640 527
rect 1334 17 1466 113
rect 1604 17 1640 181
rect 1674 51 1740 493
rect 1889 365 1923 527
rect 1973 289 2025 493
rect 1982 165 2025 289
rect 1889 17 1923 117
rect 1973 51 2025 165
rect 0 -17 2116 17
<< obsli1 >>
rect 35 393 69 493
rect 35 391 168 393
rect 35 359 129 391
rect 122 357 129 359
rect 163 357 168 391
rect 122 161 168 357
rect 35 127 168 161
rect 203 187 248 493
rect 391 393 425 493
rect 472 450 638 484
rect 203 153 213 187
rect 247 153 248 187
rect 35 69 69 127
rect 203 69 248 153
rect 286 359 425 393
rect 286 165 320 359
rect 470 357 489 391
rect 523 357 570 391
rect 470 315 570 357
rect 286 127 425 165
rect 470 141 514 315
rect 604 281 638 450
rect 798 417 832 475
rect 1022 433 1152 483
rect 1118 417 1152 433
rect 1308 417 1356 475
rect 672 367 942 417
rect 672 315 722 367
rect 824 281 874 313
rect 604 247 874 281
rect 604 239 688 247
rect 550 187 620 203
rect 550 153 581 187
rect 615 153 620 187
rect 550 129 620 153
rect 391 61 425 127
rect 654 93 688 239
rect 908 213 942 367
rect 862 145 942 213
rect 980 391 1080 393
rect 980 357 1041 391
rect 1075 357 1080 391
rect 980 331 1080 357
rect 1118 383 1356 417
rect 980 179 1014 331
rect 1048 255 1084 295
rect 1048 221 1049 255
rect 1083 221 1084 255
rect 1118 281 1152 383
rect 1502 353 1536 475
rect 1502 349 1566 353
rect 1186 315 1566 349
rect 1118 247 1494 281
rect 1048 213 1084 221
rect 1164 179 1230 203
rect 980 145 1230 179
rect 485 53 688 93
rect 862 59 912 145
rect 1264 95 1298 247
rect 1428 235 1494 247
rect 1528 136 1566 315
rect 1128 61 1298 95
rect 1502 70 1566 136
rect 1778 265 1844 493
rect 1778 199 1948 265
rect 1778 51 1844 199
<< obsli1c >>
rect 129 357 163 391
rect 213 153 247 187
rect 489 357 523 391
rect 581 153 615 187
rect 1041 357 1075 391
rect 1049 221 1083 255
<< metal1 >>
rect 0 496 2116 592
rect 753 184 811 193
rect 1397 184 1455 193
rect 753 156 1455 184
rect 753 147 811 156
rect 1397 147 1455 156
rect 0 -48 2116 48
<< obsm1 >>
rect 117 391 175 397
rect 117 357 129 391
rect 163 388 175 391
rect 477 391 535 397
rect 477 388 489 391
rect 163 360 489 388
rect 163 357 175 360
rect 117 351 175 357
rect 477 357 489 360
rect 523 388 535 391
rect 1029 391 1087 397
rect 1029 388 1041 391
rect 523 360 1041 388
rect 523 357 535 360
rect 477 351 535 357
rect 1029 357 1041 360
rect 1075 357 1087 391
rect 1029 351 1087 357
rect 1037 255 1095 261
rect 1037 252 1049 255
rect 584 224 1049 252
rect 584 193 627 224
rect 1037 221 1049 224
rect 1083 221 1095 255
rect 1037 215 1095 221
rect 201 187 259 193
rect 201 153 213 187
rect 247 184 259 187
rect 569 187 627 193
rect 569 184 581 187
rect 247 156 581 184
rect 247 153 259 156
rect 201 147 259 153
rect 569 153 581 156
rect 615 153 627 187
rect 569 147 627 153
<< labels >>
rlabel locali s 354 201 436 325 6 D
port 1 nsew signal input
rlabel locali s 1982 165 2025 289 6 Q
port 2 nsew signal output
rlabel locali s 1973 289 2025 493 6 Q
port 2 nsew signal output
rlabel locali s 1973 51 2025 165 6 Q
port 2 nsew signal output
rlabel locali s 1674 51 1740 493 6 Q_N
port 3 nsew signal output
rlabel locali s 722 147 804 213 6 SET_B
port 4 nsew signal input
rlabel locali s 1332 201 1398 213 6 SET_B
port 4 nsew signal input
rlabel locali s 1332 147 1464 201 6 SET_B
port 4 nsew signal input
rlabel metal1 s 1397 184 1455 193 6 SET_B
port 4 nsew signal input
rlabel metal1 s 1397 147 1455 156 6 SET_B
port 4 nsew signal input
rlabel metal1 s 753 184 811 193 6 SET_B
port 4 nsew signal input
rlabel metal1 s 753 156 1455 184 6 SET_B
port 4 nsew signal input
rlabel metal1 s 753 147 811 156 6 SET_B
port 4 nsew signal input
rlabel locali s 18 195 88 325 6 CLK
port 5 nsew clock input
rlabel locali s 1889 17 1923 117 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1604 17 1640 181 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1334 17 1466 113 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 948 17 1016 109 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 722 17 804 105 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 291 17 357 93 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 103 17 169 93 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 2116 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 2116 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1889 365 1923 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1604 296 1640 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1402 389 1468 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1186 451 1268 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 866 451 932 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 686 451 762 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 291 427 357 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 103 427 169 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 2116 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 2116 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2116 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3436490
string GDS_START 3418724
<< end >>
