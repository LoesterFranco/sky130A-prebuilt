magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 406 582
<< pwell >>
rect 29 -17 63 17
<< ndiode >>
rect 31 159 337 177
rect 31 125 40 159
rect 74 125 115 159
rect 149 125 219 159
rect 253 125 294 159
rect 328 125 337 159
rect 31 91 337 125
rect 31 57 40 91
rect 74 57 115 91
rect 149 57 219 91
rect 253 57 294 91
rect 328 57 337 91
rect 31 39 337 57
<< ndiodec >>
rect 40 125 74 159
rect 115 125 149 159
rect 219 125 253 159
rect 294 125 328 159
rect 40 57 74 91
rect 115 57 149 91
rect 219 57 253 91
rect 294 57 328 91
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 17 159 351 493
rect 17 125 40 159
rect 74 125 115 159
rect 149 125 219 159
rect 253 125 294 159
rect 328 125 351 159
rect 17 91 351 125
rect 17 57 40 91
rect 74 57 115 91
rect 149 57 219 91
rect 253 57 294 91
rect 328 57 351 91
rect 17 51 351 57
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
<< metal1 >>
rect 0 561 368 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 0 496 368 527
rect 0 17 368 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
rect 0 -48 368 -17
<< labels >>
flabel corelocali s 121 85 155 119 0 FreeSans 200 0 0 0 DIODE
port 1 nsew
flabel corelocali s 121 357 155 391 0 FreeSans 200 0 0 0 DIODE
port 1 nsew
flabel corelocali s 29 357 63 391 0 FreeSans 200 0 0 0 DIODE
port 1 nsew
flabel corelocali s 121 425 155 459 0 FreeSans 200 0 0 0 DIODE
port 1 nsew
flabel corelocali s 29 425 63 459 0 FreeSans 200 0 0 0 DIODE
port 1 nsew
flabel corelocali s 29 289 63 323 0 FreeSans 200 0 0 0 DIODE
port 1 nsew
flabel corelocali s 121 289 155 323 0 FreeSans 200 0 0 0 DIODE
port 1 nsew
flabel corelocali s 29 221 63 255 0 FreeSans 200 0 0 0 DIODE
port 1 nsew
flabel corelocali s 121 221 155 255 0 FreeSans 200 0 0 0 DIODE
port 1 nsew
flabel corelocali s 121 153 155 187 0 FreeSans 200 0 0 0 DIODE
port 1 nsew
flabel corelocali s 29 153 63 187 0 FreeSans 200 0 0 0 DIODE
port 1 nsew
flabel corelocali s 29 85 63 119 0 FreeSans 200 0 0 0 DIODE
port 1 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew
rlabel comment s 0 0 0 0 4 diode_4
<< properties >>
string FIXED_BBOX 0 0 368 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3598584
string GDS_START 3594578
<< end >>
