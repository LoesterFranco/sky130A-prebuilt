magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 18 299 85 493
rect 214 459 683 493
rect 18 51 69 299
rect 214 265 254 459
rect 199 199 254 265
rect 356 323 615 357
rect 356 162 390 323
rect 458 51 523 283
rect 557 51 615 323
rect 649 326 683 459
rect 649 288 799 326
rect 761 211 799 288
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 129 299 163 527
rect 103 165 137 265
rect 288 391 577 425
rect 288 165 322 391
rect 103 131 322 165
rect 287 124 322 131
rect 103 17 179 97
rect 287 51 391 124
rect 717 367 763 527
rect 797 367 877 493
rect 665 173 699 237
rect 843 173 877 367
rect 665 139 877 173
rect 650 17 753 105
rect 807 51 856 139
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
rlabel locali s 458 51 523 283 6 A0
port 1 nsew signal input
rlabel locali s 557 51 615 323 6 A1
port 2 nsew signal input
rlabel locali s 356 323 615 357 6 A1
port 2 nsew signal input
rlabel locali s 356 162 390 323 6 A1
port 2 nsew signal input
rlabel locali s 761 211 799 288 6 S
port 3 nsew signal input
rlabel locali s 649 326 683 459 6 S
port 3 nsew signal input
rlabel locali s 649 288 799 326 6 S
port 3 nsew signal input
rlabel locali s 214 459 683 493 6 S
port 3 nsew signal input
rlabel locali s 214 265 254 459 6 S
port 3 nsew signal input
rlabel locali s 199 199 254 265 6 S
port 3 nsew signal input
rlabel locali s 18 299 85 493 6 X
port 4 nsew signal output
rlabel locali s 18 51 69 299 6 X
port 4 nsew signal output
rlabel metal1 s 0 -48 920 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 920 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 920 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3276240
string GDS_START 3269040
<< end >>
