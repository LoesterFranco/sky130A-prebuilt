magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 2630 704
rect 1101 311 1309 332
<< pwell >>
rect 0 0 2592 49
<< scnmos >>
rect 84 74 114 158
rect 282 74 312 222
rect 368 74 398 222
rect 582 74 612 158
rect 702 74 732 158
rect 780 74 810 158
rect 1005 118 1035 202
rect 1083 118 1113 202
rect 1195 74 1225 202
rect 1304 74 1334 202
rect 1406 88 1436 172
rect 1484 88 1514 172
rect 1562 88 1592 172
rect 1799 88 1829 172
rect 2011 74 2041 222
rect 2111 74 2141 222
rect 2197 74 2227 222
rect 2369 74 2399 222
rect 2464 74 2494 222
<< pmoshvt >>
rect 86 504 116 588
rect 288 368 318 592
rect 378 368 408 592
rect 586 463 616 547
rect 686 463 716 547
rect 770 463 800 547
rect 957 463 987 547
rect 1047 463 1077 547
rect 1190 347 1220 547
rect 1291 392 1321 592
rect 1450 508 1480 592
rect 1534 508 1564 592
rect 1624 508 1654 592
rect 1819 508 1849 592
rect 2014 368 2044 536
rect 2104 368 2134 536
rect 2208 368 2238 592
rect 2298 368 2328 592
rect 2388 368 2418 592
rect 2478 368 2508 592
<< ndiff >>
rect 225 195 282 222
rect 225 161 237 195
rect 271 161 282 195
rect 27 133 84 158
rect 27 99 39 133
rect 73 99 84 133
rect 27 74 84 99
rect 114 133 171 158
rect 114 99 125 133
rect 159 99 171 133
rect 114 74 171 99
rect 225 120 282 161
rect 225 86 237 120
rect 271 86 282 120
rect 225 74 282 86
rect 312 186 368 222
rect 312 152 323 186
rect 357 152 368 186
rect 312 116 368 152
rect 312 82 323 116
rect 357 82 368 116
rect 312 74 368 82
rect 398 210 455 222
rect 398 176 409 210
rect 443 176 455 210
rect 398 120 455 176
rect 398 86 409 120
rect 443 86 455 120
rect 398 74 455 86
rect 509 169 567 181
rect 509 135 521 169
rect 555 158 567 169
rect 934 174 1005 202
rect 555 135 582 158
rect 509 74 582 135
rect 612 133 702 158
rect 612 99 657 133
rect 691 99 702 133
rect 612 74 702 99
rect 732 74 780 158
rect 810 120 880 158
rect 810 86 827 120
rect 861 86 880 120
rect 934 140 953 174
rect 987 140 1005 174
rect 934 118 1005 140
rect 1035 118 1083 202
rect 1113 190 1195 202
rect 1113 156 1150 190
rect 1184 156 1195 190
rect 1113 120 1195 156
rect 1113 118 1150 120
rect 810 74 880 86
rect 1138 86 1150 118
rect 1184 86 1195 120
rect 1138 74 1195 86
rect 1225 74 1304 202
rect 1334 172 1391 202
rect 1940 210 2011 222
rect 1940 176 1952 210
rect 1986 176 2011 210
rect 1334 169 1406 172
rect 1334 135 1345 169
rect 1379 135 1406 169
rect 1334 88 1406 135
rect 1436 88 1484 172
rect 1514 88 1562 172
rect 1592 134 1799 172
rect 1592 100 1603 134
rect 1637 100 1671 134
rect 1705 100 1740 134
rect 1774 100 1799 134
rect 1592 88 1799 100
rect 1829 147 1886 172
rect 1829 113 1840 147
rect 1874 113 1886 147
rect 1829 88 1886 113
rect 1940 120 2011 176
rect 1334 74 1384 88
rect 1940 86 1952 120
rect 1986 86 2011 120
rect 1940 74 2011 86
rect 2041 210 2111 222
rect 2041 176 2052 210
rect 2086 176 2111 210
rect 2041 120 2111 176
rect 2041 86 2052 120
rect 2086 86 2111 120
rect 2041 74 2111 86
rect 2141 210 2197 222
rect 2141 176 2152 210
rect 2186 176 2197 210
rect 2141 120 2197 176
rect 2141 86 2152 120
rect 2186 86 2197 120
rect 2141 74 2197 86
rect 2227 144 2369 222
rect 2227 110 2238 144
rect 2272 110 2324 144
rect 2358 110 2369 144
rect 2227 74 2369 110
rect 2399 210 2464 222
rect 2399 176 2419 210
rect 2453 176 2464 210
rect 2399 120 2464 176
rect 2399 86 2419 120
rect 2453 86 2464 120
rect 2399 74 2464 86
rect 2494 146 2565 222
rect 2494 112 2519 146
rect 2553 112 2565 146
rect 2494 74 2565 112
<< pdiff >>
rect 27 563 86 588
rect 27 529 39 563
rect 73 529 86 563
rect 27 504 86 529
rect 116 563 175 588
rect 116 529 129 563
rect 163 529 175 563
rect 116 504 175 529
rect 229 414 288 592
rect 229 380 241 414
rect 275 380 288 414
rect 229 368 288 380
rect 318 565 378 592
rect 318 531 331 565
rect 365 531 378 565
rect 318 368 378 531
rect 408 532 467 592
rect 408 498 421 532
rect 455 498 467 532
rect 408 368 467 498
rect 1238 547 1291 592
rect 527 520 586 547
rect 527 486 539 520
rect 573 486 586 520
rect 527 463 586 486
rect 616 520 686 547
rect 616 486 639 520
rect 673 486 686 520
rect 616 463 686 486
rect 716 463 770 547
rect 800 535 957 547
rect 800 501 816 535
rect 850 501 957 535
rect 800 463 957 501
rect 987 520 1047 547
rect 987 486 1000 520
rect 1034 486 1047 520
rect 987 463 1047 486
rect 1077 537 1190 547
rect 1077 503 1137 537
rect 1171 503 1190 537
rect 1077 463 1190 503
rect 1137 347 1190 463
rect 1220 392 1291 547
rect 1321 580 1450 592
rect 1321 546 1334 580
rect 1368 546 1403 580
rect 1437 546 1450 580
rect 1321 512 1450 546
rect 1321 478 1334 512
rect 1368 508 1450 512
rect 1480 508 1534 592
rect 1564 580 1624 592
rect 1564 546 1577 580
rect 1611 546 1624 580
rect 1564 508 1624 546
rect 1654 567 1709 592
rect 1654 533 1667 567
rect 1701 533 1709 567
rect 1654 508 1709 533
rect 1763 580 1819 592
rect 1763 546 1772 580
rect 1806 546 1819 580
rect 1763 508 1819 546
rect 1849 580 1904 592
rect 1849 546 1862 580
rect 1896 546 1904 580
rect 2152 580 2208 592
rect 1849 508 1904 546
rect 2152 546 2161 580
rect 2195 546 2208 580
rect 2152 536 2208 546
rect 1958 524 2014 536
rect 1368 478 1377 508
rect 1321 444 1377 478
rect 1321 410 1334 444
rect 1368 410 1377 444
rect 1321 392 1377 410
rect 1220 347 1273 392
rect 1958 490 1967 524
rect 2001 490 2014 524
rect 1958 414 2014 490
rect 1958 380 1967 414
rect 2001 380 2014 414
rect 1958 368 2014 380
rect 2044 524 2104 536
rect 2044 490 2057 524
rect 2091 490 2104 524
rect 2044 414 2104 490
rect 2044 380 2057 414
rect 2091 380 2104 414
rect 2044 368 2104 380
rect 2134 494 2208 536
rect 2134 460 2161 494
rect 2195 460 2208 494
rect 2134 414 2208 460
rect 2134 380 2161 414
rect 2195 380 2208 414
rect 2134 368 2208 380
rect 2238 580 2298 592
rect 2238 546 2251 580
rect 2285 546 2298 580
rect 2238 494 2298 546
rect 2238 460 2251 494
rect 2285 460 2298 494
rect 2238 414 2298 460
rect 2238 380 2251 414
rect 2285 380 2298 414
rect 2238 368 2298 380
rect 2328 580 2388 592
rect 2328 546 2341 580
rect 2375 546 2388 580
rect 2328 484 2388 546
rect 2328 450 2341 484
rect 2375 450 2388 484
rect 2328 368 2388 450
rect 2418 580 2478 592
rect 2418 546 2431 580
rect 2465 546 2478 580
rect 2418 494 2478 546
rect 2418 460 2431 494
rect 2465 460 2478 494
rect 2418 414 2478 460
rect 2418 380 2431 414
rect 2465 380 2478 414
rect 2418 368 2478 380
rect 2508 580 2565 592
rect 2508 546 2521 580
rect 2555 546 2565 580
rect 2508 498 2565 546
rect 2508 464 2521 498
rect 2555 464 2565 498
rect 2508 368 2565 464
<< ndiffc >>
rect 237 161 271 195
rect 39 99 73 133
rect 125 99 159 133
rect 237 86 271 120
rect 323 152 357 186
rect 323 82 357 116
rect 409 176 443 210
rect 409 86 443 120
rect 521 135 555 169
rect 657 99 691 133
rect 827 86 861 120
rect 953 140 987 174
rect 1150 156 1184 190
rect 1150 86 1184 120
rect 1952 176 1986 210
rect 1345 135 1379 169
rect 1603 100 1637 134
rect 1671 100 1705 134
rect 1740 100 1774 134
rect 1840 113 1874 147
rect 1952 86 1986 120
rect 2052 176 2086 210
rect 2052 86 2086 120
rect 2152 176 2186 210
rect 2152 86 2186 120
rect 2238 110 2272 144
rect 2324 110 2358 144
rect 2419 176 2453 210
rect 2419 86 2453 120
rect 2519 112 2553 146
<< pdiffc >>
rect 39 529 73 563
rect 129 529 163 563
rect 241 380 275 414
rect 331 531 365 565
rect 421 498 455 532
rect 539 486 573 520
rect 639 486 673 520
rect 816 501 850 535
rect 1000 486 1034 520
rect 1137 503 1171 537
rect 1334 546 1368 580
rect 1403 546 1437 580
rect 1334 478 1368 512
rect 1577 546 1611 580
rect 1667 533 1701 567
rect 1772 546 1806 580
rect 1862 546 1896 580
rect 2161 546 2195 580
rect 1334 410 1368 444
rect 1967 490 2001 524
rect 1967 380 2001 414
rect 2057 490 2091 524
rect 2057 380 2091 414
rect 2161 460 2195 494
rect 2161 380 2195 414
rect 2251 546 2285 580
rect 2251 460 2285 494
rect 2251 380 2285 414
rect 2341 546 2375 580
rect 2341 450 2375 484
rect 2431 546 2465 580
rect 2431 460 2465 494
rect 2431 380 2465 414
rect 2521 546 2555 580
rect 2521 464 2555 498
<< poly >>
rect 86 588 116 614
rect 288 592 318 618
rect 378 592 408 618
rect 482 615 1324 645
rect 86 489 116 504
rect 83 398 119 489
rect 83 382 161 398
rect 83 348 111 382
rect 145 348 161 382
rect 288 353 318 368
rect 378 353 408 368
rect 83 314 161 348
rect 83 280 111 314
rect 145 280 161 314
rect 285 310 321 353
rect 375 336 411 353
rect 482 336 512 615
rect 586 547 616 573
rect 683 562 719 615
rect 1288 607 1324 615
rect 1291 592 1321 607
rect 1450 592 1480 618
rect 1534 592 1564 618
rect 1624 592 1654 618
rect 1819 592 1849 618
rect 2208 592 2238 618
rect 2298 592 2328 618
rect 2388 592 2418 618
rect 2478 592 2508 618
rect 686 547 716 562
rect 770 547 800 573
rect 957 547 987 573
rect 1047 547 1077 573
rect 1190 547 1220 573
rect 586 448 616 463
rect 583 425 619 448
rect 686 437 716 463
rect 770 448 800 463
rect 957 448 987 463
rect 1047 448 1077 463
rect 767 432 803 448
rect 368 320 512 336
rect 83 246 161 280
rect 83 212 111 246
rect 145 212 161 246
rect 260 294 326 310
rect 260 260 276 294
rect 310 260 326 294
rect 260 244 326 260
rect 368 286 405 320
rect 439 286 512 320
rect 557 409 623 425
rect 557 375 573 409
rect 607 375 623 409
rect 767 402 889 432
rect 557 360 623 375
rect 823 390 889 402
rect 557 344 775 360
rect 557 341 725 344
rect 557 307 573 341
rect 607 310 725 341
rect 759 310 775 344
rect 823 356 839 390
rect 873 356 889 390
rect 823 340 889 356
rect 607 307 775 310
rect 557 294 775 307
rect 557 291 623 294
rect 368 270 512 286
rect 282 222 312 244
rect 368 222 398 270
rect 482 243 512 270
rect 83 196 161 212
rect 84 158 114 196
rect 482 213 612 243
rect 582 158 612 213
rect 702 158 732 294
rect 846 246 876 340
rect 954 290 990 448
rect 1044 398 1080 448
rect 1039 382 1113 398
rect 1039 348 1055 382
rect 1089 348 1113 382
rect 1039 332 1113 348
rect 2014 536 2044 562
rect 2104 536 2134 562
rect 1450 493 1480 508
rect 1534 493 1564 508
rect 1624 493 1654 508
rect 1819 493 1849 508
rect 1447 470 1483 493
rect 1409 454 1483 470
rect 1409 420 1425 454
rect 1459 420 1483 454
rect 1409 404 1483 420
rect 1291 377 1321 392
rect 1288 362 1324 377
rect 1190 332 1220 347
rect 1288 332 1436 362
rect 954 274 1035 290
rect 846 230 912 246
rect 846 210 862 230
rect 780 196 862 210
rect 896 196 912 230
rect 954 240 970 274
rect 1004 240 1035 274
rect 954 224 1035 240
rect 1005 202 1035 224
rect 1083 202 1113 332
rect 1187 306 1223 332
rect 1161 290 1227 306
rect 1161 256 1177 290
rect 1211 256 1227 290
rect 1161 240 1227 256
rect 1273 274 1339 290
rect 1273 240 1289 274
rect 1323 240 1339 274
rect 1195 202 1225 240
rect 1273 224 1339 240
rect 1304 202 1334 224
rect 780 180 912 196
rect 780 158 810 180
rect 1005 92 1035 118
rect 1083 92 1113 118
rect 1406 172 1436 332
rect 1531 331 1567 493
rect 1621 370 1657 493
rect 1816 476 1852 493
rect 1756 460 1852 476
rect 1756 426 1772 460
rect 1806 426 1852 460
rect 1756 392 1852 426
rect 1621 354 1703 370
rect 1484 315 1575 331
rect 1484 281 1525 315
rect 1559 281 1575 315
rect 1484 265 1575 281
rect 1621 320 1653 354
rect 1687 320 1703 354
rect 1621 286 1703 320
rect 1484 172 1514 265
rect 1621 252 1653 286
rect 1687 252 1703 286
rect 1756 358 1772 392
rect 1806 358 1852 392
rect 1756 324 1852 358
rect 2014 353 2044 368
rect 2104 353 2134 368
rect 2208 353 2238 368
rect 2298 353 2328 368
rect 2388 353 2418 368
rect 2478 353 2508 368
rect 1756 290 1772 324
rect 1806 323 1852 324
rect 2011 323 2137 353
rect 2205 330 2241 353
rect 2295 330 2331 353
rect 2385 330 2421 353
rect 2475 330 2511 353
rect 1806 290 2041 323
rect 1756 274 2041 290
rect 2197 314 2511 330
rect 2197 280 2213 314
rect 2247 280 2281 314
rect 2315 280 2349 314
rect 2383 300 2511 314
rect 2383 280 2494 300
rect 2197 275 2494 280
rect 1621 236 1703 252
rect 1621 217 1653 236
rect 1562 187 1653 217
rect 1562 172 1592 187
rect 1799 172 1829 274
rect 2011 222 2041 274
rect 2111 264 2494 275
rect 2111 245 2399 264
rect 2111 222 2141 245
rect 2197 222 2227 245
rect 2369 222 2399 245
rect 2464 222 2494 264
rect 84 48 114 74
rect 282 48 312 74
rect 368 48 398 74
rect 582 48 612 74
rect 702 48 732 74
rect 780 48 810 74
rect 1195 48 1225 74
rect 1304 48 1334 74
rect 1406 62 1436 88
rect 1484 62 1514 88
rect 1562 62 1592 88
rect 1799 62 1829 88
rect 2011 48 2041 74
rect 2111 48 2141 74
rect 2197 48 2227 74
rect 2369 48 2399 74
rect 2464 48 2494 74
<< polycont >>
rect 111 348 145 382
rect 111 280 145 314
rect 111 212 145 246
rect 276 260 310 294
rect 405 286 439 320
rect 573 375 607 409
rect 573 307 607 341
rect 725 310 759 344
rect 839 356 873 390
rect 1055 348 1089 382
rect 1425 420 1459 454
rect 862 196 896 230
rect 970 240 1004 274
rect 1177 256 1211 290
rect 1289 240 1323 274
rect 1772 426 1806 460
rect 1525 281 1559 315
rect 1653 320 1687 354
rect 1653 252 1687 286
rect 1772 358 1806 392
rect 1772 290 1806 324
rect 2213 280 2247 314
rect 2281 280 2315 314
rect 2349 280 2383 314
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2592 683
rect 23 563 73 592
rect 23 529 39 563
rect 23 482 73 529
rect 113 563 179 649
rect 113 529 129 563
rect 163 529 179 563
rect 113 516 179 529
rect 315 565 381 649
rect 315 531 331 565
rect 365 531 381 565
rect 315 516 381 531
rect 421 581 759 615
rect 421 532 455 581
rect 421 482 455 498
rect 489 520 589 547
rect 489 486 539 520
rect 573 486 589 520
rect 23 448 359 482
rect 489 459 589 486
rect 623 520 691 547
rect 623 486 639 520
rect 673 486 691 520
rect 623 459 691 486
rect 489 448 523 459
rect 23 162 57 448
rect 325 414 523 448
rect 95 382 161 398
rect 95 348 111 382
rect 145 348 161 382
rect 95 314 161 348
rect 95 280 111 314
rect 145 280 161 314
rect 95 246 161 280
rect 95 212 111 246
rect 145 212 161 246
rect 95 196 161 212
rect 195 380 241 414
rect 275 380 291 414
rect 195 378 291 380
rect 195 344 455 378
rect 195 202 229 344
rect 389 320 455 344
rect 263 294 355 310
rect 263 260 276 294
rect 310 260 355 294
rect 389 286 405 320
rect 439 286 455 320
rect 389 270 455 286
rect 263 236 355 260
rect 409 210 443 226
rect 195 195 287 202
rect 23 133 73 162
rect 23 99 39 133
rect 23 70 73 99
rect 109 133 159 162
rect 109 99 125 133
rect 109 17 159 99
rect 195 161 237 195
rect 271 161 287 195
rect 195 120 287 161
rect 195 86 237 120
rect 271 86 287 120
rect 195 68 287 86
rect 323 186 373 202
rect 357 152 373 186
rect 323 116 373 152
rect 357 82 373 116
rect 323 17 373 82
rect 409 120 443 176
rect 489 185 523 414
rect 557 409 623 425
rect 557 375 573 409
rect 607 375 623 409
rect 557 341 623 375
rect 557 307 573 341
rect 607 307 623 341
rect 557 291 623 307
rect 489 169 555 185
rect 489 135 521 169
rect 489 119 555 135
rect 409 85 443 86
rect 589 85 623 291
rect 409 51 623 85
rect 657 260 691 459
rect 725 467 759 581
rect 797 551 831 649
rect 903 581 1102 615
rect 797 535 869 551
rect 797 501 816 535
rect 850 501 869 535
rect 903 467 937 581
rect 725 433 937 467
rect 971 520 1034 547
rect 971 486 1000 520
rect 971 459 1034 486
rect 725 344 759 433
rect 971 399 1005 459
rect 1068 453 1102 581
rect 1136 537 1188 649
rect 1136 503 1137 537
rect 1171 503 1188 537
rect 1318 580 1453 596
rect 1318 546 1334 580
rect 1368 546 1403 580
rect 1437 546 1453 580
rect 1318 530 1453 546
rect 1577 580 1611 649
rect 1577 530 1611 546
rect 1651 567 1717 596
rect 1651 533 1667 567
rect 1701 533 1717 567
rect 1136 487 1188 503
rect 1334 512 1543 530
rect 1368 496 1543 512
rect 1651 496 1717 533
rect 1756 580 1806 649
rect 1756 546 1772 580
rect 1756 530 1806 546
rect 1846 580 1912 596
rect 1846 546 1862 580
rect 1896 546 1912 580
rect 1846 530 1912 546
rect 1068 419 1295 453
rect 823 390 1005 399
rect 823 356 839 390
rect 873 356 1005 390
rect 823 348 1005 356
rect 1039 382 1127 385
rect 1039 348 1055 382
rect 1089 350 1127 382
rect 1039 316 1087 348
rect 1121 316 1127 350
rect 725 294 759 310
rect 793 280 1005 314
rect 1039 310 1127 316
rect 793 260 827 280
rect 657 226 827 260
rect 954 274 1005 280
rect 1161 290 1227 298
rect 1161 274 1177 290
rect 861 230 918 246
rect 657 133 707 226
rect 861 196 862 230
rect 896 196 918 230
rect 954 240 970 274
rect 1004 256 1177 274
rect 1211 256 1227 290
rect 1004 240 1227 256
rect 1261 290 1295 419
rect 1334 444 1368 478
rect 1509 462 1822 496
rect 1334 358 1368 410
rect 1409 454 1475 462
rect 1409 420 1425 454
rect 1459 420 1475 454
rect 1409 404 1475 420
rect 1334 324 1407 358
rect 1261 274 1339 290
rect 1261 240 1289 274
rect 1323 240 1339 274
rect 954 224 1005 240
rect 1261 224 1339 240
rect 861 190 918 196
rect 1134 190 1200 206
rect 861 174 1010 190
rect 861 156 953 174
rect 691 99 707 133
rect 918 140 953 156
rect 987 140 1010 174
rect 918 124 1010 140
rect 1134 156 1150 190
rect 1184 156 1200 190
rect 1134 120 1200 156
rect 657 70 707 99
rect 805 86 827 120
rect 861 86 884 120
rect 805 17 884 86
rect 1134 86 1150 120
rect 1184 86 1200 120
rect 1134 17 1200 86
rect 1261 85 1295 224
rect 1373 185 1407 324
rect 1329 169 1407 185
rect 1329 135 1345 169
rect 1379 135 1407 169
rect 1329 119 1407 135
rect 1441 85 1475 404
rect 1756 460 1822 462
rect 1756 426 1772 460
rect 1806 426 1822 460
rect 1756 392 1822 426
rect 1637 354 1703 370
rect 1509 315 1575 331
rect 1509 281 1525 315
rect 1559 281 1575 315
rect 1509 202 1575 281
rect 1637 320 1653 354
rect 1687 350 1703 354
rect 1637 316 1663 320
rect 1697 316 1703 350
rect 1637 286 1703 316
rect 1637 252 1653 286
rect 1687 252 1703 286
rect 1756 358 1772 392
rect 1806 358 1822 392
rect 1756 324 1822 358
rect 1756 290 1772 324
rect 1806 290 1822 324
rect 1756 274 1822 290
rect 1637 236 1703 252
rect 1856 202 1890 530
rect 1951 524 2001 649
rect 2145 580 2201 649
rect 2145 546 2161 580
rect 2195 546 2201 580
rect 1951 490 1967 524
rect 1951 414 2001 490
rect 1951 380 1967 414
rect 1951 364 2001 380
rect 2041 524 2107 540
rect 2041 490 2057 524
rect 2091 490 2107 524
rect 2041 414 2107 490
rect 2041 380 2057 414
rect 2091 380 2107 414
rect 2041 330 2107 380
rect 2145 494 2201 546
rect 2145 460 2161 494
rect 2195 460 2201 494
rect 2145 414 2201 460
rect 2145 380 2161 414
rect 2195 380 2201 414
rect 2145 364 2201 380
rect 2235 580 2291 596
rect 2235 546 2251 580
rect 2285 546 2291 580
rect 2235 494 2291 546
rect 2235 460 2251 494
rect 2285 460 2291 494
rect 2235 416 2291 460
rect 2325 580 2391 649
rect 2325 546 2341 580
rect 2375 546 2391 580
rect 2325 484 2391 546
rect 2325 450 2341 484
rect 2375 450 2391 484
rect 2425 580 2471 596
rect 2425 546 2431 580
rect 2465 546 2471 580
rect 2425 494 2471 546
rect 2425 460 2431 494
rect 2465 460 2471 494
rect 2505 580 2571 649
rect 2505 546 2521 580
rect 2555 546 2571 580
rect 2505 498 2571 546
rect 2505 464 2521 498
rect 2555 464 2571 498
rect 2425 430 2471 460
rect 2425 416 2567 430
rect 2235 414 2567 416
rect 2235 380 2251 414
rect 2285 380 2431 414
rect 2465 380 2567 414
rect 2235 364 2567 380
rect 2041 314 2399 330
rect 2041 298 2213 314
rect 1509 168 1890 202
rect 1824 147 1890 168
rect 1261 51 1475 85
rect 1587 100 1603 134
rect 1637 100 1671 134
rect 1705 100 1740 134
rect 1774 100 1790 134
rect 1587 17 1790 100
rect 1824 113 1840 147
rect 1874 113 1890 147
rect 1824 84 1890 113
rect 1936 280 2213 298
rect 2247 280 2281 314
rect 2315 280 2349 314
rect 2383 280 2399 314
rect 1936 264 2399 280
rect 1936 210 2002 264
rect 2521 230 2567 364
rect 1936 176 1952 210
rect 1986 176 2002 210
rect 1936 120 2002 176
rect 1936 86 1952 120
rect 1986 86 2002 120
rect 1936 70 2002 86
rect 2036 210 2102 226
rect 2036 176 2052 210
rect 2086 176 2102 210
rect 2036 120 2102 176
rect 2036 86 2052 120
rect 2086 86 2102 120
rect 2036 17 2102 86
rect 2136 210 2567 230
rect 2136 176 2152 210
rect 2186 196 2419 210
rect 2186 176 2202 196
rect 2136 120 2202 176
rect 2403 176 2419 196
rect 2453 196 2567 210
rect 2453 176 2469 196
rect 2136 86 2152 120
rect 2186 86 2202 120
rect 2136 70 2202 86
rect 2236 144 2369 160
rect 2236 110 2238 144
rect 2272 110 2324 144
rect 2358 110 2369 144
rect 2236 17 2369 110
rect 2403 120 2469 176
rect 2403 86 2419 120
rect 2453 86 2469 120
rect 2403 70 2469 86
rect 2503 146 2569 162
rect 2503 112 2519 146
rect 2553 112 2569 146
rect 2503 17 2569 112
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2592 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 1087 348 1089 350
rect 1089 348 1121 350
rect 1087 316 1121 348
rect 1663 320 1687 350
rect 1687 320 1697 350
rect 1663 316 1697 320
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
<< metal1 >>
rect 0 683 2592 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2592 683
rect 0 617 2592 649
rect 1075 350 1133 356
rect 1075 316 1087 350
rect 1121 347 1133 350
rect 1651 350 1709 356
rect 1651 347 1663 350
rect 1121 319 1663 347
rect 1121 316 1133 319
rect 1075 310 1133 316
rect 1651 316 1663 319
rect 1697 316 1709 350
rect 1651 310 1709 316
rect 0 17 2592 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2592 17
rect 0 -49 2592 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dfstp_4
flabel comment s 861 265 861 265 0 FreeSans 200 0 0 0 no_jumper_check
flabel comment s 643 320 643 320 0 FreeSans 200 0 0 0 no_jumper_check
flabel pwell s 0 0 2592 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 2592 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 1663 316 1697 350 0 FreeSans 340 0 0 0 SET_B
port 3 nsew
flabel metal1 s 0 617 2592 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 2592 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 319 242 353 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 127 242 161 276 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 2527 242 2561 276 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 2527 316 2561 350 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 2527 390 2561 424 0 FreeSans 340 0 0 0 Q
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 2592 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2715150
string GDS_START 2696320
<< end >>
