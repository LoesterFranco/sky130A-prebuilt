magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1012 561
rect 103 367 169 527
rect 282 367 348 527
rect 450 367 528 527
rect 638 296 704 415
rect 806 296 872 415
rect 17 199 69 265
rect 103 17 169 97
rect 291 17 357 97
rect 459 17 525 97
rect 638 124 872 296
rect 906 124 995 265
rect 0 -17 1012 17
<< obsli1 >>
rect 17 333 69 493
rect 203 333 248 493
rect 382 333 416 493
rect 562 459 995 493
rect 562 333 604 459
rect 17 299 169 333
rect 203 299 604 333
rect 103 265 169 299
rect 738 330 772 459
rect 906 330 995 459
rect 103 199 604 265
rect 103 165 169 199
rect 17 131 169 165
rect 203 131 599 165
rect 17 51 69 131
rect 203 51 257 131
rect 391 51 425 131
rect 565 90 599 131
rect 565 51 995 90
<< metal1 >>
rect 0 496 1012 592
rect 0 -48 1012 48
<< labels >>
rlabel locali s 906 124 995 265 6 A
port 1 nsew signal input
rlabel locali s 17 199 69 265 6 TE_B
port 2 nsew signal input
rlabel locali s 806 296 872 415 6 Z
port 3 nsew signal output
rlabel locali s 638 296 704 415 6 Z
port 3 nsew signal output
rlabel locali s 638 124 872 296 6 Z
port 3 nsew signal output
rlabel locali s 459 17 525 97 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 291 17 357 97 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 103 17 169 97 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 1012 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1012 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 450 367 528 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 282 367 348 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 103 367 169 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 1012 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 1012 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1012 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2907972
string GDS_START 2900194
<< end >>
