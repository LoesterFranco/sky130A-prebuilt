magic
tech sky130A
magscale 1 2
timestamp 1604502701
<< nwell >>
rect -38 332 2630 704
<< pwell >>
rect 0 0 2592 49
<< scpmos >>
rect 104 368 134 592
rect 220 368 250 592
rect 489 463 519 547
rect 579 463 609 547
rect 683 379 713 463
rect 761 379 791 463
rect 879 379 909 547
rect 987 379 1017 547
rect 1071 379 1101 547
rect 1173 379 1203 547
rect 1281 424 1311 592
rect 1388 508 1418 592
rect 1477 508 1507 592
rect 1681 392 1711 592
rect 1784 392 1814 592
rect 1867 392 1897 592
rect 2078 368 2108 496
rect 2181 368 2211 592
rect 2375 410 2405 578
rect 2478 368 2508 592
<< nmoslvt >>
rect 84 74 114 222
rect 184 74 214 222
rect 392 125 422 209
rect 490 87 520 171
rect 576 87 606 171
rect 671 119 701 203
rect 842 119 872 229
rect 976 119 1006 229
rect 1062 119 1092 229
rect 1288 119 1318 229
rect 1360 119 1390 229
rect 1468 74 1498 158
rect 1576 74 1606 158
rect 1678 74 1708 222
rect 1778 74 1808 222
rect 1865 74 1895 222
rect 2072 74 2102 158
rect 2188 74 2218 222
rect 2386 74 2416 158
rect 2481 74 2511 222
<< ndiff >>
rect 27 202 84 222
rect 27 168 39 202
rect 73 168 84 202
rect 27 120 84 168
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 202 184 222
rect 114 168 139 202
rect 173 168 184 202
rect 114 120 184 168
rect 114 86 139 120
rect 173 86 184 120
rect 114 74 184 86
rect 214 210 271 222
rect 214 176 225 210
rect 259 176 271 210
rect 214 120 271 176
rect 214 86 225 120
rect 259 86 271 120
rect 214 74 271 86
rect 335 184 392 209
rect 335 150 347 184
rect 381 150 392 184
rect 335 125 392 150
rect 422 184 475 209
rect 422 150 433 184
rect 467 171 475 184
rect 792 203 842 229
rect 621 171 671 203
rect 467 150 490 171
rect 422 125 490 150
rect 440 87 490 125
rect 520 133 576 171
rect 520 99 531 133
rect 565 99 576 133
rect 520 87 576 99
rect 606 119 671 171
rect 701 119 842 203
rect 872 119 976 229
rect 1006 177 1062 229
rect 1006 143 1017 177
rect 1051 143 1062 177
rect 1006 119 1062 143
rect 1092 119 1163 229
rect 606 87 656 119
rect 716 112 827 119
rect 716 78 754 112
rect 788 78 827 112
rect 887 112 961 119
rect 716 66 827 78
rect 887 78 907 112
rect 941 78 961 112
rect 1107 117 1163 119
rect 887 66 961 78
rect 1107 83 1118 117
rect 1152 83 1163 117
rect 1107 71 1163 83
rect 1217 201 1288 229
rect 1217 167 1243 201
rect 1277 167 1288 201
rect 1217 119 1288 167
rect 1318 119 1360 229
rect 1390 169 1446 229
rect 1390 135 1401 169
rect 1435 158 1446 169
rect 1621 192 1678 222
rect 1621 158 1633 192
rect 1667 158 1678 192
rect 1435 135 1468 158
rect 1390 119 1468 135
rect 1217 118 1273 119
rect 1217 84 1228 118
rect 1262 84 1273 118
rect 1217 72 1273 84
rect 1418 74 1468 119
rect 1498 74 1576 158
rect 1606 116 1678 158
rect 1606 82 1633 116
rect 1667 82 1678 116
rect 1606 74 1678 82
rect 1708 192 1778 222
rect 1708 158 1733 192
rect 1767 158 1778 192
rect 1708 116 1778 158
rect 1708 82 1733 116
rect 1767 82 1778 116
rect 1708 74 1778 82
rect 1808 172 1865 222
rect 1808 138 1820 172
rect 1854 138 1865 172
rect 1808 74 1865 138
rect 1895 188 1957 222
rect 1895 154 1911 188
rect 1945 154 1957 188
rect 2138 158 2188 222
rect 1895 120 1957 154
rect 1895 86 1911 120
rect 1945 86 1957 120
rect 1895 74 1957 86
rect 2015 133 2072 158
rect 2015 99 2027 133
rect 2061 99 2072 133
rect 2015 74 2072 99
rect 2102 133 2188 158
rect 2102 99 2129 133
rect 2163 99 2188 133
rect 2102 74 2188 99
rect 2218 210 2275 222
rect 2218 176 2229 210
rect 2263 176 2275 210
rect 2218 120 2275 176
rect 2431 158 2481 222
rect 2218 86 2229 120
rect 2263 86 2275 120
rect 2218 74 2275 86
rect 2329 133 2386 158
rect 2329 99 2341 133
rect 2375 99 2386 133
rect 2329 74 2386 99
rect 2416 133 2481 158
rect 2416 99 2427 133
rect 2461 99 2481 133
rect 2416 74 2481 99
rect 2511 210 2565 222
rect 2511 176 2522 210
rect 2556 176 2565 210
rect 2511 120 2565 176
rect 2511 86 2522 120
rect 2556 86 2565 120
rect 2511 74 2565 86
<< pdiff >>
rect 45 580 104 592
rect 45 546 57 580
rect 91 546 104 580
rect 45 497 104 546
rect 45 463 57 497
rect 91 463 104 497
rect 45 414 104 463
rect 45 380 57 414
rect 91 380 104 414
rect 45 368 104 380
rect 134 582 220 592
rect 134 548 157 582
rect 191 548 220 582
rect 134 514 220 548
rect 134 480 157 514
rect 191 480 220 514
rect 134 446 220 480
rect 134 412 157 446
rect 191 412 220 446
rect 134 368 220 412
rect 250 580 305 592
rect 250 546 263 580
rect 297 546 305 580
rect 250 497 305 546
rect 250 463 263 497
rect 297 463 305 497
rect 250 414 305 463
rect 250 380 263 414
rect 297 380 305 414
rect 250 368 305 380
rect 365 535 489 547
rect 365 501 373 535
rect 407 501 441 535
rect 475 501 489 535
rect 365 463 489 501
rect 519 522 579 547
rect 519 488 532 522
rect 566 488 579 522
rect 519 463 579 488
rect 609 463 662 547
rect 1228 547 1281 592
rect 826 463 879 547
rect 627 451 683 463
rect 627 417 636 451
rect 670 417 683 451
rect 627 379 683 417
rect 713 379 761 463
rect 791 447 879 463
rect 791 413 804 447
rect 838 413 879 447
rect 791 379 879 413
rect 909 531 987 547
rect 909 497 940 531
rect 974 497 987 531
rect 909 425 987 497
rect 909 391 940 425
rect 974 391 987 425
rect 909 379 987 391
rect 1017 379 1071 547
rect 1101 535 1173 547
rect 1101 501 1120 535
rect 1154 501 1173 535
rect 1101 379 1173 501
rect 1203 424 1281 547
rect 1311 547 1388 592
rect 1311 513 1324 547
rect 1358 513 1388 547
rect 1311 508 1388 513
rect 1418 508 1477 592
rect 1507 580 1681 592
rect 1507 546 1528 580
rect 1562 546 1634 580
rect 1668 546 1681 580
rect 1507 508 1681 546
rect 1311 471 1370 508
rect 1311 437 1324 471
rect 1358 437 1370 471
rect 1311 424 1370 437
rect 1203 379 1256 424
rect 1628 392 1681 508
rect 1711 580 1784 592
rect 1711 546 1737 580
rect 1771 546 1784 580
rect 1711 512 1784 546
rect 1711 478 1737 512
rect 1771 478 1784 512
rect 1711 444 1784 478
rect 1711 410 1737 444
rect 1771 410 1784 444
rect 1711 392 1784 410
rect 1814 392 1867 592
rect 1897 573 1956 592
rect 1897 539 1910 573
rect 1944 539 1956 573
rect 1897 392 1956 539
rect 2126 566 2181 592
rect 2126 532 2134 566
rect 2168 532 2181 566
rect 2126 496 2181 532
rect 2023 414 2078 496
rect 2023 380 2031 414
rect 2065 380 2078 414
rect 2023 368 2078 380
rect 2108 368 2181 496
rect 2211 580 2266 592
rect 2211 546 2224 580
rect 2258 546 2266 580
rect 2423 580 2478 592
rect 2423 578 2431 580
rect 2211 497 2266 546
rect 2211 463 2224 497
rect 2258 463 2266 497
rect 2211 414 2266 463
rect 2211 380 2224 414
rect 2258 380 2266 414
rect 2320 566 2375 578
rect 2320 532 2328 566
rect 2362 532 2375 566
rect 2320 456 2375 532
rect 2320 422 2328 456
rect 2362 422 2375 456
rect 2320 410 2375 422
rect 2405 546 2431 578
rect 2465 546 2478 580
rect 2405 497 2478 546
rect 2405 463 2431 497
rect 2465 463 2478 497
rect 2405 414 2478 463
rect 2405 410 2431 414
rect 2211 368 2266 380
rect 2423 380 2431 410
rect 2465 380 2478 414
rect 2423 368 2478 380
rect 2508 580 2565 592
rect 2508 546 2521 580
rect 2555 546 2565 580
rect 2508 497 2565 546
rect 2508 463 2521 497
rect 2555 463 2565 497
rect 2508 414 2565 463
rect 2508 380 2521 414
rect 2555 380 2565 414
rect 2508 368 2565 380
<< ndiffc >>
rect 39 168 73 202
rect 39 86 73 120
rect 139 168 173 202
rect 139 86 173 120
rect 225 176 259 210
rect 225 86 259 120
rect 347 150 381 184
rect 433 150 467 184
rect 531 99 565 133
rect 1017 143 1051 177
rect 754 78 788 112
rect 907 78 941 112
rect 1118 83 1152 117
rect 1243 167 1277 201
rect 1401 135 1435 169
rect 1633 158 1667 192
rect 1228 84 1262 118
rect 1633 82 1667 116
rect 1733 158 1767 192
rect 1733 82 1767 116
rect 1820 138 1854 172
rect 1911 154 1945 188
rect 1911 86 1945 120
rect 2027 99 2061 133
rect 2129 99 2163 133
rect 2229 176 2263 210
rect 2229 86 2263 120
rect 2341 99 2375 133
rect 2427 99 2461 133
rect 2522 176 2556 210
rect 2522 86 2556 120
<< pdiffc >>
rect 57 546 91 580
rect 57 463 91 497
rect 57 380 91 414
rect 157 548 191 582
rect 157 480 191 514
rect 157 412 191 446
rect 263 546 297 580
rect 263 463 297 497
rect 263 380 297 414
rect 373 501 407 535
rect 441 501 475 535
rect 532 488 566 522
rect 636 417 670 451
rect 804 413 838 447
rect 940 497 974 531
rect 940 391 974 425
rect 1120 501 1154 535
rect 1324 513 1358 547
rect 1528 546 1562 580
rect 1634 546 1668 580
rect 1324 437 1358 471
rect 1737 546 1771 580
rect 1737 478 1771 512
rect 1737 410 1771 444
rect 1910 539 1944 573
rect 2134 532 2168 566
rect 2031 380 2065 414
rect 2224 546 2258 580
rect 2224 463 2258 497
rect 2224 380 2258 414
rect 2328 532 2362 566
rect 2328 422 2362 456
rect 2431 546 2465 580
rect 2431 463 2465 497
rect 2431 380 2465 414
rect 2521 546 2555 580
rect 2521 463 2555 497
rect 2521 380 2555 414
<< poly >>
rect 104 592 134 618
rect 220 592 250 618
rect 320 615 1314 645
rect 104 353 134 368
rect 220 353 250 368
rect 101 310 137 353
rect 217 326 253 353
rect 71 294 137 310
rect 71 260 87 294
rect 121 260 137 294
rect 179 310 253 326
rect 179 276 195 310
rect 229 290 253 310
rect 320 290 350 615
rect 489 547 519 573
rect 579 547 609 573
rect 680 478 716 615
rect 1278 607 1314 615
rect 1281 592 1311 607
rect 1388 592 1418 618
rect 1477 592 1507 618
rect 1681 592 1711 618
rect 1784 592 1814 618
rect 1867 592 1897 618
rect 2181 592 2211 618
rect 879 547 909 573
rect 987 547 1017 573
rect 1071 547 1101 573
rect 1173 547 1203 573
rect 683 463 713 478
rect 761 463 791 489
rect 489 448 519 463
rect 579 448 609 463
rect 486 431 522 448
rect 229 276 350 290
rect 179 260 350 276
rect 392 415 522 431
rect 392 381 408 415
rect 442 401 522 415
rect 442 381 458 401
rect 392 365 458 381
rect 71 244 137 260
rect 84 222 114 244
rect 184 222 214 260
rect 84 48 114 74
rect 184 48 214 74
rect 290 51 320 260
rect 392 209 422 365
rect 464 301 530 317
rect 464 267 480 301
rect 514 281 530 301
rect 576 281 612 448
rect 1388 493 1418 508
rect 1477 493 1507 508
rect 1385 466 1421 493
rect 1474 476 1510 493
rect 1385 436 1426 466
rect 1474 460 1590 476
rect 1474 446 1540 460
rect 1281 409 1311 424
rect 1278 388 1314 409
rect 683 353 713 379
rect 761 364 791 379
rect 879 364 909 379
rect 987 364 1017 379
rect 1071 364 1101 379
rect 1173 364 1203 379
rect 1278 372 1354 388
rect 758 291 794 364
rect 876 339 912 364
rect 514 267 612 281
rect 464 251 612 267
rect 671 275 794 291
rect 490 171 520 197
rect 576 171 606 251
rect 671 241 701 275
rect 735 261 794 275
rect 842 323 912 339
rect 842 289 862 323
rect 896 289 912 323
rect 984 317 1020 364
rect 1068 317 1104 364
rect 1170 317 1206 364
rect 1278 338 1304 372
rect 1338 338 1354 372
rect 1278 322 1354 338
rect 842 273 912 289
rect 954 301 1020 317
rect 735 241 751 261
rect 671 225 751 241
rect 842 229 872 273
rect 954 267 970 301
rect 1004 267 1020 301
rect 954 251 1020 267
rect 1062 301 1128 317
rect 1062 267 1078 301
rect 1112 267 1128 301
rect 1062 251 1128 267
rect 1170 301 1236 317
rect 1170 267 1186 301
rect 1220 274 1236 301
rect 1396 274 1426 436
rect 1524 426 1540 446
rect 1574 426 1590 460
rect 1524 410 1590 426
rect 1560 377 1590 410
rect 2078 496 2108 522
rect 1681 377 1711 392
rect 1784 377 1814 392
rect 1867 377 1897 392
rect 1560 347 1606 377
rect 1678 360 1714 377
rect 1220 267 1318 274
rect 976 229 1006 251
rect 1062 229 1092 251
rect 1170 244 1318 267
rect 1288 229 1318 244
rect 1360 244 1426 274
rect 1360 229 1390 244
rect 1468 230 1534 246
rect 671 203 701 225
rect 392 99 422 125
rect 671 93 701 119
rect 490 51 520 87
rect 290 21 520 51
rect 576 51 606 87
rect 842 93 872 119
rect 976 93 1006 119
rect 1062 93 1092 119
rect 1468 196 1484 230
rect 1518 196 1534 230
rect 1468 180 1534 196
rect 1468 158 1498 180
rect 1576 158 1606 347
rect 1648 344 1714 360
rect 1648 310 1664 344
rect 1698 310 1714 344
rect 1781 310 1817 377
rect 1648 294 1714 310
rect 1756 294 1822 310
rect 1678 222 1708 294
rect 1756 260 1772 294
rect 1806 260 1822 294
rect 1756 244 1822 260
rect 1864 274 1900 377
rect 2375 578 2405 604
rect 2478 592 2508 618
rect 2375 395 2405 410
rect 2078 353 2108 368
rect 2181 353 2211 368
rect 2327 365 2408 395
rect 2075 330 2111 353
rect 2178 330 2214 353
rect 2327 330 2357 365
rect 2478 353 2508 368
rect 2050 314 2116 330
rect 1942 294 2008 310
rect 1942 274 1958 294
rect 1864 260 1958 274
rect 1992 260 2008 294
rect 1864 244 2008 260
rect 2050 280 2066 314
rect 2100 280 2116 314
rect 2050 246 2116 280
rect 2158 314 2357 330
rect 2475 317 2511 353
rect 2158 280 2174 314
rect 2208 280 2357 314
rect 2158 264 2357 280
rect 1778 222 1808 244
rect 1865 222 1895 244
rect 1288 93 1318 119
rect 1360 51 1390 119
rect 2050 212 2066 246
rect 2100 212 2116 246
rect 2188 222 2218 264
rect 2050 196 2116 212
rect 2072 158 2102 196
rect 2327 203 2357 264
rect 2405 301 2511 317
rect 2405 267 2421 301
rect 2455 267 2511 301
rect 2405 251 2511 267
rect 2481 222 2511 251
rect 2327 173 2416 203
rect 2386 158 2416 173
rect 576 21 1390 51
rect 1468 48 1498 74
rect 1576 48 1606 74
rect 1678 48 1708 74
rect 1778 48 1808 74
rect 1865 48 1895 74
rect 2072 48 2102 74
rect 2188 48 2218 74
rect 2386 48 2416 74
rect 2481 48 2511 74
<< polycont >>
rect 87 260 121 294
rect 195 276 229 310
rect 408 381 442 415
rect 480 267 514 301
rect 701 241 735 275
rect 862 289 896 323
rect 1304 338 1338 372
rect 970 267 1004 301
rect 1078 267 1112 301
rect 1186 267 1220 301
rect 1540 426 1574 460
rect 1484 196 1518 230
rect 1664 310 1698 344
rect 1772 260 1806 294
rect 1958 260 1992 294
rect 2066 280 2100 314
rect 2174 280 2208 314
rect 2066 212 2100 246
rect 2421 267 2455 301
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2592 683
rect 17 580 107 596
rect 17 546 57 580
rect 91 546 107 580
rect 17 497 107 546
rect 17 463 57 497
rect 91 463 107 497
rect 17 414 107 463
rect 17 380 57 414
rect 91 380 107 414
rect 141 582 207 649
rect 141 548 157 582
rect 191 548 207 582
rect 141 514 207 548
rect 141 480 157 514
rect 191 480 207 514
rect 141 446 207 480
rect 141 412 157 446
rect 191 412 207 446
rect 263 580 313 596
rect 297 546 313 580
rect 263 497 313 546
rect 297 463 313 497
rect 361 535 482 649
rect 361 501 373 535
rect 407 501 441 535
rect 475 501 482 535
rect 361 485 482 501
rect 516 522 591 551
rect 516 488 532 522
rect 566 488 591 522
rect 263 414 313 463
rect 516 459 591 488
rect 17 378 107 380
rect 297 380 313 414
rect 17 344 229 378
rect 17 202 51 344
rect 195 310 229 344
rect 85 294 161 310
rect 85 260 87 294
rect 121 260 161 294
rect 195 260 229 276
rect 263 317 313 380
rect 392 415 458 431
rect 392 381 408 415
rect 442 381 458 415
rect 392 365 458 381
rect 263 301 523 317
rect 263 267 480 301
rect 514 267 523 301
rect 85 236 161 260
rect 263 251 523 267
rect 263 226 297 251
rect 225 210 297 226
rect 557 217 591 459
rect 17 168 39 202
rect 73 168 89 202
rect 17 120 89 168
rect 17 86 39 120
rect 73 86 89 120
rect 17 70 89 86
rect 123 168 139 202
rect 173 168 189 202
rect 123 120 189 168
rect 123 86 139 120
rect 173 86 189 120
rect 123 17 189 86
rect 259 176 297 210
rect 225 120 297 176
rect 259 86 297 120
rect 225 70 297 86
rect 331 184 381 213
rect 331 150 347 184
rect 331 17 381 150
rect 417 184 591 217
rect 417 150 433 184
rect 467 183 591 184
rect 625 451 686 467
rect 625 417 636 451
rect 670 417 686 451
rect 625 359 686 417
rect 788 447 838 649
rect 788 413 804 447
rect 788 393 838 413
rect 872 581 1066 615
rect 625 325 812 359
rect 872 331 906 581
rect 940 531 990 547
rect 974 497 990 531
rect 940 425 990 497
rect 1032 467 1066 581
rect 1100 535 1174 649
rect 1100 501 1120 535
rect 1154 501 1174 535
rect 1208 581 1490 615
rect 1208 467 1242 581
rect 1032 433 1242 467
rect 1308 513 1324 547
rect 1358 513 1374 547
rect 1308 471 1374 513
rect 1308 437 1324 471
rect 1358 456 1374 471
rect 1358 437 1422 456
rect 974 399 990 425
rect 1308 422 1422 437
rect 974 391 1204 399
rect 940 365 1204 391
rect 417 121 467 150
rect 625 149 659 325
rect 515 133 659 149
rect 693 275 744 291
rect 693 241 701 275
rect 735 241 744 275
rect 693 180 744 241
rect 778 248 812 325
rect 846 323 912 331
rect 846 289 862 323
rect 896 289 912 323
rect 1170 317 1204 365
rect 1288 372 1354 388
rect 1288 338 1304 372
rect 1338 338 1354 372
rect 1288 322 1354 338
rect 846 282 912 289
rect 949 301 1020 317
rect 949 267 970 301
rect 1004 267 1020 301
rect 949 251 1020 267
rect 1062 301 1128 317
rect 1062 267 1078 301
rect 1112 276 1128 301
rect 949 248 983 251
rect 778 214 983 248
rect 1062 242 1087 267
rect 1121 242 1128 276
rect 1062 236 1128 242
rect 1170 301 1236 317
rect 1170 267 1186 301
rect 1220 267 1236 301
rect 1170 251 1236 267
rect 1170 202 1204 251
rect 1017 180 1204 202
rect 693 177 1204 180
rect 693 146 1017 177
rect 515 99 531 133
rect 565 99 659 133
rect 1003 143 1017 146
rect 1051 168 1204 177
rect 1238 201 1286 217
rect 1051 143 1067 168
rect 1003 119 1067 143
rect 1238 167 1243 201
rect 1277 167 1286 201
rect 1238 134 1286 167
rect 1102 117 1168 134
rect 515 83 659 99
rect 712 78 754 112
rect 788 78 831 112
rect 712 17 831 78
rect 883 78 907 112
rect 941 85 965 112
rect 1102 85 1118 117
rect 941 83 1118 85
rect 1152 83 1168 117
rect 941 78 1168 83
rect 883 51 1168 78
rect 1212 118 1286 134
rect 1212 84 1228 118
rect 1262 84 1286 118
rect 1212 17 1286 84
rect 1320 85 1354 322
rect 1388 314 1422 422
rect 1456 382 1490 581
rect 1524 580 1684 649
rect 1524 546 1528 580
rect 1562 546 1634 580
rect 1668 546 1684 580
rect 1524 530 1684 546
rect 1737 580 1787 596
rect 1771 546 1787 580
rect 1737 512 1787 546
rect 1894 573 1960 649
rect 1894 539 1910 573
rect 1944 539 1960 573
rect 1894 516 1960 539
rect 2118 566 2184 649
rect 2118 532 2134 566
rect 2168 532 2184 566
rect 2118 516 2184 532
rect 2224 580 2292 596
rect 2258 546 2292 580
rect 1771 482 1787 512
rect 2224 497 2292 546
rect 1771 478 2190 482
rect 1737 476 2190 478
rect 1524 460 2190 476
rect 1524 426 1540 460
rect 1574 448 2190 460
rect 1574 444 1877 448
rect 1574 426 1737 444
rect 1524 416 1737 426
rect 1771 410 1877 444
rect 1737 394 1877 410
rect 1456 360 1703 382
rect 1456 348 1714 360
rect 1648 344 1714 348
rect 1388 280 1614 314
rect 1648 310 1664 344
rect 1698 310 1714 344
rect 1648 294 1714 310
rect 1756 294 1809 310
rect 1388 169 1435 280
rect 1580 260 1614 280
rect 1756 260 1772 294
rect 1806 260 1809 294
rect 1388 135 1401 169
rect 1388 119 1435 135
rect 1469 230 1534 246
rect 1469 196 1484 230
rect 1518 196 1534 230
rect 1580 226 1809 260
rect 1469 85 1534 196
rect 1843 192 1877 394
rect 1942 380 2031 414
rect 2065 380 2081 414
rect 1942 364 2081 380
rect 1942 294 2013 364
rect 2156 330 2190 448
rect 2258 463 2292 497
rect 2224 414 2292 463
rect 2258 380 2292 414
rect 2224 364 2292 380
rect 1942 276 1958 294
rect 1942 242 1951 276
rect 1992 260 2013 294
rect 1985 242 2013 260
rect 1942 238 2013 242
rect 1320 51 1534 85
rect 1617 158 1633 192
rect 1667 158 1683 192
rect 1617 116 1683 158
rect 1617 82 1633 116
rect 1667 82 1683 116
rect 1617 17 1683 82
rect 1717 158 1733 192
rect 1767 158 1783 192
rect 1717 116 1783 158
rect 1817 172 1877 192
rect 1817 138 1820 172
rect 1854 138 1877 172
rect 1817 119 1877 138
rect 1911 188 1945 204
rect 1911 120 1945 154
rect 1717 82 1733 116
rect 1767 85 1783 116
rect 1911 85 1945 86
rect 1767 82 1945 85
rect 1717 51 1945 82
rect 1979 162 2013 238
rect 2047 314 2116 330
rect 2047 280 2066 314
rect 2100 280 2116 314
rect 2047 246 2116 280
rect 2156 314 2224 330
rect 2156 280 2174 314
rect 2208 280 2224 314
rect 2156 264 2224 280
rect 2047 212 2066 246
rect 2100 212 2116 246
rect 2258 226 2292 364
rect 2047 196 2116 212
rect 2213 210 2292 226
rect 2213 176 2229 210
rect 2263 176 2292 210
rect 1979 133 2077 162
rect 1979 99 2027 133
rect 2061 99 2077 133
rect 1979 70 2077 99
rect 2113 133 2179 162
rect 2113 99 2129 133
rect 2163 99 2179 133
rect 2113 17 2179 99
rect 2213 120 2292 176
rect 2213 86 2229 120
rect 2263 86 2292 120
rect 2213 70 2292 86
rect 2328 566 2378 582
rect 2362 532 2378 566
rect 2328 456 2378 532
rect 2362 422 2378 456
rect 2328 406 2378 422
rect 2415 580 2465 649
rect 2415 546 2431 580
rect 2415 497 2465 546
rect 2415 463 2431 497
rect 2415 414 2465 463
rect 2328 317 2362 406
rect 2415 380 2431 414
rect 2415 364 2465 380
rect 2505 580 2572 596
rect 2505 546 2521 580
rect 2555 546 2572 580
rect 2505 497 2572 546
rect 2505 463 2521 497
rect 2555 463 2572 497
rect 2505 414 2572 463
rect 2505 380 2521 414
rect 2555 380 2572 414
rect 2328 301 2471 317
rect 2328 267 2421 301
rect 2455 267 2471 301
rect 2328 251 2471 267
rect 2328 133 2375 251
rect 2505 210 2572 380
rect 2505 176 2522 210
rect 2556 176 2572 210
rect 2328 99 2341 133
rect 2328 70 2375 99
rect 2411 133 2461 162
rect 2411 99 2427 133
rect 2411 17 2461 99
rect 2505 120 2572 176
rect 2505 86 2522 120
rect 2556 86 2572 120
rect 2505 70 2572 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2592 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 1087 267 1112 276
rect 1112 267 1121 276
rect 1087 242 1121 267
rect 1951 260 1958 276
rect 1958 260 1985 276
rect 1951 242 1985 260
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
<< metal1 >>
rect 0 683 2592 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2592 683
rect 0 617 2592 649
rect 1075 276 1133 282
rect 1075 242 1087 276
rect 1121 273 1133 276
rect 1939 276 1997 282
rect 1939 273 1951 276
rect 1121 245 1951 273
rect 1121 242 1133 245
rect 1075 236 1133 242
rect 1939 242 1951 245
rect 1985 242 1997 276
rect 1939 236 1997 242
rect 0 17 2592 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2592 17
rect 0 -49 2592 -17
<< labels >>
flabel comment s 640 631 640 631 0 FreeSans 200 0 0 0 no_jumper_check
rlabel comment s 0 0 0 0 4 dfbbp_1
flabel pwell s 0 0 2592 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 2592 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 2592 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 2592 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 2527 94 2561 128 0 FreeSans 340 0 0 0 Q
port 9 nsew
flabel corelocali s 2527 168 2561 202 0 FreeSans 340 0 0 0 Q
port 9 nsew
flabel corelocali s 2527 242 2561 276 0 FreeSans 340 0 0 0 Q
port 9 nsew
flabel corelocali s 2527 316 2561 350 0 FreeSans 340 0 0 0 Q
port 9 nsew
flabel corelocali s 2527 390 2561 424 0 FreeSans 340 0 0 0 Q
port 9 nsew
flabel corelocali s 2527 464 2561 498 0 FreeSans 340 0 0 0 Q
port 9 nsew
flabel corelocali s 2527 538 2561 572 0 FreeSans 340 0 0 0 Q
port 9 nsew
flabel corelocali s 127 242 161 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 415 390 449 424 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 2047 242 2081 276 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew
flabel corelocali s 2239 390 2273 424 0 FreeSans 340 0 0 0 Q_N
port 10 nsew
flabel corelocali s 2239 464 2273 498 0 FreeSans 340 0 0 0 Q_N
port 10 nsew
flabel corelocali s 2239 538 2273 572 0 FreeSans 340 0 0 0 Q_N
port 10 nsew
flabel corelocali s 1663 316 1697 350 0 FreeSans 340 0 0 0 SET_B
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 2592 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 2731958
string GDS_START 2712038
<< end >>
