magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 17 288 73 493
rect 17 70 69 288
rect 343 215 466 265
rect 1325 289 1451 323
rect 1325 199 1369 289
rect 1499 215 1643 265
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 107 443 184 527
rect 220 447 534 481
rect 685 447 751 527
rect 838 455 1497 489
rect 1583 455 1719 527
rect 220 409 264 447
rect 838 413 872 455
rect 107 375 264 409
rect 332 379 872 413
rect 107 266 151 375
rect 197 307 534 341
rect 103 173 151 266
rect 103 139 241 173
rect 103 17 163 105
rect 197 85 241 139
rect 275 119 309 307
rect 500 265 534 307
rect 578 305 655 339
rect 599 275 655 305
rect 500 199 565 265
rect 369 159 445 181
rect 599 159 633 275
rect 689 241 723 379
rect 769 289 873 343
rect 369 125 633 159
rect 667 207 723 241
rect 667 91 701 207
rect 434 85 531 91
rect 197 51 531 85
rect 575 57 701 91
rect 735 17 769 173
rect 815 83 873 289
rect 909 119 943 421
rect 977 178 1011 455
rect 1763 421 1822 493
rect 1057 323 1140 409
rect 1257 387 1822 421
rect 1057 289 1223 323
rect 1060 199 1145 254
rect 977 165 1029 178
rect 977 144 1069 165
rect 985 131 1069 144
rect 909 97 951 119
rect 909 53 991 97
rect 1035 64 1069 131
rect 1103 126 1145 199
rect 1189 85 1223 289
rect 1257 119 1291 387
rect 1715 375 1822 387
rect 1495 299 1732 341
rect 1698 265 1732 299
rect 1403 189 1465 255
rect 1698 199 1754 265
rect 1403 146 1444 189
rect 1698 181 1732 199
rect 1511 150 1732 181
rect 1503 147 1732 150
rect 1325 85 1428 93
rect 1189 51 1428 85
rect 1503 59 1561 147
rect 1788 117 1822 375
rect 1610 17 1702 113
rect 1762 51 1822 117
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
<< metal1 >>
rect 0 561 1840 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 0 496 1840 527
rect 0 17 1840 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
rect 0 -48 1840 -17
<< obsm1 >>
rect 609 320 667 329
rect 1099 320 1157 329
rect 609 292 1157 320
rect 609 283 667 292
rect 1099 283 1157 292
rect 803 184 861 193
rect 1099 184 1157 193
rect 1395 184 1453 193
rect 803 156 1453 184
rect 803 147 861 156
rect 1099 147 1157 156
rect 1395 147 1453 156
rect 905 116 963 125
rect 1497 116 1555 125
rect 905 88 1555 116
rect 905 79 963 88
rect 1497 79 1555 88
<< labels >>
rlabel locali s 1499 215 1643 265 6 A
port 1 nsew signal input
rlabel locali s 1325 289 1451 323 6 B
port 2 nsew signal input
rlabel locali s 1325 199 1369 289 6 B
port 2 nsew signal input
rlabel locali s 343 215 466 265 6 C
port 3 nsew signal input
rlabel locali s 17 288 73 493 6 X
port 4 nsew signal output
rlabel locali s 17 70 69 288 6 X
port 4 nsew signal output
rlabel metal1 s 0 -48 1840 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 1840 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1840 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 723090
string GDS_START 710828
<< end >>
