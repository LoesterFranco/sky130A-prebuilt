magic
tech sky130A
magscale 1 2
timestamp 1604502701
<< nwell >>
rect -38 332 230 704
<< pwell >>
rect 0 0 192 49
<< ndiode >>
rect 27 242 165 250
rect 27 208 39 242
rect 73 208 119 242
rect 153 208 165 242
rect 27 174 165 208
rect 27 140 39 174
rect 73 140 119 174
rect 153 140 165 174
rect 27 106 165 140
rect 27 72 39 106
rect 73 72 119 106
rect 153 72 165 106
rect 27 64 165 72
<< ndiodec >>
rect 39 208 73 242
rect 119 208 153 242
rect 39 140 73 174
rect 119 140 153 174
rect 39 72 73 106
rect 119 72 153 106
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 192 683
rect 19 242 173 613
rect 19 208 39 242
rect 73 208 119 242
rect 153 208 173 242
rect 19 174 173 208
rect 19 140 39 174
rect 73 140 119 174
rect 153 140 173 174
rect 19 106 173 140
rect 19 72 39 106
rect 73 72 119 106
rect 153 72 173 106
rect 19 53 173 72
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 192 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 31 -17 65 17
rect 127 -17 161 17
<< metal1 >>
rect 0 683 192 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 192 683
rect 0 617 192 649
rect 0 17 192 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 192 17
rect 0 -49 192 -17
<< labels >>
flabel corelocali s 31 464 65 498 0 FreeSans 200 0 0 0 DIODE
port 1 nsew
flabel corelocali s 127 168 161 202 0 FreeSans 200 0 0 0 DIODE
port 1 nsew
flabel corelocali s 127 464 161 498 0 FreeSans 200 0 0 0 DIODE
port 1 nsew
flabel corelocali s 31 94 65 128 0 FreeSans 200 0 0 0 DIODE
port 1 nsew
flabel corelocali s 127 242 161 276 0 FreeSans 200 0 0 0 DIODE
port 1 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 200 0 0 0 DIODE
port 1 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 200 0 0 0 DIODE
port 1 nsew
flabel corelocali s 31 168 65 202 0 FreeSans 200 0 0 0 DIODE
port 1 nsew
flabel corelocali s 127 94 161 128 0 FreeSans 200 0 0 0 DIODE
port 1 nsew
flabel corelocali s 31 538 65 572 0 FreeSans 200 0 0 0 DIODE
port 1 nsew
flabel corelocali s 31 390 65 424 0 FreeSans 200 0 0 0 DIODE
port 1 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 200 0 0 0 DIODE
port 1 nsew
flabel corelocali s 127 538 161 572 0 FreeSans 200 0 0 0 DIODE
port 1 nsew
flabel corelocali s 127 390 161 424 0 FreeSans 200 0 0 0 DIODE
port 1 nsew
flabel pwell s 0 0 192 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew
flabel nbase s 0 617 192 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew
rlabel comment s 0 0 0 0 4 diode_2
flabel metal1 s 0 617 192 666 0 FreeSans 200 0 0 0 VPWR
port 5 nsew
flabel metal1 s 0 0 192 49 0 FreeSans 200 0 0 0 VGND
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 192 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3006974
string GDS_START 3003156
<< end >>
