magic
tech sky130A
magscale 1 2
timestamp 1599588244
<< locali >>
rect 21 260 87 356
rect 213 364 359 430
rect 213 226 247 364
rect 395 270 461 430
rect 503 270 569 356
rect 213 192 291 226
rect 225 70 291 192
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 23 498 89 540
rect 130 532 196 649
rect 327 532 414 649
rect 23 464 529 498
rect 23 390 155 464
rect 121 226 155 390
rect 37 192 155 226
rect 281 260 359 326
rect 495 424 529 464
rect 647 458 751 572
rect 495 390 683 424
rect 617 270 683 390
rect 325 236 359 260
rect 717 236 751 458
rect 325 202 751 236
rect 37 108 121 192
rect 155 17 189 158
rect 325 17 427 156
rect 470 90 536 202
rect 570 17 636 168
rect 670 90 751 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel locali s 395 270 461 430 6 A
port 1 nsew signal input
rlabel locali s 503 270 569 356 6 B
port 2 nsew signal input
rlabel locali s 21 260 87 356 6 C_N
port 3 nsew signal input
rlabel locali s 225 70 291 192 6 X
port 4 nsew signal output
rlabel locali s 213 364 359 430 6 X
port 4 nsew signal output
rlabel locali s 213 226 247 364 6 X
port 4 nsew signal output
rlabel locali s 213 192 291 226 6 X
port 4 nsew signal output
rlabel metal1 s 0 -49 768 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 6 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 617 768 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 830120
string GDS_START 823926
<< end >>
