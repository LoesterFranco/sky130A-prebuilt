magic
tech sky130A
magscale 1 2
timestamp 1604502701
<< nwell >>
rect -38 357 1382 704
rect -38 332 534 357
rect 1007 332 1382 357
<< pwell >>
rect 0 0 1344 49
<< scpmos >>
rect 86 368 116 592
rect 228 392 258 592
rect 312 392 342 592
rect 454 508 484 592
rect 538 508 568 592
rect 647 398 677 566
rect 849 393 879 561
rect 957 393 987 561
rect 1049 393 1079 561
rect 1214 368 1244 592
<< nmoslvt >>
rect 84 74 114 222
rect 237 80 267 208
rect 315 80 345 208
rect 447 124 477 208
rect 525 124 555 208
rect 652 125 682 273
rect 852 125 882 273
rect 954 125 984 253
rect 1032 125 1062 253
rect 1230 74 1260 222
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 208 164 222
rect 602 208 652 273
rect 114 108 237 208
rect 114 74 141 108
rect 175 80 237 108
rect 267 80 315 208
rect 345 180 447 208
rect 345 146 379 180
rect 413 146 447 180
rect 345 124 447 146
rect 477 124 525 208
rect 555 171 652 208
rect 555 137 586 171
rect 620 137 652 171
rect 555 125 652 137
rect 682 250 739 273
rect 682 216 693 250
rect 727 216 739 250
rect 682 171 739 216
rect 682 137 693 171
rect 727 137 739 171
rect 682 125 739 137
rect 793 261 852 273
rect 793 227 806 261
rect 840 227 852 261
rect 793 125 852 227
rect 882 253 939 273
rect 882 245 954 253
rect 882 211 893 245
rect 927 211 954 245
rect 882 171 954 211
rect 882 137 893 171
rect 927 137 954 171
rect 882 125 954 137
rect 984 125 1032 253
rect 1062 241 1119 253
rect 1062 207 1073 241
rect 1107 207 1119 241
rect 1062 171 1119 207
rect 1062 137 1073 171
rect 1107 137 1119 171
rect 1062 125 1119 137
rect 1173 210 1230 222
rect 1173 176 1185 210
rect 1219 176 1230 210
rect 555 124 605 125
rect 345 80 395 124
rect 175 74 187 80
rect 129 62 187 74
rect 1173 120 1230 176
rect 1173 86 1185 120
rect 1219 86 1230 120
rect 1173 74 1230 86
rect 1260 210 1317 222
rect 1260 176 1271 210
rect 1305 176 1317 210
rect 1260 120 1317 176
rect 1260 86 1271 120
rect 1305 86 1317 120
rect 1260 74 1317 86
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 497 86 546
rect 27 463 39 497
rect 73 463 86 497
rect 27 414 86 463
rect 27 380 39 414
rect 73 380 86 414
rect 27 368 86 380
rect 116 580 228 592
rect 116 546 139 580
rect 173 546 228 580
rect 116 512 228 546
rect 116 478 139 512
rect 173 478 228 512
rect 116 392 228 478
rect 258 392 312 592
rect 342 560 454 592
rect 342 526 381 560
rect 415 526 454 560
rect 342 508 454 526
rect 484 508 538 592
rect 568 580 629 592
rect 568 546 583 580
rect 617 566 629 580
rect 617 546 647 566
rect 568 508 647 546
rect 342 392 395 508
rect 116 368 169 392
rect 594 398 647 508
rect 677 444 736 566
rect 1145 580 1214 592
rect 1145 561 1157 580
rect 677 410 690 444
rect 724 410 736 444
rect 677 398 736 410
rect 790 549 849 561
rect 790 515 802 549
rect 836 515 849 549
rect 790 439 849 515
rect 790 405 802 439
rect 836 405 849 439
rect 790 393 849 405
rect 879 549 957 561
rect 879 515 902 549
rect 936 515 957 549
rect 879 445 957 515
rect 879 411 902 445
rect 936 411 957 445
rect 879 393 957 411
rect 987 549 1049 561
rect 987 515 1002 549
rect 1036 515 1049 549
rect 987 445 1049 515
rect 987 411 1002 445
rect 1036 411 1049 445
rect 987 393 1049 411
rect 1079 546 1157 561
rect 1191 546 1214 580
rect 1079 509 1214 546
rect 1079 475 1157 509
rect 1191 475 1214 509
rect 1079 439 1214 475
rect 1079 405 1157 439
rect 1191 405 1214 439
rect 1079 393 1214 405
rect 1145 368 1214 393
rect 1244 580 1303 592
rect 1244 546 1257 580
rect 1291 546 1303 580
rect 1244 497 1303 546
rect 1244 463 1257 497
rect 1291 463 1303 497
rect 1244 414 1303 463
rect 1244 380 1257 414
rect 1291 380 1303 414
rect 1244 368 1303 380
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 141 74 175 108
rect 379 146 413 180
rect 586 137 620 171
rect 693 216 727 250
rect 693 137 727 171
rect 806 227 840 261
rect 893 211 927 245
rect 893 137 927 171
rect 1073 207 1107 241
rect 1073 137 1107 171
rect 1185 176 1219 210
rect 1185 86 1219 120
rect 1271 176 1305 210
rect 1271 86 1305 120
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 139 546 173 580
rect 139 478 173 512
rect 381 526 415 560
rect 583 546 617 580
rect 690 410 724 444
rect 802 515 836 549
rect 802 405 836 439
rect 902 515 936 549
rect 902 411 936 445
rect 1002 515 1036 549
rect 1002 411 1036 445
rect 1157 546 1191 580
rect 1157 475 1191 509
rect 1157 405 1191 439
rect 1257 546 1291 580
rect 1257 463 1291 497
rect 1257 380 1291 414
<< poly >>
rect 86 592 116 618
rect 228 592 258 618
rect 312 592 342 618
rect 454 592 484 618
rect 538 592 568 618
rect 1214 592 1244 618
rect 647 566 677 592
rect 454 493 484 508
rect 538 493 568 508
rect 451 476 487 493
rect 427 460 493 476
rect 427 426 443 460
rect 477 426 493 460
rect 427 410 493 426
rect 535 446 571 493
rect 535 416 579 446
rect 228 377 258 392
rect 312 377 342 392
rect 86 353 116 368
rect 225 360 261 377
rect 309 368 345 377
rect 83 326 119 353
rect 201 344 267 360
rect 83 310 153 326
rect 83 276 103 310
rect 137 276 153 310
rect 201 310 217 344
rect 251 310 267 344
rect 309 352 507 368
rect 309 338 457 352
rect 201 294 267 310
rect 441 318 457 338
rect 491 318 507 352
rect 441 302 507 318
rect 83 260 153 276
rect 84 222 114 260
rect 237 208 267 294
rect 315 280 399 296
rect 315 246 349 280
rect 383 246 399 280
rect 315 230 399 246
rect 315 208 345 230
rect 447 208 477 302
rect 549 253 579 416
rect 849 561 879 587
rect 957 561 987 587
rect 1049 561 1079 587
rect 647 383 677 398
rect 644 366 680 383
rect 849 378 879 393
rect 957 378 987 393
rect 1049 378 1079 393
rect 846 376 882 378
rect 954 376 990 378
rect 621 350 687 366
rect 621 316 637 350
rect 671 316 687 350
rect 621 300 687 316
rect 846 346 990 376
rect 846 345 984 346
rect 846 311 934 345
rect 968 311 984 345
rect 652 273 682 300
rect 846 295 984 311
rect 1046 298 1082 378
rect 1214 353 1244 368
rect 1211 326 1247 353
rect 852 273 882 295
rect 525 223 579 253
rect 525 208 555 223
rect 954 253 984 295
rect 1032 268 1082 298
rect 1141 310 1247 326
rect 1141 276 1157 310
rect 1191 290 1247 310
rect 1191 276 1260 290
rect 1032 253 1062 268
rect 1141 260 1260 276
rect 1230 222 1260 260
rect 447 98 477 124
rect 525 102 555 124
rect 525 86 591 102
rect 652 99 682 125
rect 852 99 882 125
rect 954 99 984 125
rect 84 48 114 74
rect 237 54 267 80
rect 315 54 345 80
rect 525 52 541 86
rect 575 52 591 86
rect 525 51 591 52
rect 1032 51 1062 125
rect 525 21 1062 51
rect 1230 48 1260 74
<< polycont >>
rect 443 426 477 460
rect 103 276 137 310
rect 217 310 251 344
rect 457 318 491 352
rect 349 246 383 280
rect 637 316 671 350
rect 934 311 968 345
rect 1157 276 1191 310
rect 541 52 575 86
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 19 580 89 596
rect 19 546 39 580
rect 73 546 89 580
rect 19 497 89 546
rect 19 463 39 497
rect 73 463 89 497
rect 19 414 89 463
rect 123 580 189 649
rect 123 546 139 580
rect 173 546 189 580
rect 567 580 633 649
rect 123 512 189 546
rect 123 478 139 512
rect 173 478 189 512
rect 123 462 189 478
rect 277 560 457 576
rect 277 526 381 560
rect 415 526 457 560
rect 567 546 583 580
rect 617 546 633 580
rect 789 549 852 565
rect 277 510 457 526
rect 789 515 802 549
rect 836 515 852 549
rect 789 512 852 515
rect 277 428 311 510
rect 606 478 852 512
rect 606 476 640 478
rect 19 380 39 414
rect 73 380 89 414
rect 19 364 89 380
rect 123 394 311 428
rect 345 460 640 476
rect 345 426 443 460
rect 477 426 640 460
rect 345 410 640 426
rect 674 410 690 444
rect 724 410 755 444
rect 19 226 53 364
rect 123 326 157 394
rect 87 310 157 326
rect 87 276 103 310
rect 137 276 157 310
rect 201 344 267 360
rect 201 310 217 344
rect 251 310 267 344
rect 201 294 267 310
rect 87 260 157 276
rect 345 280 399 410
rect 123 226 311 260
rect 345 246 349 280
rect 383 246 399 280
rect 345 230 399 246
rect 441 352 507 368
rect 441 318 457 352
rect 491 318 507 352
rect 441 266 507 318
rect 606 366 640 410
rect 606 350 687 366
rect 606 316 637 350
rect 671 316 687 350
rect 606 300 687 316
rect 721 266 755 410
rect 441 250 755 266
rect 441 232 693 250
rect 19 210 89 226
rect 19 176 39 210
rect 73 192 89 210
rect 277 196 311 226
rect 727 216 755 250
rect 73 176 243 192
rect 19 158 243 176
rect 19 120 89 158
rect 19 86 39 120
rect 73 86 89 120
rect 19 70 89 86
rect 125 108 175 124
rect 125 74 141 108
rect 125 17 175 74
rect 209 85 243 158
rect 277 180 452 196
rect 277 146 379 180
rect 413 146 452 180
rect 277 130 452 146
rect 550 171 659 187
rect 550 137 586 171
rect 620 137 659 171
rect 525 86 591 102
rect 525 85 541 86
rect 209 52 541 85
rect 575 52 591 86
rect 209 51 591 52
rect 625 17 659 137
rect 693 171 755 216
rect 789 439 852 478
rect 789 405 802 439
rect 836 405 852 439
rect 789 389 852 405
rect 886 549 952 649
rect 1141 580 1207 649
rect 886 515 902 549
rect 936 515 952 549
rect 886 445 952 515
rect 886 411 902 445
rect 936 411 952 445
rect 886 395 952 411
rect 986 549 1052 565
rect 986 515 1002 549
rect 1036 515 1052 549
rect 986 445 1052 515
rect 986 411 1002 445
rect 1036 429 1052 445
rect 1141 546 1157 580
rect 1191 546 1207 580
rect 1141 509 1207 546
rect 1141 475 1157 509
rect 1191 475 1207 509
rect 1141 439 1207 475
rect 1036 411 1107 429
rect 986 395 1107 411
rect 789 261 841 389
rect 889 345 1031 361
rect 889 311 934 345
rect 968 311 1031 345
rect 889 295 1031 311
rect 1073 326 1107 395
rect 1141 405 1157 439
rect 1191 405 1207 439
rect 1141 389 1207 405
rect 1241 580 1321 596
rect 1241 546 1257 580
rect 1291 546 1321 580
rect 1241 497 1321 546
rect 1241 463 1257 497
rect 1291 463 1321 497
rect 1241 414 1321 463
rect 1241 380 1257 414
rect 1291 380 1321 414
rect 1073 310 1207 326
rect 1241 310 1321 380
rect 1073 276 1157 310
rect 1191 276 1207 310
rect 789 227 806 261
rect 840 227 841 261
rect 789 211 841 227
rect 877 245 943 261
rect 1073 260 1207 276
rect 1073 257 1123 260
rect 877 211 893 245
rect 927 211 943 245
rect 727 137 755 171
rect 693 121 755 137
rect 877 171 943 211
rect 877 137 893 171
rect 927 137 943 171
rect 877 17 943 137
rect 1057 241 1123 257
rect 1057 207 1073 241
rect 1107 207 1123 241
rect 1057 171 1123 207
rect 1057 137 1073 171
rect 1107 137 1123 171
rect 1057 121 1123 137
rect 1169 210 1219 226
rect 1169 176 1185 210
rect 1169 120 1219 176
rect 1169 86 1185 120
rect 1169 17 1219 86
rect 1255 210 1321 310
rect 1255 176 1271 210
rect 1305 176 1321 210
rect 1255 120 1321 176
rect 1255 86 1271 120
rect 1305 86 1321 120
rect 1255 70 1321 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
<< metal1 >>
rect 0 683 1344 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 0 617 1344 649
rect 0 17 1344 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
rect 0 -49 1344 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dlclkp_1
flabel pwell s 0 0 1344 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 0 617 1344 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 0 617 1344 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 1344 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 1279 316 1313 350 0 FreeSans 340 0 0 0 GCLK
port 7 nsew
flabel corelocali s 1279 390 1313 424 0 FreeSans 340 0 0 0 GCLK
port 7 nsew
flabel corelocali s 1279 464 1313 498 0 FreeSans 340 0 0 0 GCLK
port 7 nsew
flabel corelocali s 1279 538 1313 572 0 FreeSans 340 0 0 0 GCLK
port 7 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 GATE
port 2 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 1344 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3017798
string GDS_START 3007032
<< end >>
