magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 1694 582
<< pwell >>
rect 124 -17 158 17
<< scnmos >>
rect 89 47 119 177
rect 183 47 213 177
rect 277 47 307 177
rect 371 47 401 177
rect 455 47 485 177
rect 549 47 579 177
rect 643 47 673 177
rect 737 47 767 177
rect 831 47 861 177
rect 925 47 955 177
rect 1019 47 1049 177
rect 1113 47 1143 177
rect 1207 47 1237 177
rect 1301 47 1331 177
rect 1395 47 1425 177
rect 1499 47 1529 177
<< pmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 457 297 493 497
rect 551 297 587 497
rect 645 297 681 497
rect 739 297 775 497
rect 833 297 869 497
rect 927 297 963 497
rect 1021 297 1057 497
rect 1115 297 1151 497
rect 1209 297 1245 497
rect 1303 297 1339 497
rect 1397 297 1433 497
rect 1491 297 1527 497
<< ndiff >>
rect 27 97 89 177
rect 27 63 35 97
rect 69 63 89 97
rect 27 47 89 63
rect 119 129 183 177
rect 119 95 129 129
rect 163 95 183 129
rect 119 47 183 95
rect 213 97 277 177
rect 213 63 223 97
rect 257 63 277 97
rect 213 47 277 63
rect 307 129 371 177
rect 307 95 317 129
rect 351 95 371 129
rect 307 47 371 95
rect 401 97 455 177
rect 401 63 411 97
rect 445 63 455 97
rect 401 47 455 63
rect 485 129 549 177
rect 485 95 505 129
rect 539 95 549 129
rect 485 47 549 95
rect 579 97 643 177
rect 579 63 599 97
rect 633 63 643 97
rect 579 47 643 63
rect 673 129 737 177
rect 673 95 693 129
rect 727 95 737 129
rect 673 47 737 95
rect 767 97 831 177
rect 767 63 787 97
rect 821 63 831 97
rect 767 47 831 63
rect 861 129 925 177
rect 861 95 881 129
rect 915 95 925 129
rect 861 47 925 95
rect 955 97 1019 177
rect 955 63 975 97
rect 1009 63 1019 97
rect 955 47 1019 63
rect 1049 129 1113 177
rect 1049 95 1069 129
rect 1103 95 1113 129
rect 1049 47 1113 95
rect 1143 97 1207 177
rect 1143 63 1163 97
rect 1197 63 1207 97
rect 1143 47 1207 63
rect 1237 129 1301 177
rect 1237 95 1257 129
rect 1291 95 1301 129
rect 1237 47 1301 95
rect 1331 97 1395 177
rect 1331 63 1351 97
rect 1385 63 1395 97
rect 1331 47 1395 63
rect 1425 129 1499 177
rect 1425 95 1445 129
rect 1479 95 1499 129
rect 1425 47 1499 95
rect 1529 161 1589 177
rect 1529 127 1539 161
rect 1573 127 1589 161
rect 1529 93 1589 127
rect 1529 59 1539 93
rect 1573 59 1589 93
rect 1529 47 1589 59
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 297 81 383
rect 117 479 175 497
rect 117 445 129 479
rect 163 445 175 479
rect 117 411 175 445
rect 117 377 129 411
rect 163 377 175 411
rect 117 343 175 377
rect 117 309 129 343
rect 163 309 175 343
rect 117 297 175 309
rect 211 485 269 497
rect 211 451 223 485
rect 257 451 269 485
rect 211 417 269 451
rect 211 383 223 417
rect 257 383 269 417
rect 211 297 269 383
rect 305 479 363 497
rect 305 445 317 479
rect 351 445 363 479
rect 305 411 363 445
rect 305 377 317 411
rect 351 377 363 411
rect 305 343 363 377
rect 305 309 317 343
rect 351 309 363 343
rect 305 297 363 309
rect 399 485 457 497
rect 399 451 411 485
rect 445 451 457 485
rect 399 417 457 451
rect 399 383 411 417
rect 445 383 457 417
rect 399 297 457 383
rect 493 463 551 497
rect 493 429 505 463
rect 539 429 551 463
rect 493 368 551 429
rect 493 334 505 368
rect 539 334 551 368
rect 493 297 551 334
rect 587 485 645 497
rect 587 451 599 485
rect 633 451 645 485
rect 587 417 645 451
rect 587 383 599 417
rect 633 383 645 417
rect 587 297 645 383
rect 681 463 739 497
rect 681 429 693 463
rect 727 429 739 463
rect 681 368 739 429
rect 681 334 693 368
rect 727 334 739 368
rect 681 297 739 334
rect 775 485 833 497
rect 775 451 787 485
rect 821 451 833 485
rect 775 417 833 451
rect 775 383 787 417
rect 821 383 833 417
rect 775 297 833 383
rect 869 463 927 497
rect 869 429 881 463
rect 915 429 927 463
rect 869 368 927 429
rect 869 334 881 368
rect 915 334 927 368
rect 869 297 927 334
rect 963 485 1021 497
rect 963 451 975 485
rect 1009 451 1021 485
rect 963 417 1021 451
rect 963 383 975 417
rect 1009 383 1021 417
rect 963 297 1021 383
rect 1057 463 1115 497
rect 1057 429 1069 463
rect 1103 429 1115 463
rect 1057 368 1115 429
rect 1057 334 1069 368
rect 1103 334 1115 368
rect 1057 297 1115 334
rect 1151 485 1209 497
rect 1151 451 1163 485
rect 1197 451 1209 485
rect 1151 417 1209 451
rect 1151 383 1163 417
rect 1197 383 1209 417
rect 1151 297 1209 383
rect 1245 463 1303 497
rect 1245 429 1257 463
rect 1291 429 1303 463
rect 1245 368 1303 429
rect 1245 334 1257 368
rect 1291 334 1303 368
rect 1245 297 1303 334
rect 1339 485 1397 497
rect 1339 451 1351 485
rect 1385 451 1397 485
rect 1339 417 1397 451
rect 1339 383 1351 417
rect 1385 383 1397 417
rect 1339 297 1397 383
rect 1433 463 1491 497
rect 1433 429 1445 463
rect 1479 429 1491 463
rect 1433 368 1491 429
rect 1433 334 1445 368
rect 1479 334 1491 368
rect 1433 297 1491 334
rect 1527 485 1589 497
rect 1527 451 1539 485
rect 1573 451 1589 485
rect 1527 417 1589 451
rect 1527 383 1539 417
rect 1573 383 1589 417
rect 1527 349 1589 383
rect 1527 315 1539 349
rect 1573 315 1589 349
rect 1527 297 1589 315
<< ndiffc >>
rect 35 63 69 97
rect 129 95 163 129
rect 223 63 257 97
rect 317 95 351 129
rect 411 63 445 97
rect 505 95 539 129
rect 599 63 633 97
rect 693 95 727 129
rect 787 63 821 97
rect 881 95 915 129
rect 975 63 1009 97
rect 1069 95 1103 129
rect 1163 63 1197 97
rect 1257 95 1291 129
rect 1351 63 1385 97
rect 1445 95 1479 129
rect 1539 127 1573 161
rect 1539 59 1573 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 129 445 163 479
rect 129 377 163 411
rect 129 309 163 343
rect 223 451 257 485
rect 223 383 257 417
rect 317 445 351 479
rect 317 377 351 411
rect 317 309 351 343
rect 411 451 445 485
rect 411 383 445 417
rect 505 429 539 463
rect 505 334 539 368
rect 599 451 633 485
rect 599 383 633 417
rect 693 429 727 463
rect 693 334 727 368
rect 787 451 821 485
rect 787 383 821 417
rect 881 429 915 463
rect 881 334 915 368
rect 975 451 1009 485
rect 975 383 1009 417
rect 1069 429 1103 463
rect 1069 334 1103 368
rect 1163 451 1197 485
rect 1163 383 1197 417
rect 1257 429 1291 463
rect 1257 334 1291 368
rect 1351 451 1385 485
rect 1351 383 1385 417
rect 1445 429 1479 463
rect 1445 334 1479 368
rect 1539 451 1573 485
rect 1539 383 1573 417
rect 1539 315 1573 349
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 457 497 493 523
rect 551 497 587 523
rect 645 497 681 523
rect 739 497 775 523
rect 833 497 869 523
rect 927 497 963 523
rect 1021 497 1057 523
rect 1115 497 1151 523
rect 1209 497 1245 523
rect 1303 497 1339 523
rect 1397 497 1433 523
rect 1491 497 1527 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 457 282 493 297
rect 551 282 587 297
rect 645 282 681 297
rect 739 282 775 297
rect 833 282 869 297
rect 927 282 963 297
rect 1021 282 1057 297
rect 1115 282 1151 297
rect 1209 282 1245 297
rect 1303 282 1339 297
rect 1397 282 1433 297
rect 1491 282 1527 297
rect 79 261 119 282
rect 27 259 119 261
rect 173 259 213 282
rect 267 259 307 282
rect 361 259 401 282
rect 27 249 401 259
rect 27 215 60 249
rect 94 215 138 249
rect 172 215 216 249
rect 250 215 284 249
rect 318 215 401 249
rect 27 205 401 215
rect 27 203 119 205
rect 89 177 119 203
rect 183 177 213 205
rect 277 177 307 205
rect 371 177 401 205
rect 455 259 495 282
rect 549 259 589 282
rect 643 259 683 282
rect 737 259 777 282
rect 831 259 871 282
rect 925 259 965 282
rect 1019 259 1059 282
rect 1113 259 1153 282
rect 1207 259 1247 282
rect 1301 259 1341 282
rect 1395 259 1435 282
rect 1489 259 1529 282
rect 455 249 1529 259
rect 455 215 475 249
rect 509 215 553 249
rect 587 215 631 249
rect 665 215 709 249
rect 743 215 787 249
rect 821 215 855 249
rect 889 215 933 249
rect 967 215 1529 249
rect 455 205 1529 215
rect 455 177 485 205
rect 549 177 579 205
rect 643 177 673 205
rect 737 177 767 205
rect 831 177 861 205
rect 925 177 955 205
rect 1019 177 1049 205
rect 1113 177 1143 205
rect 1207 177 1237 205
rect 1301 177 1331 205
rect 1395 177 1425 205
rect 1499 177 1529 205
rect 89 21 119 47
rect 183 21 213 47
rect 277 21 307 47
rect 371 21 401 47
rect 455 21 485 47
rect 549 21 579 47
rect 643 21 673 47
rect 737 21 767 47
rect 831 21 861 47
rect 925 21 955 47
rect 1019 21 1049 47
rect 1113 21 1143 47
rect 1207 21 1237 47
rect 1301 21 1331 47
rect 1395 21 1425 47
rect 1499 21 1529 47
<< polycont >>
rect 60 215 94 249
rect 138 215 172 249
rect 216 215 250 249
rect 284 215 318 249
rect 475 215 509 249
rect 553 215 587 249
rect 631 215 665 249
rect 709 215 743 249
rect 787 215 821 249
rect 855 215 889 249
rect 933 215 967 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 35 485 69 527
rect 35 417 69 451
rect 35 367 69 383
rect 103 479 179 493
rect 103 445 129 479
rect 163 445 179 479
rect 103 411 179 445
rect 103 377 129 411
rect 163 377 179 411
rect 103 343 179 377
rect 223 485 257 527
rect 223 417 257 451
rect 223 367 257 383
rect 291 479 367 493
rect 291 445 317 479
rect 351 445 367 479
rect 291 411 367 445
rect 291 377 317 411
rect 351 377 367 411
rect 103 309 129 343
rect 163 323 179 343
rect 291 343 367 377
rect 411 485 445 527
rect 411 417 445 451
rect 411 367 445 383
rect 505 463 539 493
rect 505 368 539 429
rect 291 323 317 343
rect 163 309 317 323
rect 351 323 367 343
rect 573 485 649 527
rect 573 451 599 485
rect 633 451 649 485
rect 573 417 649 451
rect 573 383 599 417
rect 633 383 649 417
rect 573 367 649 383
rect 693 463 727 493
rect 693 368 727 429
rect 505 323 539 334
rect 761 485 837 527
rect 761 451 787 485
rect 821 451 837 485
rect 761 417 837 451
rect 761 383 787 417
rect 821 383 837 417
rect 761 367 837 383
rect 881 463 915 493
rect 881 368 915 429
rect 693 323 727 334
rect 949 485 1025 527
rect 949 451 975 485
rect 1009 451 1025 485
rect 949 417 1025 451
rect 949 383 975 417
rect 1009 383 1025 417
rect 949 367 1025 383
rect 1069 463 1103 493
rect 1069 368 1103 429
rect 881 323 915 334
rect 1137 485 1213 527
rect 1137 451 1163 485
rect 1197 451 1213 485
rect 1137 417 1213 451
rect 1137 383 1163 417
rect 1197 383 1213 417
rect 1137 367 1213 383
rect 1257 463 1291 493
rect 1257 368 1291 429
rect 1069 323 1103 334
rect 1325 485 1401 527
rect 1325 451 1351 485
rect 1385 451 1401 485
rect 1325 417 1401 451
rect 1325 383 1351 417
rect 1385 383 1401 417
rect 1325 367 1401 383
rect 1445 463 1479 493
rect 1445 368 1479 429
rect 1257 323 1291 334
rect 1445 323 1479 334
rect 351 309 443 323
rect 103 289 443 309
rect 505 289 1479 323
rect 1513 485 1589 527
rect 1513 451 1539 485
rect 1573 451 1589 485
rect 1513 417 1589 451
rect 1513 383 1539 417
rect 1573 383 1589 417
rect 1513 349 1589 383
rect 1513 315 1539 349
rect 1573 315 1589 349
rect 1513 297 1589 315
rect 27 249 362 255
rect 27 215 60 249
rect 94 215 138 249
rect 172 215 216 249
rect 250 215 284 249
rect 318 215 362 249
rect 408 249 443 289
rect 408 215 475 249
rect 509 215 553 249
rect 587 215 631 249
rect 665 215 709 249
rect 743 215 787 249
rect 821 215 855 249
rect 889 215 933 249
rect 967 215 993 249
rect 408 181 443 215
rect 1042 181 1479 289
rect 129 147 443 181
rect 505 147 1479 181
rect 129 129 163 147
rect 19 97 85 113
rect 19 63 35 97
rect 69 63 85 97
rect 19 17 85 63
rect 317 129 351 147
rect 129 51 163 95
rect 197 97 273 113
rect 197 63 223 97
rect 257 63 273 97
rect 197 17 273 63
rect 505 129 539 147
rect 317 52 351 95
rect 385 97 461 113
rect 385 63 411 97
rect 445 63 461 97
rect 385 17 461 63
rect 693 129 727 147
rect 505 51 539 95
rect 573 97 649 113
rect 573 63 599 97
rect 633 63 649 97
rect 573 17 649 63
rect 881 129 915 147
rect 693 51 727 95
rect 761 97 837 113
rect 761 63 787 97
rect 821 63 837 97
rect 761 17 837 63
rect 1069 129 1103 147
rect 881 51 915 95
rect 949 97 1025 113
rect 949 63 975 97
rect 1009 63 1025 97
rect 949 17 1025 63
rect 1257 129 1291 147
rect 1069 51 1103 95
rect 1137 97 1213 113
rect 1137 63 1163 97
rect 1197 63 1213 97
rect 1137 17 1213 63
rect 1445 129 1479 147
rect 1257 51 1291 95
rect 1325 97 1401 113
rect 1325 63 1351 97
rect 1385 63 1401 97
rect 1325 17 1401 63
rect 1445 51 1479 95
rect 1513 161 1589 177
rect 1513 127 1539 161
rect 1573 127 1589 161
rect 1513 93 1589 127
rect 1513 59 1539 93
rect 1573 59 1589 93
rect 1513 17 1589 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
<< metal1 >>
rect 0 561 1656 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 0 496 1656 527
rect 0 17 1656 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
rect 0 -48 1656 -17
<< labels >>
flabel corelocali s 304 221 338 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 1052 153 1086 187 0 FreeSans 200 0 0 0 X
port 6 nsew
flabel corelocali s 1052 221 1086 255 0 FreeSans 200 0 0 0 X
port 6 nsew
flabel corelocali s 215 221 249 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 124 -17 158 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel corelocali s 124 527 158 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew
flabel corelocali s 1052 289 1086 323 0 FreeSans 200 0 0 0 X
port 6 nsew
flabel corelocali s 124 221 158 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 39 221 73 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel nwell s 124 527 158 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew
flabel pwell s 124 -17 158 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew
flabel metal1 s 124 -17 158 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 124 527 158 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 1656 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1639512
string GDS_START 1627650
<< end >>
