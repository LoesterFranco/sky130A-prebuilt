magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 2054 704
<< pwell >>
rect 0 0 2016 49
<< scnmos >>
rect 84 84 114 232
rect 170 84 200 232
rect 256 84 286 232
rect 342 84 372 232
rect 540 74 570 222
rect 626 74 656 222
rect 712 74 742 222
rect 798 74 828 222
rect 884 74 914 222
rect 970 74 1000 222
rect 1056 74 1086 222
rect 1142 74 1172 222
rect 1242 74 1272 222
rect 1356 74 1386 222
rect 1442 74 1472 222
rect 1542 74 1572 222
rect 1628 74 1658 222
rect 1716 74 1746 222
rect 1816 74 1846 222
rect 1902 74 1932 222
<< pmoshvt >>
rect 86 368 116 592
rect 176 368 206 592
rect 283 368 313 592
rect 378 368 408 592
rect 478 368 508 592
rect 568 368 598 592
rect 678 368 708 592
rect 768 368 798 592
rect 858 368 888 592
rect 948 368 978 592
rect 1048 368 1078 592
rect 1148 368 1178 592
rect 1258 368 1288 592
rect 1359 368 1389 592
rect 1449 368 1479 592
rect 1539 368 1569 592
rect 1629 368 1659 592
rect 1719 368 1749 592
rect 1809 368 1839 592
rect 1899 368 1929 592
<< ndiff >>
rect 27 220 84 232
rect 27 186 39 220
rect 73 186 84 220
rect 27 130 84 186
rect 27 96 39 130
rect 73 96 84 130
rect 27 84 84 96
rect 114 221 170 232
rect 114 187 125 221
rect 159 187 170 221
rect 114 153 170 187
rect 114 119 125 153
rect 159 119 170 153
rect 114 84 170 119
rect 200 149 256 232
rect 200 115 211 149
rect 245 115 256 149
rect 200 84 256 115
rect 286 221 342 232
rect 286 187 297 221
rect 331 187 342 221
rect 286 153 342 187
rect 286 119 297 153
rect 331 119 342 153
rect 286 84 342 119
rect 372 220 429 232
rect 372 186 383 220
rect 417 186 429 220
rect 372 130 429 186
rect 372 96 383 130
rect 417 96 429 130
rect 372 84 429 96
rect 483 120 540 222
rect 483 86 495 120
rect 529 86 540 120
rect 483 74 540 86
rect 570 207 626 222
rect 570 173 581 207
rect 615 173 626 207
rect 570 74 626 173
rect 656 136 712 222
rect 656 102 667 136
rect 701 102 712 136
rect 656 74 712 102
rect 742 207 798 222
rect 742 173 753 207
rect 787 173 798 207
rect 742 74 798 173
rect 828 120 884 222
rect 828 86 839 120
rect 873 86 884 120
rect 828 74 884 86
rect 914 195 970 222
rect 914 161 925 195
rect 959 161 970 195
rect 914 74 970 161
rect 1000 120 1056 222
rect 1000 86 1011 120
rect 1045 86 1056 120
rect 1000 74 1056 86
rect 1086 199 1142 222
rect 1086 165 1097 199
rect 1131 165 1142 199
rect 1086 74 1142 165
rect 1172 202 1242 222
rect 1172 168 1197 202
rect 1231 168 1242 202
rect 1172 120 1242 168
rect 1172 86 1197 120
rect 1231 86 1242 120
rect 1172 74 1242 86
rect 1272 116 1356 222
rect 1272 82 1297 116
rect 1331 82 1356 116
rect 1272 74 1356 82
rect 1386 144 1442 222
rect 1386 110 1397 144
rect 1431 110 1442 144
rect 1386 74 1442 110
rect 1472 116 1542 222
rect 1472 82 1483 116
rect 1517 82 1542 116
rect 1472 74 1542 82
rect 1572 144 1628 222
rect 1572 110 1583 144
rect 1617 110 1628 144
rect 1572 74 1628 110
rect 1658 116 1716 222
rect 1658 82 1670 116
rect 1704 82 1716 116
rect 1658 74 1716 82
rect 1746 202 1816 222
rect 1746 168 1771 202
rect 1805 168 1816 202
rect 1746 120 1816 168
rect 1746 86 1771 120
rect 1805 86 1816 120
rect 1746 74 1816 86
rect 1846 127 1902 222
rect 1846 93 1857 127
rect 1891 93 1902 127
rect 1846 74 1902 93
rect 1932 202 1989 222
rect 1932 168 1943 202
rect 1977 168 1989 202
rect 1932 120 1989 168
rect 1932 86 1943 120
rect 1977 86 1989 120
rect 1932 74 1989 86
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 510 86 546
rect 27 476 39 510
rect 73 476 86 510
rect 27 440 86 476
rect 27 406 39 440
rect 73 406 86 440
rect 27 368 86 406
rect 116 580 176 592
rect 116 546 129 580
rect 163 546 176 580
rect 116 510 176 546
rect 116 476 129 510
rect 163 476 176 510
rect 116 440 176 476
rect 116 406 129 440
rect 163 406 176 440
rect 116 368 176 406
rect 206 580 283 592
rect 206 546 229 580
rect 263 546 283 580
rect 206 508 283 546
rect 206 474 229 508
rect 263 474 283 508
rect 206 368 283 474
rect 313 580 378 592
rect 313 546 331 580
rect 365 546 378 580
rect 313 497 378 546
rect 313 463 331 497
rect 365 463 378 497
rect 313 414 378 463
rect 313 380 331 414
rect 365 380 378 414
rect 313 368 378 380
rect 408 580 478 592
rect 408 546 421 580
rect 455 546 478 580
rect 408 512 478 546
rect 408 478 421 512
rect 455 478 478 512
rect 408 368 478 478
rect 508 580 568 592
rect 508 546 521 580
rect 555 546 568 580
rect 508 512 568 546
rect 508 478 521 512
rect 555 478 568 512
rect 508 368 568 478
rect 598 580 678 592
rect 598 546 621 580
rect 655 546 678 580
rect 598 368 678 546
rect 708 580 768 592
rect 708 546 721 580
rect 755 546 768 580
rect 708 512 768 546
rect 708 478 721 512
rect 755 478 768 512
rect 708 368 768 478
rect 798 531 858 592
rect 798 497 811 531
rect 845 497 858 531
rect 798 444 858 497
rect 798 410 811 444
rect 845 410 858 444
rect 798 368 858 410
rect 888 580 948 592
rect 888 546 901 580
rect 935 546 948 580
rect 888 512 948 546
rect 888 478 901 512
rect 935 478 948 512
rect 888 368 948 478
rect 978 531 1048 592
rect 978 497 1001 531
rect 1035 497 1048 531
rect 978 444 1048 497
rect 978 410 1001 444
rect 1035 410 1048 444
rect 978 368 1048 410
rect 1078 580 1148 592
rect 1078 546 1101 580
rect 1135 546 1148 580
rect 1078 512 1148 546
rect 1078 478 1101 512
rect 1135 478 1148 512
rect 1078 368 1148 478
rect 1178 580 1258 592
rect 1178 546 1201 580
rect 1235 546 1258 580
rect 1178 512 1258 546
rect 1178 478 1201 512
rect 1235 478 1258 512
rect 1178 368 1258 478
rect 1288 580 1359 592
rect 1288 546 1301 580
rect 1335 546 1359 580
rect 1288 368 1359 546
rect 1389 531 1449 592
rect 1389 497 1402 531
rect 1436 497 1449 531
rect 1389 440 1449 497
rect 1389 406 1402 440
rect 1436 406 1449 440
rect 1389 368 1449 406
rect 1479 580 1539 592
rect 1479 546 1492 580
rect 1526 546 1539 580
rect 1479 508 1539 546
rect 1479 474 1492 508
rect 1526 474 1539 508
rect 1479 368 1539 474
rect 1569 531 1629 592
rect 1569 497 1582 531
rect 1616 497 1629 531
rect 1569 440 1629 497
rect 1569 406 1582 440
rect 1616 406 1629 440
rect 1569 368 1629 406
rect 1659 580 1719 592
rect 1659 546 1672 580
rect 1706 546 1719 580
rect 1659 510 1719 546
rect 1659 476 1672 510
rect 1706 476 1719 510
rect 1659 440 1719 476
rect 1659 406 1672 440
rect 1706 406 1719 440
rect 1659 368 1719 406
rect 1749 580 1809 592
rect 1749 546 1762 580
rect 1796 546 1809 580
rect 1749 508 1809 546
rect 1749 474 1762 508
rect 1796 474 1809 508
rect 1749 368 1809 474
rect 1839 580 1899 592
rect 1839 546 1852 580
rect 1886 546 1899 580
rect 1839 510 1899 546
rect 1839 476 1852 510
rect 1886 476 1899 510
rect 1839 440 1899 476
rect 1839 406 1852 440
rect 1886 406 1899 440
rect 1839 368 1899 406
rect 1929 580 1988 592
rect 1929 546 1942 580
rect 1976 546 1988 580
rect 1929 510 1988 546
rect 1929 476 1942 510
rect 1976 476 1988 510
rect 1929 440 1988 476
rect 1929 406 1942 440
rect 1976 406 1988 440
rect 1929 368 1988 406
<< ndiffc >>
rect 39 186 73 220
rect 39 96 73 130
rect 125 187 159 221
rect 125 119 159 153
rect 211 115 245 149
rect 297 187 331 221
rect 297 119 331 153
rect 383 186 417 220
rect 383 96 417 130
rect 495 86 529 120
rect 581 173 615 207
rect 667 102 701 136
rect 753 173 787 207
rect 839 86 873 120
rect 925 161 959 195
rect 1011 86 1045 120
rect 1097 165 1131 199
rect 1197 168 1231 202
rect 1197 86 1231 120
rect 1297 82 1331 116
rect 1397 110 1431 144
rect 1483 82 1517 116
rect 1583 110 1617 144
rect 1670 82 1704 116
rect 1771 168 1805 202
rect 1771 86 1805 120
rect 1857 93 1891 127
rect 1943 168 1977 202
rect 1943 86 1977 120
<< pdiffc >>
rect 39 546 73 580
rect 39 476 73 510
rect 39 406 73 440
rect 129 546 163 580
rect 129 476 163 510
rect 129 406 163 440
rect 229 546 263 580
rect 229 474 263 508
rect 331 546 365 580
rect 331 463 365 497
rect 331 380 365 414
rect 421 546 455 580
rect 421 478 455 512
rect 521 546 555 580
rect 521 478 555 512
rect 621 546 655 580
rect 721 546 755 580
rect 721 478 755 512
rect 811 497 845 531
rect 811 410 845 444
rect 901 546 935 580
rect 901 478 935 512
rect 1001 497 1035 531
rect 1001 410 1035 444
rect 1101 546 1135 580
rect 1101 478 1135 512
rect 1201 546 1235 580
rect 1201 478 1235 512
rect 1301 546 1335 580
rect 1402 497 1436 531
rect 1402 406 1436 440
rect 1492 546 1526 580
rect 1492 474 1526 508
rect 1582 497 1616 531
rect 1582 406 1616 440
rect 1672 546 1706 580
rect 1672 476 1706 510
rect 1672 406 1706 440
rect 1762 546 1796 580
rect 1762 474 1796 508
rect 1852 546 1886 580
rect 1852 476 1886 510
rect 1852 406 1886 440
rect 1942 546 1976 580
rect 1942 476 1976 510
rect 1942 406 1976 440
<< poly >>
rect 86 592 116 618
rect 176 592 206 618
rect 283 592 313 618
rect 378 592 408 618
rect 478 592 508 618
rect 568 592 598 618
rect 678 592 708 618
rect 768 592 798 618
rect 858 592 888 618
rect 948 592 978 618
rect 1048 592 1078 618
rect 1148 592 1178 618
rect 1258 592 1288 618
rect 1359 592 1389 618
rect 1449 592 1479 618
rect 1539 592 1569 618
rect 1629 592 1659 618
rect 1719 592 1749 618
rect 1809 592 1839 618
rect 1899 592 1929 618
rect 86 353 116 368
rect 176 353 206 368
rect 283 353 313 368
rect 378 353 408 368
rect 478 353 508 368
rect 568 353 598 368
rect 678 353 708 368
rect 768 353 798 368
rect 858 353 888 368
rect 948 353 978 368
rect 1048 353 1078 368
rect 1148 353 1178 368
rect 1258 353 1288 368
rect 1359 353 1389 368
rect 1449 353 1479 368
rect 1539 353 1569 368
rect 1629 353 1659 368
rect 1719 353 1749 368
rect 1809 353 1839 368
rect 1899 353 1929 368
rect 83 336 119 353
rect 173 336 209 353
rect 280 336 316 353
rect 375 336 411 353
rect 79 320 411 336
rect 79 286 95 320
rect 129 286 163 320
rect 197 286 231 320
rect 265 306 411 320
rect 475 336 511 353
rect 565 336 601 353
rect 675 336 711 353
rect 475 320 711 336
rect 265 286 372 306
rect 79 270 372 286
rect 475 286 525 320
rect 559 286 593 320
rect 627 286 661 320
rect 695 286 711 320
rect 765 345 801 353
rect 855 345 891 353
rect 765 315 891 345
rect 475 270 711 286
rect 84 232 114 270
rect 170 232 200 270
rect 256 232 286 270
rect 342 232 372 270
rect 540 222 570 270
rect 626 267 711 270
rect 798 310 891 315
rect 945 310 981 353
rect 1045 310 1081 353
rect 1145 336 1181 353
rect 1134 320 1200 336
rect 798 294 1086 310
rect 626 237 742 267
rect 626 222 656 237
rect 712 222 742 237
rect 798 260 853 294
rect 887 260 921 294
rect 955 260 989 294
rect 1023 260 1086 294
rect 1134 286 1150 320
rect 1184 286 1200 320
rect 1255 318 1291 353
rect 1356 336 1392 353
rect 1446 336 1482 353
rect 1536 336 1572 353
rect 1626 336 1662 353
rect 1356 320 1662 336
rect 1134 270 1200 286
rect 1242 302 1308 318
rect 798 244 1086 260
rect 798 222 828 244
rect 884 222 914 244
rect 970 222 1000 244
rect 1056 222 1086 244
rect 1142 222 1172 270
rect 1242 268 1258 302
rect 1292 268 1308 302
rect 1242 252 1308 268
rect 1356 286 1385 320
rect 1419 286 1453 320
rect 1487 286 1521 320
rect 1555 306 1662 320
rect 1716 318 1752 353
rect 1806 318 1842 353
rect 1896 318 1932 353
rect 1555 286 1658 306
rect 1356 270 1658 286
rect 1242 222 1272 252
rect 1356 222 1386 270
rect 1442 222 1472 270
rect 1542 222 1572 270
rect 1628 222 1658 270
rect 1716 302 1932 318
rect 1716 268 1732 302
rect 1766 268 1800 302
rect 1834 268 1868 302
rect 1902 268 1932 302
rect 1716 252 1932 268
rect 1716 222 1746 252
rect 1816 222 1846 252
rect 1902 222 1932 252
rect 84 58 114 84
rect 170 58 200 84
rect 256 58 286 84
rect 342 58 372 84
rect 540 48 570 74
rect 626 48 656 74
rect 712 48 742 74
rect 798 48 828 74
rect 884 48 914 74
rect 970 48 1000 74
rect 1056 48 1086 74
rect 1142 48 1172 74
rect 1242 48 1272 74
rect 1356 48 1386 74
rect 1442 48 1472 74
rect 1542 48 1572 74
rect 1628 48 1658 74
rect 1716 48 1746 74
rect 1816 48 1846 74
rect 1902 48 1932 74
<< polycont >>
rect 95 286 129 320
rect 163 286 197 320
rect 231 286 265 320
rect 525 286 559 320
rect 593 286 627 320
rect 661 286 695 320
rect 853 260 887 294
rect 921 260 955 294
rect 989 260 1023 294
rect 1150 286 1184 320
rect 1258 268 1292 302
rect 1385 286 1419 320
rect 1453 286 1487 320
rect 1521 286 1555 320
rect 1732 268 1766 302
rect 1800 268 1834 302
rect 1868 268 1902 302
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 23 580 73 649
rect 23 546 39 580
rect 23 510 73 546
rect 23 476 39 510
rect 23 440 73 476
rect 23 406 39 440
rect 23 390 73 406
rect 113 580 179 596
rect 113 546 129 580
rect 163 546 179 580
rect 113 510 179 546
rect 113 476 129 510
rect 163 476 179 510
rect 113 440 179 476
rect 213 580 279 649
rect 213 546 229 580
rect 263 546 279 580
rect 213 508 279 546
rect 213 474 229 508
rect 263 474 279 508
rect 213 458 279 474
rect 315 580 365 596
rect 315 546 331 580
rect 315 497 365 546
rect 315 463 331 497
rect 405 580 471 649
rect 405 546 421 580
rect 455 546 471 580
rect 405 512 471 546
rect 405 478 421 512
rect 455 478 471 512
rect 505 580 571 596
rect 505 546 521 580
rect 555 546 571 580
rect 605 580 671 649
rect 605 546 621 580
rect 655 546 671 580
rect 705 581 1151 615
rect 705 580 771 581
rect 705 546 721 580
rect 755 546 771 580
rect 885 580 951 581
rect 505 512 571 546
rect 705 512 771 546
rect 505 478 521 512
rect 555 478 721 512
rect 755 478 771 512
rect 811 531 845 547
rect 113 406 129 440
rect 163 424 179 440
rect 315 444 365 463
rect 811 444 845 497
rect 885 546 901 580
rect 935 546 951 580
rect 1085 580 1151 581
rect 885 512 951 546
rect 885 478 901 512
rect 935 478 951 512
rect 985 531 1051 547
rect 985 497 1001 531
rect 1035 497 1051 531
rect 985 444 1051 497
rect 1085 546 1101 580
rect 1135 546 1151 580
rect 1085 512 1151 546
rect 1085 478 1101 512
rect 1135 478 1151 512
rect 1185 580 1251 649
rect 1185 546 1201 580
rect 1235 546 1251 580
rect 1185 512 1251 546
rect 1285 581 1706 615
rect 1285 580 1352 581
rect 1285 546 1301 580
rect 1335 546 1352 580
rect 1492 580 1526 581
rect 1285 530 1335 546
rect 1386 531 1452 547
rect 1185 478 1201 512
rect 1235 478 1251 512
rect 1386 504 1402 531
rect 1369 497 1402 504
rect 1436 497 1452 531
rect 1369 444 1452 497
rect 1672 580 1706 581
rect 1492 508 1526 546
rect 1492 458 1526 474
rect 1566 531 1632 547
rect 1566 497 1582 531
rect 1616 497 1632 531
rect 315 424 811 444
rect 163 414 811 424
rect 163 406 331 414
rect 113 390 331 406
rect 315 380 331 390
rect 365 410 811 414
rect 845 410 1001 444
rect 1035 440 1452 444
rect 1035 410 1402 440
rect 1369 406 1402 410
rect 1436 424 1452 440
rect 1566 440 1632 497
rect 1566 424 1582 440
rect 1436 406 1582 424
rect 1616 406 1632 440
rect 1369 390 1632 406
rect 1672 510 1706 546
rect 1672 440 1706 476
rect 1746 580 1796 649
rect 1746 546 1762 580
rect 1746 508 1796 546
rect 1746 474 1762 508
rect 1746 458 1796 474
rect 1836 580 1902 596
rect 1836 546 1852 580
rect 1886 546 1902 580
rect 1836 510 1902 546
rect 1836 476 1852 510
rect 1886 476 1902 510
rect 1836 440 1902 476
rect 1836 424 1852 440
rect 1706 406 1852 424
rect 1886 406 1902 440
rect 1672 390 1902 406
rect 1942 580 1992 649
rect 1976 546 1992 580
rect 1942 510 1992 546
rect 1976 476 1992 510
rect 1942 440 1992 476
rect 1976 406 1992 440
rect 1942 390 1992 406
rect 315 364 365 380
rect 25 320 281 356
rect 25 286 95 320
rect 129 286 163 320
rect 197 286 231 320
rect 265 286 281 320
rect 25 270 281 286
rect 315 236 349 364
rect 509 342 1200 376
rect 509 320 711 342
rect 509 286 525 320
rect 559 286 593 320
rect 627 286 661 320
rect 695 286 711 320
rect 1081 320 1200 342
rect 509 270 711 286
rect 837 294 1039 308
rect 837 260 853 294
rect 887 260 921 294
rect 955 260 989 294
rect 1023 260 1039 294
rect 1081 286 1150 320
rect 1184 286 1200 320
rect 1369 320 1607 356
rect 1081 270 1200 286
rect 1242 302 1315 318
rect 837 236 1039 260
rect 1242 268 1258 302
rect 1292 268 1315 302
rect 1369 286 1385 320
rect 1419 286 1453 320
rect 1487 286 1521 320
rect 1555 286 1607 320
rect 1657 302 1991 356
rect 1242 252 1315 268
rect 1657 268 1732 302
rect 1766 268 1800 302
rect 1834 268 1868 302
rect 1902 268 1991 302
rect 1657 252 1991 268
rect 23 220 75 236
rect 23 186 39 220
rect 73 186 75 220
rect 23 130 75 186
rect 23 96 39 130
rect 73 96 75 130
rect 109 221 349 236
rect 109 187 125 221
rect 159 202 297 221
rect 159 187 175 202
rect 109 153 175 187
rect 281 187 297 202
rect 331 187 349 221
rect 109 119 125 153
rect 159 119 175 153
rect 209 149 247 168
rect 23 85 75 96
rect 209 115 211 149
rect 245 115 247 149
rect 281 153 349 187
rect 281 119 297 153
rect 331 119 349 153
rect 383 220 803 236
rect 417 207 803 220
rect 1281 218 1691 252
rect 417 186 581 207
rect 383 173 581 186
rect 615 202 753 207
rect 615 173 631 202
rect 383 154 631 173
rect 737 173 753 202
rect 787 202 803 207
rect 1081 202 1147 210
rect 787 199 1147 202
rect 787 195 1097 199
rect 787 173 925 195
rect 383 130 433 154
rect 209 85 247 115
rect 417 96 433 130
rect 667 136 701 168
rect 737 161 925 173
rect 959 165 1097 195
rect 1131 165 1147 199
rect 959 161 1147 165
rect 737 154 1147 161
rect 1181 202 1247 218
rect 1181 168 1197 202
rect 1231 184 1247 202
rect 1755 202 1993 218
rect 1755 184 1771 202
rect 1231 168 1771 184
rect 1805 184 1943 202
rect 383 85 433 96
rect 23 51 433 85
rect 479 86 495 120
rect 529 102 667 120
rect 1181 150 1805 168
rect 1977 168 1993 202
rect 1181 120 1247 150
rect 701 102 839 120
rect 529 86 839 102
rect 873 86 1011 120
rect 1045 86 1197 120
rect 1231 86 1247 120
rect 1381 144 1431 150
rect 479 70 1247 86
rect 1281 82 1297 116
rect 1331 82 1347 116
rect 1281 17 1347 82
rect 1381 110 1397 144
rect 1567 144 1617 150
rect 1381 70 1431 110
rect 1467 82 1483 116
rect 1517 82 1533 116
rect 1467 17 1533 82
rect 1567 110 1583 144
rect 1755 120 1805 150
rect 1567 70 1617 110
rect 1653 82 1670 116
rect 1704 82 1721 116
rect 1653 17 1721 82
rect 1755 86 1771 120
rect 1755 70 1805 86
rect 1841 127 1907 150
rect 1841 93 1857 127
rect 1891 93 1907 127
rect 1841 17 1907 93
rect 1943 120 1993 168
rect 1977 86 1993 120
rect 1943 70 1993 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o221ai_4
flabel pwell s 0 0 2016 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 0 617 2016 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 0 617 2016 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 2016 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 1087 316 1121 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 1375 316 1409 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 1471 316 1505 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 1567 316 1601 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 C1
port 5 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 C1
port 5 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 C1
port 5 nsew
flabel corelocali s 895 242 929 276 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 991 242 1025 276 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 1375 464 1409 498 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 1663 316 1697 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 1759 316 1793 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 1855 316 1889 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 1951 316 1985 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 2016 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1473812
string GDS_START 1457730
<< end >>
