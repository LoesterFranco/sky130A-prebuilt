magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 17 296 85 493
rect 17 165 68 296
rect 206 199 276 265
rect 17 90 89 165
rect 446 215 570 257
rect 604 215 714 257
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 119 441 201 527
rect 354 443 420 527
rect 456 407 517 493
rect 129 373 517 407
rect 129 265 172 373
rect 215 305 344 339
rect 102 199 172 265
rect 310 165 344 305
rect 135 17 169 165
rect 242 131 344 165
rect 378 291 517 373
rect 634 307 710 527
rect 242 90 276 131
rect 378 51 412 291
rect 456 147 713 181
rect 456 51 522 147
rect 566 17 600 111
rect 647 54 713 147
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel locali s 604 215 714 257 6 A1
port 1 nsew signal input
rlabel locali s 446 215 570 257 6 A2
port 2 nsew signal input
rlabel locali s 206 199 276 265 6 B1_N
port 3 nsew signal input
rlabel locali s 17 296 85 493 6 X
port 4 nsew signal output
rlabel locali s 17 165 68 296 6 X
port 4 nsew signal output
rlabel locali s 17 90 89 165 6 X
port 4 nsew signal output
rlabel metal1 s 0 -48 736 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 736 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 994076
string GDS_START 987844
<< end >>
