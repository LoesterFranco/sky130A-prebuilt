magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 92 561
rect 0 -17 92 17
<< metal1 >>
rect 0 496 92 592
rect 0 -48 92 48
<< labels >>
rlabel locali s 0 -17 92 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 92 48 8 VGND
port 1 nsew ground bidirectional abutment
rlabel locali s 0 527 92 561 6 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 0 496 92 592 6 VPWR
port 2 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE SPACER
string FIXED_BBOX 0 0 92 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2107444
string GDS_START 2106216
<< end >>
