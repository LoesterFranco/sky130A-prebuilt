magic
tech sky130A
magscale 1 2
timestamp 1601050082
<< locali >>
rect 121 332 359 367
rect 121 298 547 332
rect 313 162 420 253
rect 481 252 547 298
rect 589 288 655 430
rect 768 252 927 318
rect 768 236 839 252
rect 2617 388 2683 596
rect 2813 388 2856 596
rect 2617 354 2951 388
rect 2817 260 2951 354
rect 2817 220 2851 260
rect 2507 186 2851 220
rect 2507 70 2573 186
rect 2817 70 2851 186
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 2976 683
rect 23 435 89 596
rect 123 469 313 649
rect 421 503 487 596
rect 619 537 685 649
rect 723 518 799 596
rect 941 550 1007 649
rect 723 516 929 518
rect 1149 516 1215 551
rect 723 503 1215 516
rect 421 484 1215 503
rect 1249 498 1377 551
rect 1434 532 1504 649
rect 1545 498 1611 551
rect 1249 485 1611 498
rect 421 469 799 484
rect 916 482 1215 484
rect 689 466 799 469
rect 23 401 541 435
rect 23 253 57 401
rect 475 366 541 401
rect 23 187 228 253
rect 23 70 73 187
rect 689 218 723 466
rect 1165 451 1215 482
rect 1343 464 1611 485
rect 757 424 833 432
rect 757 390 799 424
rect 757 366 833 390
rect 867 398 903 450
rect 867 364 995 398
rect 1031 383 1131 448
rect 1165 417 1309 451
rect 1031 382 1241 383
rect 961 348 995 364
rect 961 282 1056 348
rect 1090 317 1241 382
rect 961 218 995 282
rect 1090 248 1124 317
rect 1275 283 1309 417
rect 513 184 723 218
rect 873 184 995 218
rect 1039 184 1124 248
rect 513 169 547 184
rect 109 17 175 153
rect 221 85 287 128
rect 454 119 547 169
rect 873 150 907 184
rect 645 85 700 150
rect 221 51 700 85
rect 734 17 799 150
rect 833 110 907 150
rect 943 17 1009 150
rect 1043 100 1124 184
rect 1158 249 1309 283
rect 1158 134 1198 249
rect 1343 215 1377 464
rect 1232 181 1377 215
rect 1411 218 1465 389
rect 1499 315 1533 464
rect 1567 424 1629 430
rect 1601 390 1629 424
rect 1567 364 1629 390
rect 1673 349 1707 649
rect 1747 315 1813 551
rect 1854 510 2059 576
rect 1499 252 1663 315
rect 1697 281 1813 315
rect 1849 413 1991 476
rect 1697 218 1731 281
rect 1849 247 1883 413
rect 2025 379 2059 510
rect 2093 504 2159 649
rect 2200 504 2266 596
rect 1411 184 1731 218
rect 1232 134 1294 181
rect 1411 116 1620 150
rect 1654 119 1731 184
rect 1765 181 1883 247
rect 1917 345 2059 379
rect 2117 424 2183 430
rect 2117 390 2143 424
rect 2177 390 2183 424
rect 2117 364 2183 390
rect 1917 211 1951 345
rect 2232 311 2266 504
rect 2330 364 2380 649
rect 2420 320 2486 540
rect 2527 364 2577 649
rect 2723 422 2773 649
rect 2894 422 2953 649
rect 2003 277 2317 311
rect 2003 245 2069 277
rect 2183 211 2249 243
rect 1411 100 1445 116
rect 1043 66 1445 100
rect 1586 85 1620 116
rect 1765 85 1799 181
rect 1917 177 2249 211
rect 1917 147 1951 177
rect 1486 17 1552 82
rect 1586 51 1799 85
rect 1833 81 1951 147
rect 2283 143 2317 277
rect 2028 17 2116 136
rect 2208 77 2317 143
rect 2351 254 2770 320
rect 2351 70 2385 254
rect 2421 17 2473 220
rect 2607 17 2781 152
rect 2887 17 2953 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 2976 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 799 390 833 424
rect 1567 390 1601 424
rect 2143 390 2177 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
<< metal1 >>
rect 0 683 2976 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 2976 683
rect 0 617 2976 649
rect 787 424 845 430
rect 787 390 799 424
rect 833 421 845 424
rect 1555 424 1613 430
rect 1555 421 1567 424
rect 833 393 1567 421
rect 833 390 845 393
rect 787 384 845 390
rect 1555 390 1567 393
rect 1601 421 1613 424
rect 2131 424 2189 430
rect 2131 421 2143 424
rect 1601 393 2143 421
rect 1601 390 1613 393
rect 1555 384 1613 390
rect 2131 390 2143 393
rect 2177 390 2189 424
rect 2131 384 2189 390
rect 0 17 2976 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 2976 17
rect 0 -49 2976 -17
<< labels >>
rlabel locali s 313 162 420 253 6 D
port 1 nsew signal input
rlabel locali s 2817 260 2951 354 6 Q
port 2 nsew signal output
rlabel locali s 2817 220 2851 260 6 Q
port 2 nsew signal output
rlabel locali s 2817 70 2851 186 6 Q
port 2 nsew signal output
rlabel locali s 2813 388 2856 596 6 Q
port 2 nsew signal output
rlabel locali s 2617 388 2683 596 6 Q
port 2 nsew signal output
rlabel locali s 2617 354 2951 388 6 Q
port 2 nsew signal output
rlabel locali s 2507 186 2851 220 6 Q
port 2 nsew signal output
rlabel locali s 2507 70 2573 186 6 Q
port 2 nsew signal output
rlabel metal1 s 2131 421 2189 430 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 2131 384 2189 393 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 1555 421 1613 430 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 1555 384 1613 393 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 787 421 845 430 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 787 393 2189 421 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 787 384 845 393 6 RESET_B
port 3 nsew signal input
rlabel locali s 589 288 655 430 6 SCD
port 4 nsew signal input
rlabel locali s 481 252 547 298 6 SCE
port 5 nsew signal input
rlabel locali s 121 332 359 367 6 SCE
port 5 nsew signal input
rlabel locali s 121 298 547 332 6 SCE
port 5 nsew signal input
rlabel locali s 768 252 927 318 6 CLK
port 6 nsew clock input
rlabel locali s 768 236 839 252 6 CLK
port 6 nsew clock input
rlabel metal1 s 0 -49 2976 49 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 617 2976 715 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2976 666
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 206836
string GDS_START 184766
<< end >>
