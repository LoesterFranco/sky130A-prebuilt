magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 276 561
rect 105 375 171 527
rect 205 312 259 493
rect 21 197 89 271
rect 223 152 259 312
rect 105 17 171 93
rect 207 51 259 152
rect 0 -17 276 17
<< obsli1 >>
rect 33 341 69 493
rect 33 307 168 341
rect 134 278 168 307
rect 134 212 189 278
rect 134 161 168 212
rect 35 127 168 161
rect 35 51 69 127
<< metal1 >>
rect 0 496 276 592
rect 0 -48 276 48
<< labels >>
rlabel locali s 21 197 89 271 6 A
port 1 nsew signal input
rlabel locali s 223 152 259 312 6 X
port 2 nsew signal output
rlabel locali s 207 51 259 152 6 X
port 2 nsew signal output
rlabel locali s 205 312 259 493 6 X
port 2 nsew signal output
rlabel locali s 105 17 171 93 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 0 -17 276 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 276 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 105 375 171 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 0 527 276 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 496 276 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 276 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3004728
string GDS_START 3000820
<< end >>
