magic
tech sky130A
magscale 1 2
timestamp 1601050056
<< nwell >>
rect -38 332 1574 704
<< pwell >>
rect 0 0 1536 49
<< scpmos >>
rect 83 387 119 587
rect 173 387 209 587
rect 264 387 300 587
rect 363 387 399 587
rect 453 387 489 587
rect 543 387 579 587
rect 730 387 766 587
rect 825 387 861 587
rect 920 387 956 587
rect 1020 387 1056 587
rect 1121 368 1157 592
rect 1226 368 1262 592
rect 1316 368 1352 592
rect 1417 368 1453 592
<< nmoslvt >>
rect 84 125 114 253
rect 170 125 200 253
rect 270 125 300 253
rect 363 125 393 253
rect 456 125 486 253
rect 543 125 573 253
rect 747 119 777 247
rect 834 119 864 247
rect 920 119 950 247
rect 1006 119 1036 247
rect 1121 99 1151 247
rect 1208 99 1238 247
rect 1322 99 1352 247
rect 1408 99 1438 247
<< ndiff >>
rect 27 239 84 253
rect 27 205 39 239
rect 73 205 84 239
rect 27 171 84 205
rect 27 137 39 171
rect 73 137 84 171
rect 27 125 84 137
rect 114 239 170 253
rect 114 205 125 239
rect 159 205 170 239
rect 114 171 170 205
rect 114 137 125 171
rect 159 137 170 171
rect 114 125 170 137
rect 200 171 270 253
rect 200 137 211 171
rect 245 137 270 171
rect 200 125 270 137
rect 300 241 363 253
rect 300 207 311 241
rect 345 207 363 241
rect 300 171 363 207
rect 300 137 311 171
rect 345 137 363 171
rect 300 125 363 137
rect 393 171 456 253
rect 393 137 411 171
rect 445 137 456 171
rect 393 125 456 137
rect 486 245 543 253
rect 486 211 497 245
rect 531 211 543 245
rect 486 177 543 211
rect 486 143 497 177
rect 531 143 543 177
rect 486 125 543 143
rect 573 171 630 253
rect 573 137 584 171
rect 618 137 630 171
rect 573 125 630 137
rect 690 168 747 247
rect 690 134 702 168
rect 736 134 747 168
rect 690 119 747 134
rect 777 235 834 247
rect 777 201 788 235
rect 822 201 834 235
rect 777 167 834 201
rect 777 133 788 167
rect 822 133 834 167
rect 777 119 834 133
rect 864 166 920 247
rect 864 132 875 166
rect 909 132 920 166
rect 864 119 920 132
rect 950 236 1006 247
rect 950 202 961 236
rect 995 202 1006 236
rect 950 168 1006 202
rect 950 134 961 168
rect 995 134 1006 168
rect 950 119 1006 134
rect 1036 228 1121 247
rect 1036 194 1063 228
rect 1097 194 1121 228
rect 1036 145 1121 194
rect 1036 119 1063 145
rect 1051 111 1063 119
rect 1097 111 1121 145
rect 1051 99 1121 111
rect 1151 220 1208 247
rect 1151 186 1163 220
rect 1197 186 1208 220
rect 1151 145 1208 186
rect 1151 111 1163 145
rect 1197 111 1208 145
rect 1151 99 1208 111
rect 1238 145 1322 247
rect 1238 111 1256 145
rect 1290 111 1322 145
rect 1238 99 1322 111
rect 1352 220 1408 247
rect 1352 186 1363 220
rect 1397 186 1408 220
rect 1352 145 1408 186
rect 1352 111 1363 145
rect 1397 111 1408 145
rect 1352 99 1408 111
rect 1438 235 1509 247
rect 1438 201 1463 235
rect 1497 201 1509 235
rect 1438 145 1509 201
rect 1438 111 1463 145
rect 1497 111 1509 145
rect 1438 99 1509 111
<< pdiff >>
rect 1071 587 1121 592
rect 27 576 83 587
rect 27 542 39 576
rect 73 542 83 576
rect 27 508 83 542
rect 27 474 39 508
rect 73 474 83 508
rect 27 440 83 474
rect 27 406 39 440
rect 73 406 83 440
rect 27 387 83 406
rect 119 575 173 587
rect 119 541 129 575
rect 163 541 173 575
rect 119 507 173 541
rect 119 473 129 507
rect 163 473 173 507
rect 119 439 173 473
rect 119 405 129 439
rect 163 405 173 439
rect 119 387 173 405
rect 209 576 264 587
rect 209 542 219 576
rect 253 542 264 576
rect 209 508 264 542
rect 209 474 219 508
rect 253 474 264 508
rect 209 387 264 474
rect 300 575 363 587
rect 300 541 319 575
rect 353 541 363 575
rect 300 500 363 541
rect 300 466 319 500
rect 353 466 363 500
rect 300 387 363 466
rect 399 531 453 587
rect 399 497 409 531
rect 443 497 453 531
rect 399 440 453 497
rect 399 406 409 440
rect 443 406 453 440
rect 399 387 453 406
rect 489 575 543 587
rect 489 541 499 575
rect 533 541 543 575
rect 489 500 543 541
rect 489 466 499 500
rect 533 466 543 500
rect 489 387 543 466
rect 579 576 730 587
rect 579 542 589 576
rect 623 542 686 576
rect 720 542 730 576
rect 579 508 730 542
rect 579 474 589 508
rect 623 474 686 508
rect 720 474 730 508
rect 579 387 730 474
rect 766 575 825 587
rect 766 541 776 575
rect 810 541 825 575
rect 766 500 825 541
rect 766 466 776 500
rect 810 466 825 500
rect 766 387 825 466
rect 861 543 920 587
rect 861 509 876 543
rect 910 509 920 543
rect 861 440 920 509
rect 861 406 876 440
rect 910 406 920 440
rect 861 387 920 406
rect 956 575 1020 587
rect 956 541 976 575
rect 1010 541 1020 575
rect 956 500 1020 541
rect 956 466 976 500
rect 1010 466 1020 500
rect 956 387 1020 466
rect 1056 575 1121 587
rect 1056 541 1076 575
rect 1110 541 1121 575
rect 1056 500 1121 541
rect 1056 466 1076 500
rect 1110 466 1121 500
rect 1056 387 1121 466
rect 1071 368 1121 387
rect 1157 580 1226 592
rect 1157 546 1182 580
rect 1216 546 1226 580
rect 1157 500 1226 546
rect 1157 466 1182 500
rect 1216 466 1226 500
rect 1157 420 1226 466
rect 1157 386 1182 420
rect 1216 386 1226 420
rect 1157 368 1226 386
rect 1262 580 1316 592
rect 1262 546 1272 580
rect 1306 546 1316 580
rect 1262 488 1316 546
rect 1262 454 1272 488
rect 1306 454 1316 488
rect 1262 368 1316 454
rect 1352 580 1417 592
rect 1352 546 1373 580
rect 1407 546 1417 580
rect 1352 497 1417 546
rect 1352 463 1373 497
rect 1407 463 1417 497
rect 1352 414 1417 463
rect 1352 380 1373 414
rect 1407 380 1417 414
rect 1352 368 1417 380
rect 1453 580 1509 592
rect 1453 546 1463 580
rect 1497 546 1509 580
rect 1453 510 1509 546
rect 1453 476 1463 510
rect 1497 476 1509 510
rect 1453 440 1509 476
rect 1453 406 1463 440
rect 1497 406 1509 440
rect 1453 368 1509 406
<< ndiffc >>
rect 39 205 73 239
rect 39 137 73 171
rect 125 205 159 239
rect 125 137 159 171
rect 211 137 245 171
rect 311 207 345 241
rect 311 137 345 171
rect 411 137 445 171
rect 497 211 531 245
rect 497 143 531 177
rect 584 137 618 171
rect 702 134 736 168
rect 788 201 822 235
rect 788 133 822 167
rect 875 132 909 166
rect 961 202 995 236
rect 961 134 995 168
rect 1063 194 1097 228
rect 1063 111 1097 145
rect 1163 186 1197 220
rect 1163 111 1197 145
rect 1256 111 1290 145
rect 1363 186 1397 220
rect 1363 111 1397 145
rect 1463 201 1497 235
rect 1463 111 1497 145
<< pdiffc >>
rect 39 542 73 576
rect 39 474 73 508
rect 39 406 73 440
rect 129 541 163 575
rect 129 473 163 507
rect 129 405 163 439
rect 219 542 253 576
rect 219 474 253 508
rect 319 541 353 575
rect 319 466 353 500
rect 409 497 443 531
rect 409 406 443 440
rect 499 541 533 575
rect 499 466 533 500
rect 589 542 623 576
rect 686 542 720 576
rect 589 474 623 508
rect 686 474 720 508
rect 776 541 810 575
rect 776 466 810 500
rect 876 509 910 543
rect 876 406 910 440
rect 976 541 1010 575
rect 976 466 1010 500
rect 1076 541 1110 575
rect 1076 466 1110 500
rect 1182 546 1216 580
rect 1182 466 1216 500
rect 1182 386 1216 420
rect 1272 546 1306 580
rect 1272 454 1306 488
rect 1373 546 1407 580
rect 1373 463 1407 497
rect 1373 380 1407 414
rect 1463 546 1497 580
rect 1463 476 1497 510
rect 1463 406 1497 440
<< poly >>
rect 83 587 119 613
rect 173 587 209 613
rect 264 587 300 613
rect 363 587 399 613
rect 453 587 489 613
rect 543 587 579 613
rect 730 587 766 613
rect 825 587 861 613
rect 920 587 956 613
rect 1020 587 1056 613
rect 1121 592 1157 618
rect 1226 592 1262 618
rect 1316 592 1352 618
rect 1417 592 1453 618
rect 83 355 119 387
rect 173 355 209 387
rect 44 339 209 355
rect 44 305 60 339
rect 94 305 128 339
rect 162 305 209 339
rect 44 289 209 305
rect 84 253 114 289
rect 170 253 200 289
rect 264 268 300 387
rect 270 253 300 268
rect 363 355 399 387
rect 453 355 489 387
rect 363 339 489 355
rect 363 305 439 339
rect 473 305 489 339
rect 363 289 489 305
rect 543 319 579 387
rect 621 339 687 355
rect 621 319 637 339
rect 543 305 637 319
rect 671 305 687 339
rect 543 289 687 305
rect 730 292 766 387
rect 825 355 861 387
rect 920 355 956 387
rect 825 339 956 355
rect 825 305 889 339
rect 923 319 956 339
rect 1020 336 1056 387
rect 1121 336 1157 368
rect 1226 336 1262 368
rect 1316 336 1352 368
rect 998 320 1064 336
rect 923 305 950 319
rect 363 253 393 289
rect 456 253 486 289
rect 543 253 573 289
rect 84 99 114 125
rect 170 99 200 125
rect 270 51 300 125
rect 363 99 393 125
rect 456 99 486 125
rect 543 99 573 125
rect 645 51 675 289
rect 730 262 777 292
rect 825 289 950 305
rect 747 247 777 262
rect 834 247 864 289
rect 920 247 950 289
rect 998 286 1014 320
rect 1048 286 1064 320
rect 998 270 1064 286
rect 1121 325 1352 336
rect 1417 325 1453 368
rect 1121 320 1453 325
rect 1121 286 1137 320
rect 1171 286 1205 320
rect 1239 286 1273 320
rect 1307 286 1453 320
rect 1121 270 1453 286
rect 1006 247 1036 270
rect 1121 247 1151 270
rect 1208 247 1238 270
rect 1322 247 1352 270
rect 1408 247 1438 270
rect 270 21 675 51
rect 747 51 777 119
rect 834 93 864 119
rect 920 93 950 119
rect 1006 51 1036 119
rect 1121 73 1151 99
rect 1208 73 1238 99
rect 1322 73 1352 99
rect 1408 73 1438 99
rect 747 21 1036 51
<< polycont >>
rect 60 305 94 339
rect 128 305 162 339
rect 439 305 473 339
rect 637 305 671 339
rect 889 305 923 339
rect 1014 286 1048 320
rect 1137 286 1171 320
rect 1205 286 1239 320
rect 1273 286 1307 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 23 576 73 649
rect 23 542 39 576
rect 23 508 73 542
rect 23 474 39 508
rect 23 440 73 474
rect 23 406 39 440
rect 23 390 73 406
rect 113 575 179 591
rect 113 541 129 575
rect 163 541 179 575
rect 113 507 179 541
rect 113 473 129 507
rect 163 473 179 507
rect 113 439 179 473
rect 219 576 269 649
rect 253 542 269 576
rect 219 508 269 542
rect 253 474 269 508
rect 219 458 269 474
rect 303 581 549 615
rect 303 575 369 581
rect 303 541 319 575
rect 353 541 369 575
rect 483 575 549 581
rect 303 500 369 541
rect 303 466 319 500
rect 353 466 369 500
rect 303 458 369 466
rect 409 531 443 547
rect 113 405 129 439
rect 163 424 179 439
rect 409 440 443 497
rect 483 541 499 575
rect 533 541 549 575
rect 483 500 549 541
rect 483 466 499 500
rect 533 466 549 500
rect 483 458 549 466
rect 583 576 726 649
rect 583 542 589 576
rect 623 542 686 576
rect 720 542 726 576
rect 583 508 726 542
rect 583 474 589 508
rect 623 474 686 508
rect 720 474 726 508
rect 583 458 726 474
rect 760 581 1026 615
rect 760 575 826 581
rect 760 541 776 575
rect 810 541 826 575
rect 960 575 1026 581
rect 760 500 826 541
rect 760 466 776 500
rect 810 466 826 500
rect 760 458 826 466
rect 860 543 926 547
rect 860 509 876 543
rect 910 509 926 543
rect 163 406 409 424
rect 860 440 926 509
rect 960 541 976 575
rect 1010 541 1026 575
rect 960 500 1026 541
rect 960 466 976 500
rect 1010 466 1026 500
rect 960 458 1026 466
rect 1060 575 1126 649
rect 1060 541 1076 575
rect 1110 541 1126 575
rect 1060 500 1126 541
rect 1060 466 1076 500
rect 1110 466 1126 500
rect 1060 458 1126 466
rect 1166 580 1232 596
rect 1166 546 1182 580
rect 1216 546 1232 580
rect 1166 500 1232 546
rect 1166 466 1182 500
rect 1216 466 1232 500
rect 860 424 876 440
rect 443 406 876 424
rect 910 424 926 440
rect 910 406 1132 424
rect 163 405 1132 406
rect 113 390 1132 405
rect 25 339 178 356
rect 25 305 60 339
rect 94 305 128 339
rect 162 305 178 339
rect 25 289 178 305
rect 212 255 246 390
rect 409 339 551 356
rect 409 305 439 339
rect 473 305 551 339
rect 409 289 551 305
rect 601 339 839 356
rect 601 305 637 339
rect 671 305 839 339
rect 601 289 839 305
rect 873 339 939 356
rect 873 305 889 339
rect 923 305 939 339
rect 873 289 939 305
rect 985 320 1064 356
rect 985 286 1014 320
rect 1048 286 1064 320
rect 985 270 1064 286
rect 1098 336 1132 390
rect 1166 420 1232 466
rect 1272 580 1322 649
rect 1306 546 1322 580
rect 1272 488 1322 546
rect 1306 454 1322 488
rect 1272 438 1322 454
rect 1357 580 1423 596
rect 1357 546 1373 580
rect 1407 546 1423 580
rect 1357 497 1423 546
rect 1357 463 1373 497
rect 1407 463 1423 497
rect 1166 386 1182 420
rect 1216 404 1232 420
rect 1357 414 1423 463
rect 1357 404 1373 414
rect 1216 386 1373 404
rect 1166 380 1373 386
rect 1407 380 1423 414
rect 1463 580 1513 649
rect 1497 546 1513 580
rect 1463 510 1513 546
rect 1497 476 1513 510
rect 1463 440 1513 476
rect 1497 406 1513 440
rect 1463 390 1513 406
rect 1166 370 1423 380
rect 1357 356 1423 370
rect 1098 320 1323 336
rect 1098 286 1137 320
rect 1171 286 1205 320
rect 1239 286 1273 320
rect 1307 286 1323 320
rect 1098 270 1323 286
rect 1357 310 1511 356
rect 23 239 73 255
rect 23 205 39 239
rect 23 171 73 205
rect 23 137 39 171
rect 23 87 73 137
rect 109 239 246 255
rect 109 205 125 239
rect 159 221 246 239
rect 295 255 361 257
rect 295 245 823 255
rect 295 241 497 245
rect 109 171 159 205
rect 295 207 311 241
rect 345 211 497 241
rect 531 236 823 245
rect 1357 236 1413 310
rect 531 235 961 236
rect 531 221 788 235
rect 531 211 548 221
rect 345 207 548 211
rect 295 205 548 207
rect 109 137 125 171
rect 109 121 159 137
rect 195 171 261 187
rect 195 137 211 171
rect 245 137 261 171
rect 195 87 261 137
rect 295 171 361 205
rect 495 177 534 205
rect 822 202 961 235
rect 995 202 1011 236
rect 822 201 823 202
rect 295 137 311 171
rect 345 137 361 171
rect 295 121 361 137
rect 395 137 411 171
rect 445 137 461 171
rect 395 91 461 137
rect 495 143 497 177
rect 531 143 534 177
rect 495 127 534 143
rect 568 137 584 171
rect 618 137 634 171
rect 568 91 634 137
rect 395 87 634 91
rect 23 57 634 87
rect 686 168 752 187
rect 686 134 702 168
rect 736 134 752 168
rect 23 53 461 57
rect 686 17 752 134
rect 788 167 823 201
rect 961 168 1011 202
rect 822 133 823 167
rect 788 117 823 133
rect 859 166 925 168
rect 859 132 875 166
rect 909 132 925 166
rect 859 17 925 132
rect 995 134 1011 168
rect 961 118 1011 134
rect 1047 228 1113 236
rect 1047 194 1063 228
rect 1097 194 1113 228
rect 1047 145 1113 194
rect 1047 111 1063 145
rect 1097 111 1113 145
rect 1047 17 1113 111
rect 1147 220 1413 236
rect 1147 186 1163 220
rect 1197 202 1363 220
rect 1147 145 1197 186
rect 1347 186 1363 202
rect 1397 186 1413 220
rect 1147 111 1163 145
rect 1147 95 1197 111
rect 1233 145 1313 161
rect 1233 111 1256 145
rect 1290 111 1313 145
rect 1233 17 1313 111
rect 1347 145 1413 186
rect 1347 111 1363 145
rect 1397 111 1413 145
rect 1347 95 1413 111
rect 1447 235 1513 251
rect 1447 201 1463 235
rect 1497 201 1513 235
rect 1447 145 1513 201
rect 1447 111 1463 145
rect 1497 111 1513 145
rect 1447 17 1513 111
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
flabel pwell s 0 0 1536 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 0 617 1536 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
rlabel comment s 0 0 0 0 4 o221a_4
flabel metal1 s 0 617 1536 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 1536 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 1471 316 1505 350 0 FreeSans 340 0 0 0 X
port 10 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 C1
port 5 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 C1
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 1536 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1155656
string GDS_START 1143054
<< end >>
