magic
tech sky130A
magscale 1 2
timestamp 1601050056
<< nwell >>
rect -38 332 806 704
<< pwell >>
rect 0 0 768 49
<< scpmos >>
rect 83 368 119 592
rect 184 368 220 592
rect 313 392 349 592
rect 397 392 433 592
rect 511 392 547 592
rect 619 392 655 592
<< nmoslvt >>
rect 98 74 128 222
rect 184 74 214 222
rect 298 74 328 222
rect 397 74 427 222
rect 511 74 541 222
rect 640 74 670 222
<< ndiff >>
rect 27 210 98 222
rect 27 176 39 210
rect 73 176 98 210
rect 27 120 98 176
rect 27 86 39 120
rect 73 86 98 120
rect 27 74 98 86
rect 128 210 184 222
rect 128 176 139 210
rect 173 176 184 210
rect 128 120 184 176
rect 128 86 139 120
rect 173 86 184 120
rect 128 74 184 86
rect 214 210 298 222
rect 214 176 239 210
rect 273 176 298 210
rect 214 120 298 176
rect 214 86 239 120
rect 273 86 298 120
rect 214 74 298 86
rect 328 210 397 222
rect 328 176 339 210
rect 373 176 397 210
rect 328 120 397 176
rect 328 86 339 120
rect 373 86 397 120
rect 328 74 397 86
rect 427 120 511 222
rect 427 86 445 120
rect 479 86 511 120
rect 427 74 511 86
rect 541 142 640 222
rect 541 108 573 142
rect 607 108 640 142
rect 541 74 640 108
rect 670 210 741 222
rect 670 176 695 210
rect 729 176 741 210
rect 670 120 741 176
rect 670 86 695 120
rect 729 86 741 120
rect 670 74 741 86
<< pdiff >>
rect 27 573 83 592
rect 27 539 39 573
rect 73 539 83 573
rect 27 368 83 539
rect 119 414 184 592
rect 119 380 134 414
rect 168 380 184 414
rect 119 368 184 380
rect 220 580 313 592
rect 220 546 249 580
rect 283 546 313 580
rect 220 392 313 546
rect 349 392 397 592
rect 433 392 511 592
rect 547 580 619 592
rect 547 546 569 580
rect 603 546 619 580
rect 547 509 619 546
rect 547 475 569 509
rect 603 475 619 509
rect 547 438 619 475
rect 547 404 569 438
rect 603 404 619 438
rect 547 392 619 404
rect 655 580 741 592
rect 655 546 695 580
rect 729 546 741 580
rect 655 510 741 546
rect 655 476 695 510
rect 729 476 741 510
rect 655 440 741 476
rect 655 406 695 440
rect 729 406 741 440
rect 655 392 741 406
rect 220 368 270 392
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 139 176 173 210
rect 139 86 173 120
rect 239 176 273 210
rect 239 86 273 120
rect 339 176 373 210
rect 339 86 373 120
rect 445 86 479 120
rect 573 108 607 142
rect 695 176 729 210
rect 695 86 729 120
<< pdiffc >>
rect 39 539 73 573
rect 134 380 168 414
rect 249 546 283 580
rect 569 546 603 580
rect 569 475 603 509
rect 569 404 603 438
rect 695 546 729 580
rect 695 476 729 510
rect 695 406 729 440
<< poly >>
rect 83 592 119 618
rect 184 592 220 618
rect 313 592 349 618
rect 397 592 433 618
rect 511 592 547 618
rect 619 592 655 618
rect 83 330 119 368
rect 55 314 128 330
rect 55 280 71 314
rect 105 294 128 314
rect 184 294 220 368
rect 313 336 349 392
rect 105 280 220 294
rect 55 264 220 280
rect 283 320 349 336
rect 283 286 299 320
rect 333 286 349 320
rect 283 270 349 286
rect 397 360 433 392
rect 397 344 463 360
rect 397 310 413 344
rect 447 310 463 344
rect 397 294 463 310
rect 511 310 547 392
rect 619 358 655 392
rect 625 326 655 358
rect 625 310 745 326
rect 511 294 577 310
rect 98 222 128 264
rect 184 222 214 264
rect 298 222 328 270
rect 397 222 427 294
rect 511 260 527 294
rect 561 260 577 294
rect 625 276 695 310
rect 729 276 745 310
rect 625 260 745 276
rect 511 244 577 260
rect 511 222 541 244
rect 640 222 670 260
rect 98 48 128 74
rect 184 48 214 74
rect 298 48 328 74
rect 397 48 427 74
rect 511 48 541 74
rect 640 48 670 74
<< polycont >>
rect 71 280 105 314
rect 299 286 333 320
rect 413 310 447 344
rect 527 260 561 294
rect 695 276 729 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 23 573 89 649
rect 23 539 39 573
rect 73 539 89 573
rect 23 532 89 539
rect 214 580 319 649
rect 214 546 249 580
rect 283 546 319 580
rect 214 532 319 546
rect 553 580 645 596
rect 553 546 569 580
rect 603 546 645 580
rect 553 509 645 546
rect 553 498 569 509
rect 45 475 569 498
rect 603 475 645 509
rect 45 464 645 475
rect 45 330 79 464
rect 553 438 645 464
rect 113 414 190 430
rect 113 380 134 414
rect 168 380 190 414
rect 113 364 190 380
rect 45 314 121 330
rect 45 280 71 314
rect 105 280 121 314
rect 45 264 121 280
rect 155 226 189 364
rect 283 320 359 430
rect 283 286 299 320
rect 333 286 359 320
rect 397 344 463 430
rect 553 404 569 438
rect 603 404 645 438
rect 553 388 645 404
rect 679 580 745 649
rect 679 546 695 580
rect 729 546 745 580
rect 679 510 745 546
rect 679 476 695 510
rect 729 476 745 510
rect 679 440 745 476
rect 679 406 695 440
rect 729 406 745 440
rect 679 390 745 406
rect 397 310 413 344
rect 447 310 463 344
rect 397 294 463 310
rect 505 294 577 310
rect 283 270 359 286
rect 505 260 527 294
rect 561 260 577 294
rect 505 236 577 260
rect 611 226 645 388
rect 679 310 745 356
rect 679 276 695 310
rect 729 276 745 310
rect 679 260 745 276
rect 23 210 89 226
rect 23 176 39 210
rect 73 176 89 210
rect 23 120 89 176
rect 23 86 39 120
rect 73 86 89 120
rect 23 17 89 86
rect 123 210 189 226
rect 123 176 139 210
rect 173 176 189 210
rect 123 120 189 176
rect 123 86 139 120
rect 173 86 189 120
rect 123 70 189 86
rect 223 210 289 226
rect 223 176 239 210
rect 273 176 289 210
rect 223 120 289 176
rect 223 86 239 120
rect 273 86 289 120
rect 223 17 289 86
rect 323 210 389 226
rect 323 176 339 210
rect 373 188 389 210
rect 611 210 745 226
rect 611 192 695 210
rect 373 176 570 188
rect 323 158 570 176
rect 679 176 695 192
rect 729 176 745 210
rect 323 154 645 158
rect 323 120 389 154
rect 536 142 645 154
rect 323 86 339 120
rect 373 86 389 120
rect 323 70 389 86
rect 423 86 445 120
rect 479 86 502 120
rect 536 108 573 142
rect 607 108 645 142
rect 536 92 645 108
rect 679 120 745 176
rect 423 17 502 86
rect 679 86 695 120
rect 729 86 745 120
rect 679 70 745 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
rlabel comment s 0 0 0 0 4 o31a_2
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 B1
port 4 nsew
flabel corelocali s 511 242 545 276 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 415 390 449 424 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 319 390 353 424 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 127 390 161 424 0 FreeSans 340 0 0 0 X
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 768 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1341732
string GDS_START 1335094
<< end >>
