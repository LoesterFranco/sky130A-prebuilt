magic
tech sky130A
magscale 1 2
timestamp 1604502741
<< locali >>
rect 21 236 87 310
rect 121 270 225 356
rect 267 270 359 356
rect 393 270 459 356
rect 579 364 645 596
rect 601 282 645 364
rect 601 226 647 282
rect 596 70 647 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 21 424 87 572
rect 121 458 187 649
rect 221 424 287 572
rect 405 458 545 649
rect 21 390 535 424
rect 21 364 87 390
rect 501 326 535 390
rect 679 364 745 649
rect 501 260 567 326
rect 501 236 535 260
rect 121 202 535 236
rect 26 70 155 202
rect 205 134 470 168
rect 205 70 271 134
rect 305 17 355 100
rect 404 70 470 134
rect 510 17 560 168
rect 682 17 748 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel locali s 393 270 459 356 6 A1
port 1 nsew signal input
rlabel locali s 267 270 359 356 6 A2
port 2 nsew signal input
rlabel locali s 121 270 225 356 6 B1
port 3 nsew signal input
rlabel locali s 21 236 87 310 6 C1
port 4 nsew signal input
rlabel locali s 601 282 645 364 6 X
port 5 nsew signal output
rlabel locali s 601 226 647 282 6 X
port 5 nsew signal output
rlabel locali s 596 70 647 226 6 X
port 5 nsew signal output
rlabel locali s 579 364 645 596 6 X
port 5 nsew signal output
rlabel metal1 s 0 -49 768 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 768 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1720268
string GDS_START 1713180
<< end >>
