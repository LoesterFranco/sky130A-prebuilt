magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 89 93 119 177
rect 196 47 226 177
rect 280 47 310 177
<< pmoshvt >>
rect 81 297 117 381
rect 188 297 224 497
rect 282 297 318 497
<< ndiff >>
rect 27 155 89 177
rect 27 121 35 155
rect 69 121 89 155
rect 27 93 89 121
rect 119 93 196 177
rect 134 59 142 93
rect 176 59 196 93
rect 134 47 196 59
rect 226 47 280 177
rect 310 93 372 177
rect 310 59 330 93
rect 364 59 372 93
rect 310 47 372 59
<< pdiff >>
rect 134 485 188 497
rect 134 451 142 485
rect 176 451 188 485
rect 134 417 188 451
rect 134 383 142 417
rect 176 383 188 417
rect 134 381 188 383
rect 27 349 81 381
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 297 188 381
rect 224 485 282 497
rect 224 451 236 485
rect 270 451 282 485
rect 224 417 282 451
rect 224 383 236 417
rect 270 383 282 417
rect 224 297 282 383
rect 318 485 372 497
rect 318 451 330 485
rect 364 451 372 485
rect 318 297 372 451
<< ndiffc >>
rect 35 121 69 155
rect 142 59 176 93
rect 330 59 364 93
<< pdiffc >>
rect 142 451 176 485
rect 142 383 176 417
rect 35 315 69 349
rect 236 451 270 485
rect 236 383 270 417
rect 330 451 364 485
<< poly >>
rect 188 497 224 523
rect 282 497 318 523
rect 81 381 117 407
rect 81 282 117 297
rect 188 282 224 297
rect 282 282 318 297
rect 79 265 119 282
rect 186 265 226 282
rect 22 249 119 265
rect 22 215 34 249
rect 68 215 119 249
rect 22 199 119 215
rect 172 249 226 265
rect 172 215 182 249
rect 216 215 226 249
rect 172 199 226 215
rect 89 177 119 199
rect 196 177 226 199
rect 280 265 320 282
rect 280 249 334 265
rect 280 215 290 249
rect 324 215 334 249
rect 280 199 334 215
rect 280 177 310 199
rect 89 67 119 93
rect 196 21 226 47
rect 280 21 310 47
<< polycont >>
rect 34 215 68 249
rect 182 215 216 249
rect 290 215 324 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 126 485 176 527
rect 126 451 142 485
rect 126 417 176 451
rect 126 383 142 417
rect 126 367 176 383
rect 210 485 286 493
rect 210 451 236 485
rect 270 451 286 485
rect 210 417 286 451
rect 330 485 373 527
rect 364 451 373 485
rect 330 435 373 451
rect 210 383 236 417
rect 270 401 286 417
rect 270 383 438 401
rect 210 367 438 383
rect 18 349 74 365
rect 18 315 35 349
rect 69 333 74 349
rect 69 315 324 333
rect 18 299 324 315
rect 18 249 84 263
rect 18 215 34 249
rect 68 215 84 249
rect 118 249 237 263
rect 118 215 182 249
rect 216 215 237 249
rect 290 249 324 299
rect 290 181 324 215
rect 18 155 324 181
rect 18 121 35 155
rect 69 147 324 155
rect 69 121 72 147
rect 18 105 72 121
rect 364 109 438 367
rect 126 93 192 109
rect 126 59 142 93
rect 176 59 192 93
rect 126 17 192 59
rect 272 93 438 109
rect 272 59 330 93
rect 364 59 438 93
rect 272 51 438 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
flabel corelocali s 379 374 379 374 0 FreeSans 250 0 0 0 Y
port 7 nsew
flabel corelocali s 379 306 379 306 0 FreeSans 250 0 0 0 Y
port 7 nsew
flabel corelocali s 379 102 379 102 0 FreeSans 250 0 0 0 Y
port 7 nsew
flabel corelocali s 379 238 379 238 0 FreeSans 250 0 0 0 Y
port 7 nsew
flabel corelocali s 379 170 379 170 0 FreeSans 250 0 0 0 Y
port 7 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 250 0 0 0 A_N
port 1 nsew
flabel corelocali s 132 221 166 255 0 FreeSans 250 0 0 0 B
port 2 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew
rlabel comment s 0 0 0 0 4 nand2b_1
<< properties >>
string FIXED_BBOX 0 0 460 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2222346
string GDS_START 2217752
<< end >>
