magic
tech sky130A
magscale 1 2
timestamp 1604502705
<< nwell >>
rect -38 332 1862 704
<< pwell >>
rect 0 0 1824 49
<< scnmos >>
rect 84 74 114 222
rect 170 74 200 222
rect 270 74 300 222
rect 370 74 400 222
rect 470 74 500 222
rect 570 74 600 222
rect 670 74 700 222
rect 770 74 800 222
rect 856 74 886 222
rect 956 74 986 222
rect 1042 74 1072 222
rect 1128 74 1158 222
rect 1214 74 1244 222
rect 1300 74 1330 222
rect 1386 74 1416 222
rect 1486 74 1516 222
rect 1696 74 1726 222
<< pmoshvt >>
rect 85 368 115 592
rect 175 368 205 592
rect 265 368 295 592
rect 355 368 385 592
rect 445 368 475 592
rect 535 368 565 592
rect 625 368 655 592
rect 715 368 745 592
rect 805 368 835 592
rect 895 368 925 592
rect 985 368 1015 592
rect 1075 368 1105 592
rect 1165 368 1195 592
rect 1255 368 1285 592
rect 1345 368 1375 592
rect 1435 368 1465 592
rect 1710 368 1740 592
<< ndiff >>
rect 27 202 84 222
rect 27 168 39 202
rect 73 168 84 202
rect 27 127 84 168
rect 27 93 39 127
rect 73 93 84 127
rect 27 74 84 93
rect 114 173 170 222
rect 114 139 125 173
rect 159 139 170 173
rect 114 74 170 139
rect 200 127 270 222
rect 200 93 225 127
rect 259 93 270 127
rect 200 74 270 93
rect 300 173 370 222
rect 300 139 325 173
rect 359 139 370 173
rect 300 74 370 139
rect 400 127 470 222
rect 400 93 425 127
rect 459 93 470 127
rect 400 74 470 93
rect 500 173 570 222
rect 500 139 525 173
rect 559 139 570 173
rect 500 74 570 139
rect 600 127 670 222
rect 600 93 625 127
rect 659 93 670 127
rect 600 74 670 93
rect 700 169 770 222
rect 700 135 725 169
rect 759 135 770 169
rect 700 74 770 135
rect 800 210 856 222
rect 800 176 811 210
rect 845 176 856 210
rect 800 120 856 176
rect 800 86 811 120
rect 845 86 856 120
rect 800 74 856 86
rect 886 203 956 222
rect 886 169 897 203
rect 931 169 956 203
rect 886 120 956 169
rect 886 86 897 120
rect 931 86 956 120
rect 886 74 956 86
rect 986 210 1042 222
rect 986 176 997 210
rect 1031 176 1042 210
rect 986 120 1042 176
rect 986 86 997 120
rect 1031 86 1042 120
rect 986 74 1042 86
rect 1072 203 1128 222
rect 1072 169 1083 203
rect 1117 169 1128 203
rect 1072 120 1128 169
rect 1072 86 1083 120
rect 1117 86 1128 120
rect 1072 74 1128 86
rect 1158 210 1214 222
rect 1158 176 1169 210
rect 1203 176 1214 210
rect 1158 120 1214 176
rect 1158 86 1169 120
rect 1203 86 1214 120
rect 1158 74 1214 86
rect 1244 203 1300 222
rect 1244 169 1255 203
rect 1289 169 1300 203
rect 1244 120 1300 169
rect 1244 86 1255 120
rect 1289 86 1300 120
rect 1244 74 1300 86
rect 1330 210 1386 222
rect 1330 176 1341 210
rect 1375 176 1386 210
rect 1330 120 1386 176
rect 1330 86 1341 120
rect 1375 86 1386 120
rect 1330 74 1386 86
rect 1416 203 1486 222
rect 1416 169 1441 203
rect 1475 169 1486 203
rect 1416 120 1486 169
rect 1416 86 1441 120
rect 1475 86 1486 120
rect 1416 74 1486 86
rect 1516 210 1573 222
rect 1516 176 1527 210
rect 1561 176 1573 210
rect 1516 120 1573 176
rect 1516 86 1527 120
rect 1561 86 1573 120
rect 1516 74 1573 86
rect 1638 198 1696 222
rect 1638 164 1651 198
rect 1685 164 1696 198
rect 1638 120 1696 164
rect 1638 86 1651 120
rect 1685 86 1696 120
rect 1638 74 1696 86
rect 1726 186 1783 222
rect 1726 152 1737 186
rect 1771 152 1783 186
rect 1726 118 1783 152
rect 1726 84 1737 118
rect 1771 84 1783 118
rect 1726 74 1783 84
<< pdiff >>
rect 27 580 85 592
rect 27 546 38 580
rect 72 546 85 580
rect 27 497 85 546
rect 27 463 38 497
rect 72 463 85 497
rect 27 414 85 463
rect 27 380 38 414
rect 72 380 85 414
rect 27 368 85 380
rect 115 547 175 592
rect 115 513 128 547
rect 162 513 175 547
rect 115 479 175 513
rect 115 445 128 479
rect 162 445 175 479
rect 115 411 175 445
rect 115 377 128 411
rect 162 377 175 411
rect 115 368 175 377
rect 205 580 265 592
rect 205 546 218 580
rect 252 546 265 580
rect 205 462 265 546
rect 205 428 218 462
rect 252 428 265 462
rect 205 368 265 428
rect 295 547 355 592
rect 295 513 308 547
rect 342 513 355 547
rect 295 479 355 513
rect 295 445 308 479
rect 342 445 355 479
rect 295 411 355 445
rect 295 377 308 411
rect 342 377 355 411
rect 295 368 355 377
rect 385 580 445 592
rect 385 546 398 580
rect 432 546 445 580
rect 385 462 445 546
rect 385 428 398 462
rect 432 428 445 462
rect 385 368 445 428
rect 475 547 535 592
rect 475 513 488 547
rect 522 513 535 547
rect 475 479 535 513
rect 475 445 488 479
rect 522 445 535 479
rect 475 411 535 445
rect 475 377 488 411
rect 522 377 535 411
rect 475 368 535 377
rect 565 580 625 592
rect 565 546 578 580
rect 612 546 625 580
rect 565 462 625 546
rect 565 428 578 462
rect 612 428 625 462
rect 565 368 625 428
rect 655 547 715 592
rect 655 513 668 547
rect 702 513 715 547
rect 655 479 715 513
rect 655 445 668 479
rect 702 445 715 479
rect 655 411 715 445
rect 655 377 668 411
rect 702 377 715 411
rect 655 368 715 377
rect 745 580 805 592
rect 745 546 758 580
rect 792 546 805 580
rect 745 462 805 546
rect 745 428 758 462
rect 792 428 805 462
rect 745 368 805 428
rect 835 582 895 592
rect 835 548 848 582
rect 882 548 895 582
rect 835 514 895 548
rect 835 480 848 514
rect 882 480 895 514
rect 835 368 895 480
rect 925 580 985 592
rect 925 546 938 580
rect 972 546 985 580
rect 925 497 985 546
rect 925 463 938 497
rect 972 463 985 497
rect 925 414 985 463
rect 925 380 938 414
rect 972 380 985 414
rect 925 368 985 380
rect 1015 580 1075 592
rect 1015 546 1028 580
rect 1062 546 1075 580
rect 1015 504 1075 546
rect 1015 470 1028 504
rect 1062 470 1075 504
rect 1015 428 1075 470
rect 1015 394 1028 428
rect 1062 394 1075 428
rect 1015 368 1075 394
rect 1105 580 1165 592
rect 1105 546 1118 580
rect 1152 546 1165 580
rect 1105 497 1165 546
rect 1105 463 1118 497
rect 1152 463 1165 497
rect 1105 414 1165 463
rect 1105 380 1118 414
rect 1152 380 1165 414
rect 1105 368 1165 380
rect 1195 580 1255 592
rect 1195 546 1208 580
rect 1242 546 1255 580
rect 1195 504 1255 546
rect 1195 470 1208 504
rect 1242 470 1255 504
rect 1195 428 1255 470
rect 1195 394 1208 428
rect 1242 394 1255 428
rect 1195 368 1255 394
rect 1285 580 1345 592
rect 1285 546 1298 580
rect 1332 546 1345 580
rect 1285 497 1345 546
rect 1285 463 1298 497
rect 1332 463 1345 497
rect 1285 414 1345 463
rect 1285 380 1298 414
rect 1332 380 1345 414
rect 1285 368 1345 380
rect 1375 580 1435 592
rect 1375 546 1388 580
rect 1422 546 1435 580
rect 1375 504 1435 546
rect 1375 470 1388 504
rect 1422 470 1435 504
rect 1375 428 1435 470
rect 1375 394 1388 428
rect 1422 394 1435 428
rect 1375 368 1435 394
rect 1465 580 1523 592
rect 1465 546 1478 580
rect 1512 546 1523 580
rect 1465 497 1523 546
rect 1465 463 1478 497
rect 1512 463 1523 497
rect 1465 414 1523 463
rect 1465 380 1478 414
rect 1512 380 1523 414
rect 1465 368 1523 380
rect 1653 580 1710 592
rect 1653 546 1663 580
rect 1697 546 1710 580
rect 1653 497 1710 546
rect 1653 463 1663 497
rect 1697 463 1710 497
rect 1653 414 1710 463
rect 1653 380 1663 414
rect 1697 380 1710 414
rect 1653 368 1710 380
rect 1740 580 1797 592
rect 1740 546 1753 580
rect 1787 546 1797 580
rect 1740 497 1797 546
rect 1740 463 1753 497
rect 1787 463 1797 497
rect 1740 414 1797 463
rect 1740 380 1753 414
rect 1787 380 1797 414
rect 1740 368 1797 380
<< ndiffc >>
rect 39 168 73 202
rect 39 93 73 127
rect 125 139 159 173
rect 225 93 259 127
rect 325 139 359 173
rect 425 93 459 127
rect 525 139 559 173
rect 625 93 659 127
rect 725 135 759 169
rect 811 176 845 210
rect 811 86 845 120
rect 897 169 931 203
rect 897 86 931 120
rect 997 176 1031 210
rect 997 86 1031 120
rect 1083 169 1117 203
rect 1083 86 1117 120
rect 1169 176 1203 210
rect 1169 86 1203 120
rect 1255 169 1289 203
rect 1255 86 1289 120
rect 1341 176 1375 210
rect 1341 86 1375 120
rect 1441 169 1475 203
rect 1441 86 1475 120
rect 1527 176 1561 210
rect 1527 86 1561 120
rect 1651 164 1685 198
rect 1651 86 1685 120
rect 1737 152 1771 186
rect 1737 84 1771 118
<< pdiffc >>
rect 38 546 72 580
rect 38 463 72 497
rect 38 380 72 414
rect 128 513 162 547
rect 128 445 162 479
rect 128 377 162 411
rect 218 546 252 580
rect 218 428 252 462
rect 308 513 342 547
rect 308 445 342 479
rect 308 377 342 411
rect 398 546 432 580
rect 398 428 432 462
rect 488 513 522 547
rect 488 445 522 479
rect 488 377 522 411
rect 578 546 612 580
rect 578 428 612 462
rect 668 513 702 547
rect 668 445 702 479
rect 668 377 702 411
rect 758 546 792 580
rect 758 428 792 462
rect 848 548 882 582
rect 848 480 882 514
rect 938 546 972 580
rect 938 463 972 497
rect 938 380 972 414
rect 1028 546 1062 580
rect 1028 470 1062 504
rect 1028 394 1062 428
rect 1118 546 1152 580
rect 1118 463 1152 497
rect 1118 380 1152 414
rect 1208 546 1242 580
rect 1208 470 1242 504
rect 1208 394 1242 428
rect 1298 546 1332 580
rect 1298 463 1332 497
rect 1298 380 1332 414
rect 1388 546 1422 580
rect 1388 470 1422 504
rect 1388 394 1422 428
rect 1478 546 1512 580
rect 1478 463 1512 497
rect 1478 380 1512 414
rect 1663 546 1697 580
rect 1663 463 1697 497
rect 1663 380 1697 414
rect 1753 546 1787 580
rect 1753 463 1787 497
rect 1753 380 1787 414
<< poly >>
rect 85 592 115 618
rect 175 592 205 618
rect 265 592 295 618
rect 355 592 385 618
rect 445 592 475 618
rect 535 592 565 618
rect 625 592 655 618
rect 715 592 745 618
rect 805 592 835 618
rect 895 592 925 618
rect 985 592 1015 618
rect 1075 592 1105 618
rect 1165 592 1195 618
rect 1255 592 1285 618
rect 1345 592 1375 618
rect 1435 592 1465 618
rect 1555 577 1621 593
rect 1710 592 1740 618
rect 1555 543 1571 577
rect 1605 543 1621 577
rect 1555 509 1621 543
rect 1555 475 1571 509
rect 1605 475 1621 509
rect 1555 441 1621 475
rect 1555 407 1571 441
rect 1605 407 1621 441
rect 1555 373 1621 407
rect 85 353 115 368
rect 175 353 205 368
rect 265 353 295 368
rect 355 353 385 368
rect 445 353 475 368
rect 535 353 565 368
rect 625 353 655 368
rect 715 353 745 368
rect 805 353 835 368
rect 895 353 925 368
rect 985 353 1015 368
rect 1075 353 1105 368
rect 1165 353 1195 368
rect 1255 353 1285 368
rect 1345 353 1375 368
rect 1435 353 1465 368
rect 1555 353 1571 373
rect 82 310 118 353
rect 172 310 208 353
rect 262 310 298 353
rect 352 310 388 353
rect 442 310 478 353
rect 532 310 568 353
rect 622 310 658 353
rect 712 310 748 353
rect 802 339 1571 353
rect 1605 339 1621 373
rect 1710 353 1740 368
rect 802 323 1621 339
rect 1707 310 1743 353
rect 82 294 748 310
rect 82 260 98 294
rect 132 260 166 294
rect 200 260 234 294
rect 268 260 302 294
rect 336 260 370 294
rect 404 260 438 294
rect 472 260 506 294
rect 540 260 574 294
rect 608 260 642 294
rect 676 274 748 294
rect 1687 294 1753 310
rect 1687 274 1703 294
rect 676 260 800 274
rect 82 244 800 260
rect 84 222 114 244
rect 170 222 200 244
rect 270 222 300 244
rect 370 222 400 244
rect 470 222 500 244
rect 570 222 600 244
rect 670 222 700 244
rect 770 222 800 244
rect 856 260 1703 274
rect 1737 260 1753 294
rect 856 244 1753 260
rect 856 222 886 244
rect 956 222 986 244
rect 1042 222 1072 244
rect 1128 222 1158 244
rect 1214 222 1244 244
rect 1300 222 1330 244
rect 1386 222 1416 244
rect 1486 222 1516 244
rect 1696 222 1726 244
rect 84 48 114 74
rect 170 48 200 74
rect 270 48 300 74
rect 370 48 400 74
rect 470 48 500 74
rect 570 48 600 74
rect 670 48 700 74
rect 770 48 800 74
rect 856 48 886 74
rect 956 48 986 74
rect 1042 48 1072 74
rect 1128 48 1158 74
rect 1214 48 1244 74
rect 1300 48 1330 74
rect 1386 48 1416 74
rect 1486 48 1516 74
rect 1696 48 1726 74
<< polycont >>
rect 1571 543 1605 577
rect 1571 475 1605 509
rect 1571 407 1605 441
rect 1571 339 1605 373
rect 98 260 132 294
rect 166 260 200 294
rect 234 260 268 294
rect 302 260 336 294
rect 370 260 404 294
rect 438 260 472 294
rect 506 260 540 294
rect 574 260 608 294
rect 642 260 676 294
rect 1703 260 1737 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 22 581 792 615
rect 22 580 75 581
rect 22 546 38 580
rect 72 546 75 580
rect 214 580 255 581
rect 22 497 75 546
rect 22 463 38 497
rect 72 463 75 497
rect 22 414 75 463
rect 22 380 38 414
rect 72 380 75 414
rect 22 364 75 380
rect 112 513 128 547
rect 162 513 178 547
rect 112 479 178 513
rect 112 445 128 479
rect 162 445 178 479
rect 112 411 178 445
rect 214 546 218 580
rect 252 546 255 580
rect 394 580 438 581
rect 214 462 255 546
rect 214 428 218 462
rect 252 428 255 462
rect 214 412 255 428
rect 292 513 308 547
rect 342 513 358 547
rect 292 479 358 513
rect 292 445 308 479
rect 342 445 358 479
rect 112 377 128 411
rect 162 378 178 411
rect 292 411 358 445
rect 394 546 398 580
rect 432 546 438 580
rect 575 580 615 581
rect 394 462 438 546
rect 394 428 398 462
rect 432 428 438 462
rect 394 412 438 428
rect 472 513 488 547
rect 522 513 538 547
rect 472 479 538 513
rect 472 445 488 479
rect 522 445 538 479
rect 292 378 308 411
rect 162 377 308 378
rect 342 378 358 411
rect 472 411 538 445
rect 575 546 578 580
rect 612 546 615 580
rect 758 580 792 581
rect 575 462 615 546
rect 575 428 578 462
rect 612 428 615 462
rect 575 412 615 428
rect 652 513 668 547
rect 702 513 718 547
rect 652 479 718 513
rect 652 445 668 479
rect 702 445 718 479
rect 472 378 488 411
rect 342 377 488 378
rect 522 378 538 411
rect 652 411 718 445
rect 758 462 792 546
rect 832 582 898 649
rect 832 548 848 582
rect 882 548 898 582
rect 832 514 898 548
rect 832 480 848 514
rect 882 480 898 514
rect 938 580 988 596
rect 972 546 988 580
rect 938 497 988 546
rect 972 463 988 497
rect 938 446 988 463
rect 792 428 988 446
rect 758 414 988 428
rect 758 412 938 414
rect 652 378 668 411
rect 522 377 668 378
rect 702 378 718 411
rect 972 380 988 414
rect 702 377 839 378
rect 112 344 839 377
rect 741 310 839 344
rect 938 344 988 380
rect 1028 580 1062 649
rect 1028 504 1062 546
rect 1028 428 1062 470
rect 1028 378 1062 394
rect 1102 580 1152 596
rect 1102 546 1118 580
rect 1102 497 1152 546
rect 1102 463 1118 497
rect 1102 414 1152 463
rect 1102 380 1118 414
rect 1102 344 1152 380
rect 1192 580 1242 649
rect 1192 546 1208 580
rect 1192 504 1242 546
rect 1192 470 1208 504
rect 1192 428 1242 470
rect 1192 394 1208 428
rect 1192 378 1242 394
rect 1282 580 1332 596
rect 1282 546 1298 580
rect 1282 497 1332 546
rect 1282 463 1298 497
rect 1282 414 1332 463
rect 1282 380 1298 414
rect 1282 344 1332 380
rect 1372 580 1422 649
rect 1372 546 1388 580
rect 1372 504 1422 546
rect 1372 470 1388 504
rect 1372 428 1422 470
rect 1372 394 1388 428
rect 1372 378 1422 394
rect 1462 580 1512 596
rect 1647 593 1713 596
rect 1462 546 1478 580
rect 1462 497 1512 546
rect 1462 463 1478 497
rect 1462 414 1512 463
rect 1462 380 1478 414
rect 1462 344 1512 380
rect 938 310 1512 344
rect 1555 580 1713 593
rect 1555 577 1663 580
rect 1555 543 1571 577
rect 1605 546 1663 577
rect 1697 546 1713 580
rect 1605 543 1713 546
rect 1555 509 1713 543
rect 1555 475 1571 509
rect 1605 497 1713 509
rect 1605 475 1663 497
rect 1555 463 1663 475
rect 1697 463 1713 497
rect 1555 441 1713 463
rect 1555 407 1571 441
rect 1605 414 1713 441
rect 1605 407 1663 414
rect 1555 380 1663 407
rect 1697 380 1713 414
rect 1555 373 1713 380
rect 1555 339 1571 373
rect 1605 364 1713 373
rect 1753 580 1803 649
rect 1787 546 1803 580
rect 1753 497 1803 546
rect 1787 463 1803 497
rect 1753 414 1803 463
rect 1787 380 1803 414
rect 1753 364 1803 380
rect 1605 339 1645 364
rect 1555 323 1645 339
rect 82 294 692 310
rect 82 260 98 294
rect 132 260 166 294
rect 200 260 234 294
rect 268 260 302 294
rect 336 260 370 294
rect 404 260 438 294
rect 472 260 506 294
rect 540 260 574 294
rect 608 260 642 294
rect 676 260 692 294
rect 82 236 692 260
rect 741 202 775 310
rect 23 168 39 202
rect 73 168 89 202
rect 23 127 89 168
rect 23 93 39 127
rect 73 93 89 127
rect 125 173 775 202
rect 159 168 325 173
rect 159 139 175 168
rect 125 123 175 139
rect 309 139 325 168
rect 359 168 525 173
rect 359 139 375 168
rect 209 127 275 134
rect 23 85 89 93
rect 209 93 225 127
rect 259 93 275 127
rect 309 123 375 139
rect 509 139 525 168
rect 559 169 775 173
rect 559 168 725 169
rect 559 139 575 168
rect 409 127 475 134
rect 209 85 275 93
rect 409 93 425 127
rect 459 93 475 127
rect 509 123 575 139
rect 709 135 725 168
rect 759 135 775 169
rect 609 127 675 134
rect 409 85 475 93
rect 609 93 625 127
rect 659 93 675 127
rect 709 119 775 135
rect 811 242 1577 276
rect 811 210 845 242
rect 981 210 1031 242
rect 811 120 845 176
rect 609 85 675 93
rect 811 85 845 86
rect 23 51 845 85
rect 881 203 947 208
rect 881 169 897 203
rect 931 169 947 203
rect 881 120 947 169
rect 881 86 897 120
rect 931 86 947 120
rect 881 17 947 86
rect 981 176 997 210
rect 1169 210 1203 242
rect 981 120 1031 176
rect 981 86 997 120
rect 981 70 1031 86
rect 1067 203 1133 208
rect 1067 169 1083 203
rect 1117 169 1133 203
rect 1067 120 1133 169
rect 1067 86 1083 120
rect 1117 86 1133 120
rect 1067 17 1133 86
rect 1341 210 1391 242
rect 1169 120 1203 176
rect 1169 70 1203 86
rect 1239 203 1305 208
rect 1239 169 1255 203
rect 1289 169 1305 203
rect 1239 120 1305 169
rect 1239 86 1255 120
rect 1289 86 1305 120
rect 1239 17 1305 86
rect 1375 176 1391 210
rect 1527 210 1577 242
rect 1341 120 1391 176
rect 1375 86 1391 120
rect 1341 70 1391 86
rect 1425 203 1491 208
rect 1425 169 1441 203
rect 1475 169 1491 203
rect 1425 120 1491 169
rect 1425 86 1441 120
rect 1475 86 1491 120
rect 1425 17 1491 86
rect 1561 176 1577 210
rect 1527 120 1577 176
rect 1561 86 1577 120
rect 1527 70 1577 86
rect 1611 202 1645 323
rect 1687 294 1753 310
rect 1687 260 1703 294
rect 1737 282 1753 294
rect 1737 260 1799 282
rect 1687 236 1799 260
rect 1611 198 1701 202
rect 1611 164 1651 198
rect 1685 164 1701 198
rect 1611 120 1701 164
rect 1611 86 1651 120
rect 1685 86 1701 120
rect 1611 70 1701 86
rect 1735 186 1787 202
rect 1735 152 1737 186
rect 1771 152 1787 186
rect 1735 118 1787 152
rect 1735 84 1737 118
rect 1771 84 1787 118
rect 1735 17 1787 84
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
<< metal1 >>
rect 0 683 1824 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 0 617 1824 649
rect 0 17 1824 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
rect 0 -49 1824 -17
<< labels >>
rlabel comment s 0 0 0 0 4 einvp_8
flabel pwell s 0 0 1824 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 0 617 1824 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 0 617 1824 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 1824 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 Z
port 7 nsew
flabel corelocali s 1759 242 1793 276 0 FreeSans 340 0 0 0 TE
port 2 nsew
flabel corelocali s 223 242 257 276 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 319 242 353 276 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 415 242 449 276 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 511 242 545 276 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 607 242 641 276 0 FreeSans 340 0 0 0 A
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 1824 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2074716
string GDS_START 2060396
<< end >>
