magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3128 561
rect 103 427 179 527
rect 17 195 87 325
rect 311 377 377 527
rect 702 443 778 527
rect 298 205 353 337
rect 103 17 179 93
rect 387 203 451 339
rect 831 265 895 475
rect 387 153 521 203
rect 387 152 451 153
rect 311 17 361 127
rect 395 69 451 152
rect 724 17 790 89
rect 1241 441 1317 527
rect 1565 383 1631 527
rect 2104 451 2180 527
rect 2388 451 2686 527
rect 1277 17 1311 105
rect 2743 326 2819 493
rect 2949 353 3008 527
rect 2764 304 2819 326
rect 2503 219 2618 265
rect 1658 17 1735 93
rect 2082 17 2144 105
rect 2620 17 2686 161
rect 2764 143 2823 304
rect 2743 51 2823 143
rect 3052 321 3109 493
rect 3062 165 3109 321
rect 2950 17 3008 109
rect 3052 51 3109 165
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3128 17
<< obsli1 >>
rect 34 393 69 493
rect 34 391 177 393
rect 34 359 131 391
rect 165 357 177 391
rect 131 161 177 357
rect 34 127 177 161
rect 223 187 264 493
rect 477 375 553 477
rect 619 381 653 493
rect 223 153 230 187
rect 34 69 69 127
rect 223 69 264 153
rect 510 273 553 375
rect 589 349 653 381
rect 589 315 779 349
rect 510 255 655 273
rect 510 237 621 255
rect 557 221 621 237
rect 557 215 655 221
rect 745 219 779 315
rect 929 255 963 493
rect 1007 450 1183 484
rect 557 119 591 215
rect 745 159 814 219
rect 510 53 591 119
rect 625 153 814 159
rect 625 125 779 153
rect 625 61 665 125
rect 929 61 963 221
rect 997 357 1029 391
rect 1063 357 1115 391
rect 997 315 1115 357
rect 997 141 1049 315
rect 1149 281 1183 450
rect 1387 407 1421 475
rect 1217 357 1517 407
rect 1860 450 2046 484
rect 1822 391 1869 397
rect 1217 315 1277 357
rect 1389 281 1439 297
rect 1149 247 1439 281
rect 1149 239 1243 247
rect 1085 187 1165 203
rect 1085 153 1131 187
rect 1085 129 1165 153
rect 1199 93 1243 239
rect 1395 231 1439 247
rect 1483 213 1517 357
rect 1822 357 1835 391
rect 1561 323 1782 331
rect 1561 289 1743 323
rect 1777 289 1782 323
rect 1822 315 1869 357
rect 1561 283 1782 289
rect 1561 247 1627 283
rect 1927 261 1978 381
rect 1834 255 1978 261
rect 1689 213 1775 247
rect 1277 187 1359 213
rect 1277 153 1317 187
rect 1351 153 1359 187
rect 1483 179 1775 213
rect 1834 221 1835 255
rect 1869 225 1978 255
rect 2012 281 2046 450
rect 2238 417 2272 475
rect 2080 383 2686 417
rect 2080 315 2140 383
rect 2012 247 2302 281
rect 1869 221 1902 225
rect 1483 153 1531 179
rect 1277 147 1359 153
rect 1455 119 1531 153
rect 1020 53 1243 93
rect 1355 85 1421 93
rect 1570 85 1609 143
rect 1834 141 1902 221
rect 2012 93 2046 247
rect 2258 215 2302 247
rect 2131 187 2216 213
rect 2131 153 2143 187
rect 2177 153 2216 187
rect 2346 163 2383 383
rect 2131 147 2216 153
rect 2307 129 2383 163
rect 2426 323 2581 349
rect 2426 289 2433 323
rect 2467 315 2581 323
rect 2467 289 2469 315
rect 2426 185 2469 289
rect 2652 265 2686 383
rect 2853 345 2904 483
rect 2652 199 2705 265
rect 2426 151 2563 185
rect 1355 51 1609 85
rect 1883 53 2046 93
rect 2196 85 2276 93
rect 2425 85 2460 117
rect 2196 51 2460 85
rect 2523 53 2563 151
rect 2863 265 2904 345
rect 2863 199 3018 265
rect 2863 51 2904 199
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 2881 527 2915 561
rect 2973 527 3007 561
rect 3065 527 3099 561
rect 131 357 165 391
rect 230 153 264 187
rect 621 221 655 255
rect 929 221 963 255
rect 1029 357 1063 391
rect 1131 153 1165 187
rect 1835 357 1869 391
rect 1743 289 1777 323
rect 1317 153 1351 187
rect 1835 221 1869 255
rect 2143 153 2177 187
rect 2433 289 2467 323
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
rect 2881 -17 2915 17
rect 2973 -17 3007 17
rect 3065 -17 3099 17
<< metal1 >>
rect 0 561 3128 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3128 561
rect 0 496 3128 527
rect 1305 187 1363 193
rect 1305 153 1317 187
rect 1351 184 1363 187
rect 2131 187 2189 193
rect 2131 184 2143 187
rect 1351 156 2143 184
rect 1351 153 1363 156
rect 1305 147 1363 153
rect 2131 153 2143 156
rect 2177 153 2189 187
rect 2131 147 2189 153
rect 0 17 3128 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3128 17
rect 0 -48 3128 -17
<< obsm1 >>
rect 119 391 177 397
rect 119 357 131 391
rect 165 388 177 391
rect 1017 391 1075 397
rect 1017 388 1029 391
rect 165 360 1029 388
rect 165 357 177 360
rect 119 351 177 357
rect 1017 357 1029 360
rect 1063 388 1075 391
rect 1823 391 1881 397
rect 1823 388 1835 391
rect 1063 360 1835 388
rect 1063 357 1075 360
rect 1017 351 1075 357
rect 1823 357 1835 360
rect 1869 357 1881 391
rect 1823 351 1881 357
rect 1731 323 1789 329
rect 1731 289 1743 323
rect 1777 320 1789 323
rect 2421 323 2479 329
rect 2421 320 2433 323
rect 1777 292 2433 320
rect 1777 289 1789 292
rect 1731 283 1789 289
rect 2421 289 2433 292
rect 2467 289 2479 323
rect 2421 283 2479 289
rect 609 255 667 261
rect 609 221 621 255
rect 655 252 667 255
rect 917 255 975 261
rect 917 252 929 255
rect 655 224 929 252
rect 655 221 667 224
rect 609 215 667 221
rect 917 221 929 224
rect 963 221 975 255
rect 1823 255 1881 261
rect 1823 252 1835 255
rect 917 215 975 221
rect 1134 224 1835 252
rect 1134 193 1177 224
rect 1823 221 1835 224
rect 1869 221 1881 255
rect 1823 215 1881 221
rect 218 187 276 193
rect 218 153 230 187
rect 264 184 276 187
rect 1119 187 1177 193
rect 1119 184 1131 187
rect 264 156 1131 184
rect 264 153 276 156
rect 218 147 276 153
rect 1119 153 1131 156
rect 1165 153 1177 187
rect 1119 147 1177 153
<< labels >>
rlabel locali s 17 195 87 325 6 CLK
port 1 nsew signal input
rlabel locali s 831 265 895 475 6 D
port 2 nsew signal input
rlabel locali s 3062 165 3109 321 6 Q
port 3 nsew signal output
rlabel locali s 3052 321 3109 493 6 Q
port 3 nsew signal output
rlabel locali s 3052 51 3109 165 6 Q
port 3 nsew signal output
rlabel locali s 2764 304 2819 326 6 Q_N
port 4 nsew signal output
rlabel locali s 2764 143 2823 304 6 Q_N
port 4 nsew signal output
rlabel locali s 2743 326 2819 493 6 Q_N
port 4 nsew signal output
rlabel locali s 2743 51 2823 143 6 Q_N
port 4 nsew signal output
rlabel locali s 2503 219 2618 265 6 RESET_B
port 5 nsew signal input
rlabel locali s 298 205 353 337 6 SCD
port 6 nsew signal input
rlabel locali s 395 69 451 152 6 SCE
port 7 nsew signal input
rlabel locali s 387 203 451 339 6 SCE
port 7 nsew signal input
rlabel locali s 387 153 521 203 6 SCE
port 7 nsew signal input
rlabel locali s 387 152 451 153 6 SCE
port 7 nsew signal input
rlabel metal1 s 2131 184 2189 193 6 SET_B
port 8 nsew signal input
rlabel metal1 s 2131 147 2189 156 6 SET_B
port 8 nsew signal input
rlabel metal1 s 1305 184 1363 193 6 SET_B
port 8 nsew signal input
rlabel metal1 s 1305 156 2189 184 6 SET_B
port 8 nsew signal input
rlabel metal1 s 1305 147 1363 156 6 SET_B
port 8 nsew signal input
rlabel metal1 s 0 -48 3128 48 8 VGND
port 9 nsew ground bidirectional
rlabel locali s 2950 17 3008 109 6 VGND
port 9 nsew ground bidirectional
rlabel locali s 2620 17 2686 161 6 VGND
port 9 nsew ground bidirectional
rlabel locali s 2082 17 2144 105 6 VGND
port 9 nsew ground bidirectional
rlabel locali s 1658 17 1735 93 6 VGND
port 9 nsew ground bidirectional
rlabel locali s 1277 17 1311 105 6 VGND
port 9 nsew ground bidirectional
rlabel locali s 724 17 790 89 6 VGND
port 9 nsew ground bidirectional
rlabel locali s 311 17 361 127 6 VGND
port 9 nsew ground bidirectional
rlabel locali s 103 17 179 93 6 VGND
port 9 nsew ground bidirectional
rlabel locali s 0 -17 3128 17 8 VGND
port 9 nsew ground bidirectional
rlabel metal1 s 0 496 3128 592 6 VPWR
port 10 nsew power bidirectional
rlabel locali s 2949 353 3008 527 6 VPWR
port 10 nsew power bidirectional
rlabel locali s 2388 451 2686 527 6 VPWR
port 10 nsew power bidirectional
rlabel locali s 2104 451 2180 527 6 VPWR
port 10 nsew power bidirectional
rlabel locali s 1565 383 1631 527 6 VPWR
port 10 nsew power bidirectional
rlabel locali s 1241 441 1317 527 6 VPWR
port 10 nsew power bidirectional
rlabel locali s 702 443 778 527 6 VPWR
port 10 nsew power bidirectional
rlabel locali s 311 377 377 527 6 VPWR
port 10 nsew power bidirectional
rlabel locali s 103 427 179 527 6 VPWR
port 10 nsew power bidirectional
rlabel locali s 0 527 3128 561 6 VPWR
port 10 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 3128 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 146246
string GDS_START 122988
<< end >>
