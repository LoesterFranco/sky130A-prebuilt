magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 920 561
rect 23 435 75 527
rect 17 199 75 394
rect 109 342 161 493
rect 195 383 261 527
rect 295 342 333 493
rect 367 383 433 527
rect 565 342 631 425
rect 109 308 631 342
rect 737 373 803 527
rect 109 134 175 308
rect 209 215 381 273
rect 473 215 667 271
rect 712 249 891 259
rect 701 215 891 249
rect 823 153 891 215
rect 479 17 545 89
rect 651 17 717 89
rect 823 17 889 89
rect 0 -17 920 17
<< obsli1 >>
rect 479 459 703 493
rect 479 420 531 459
rect 665 339 703 459
rect 837 339 889 493
rect 665 305 889 339
rect 209 93 247 178
rect 281 127 789 169
rect 751 103 789 127
rect 209 89 433 93
rect 19 51 433 89
<< metal1 >>
rect 0 496 920 592
rect 0 -48 920 48
<< labels >>
rlabel locali s 823 153 891 215 6 A1
port 1 nsew signal input
rlabel locali s 712 249 891 259 6 A1
port 1 nsew signal input
rlabel locali s 701 215 891 249 6 A1
port 1 nsew signal input
rlabel locali s 473 215 667 271 6 A2
port 2 nsew signal input
rlabel locali s 209 215 381 273 6 B1
port 3 nsew signal input
rlabel locali s 17 199 75 394 6 C1
port 4 nsew signal input
rlabel locali s 565 342 631 425 6 Y
port 5 nsew signal output
rlabel locali s 295 342 333 493 6 Y
port 5 nsew signal output
rlabel locali s 109 342 161 493 6 Y
port 5 nsew signal output
rlabel locali s 109 308 631 342 6 Y
port 5 nsew signal output
rlabel locali s 109 134 175 308 6 Y
port 5 nsew signal output
rlabel locali s 823 17 889 89 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 651 17 717 89 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 479 17 545 89 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 920 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 920 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 737 373 803 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 367 383 433 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 195 383 261 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 23 435 75 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 920 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 920 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 920 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1315528
string GDS_START 1308132
<< end >>
