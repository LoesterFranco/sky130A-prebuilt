magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1748 561
rect 119 367 257 527
rect 199 299 257 367
rect 291 333 357 493
rect 391 367 425 527
rect 459 333 525 493
rect 559 367 593 527
rect 627 333 693 493
rect 727 367 761 527
rect 795 333 861 493
rect 895 367 1033 527
rect 1067 333 1133 493
rect 1167 367 1201 527
rect 1235 333 1301 493
rect 1335 367 1369 527
rect 1403 333 1469 493
rect 1503 367 1537 527
rect 1571 333 1637 493
rect 291 289 1637 333
rect 1671 289 1722 527
rect 22 215 88 255
rect 475 181 528 289
rect 586 215 918 255
rect 958 215 1302 255
rect 1403 215 1731 255
rect 119 17 169 109
rect 291 127 528 181
rect 1419 17 1453 109
rect 1587 17 1621 109
rect 0 -17 1748 17
<< obsli1 >>
rect 18 333 85 493
rect 18 299 161 333
rect 122 255 161 299
rect 122 215 441 255
rect 122 181 161 215
rect 18 147 161 181
rect 18 51 85 147
rect 207 93 257 181
rect 627 127 1301 181
rect 1335 147 1722 181
rect 1335 93 1385 147
rect 207 51 945 93
rect 983 51 1385 93
rect 1487 51 1553 147
rect 1655 51 1722 147
<< metal1 >>
rect 0 496 1748 592
rect 0 -48 1748 48
<< labels >>
rlabel locali s 22 215 88 255 6 A_N
port 1 nsew signal input
rlabel locali s 586 215 918 255 6 B
port 2 nsew signal input
rlabel locali s 958 215 1302 255 6 C
port 3 nsew signal input
rlabel locali s 1403 215 1731 255 6 D
port 4 nsew signal input
rlabel locali s 1571 333 1637 493 6 Y
port 5 nsew signal output
rlabel locali s 1403 333 1469 493 6 Y
port 5 nsew signal output
rlabel locali s 1235 333 1301 493 6 Y
port 5 nsew signal output
rlabel locali s 1067 333 1133 493 6 Y
port 5 nsew signal output
rlabel locali s 795 333 861 493 6 Y
port 5 nsew signal output
rlabel locali s 627 333 693 493 6 Y
port 5 nsew signal output
rlabel locali s 475 181 528 289 6 Y
port 5 nsew signal output
rlabel locali s 459 333 525 493 6 Y
port 5 nsew signal output
rlabel locali s 291 333 357 493 6 Y
port 5 nsew signal output
rlabel locali s 291 289 1637 333 6 Y
port 5 nsew signal output
rlabel locali s 291 127 528 181 6 Y
port 5 nsew signal output
rlabel locali s 1587 17 1621 109 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1419 17 1453 109 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 119 17 169 109 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 1748 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1748 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1671 289 1722 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1503 367 1537 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1335 367 1369 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1167 367 1201 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 895 367 1033 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 727 367 761 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 559 367 593 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 391 367 425 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 199 299 257 367 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 119 367 257 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 1748 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 1748 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1748 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1894594
string GDS_START 1879666
<< end >>
