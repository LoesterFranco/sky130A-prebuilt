magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 736 561
rect 103 448 169 527
rect 294 391 411 425
rect 86 199 156 339
rect 190 199 248 265
rect 131 17 165 165
rect 371 165 411 391
rect 565 326 617 482
rect 651 375 717 527
rect 523 289 617 326
rect 523 199 589 289
rect 659 255 719 341
rect 623 199 719 255
rect 371 131 617 165
rect 303 17 369 96
rect 403 60 443 131
rect 477 17 543 97
rect 577 62 617 131
rect 651 17 717 165
rect 0 -17 736 17
<< obsli1 >>
rect 17 414 69 491
rect 207 459 479 493
rect 207 414 241 459
rect 17 377 241 414
rect 17 165 52 377
rect 199 305 318 343
rect 282 265 318 305
rect 282 199 337 265
rect 282 165 318 199
rect 17 90 81 165
rect 215 131 318 165
rect 445 199 479 459
rect 215 90 249 131
<< metal1 >>
rect 0 496 736 592
rect 0 -48 736 48
<< labels >>
rlabel locali s 659 255 719 341 6 A
port 1 nsew signal input
rlabel locali s 623 199 719 255 6 A
port 1 nsew signal input
rlabel locali s 565 326 617 482 6 B
port 2 nsew signal input
rlabel locali s 523 289 617 326 6 B
port 2 nsew signal input
rlabel locali s 523 199 589 289 6 B
port 2 nsew signal input
rlabel locali s 86 199 156 339 6 C_N
port 3 nsew signal input
rlabel locali s 190 199 248 265 6 D_N
port 4 nsew signal input
rlabel locali s 577 62 617 131 6 Y
port 5 nsew signal output
rlabel locali s 403 60 443 131 6 Y
port 5 nsew signal output
rlabel locali s 371 165 411 391 6 Y
port 5 nsew signal output
rlabel locali s 371 131 617 165 6 Y
port 5 nsew signal output
rlabel locali s 294 391 411 425 6 Y
port 5 nsew signal output
rlabel locali s 651 17 717 165 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 477 17 543 97 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 303 17 369 96 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 131 17 165 165 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 736 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 736 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 651 375 717 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 103 448 169 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 736 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 736 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1197490
string GDS_START 1191130
<< end >>
