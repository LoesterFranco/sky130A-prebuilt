magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 828 561
rect 18 299 69 527
rect 103 319 165 493
rect 205 435 263 527
rect 665 435 709 527
rect 18 17 69 177
rect 103 150 137 319
rect 455 263 618 325
rect 455 256 489 263
rect 103 51 153 150
rect 363 153 489 256
rect 525 147 618 205
rect 672 151 710 325
rect 187 17 253 93
rect 580 84 618 147
rect 670 17 710 117
rect 0 -17 828 17
<< obsli1 >>
rect 297 451 559 485
rect 297 401 331 451
rect 743 401 810 493
rect 199 367 331 401
rect 365 367 810 401
rect 199 265 233 367
rect 365 333 399 367
rect 171 199 233 265
rect 267 299 399 333
rect 267 199 301 299
rect 199 161 233 199
rect 199 127 321 161
rect 287 93 321 127
rect 287 59 546 93
rect 744 51 810 367
<< metal1 >>
rect 0 496 828 592
rect 0 -48 828 48
<< labels >>
rlabel locali s 455 263 618 325 6 A0
port 1 nsew signal input
rlabel locali s 455 256 489 263 6 A0
port 1 nsew signal input
rlabel locali s 363 153 489 256 6 A0
port 1 nsew signal input
rlabel locali s 580 84 618 147 6 A1
port 2 nsew signal input
rlabel locali s 525 147 618 205 6 A1
port 2 nsew signal input
rlabel locali s 672 151 710 325 6 S
port 3 nsew signal input
rlabel locali s 103 319 165 493 6 X
port 4 nsew signal output
rlabel locali s 103 150 137 319 6 X
port 4 nsew signal output
rlabel locali s 103 51 153 150 6 X
port 4 nsew signal output
rlabel locali s 670 17 710 117 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 187 17 253 93 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 18 17 69 177 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 828 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 828 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 665 435 709 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 205 435 263 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 18 299 69 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 828 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 828 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1650730
string GDS_START 1643540
<< end >>
