magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 736 561
rect 120 360 186 527
rect 17 215 112 258
rect 426 360 509 527
rect 543 305 630 493
rect 664 325 719 527
rect 543 284 636 305
rect 602 189 636 284
rect 117 17 183 113
rect 593 156 636 189
rect 593 128 630 156
rect 433 17 507 113
rect 541 54 630 128
rect 664 17 719 129
rect 0 -17 736 17
<< obsli1 >>
rect 17 326 86 493
rect 222 360 288 493
rect 17 292 211 326
rect 146 181 211 292
rect 17 147 211 181
rect 254 251 288 360
rect 326 326 392 493
rect 326 292 509 326
rect 254 215 441 251
rect 475 249 509 292
rect 475 215 568 249
rect 17 54 83 147
rect 254 120 288 215
rect 475 181 509 215
rect 232 54 288 120
rect 326 147 509 181
rect 326 54 392 147
<< metal1 >>
rect 0 496 736 592
rect 0 -48 736 48
<< labels >>
rlabel locali s 17 215 112 258 6 A
port 1 nsew signal input
rlabel locali s 602 189 636 284 6 X
port 2 nsew signal output
rlabel locali s 593 156 636 189 6 X
port 2 nsew signal output
rlabel locali s 593 128 630 156 6 X
port 2 nsew signal output
rlabel locali s 543 305 630 493 6 X
port 2 nsew signal output
rlabel locali s 543 284 636 305 6 X
port 2 nsew signal output
rlabel locali s 541 54 630 128 6 X
port 2 nsew signal output
rlabel locali s 664 17 719 129 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 433 17 507 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 117 17 183 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 0 -17 736 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 736 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 664 325 719 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 426 360 509 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 120 360 186 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 0 527 736 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 496 736 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3135986
string GDS_START 3129876
<< end >>
