magic
tech sky130A
magscale 1 2
timestamp 1604502697
<< nwell >>
rect -38 261 2338 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 79 47 109 177
rect 173 47 203 177
rect 267 47 297 177
rect 361 47 391 177
rect 455 47 485 177
rect 559 47 589 177
rect 643 47 673 177
rect 737 47 767 177
rect 831 47 861 177
rect 925 47 955 177
rect 1019 47 1049 177
rect 1113 47 1143 177
rect 1207 47 1237 177
rect 1301 47 1331 177
rect 1395 47 1425 177
rect 1489 47 1519 177
rect 1583 47 1613 177
rect 1677 47 1707 177
rect 1771 47 1801 177
rect 1865 47 1895 177
rect 1959 47 1989 177
rect 2063 47 2093 177
<< pmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 457 297 493 497
rect 551 297 587 497
rect 645 297 681 497
rect 739 297 775 497
rect 833 297 869 497
rect 927 297 963 497
rect 1021 297 1057 497
rect 1115 297 1151 497
rect 1209 297 1245 497
rect 1303 297 1339 497
rect 1397 297 1433 497
rect 1491 297 1527 497
rect 1585 297 1621 497
rect 1679 297 1715 497
rect 1773 297 1809 497
rect 1867 297 1903 497
rect 1961 297 1997 497
rect 2055 297 2091 497
<< ndiff >>
rect 27 165 79 177
rect 27 131 35 165
rect 69 131 79 165
rect 27 97 79 131
rect 27 63 35 97
rect 69 63 79 97
rect 27 47 79 63
rect 109 165 173 177
rect 109 131 129 165
rect 163 131 173 165
rect 109 97 173 131
rect 109 63 129 97
rect 163 63 173 97
rect 109 47 173 63
rect 203 97 267 177
rect 203 63 223 97
rect 257 63 267 97
rect 203 47 267 63
rect 297 165 361 177
rect 297 131 317 165
rect 351 131 361 165
rect 297 97 361 131
rect 297 63 317 97
rect 351 63 361 97
rect 297 47 361 63
rect 391 97 455 177
rect 391 63 411 97
rect 445 63 455 97
rect 391 47 455 63
rect 485 165 559 177
rect 485 131 505 165
rect 539 131 559 165
rect 485 97 559 131
rect 485 63 505 97
rect 539 63 559 97
rect 485 47 559 63
rect 589 97 643 177
rect 589 63 599 97
rect 633 63 643 97
rect 589 47 643 63
rect 673 165 737 177
rect 673 131 693 165
rect 727 131 737 165
rect 673 97 737 131
rect 673 63 693 97
rect 727 63 737 97
rect 673 47 737 63
rect 767 97 831 177
rect 767 63 787 97
rect 821 63 831 97
rect 767 47 831 63
rect 861 165 925 177
rect 861 131 881 165
rect 915 131 925 165
rect 861 97 925 131
rect 861 63 881 97
rect 915 63 925 97
rect 861 47 925 63
rect 955 97 1019 177
rect 955 63 975 97
rect 1009 63 1019 97
rect 955 47 1019 63
rect 1049 165 1113 177
rect 1049 131 1069 165
rect 1103 131 1113 165
rect 1049 97 1113 131
rect 1049 63 1069 97
rect 1103 63 1113 97
rect 1049 47 1113 63
rect 1143 97 1207 177
rect 1143 63 1163 97
rect 1197 63 1207 97
rect 1143 47 1207 63
rect 1237 165 1301 177
rect 1237 131 1257 165
rect 1291 131 1301 165
rect 1237 97 1301 131
rect 1237 63 1257 97
rect 1291 63 1301 97
rect 1237 47 1301 63
rect 1331 97 1395 177
rect 1331 63 1351 97
rect 1385 63 1395 97
rect 1331 47 1395 63
rect 1425 165 1489 177
rect 1425 131 1445 165
rect 1479 131 1489 165
rect 1425 97 1489 131
rect 1425 63 1445 97
rect 1479 63 1489 97
rect 1425 47 1489 63
rect 1519 97 1583 177
rect 1519 63 1539 97
rect 1573 63 1583 97
rect 1519 47 1583 63
rect 1613 165 1677 177
rect 1613 131 1633 165
rect 1667 131 1677 165
rect 1613 97 1677 131
rect 1613 63 1633 97
rect 1667 63 1677 97
rect 1613 47 1677 63
rect 1707 97 1771 177
rect 1707 63 1727 97
rect 1761 63 1771 97
rect 1707 47 1771 63
rect 1801 165 1865 177
rect 1801 131 1821 165
rect 1855 131 1865 165
rect 1801 97 1865 131
rect 1801 63 1821 97
rect 1855 63 1865 97
rect 1801 47 1865 63
rect 1895 97 1959 177
rect 1895 63 1915 97
rect 1949 63 1959 97
rect 1895 47 1959 63
rect 1989 165 2063 177
rect 1989 131 2009 165
rect 2043 131 2063 165
rect 1989 97 2063 131
rect 1989 63 2009 97
rect 2043 63 2063 97
rect 1989 47 2063 63
rect 2093 97 2145 177
rect 2093 63 2103 97
rect 2137 63 2145 97
rect 2093 47 2145 63
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 479 175 497
rect 117 445 129 479
rect 163 445 175 479
rect 117 411 175 445
rect 117 377 129 411
rect 163 377 175 411
rect 117 343 175 377
rect 117 309 129 343
rect 163 309 175 343
rect 117 297 175 309
rect 211 485 269 497
rect 211 451 223 485
rect 257 451 269 485
rect 211 417 269 451
rect 211 383 223 417
rect 257 383 269 417
rect 211 297 269 383
rect 305 479 363 497
rect 305 445 317 479
rect 351 445 363 479
rect 305 411 363 445
rect 305 377 317 411
rect 351 377 363 411
rect 305 343 363 377
rect 305 309 317 343
rect 351 309 363 343
rect 305 297 363 309
rect 399 485 457 497
rect 399 451 411 485
rect 445 451 457 485
rect 399 417 457 451
rect 399 383 411 417
rect 445 383 457 417
rect 399 297 457 383
rect 493 479 551 497
rect 493 445 505 479
rect 539 445 551 479
rect 493 411 551 445
rect 493 377 505 411
rect 539 377 551 411
rect 493 343 551 377
rect 493 309 505 343
rect 539 309 551 343
rect 493 297 551 309
rect 587 485 645 497
rect 587 451 599 485
rect 633 451 645 485
rect 587 417 645 451
rect 587 383 599 417
rect 633 383 645 417
rect 587 297 645 383
rect 681 479 739 497
rect 681 445 693 479
rect 727 445 739 479
rect 681 411 739 445
rect 681 377 693 411
rect 727 377 739 411
rect 681 343 739 377
rect 681 309 693 343
rect 727 309 739 343
rect 681 297 739 309
rect 775 485 833 497
rect 775 451 787 485
rect 821 451 833 485
rect 775 417 833 451
rect 775 383 787 417
rect 821 383 833 417
rect 775 297 833 383
rect 869 479 927 497
rect 869 445 881 479
rect 915 445 927 479
rect 869 411 927 445
rect 869 377 881 411
rect 915 377 927 411
rect 869 343 927 377
rect 869 309 881 343
rect 915 309 927 343
rect 869 297 927 309
rect 963 485 1021 497
rect 963 451 975 485
rect 1009 451 1021 485
rect 963 417 1021 451
rect 963 383 975 417
rect 1009 383 1021 417
rect 963 297 1021 383
rect 1057 479 1115 497
rect 1057 445 1069 479
rect 1103 445 1115 479
rect 1057 411 1115 445
rect 1057 377 1069 411
rect 1103 377 1115 411
rect 1057 343 1115 377
rect 1057 309 1069 343
rect 1103 309 1115 343
rect 1057 297 1115 309
rect 1151 485 1209 497
rect 1151 451 1163 485
rect 1197 451 1209 485
rect 1151 417 1209 451
rect 1151 383 1163 417
rect 1197 383 1209 417
rect 1151 297 1209 383
rect 1245 479 1303 497
rect 1245 445 1257 479
rect 1291 445 1303 479
rect 1245 411 1303 445
rect 1245 377 1257 411
rect 1291 377 1303 411
rect 1245 343 1303 377
rect 1245 309 1257 343
rect 1291 309 1303 343
rect 1245 297 1303 309
rect 1339 485 1397 497
rect 1339 451 1351 485
rect 1385 451 1397 485
rect 1339 417 1397 451
rect 1339 383 1351 417
rect 1385 383 1397 417
rect 1339 297 1397 383
rect 1433 479 1491 497
rect 1433 445 1445 479
rect 1479 445 1491 479
rect 1433 411 1491 445
rect 1433 377 1445 411
rect 1479 377 1491 411
rect 1433 343 1491 377
rect 1433 309 1445 343
rect 1479 309 1491 343
rect 1433 297 1491 309
rect 1527 485 1585 497
rect 1527 451 1539 485
rect 1573 451 1585 485
rect 1527 417 1585 451
rect 1527 383 1539 417
rect 1573 383 1585 417
rect 1527 297 1585 383
rect 1621 479 1679 497
rect 1621 445 1633 479
rect 1667 445 1679 479
rect 1621 411 1679 445
rect 1621 377 1633 411
rect 1667 377 1679 411
rect 1621 343 1679 377
rect 1621 309 1633 343
rect 1667 309 1679 343
rect 1621 297 1679 309
rect 1715 485 1773 497
rect 1715 451 1727 485
rect 1761 451 1773 485
rect 1715 417 1773 451
rect 1715 383 1727 417
rect 1761 383 1773 417
rect 1715 297 1773 383
rect 1809 479 1867 497
rect 1809 445 1821 479
rect 1855 445 1867 479
rect 1809 411 1867 445
rect 1809 377 1821 411
rect 1855 377 1867 411
rect 1809 343 1867 377
rect 1809 309 1821 343
rect 1855 309 1867 343
rect 1809 297 1867 309
rect 1903 485 1961 497
rect 1903 451 1915 485
rect 1949 451 1961 485
rect 1903 417 1961 451
rect 1903 383 1915 417
rect 1949 383 1961 417
rect 1903 297 1961 383
rect 1997 479 2055 497
rect 1997 445 2009 479
rect 2043 445 2055 479
rect 1997 411 2055 445
rect 1997 377 2009 411
rect 2043 377 2055 411
rect 1997 343 2055 377
rect 1997 309 2009 343
rect 2043 309 2055 343
rect 1997 297 2055 309
rect 2091 485 2145 497
rect 2091 451 2103 485
rect 2137 451 2145 485
rect 2091 417 2145 451
rect 2091 383 2103 417
rect 2137 383 2145 417
rect 2091 297 2145 383
<< ndiffc >>
rect 35 131 69 165
rect 35 63 69 97
rect 129 131 163 165
rect 129 63 163 97
rect 223 63 257 97
rect 317 131 351 165
rect 317 63 351 97
rect 411 63 445 97
rect 505 131 539 165
rect 505 63 539 97
rect 599 63 633 97
rect 693 131 727 165
rect 693 63 727 97
rect 787 63 821 97
rect 881 131 915 165
rect 881 63 915 97
rect 975 63 1009 97
rect 1069 131 1103 165
rect 1069 63 1103 97
rect 1163 63 1197 97
rect 1257 131 1291 165
rect 1257 63 1291 97
rect 1351 63 1385 97
rect 1445 131 1479 165
rect 1445 63 1479 97
rect 1539 63 1573 97
rect 1633 131 1667 165
rect 1633 63 1667 97
rect 1727 63 1761 97
rect 1821 131 1855 165
rect 1821 63 1855 97
rect 1915 63 1949 97
rect 2009 131 2043 165
rect 2009 63 2043 97
rect 2103 63 2137 97
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 445 163 479
rect 129 377 163 411
rect 129 309 163 343
rect 223 451 257 485
rect 223 383 257 417
rect 317 445 351 479
rect 317 377 351 411
rect 317 309 351 343
rect 411 451 445 485
rect 411 383 445 417
rect 505 445 539 479
rect 505 377 539 411
rect 505 309 539 343
rect 599 451 633 485
rect 599 383 633 417
rect 693 445 727 479
rect 693 377 727 411
rect 693 309 727 343
rect 787 451 821 485
rect 787 383 821 417
rect 881 445 915 479
rect 881 377 915 411
rect 881 309 915 343
rect 975 451 1009 485
rect 975 383 1009 417
rect 1069 445 1103 479
rect 1069 377 1103 411
rect 1069 309 1103 343
rect 1163 451 1197 485
rect 1163 383 1197 417
rect 1257 445 1291 479
rect 1257 377 1291 411
rect 1257 309 1291 343
rect 1351 451 1385 485
rect 1351 383 1385 417
rect 1445 445 1479 479
rect 1445 377 1479 411
rect 1445 309 1479 343
rect 1539 451 1573 485
rect 1539 383 1573 417
rect 1633 445 1667 479
rect 1633 377 1667 411
rect 1633 309 1667 343
rect 1727 451 1761 485
rect 1727 383 1761 417
rect 1821 445 1855 479
rect 1821 377 1855 411
rect 1821 309 1855 343
rect 1915 451 1949 485
rect 1915 383 1949 417
rect 2009 445 2043 479
rect 2009 377 2043 411
rect 2009 309 2043 343
rect 2103 451 2137 485
rect 2103 383 2137 417
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 457 497 493 523
rect 551 497 587 523
rect 645 497 681 523
rect 739 497 775 523
rect 833 497 869 523
rect 927 497 963 523
rect 1021 497 1057 523
rect 1115 497 1151 523
rect 1209 497 1245 523
rect 1303 497 1339 523
rect 1397 497 1433 523
rect 1491 497 1527 523
rect 1585 497 1621 523
rect 1679 497 1715 523
rect 1773 497 1809 523
rect 1867 497 1903 523
rect 1961 497 1997 523
rect 2055 497 2091 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 457 282 493 297
rect 551 282 587 297
rect 645 282 681 297
rect 739 282 775 297
rect 833 282 869 297
rect 927 282 963 297
rect 1021 282 1057 297
rect 1115 282 1151 297
rect 1209 282 1245 297
rect 1303 282 1339 297
rect 1397 282 1433 297
rect 1491 282 1527 297
rect 1585 282 1621 297
rect 1679 282 1715 297
rect 1773 282 1809 297
rect 1867 282 1903 297
rect 1961 282 1997 297
rect 2055 282 2091 297
rect 79 259 119 282
rect 173 259 213 282
rect 267 259 307 282
rect 361 259 401 282
rect 455 259 495 282
rect 549 259 589 282
rect 79 249 589 259
rect 79 215 103 249
rect 137 215 181 249
rect 215 215 259 249
rect 293 215 337 249
rect 371 215 415 249
rect 449 215 483 249
rect 517 215 589 249
rect 79 205 589 215
rect 79 177 109 205
rect 173 177 203 205
rect 267 177 297 205
rect 361 177 391 205
rect 455 177 485 205
rect 559 177 589 205
rect 643 259 683 282
rect 737 259 777 282
rect 831 259 871 282
rect 925 259 965 282
rect 1019 259 1059 282
rect 1113 259 1153 282
rect 1207 259 1247 282
rect 1301 259 1341 282
rect 1395 259 1435 282
rect 1489 259 1529 282
rect 1583 259 1623 282
rect 1677 259 1717 282
rect 1771 259 1811 282
rect 1865 259 1905 282
rect 1959 259 1999 282
rect 2053 259 2093 282
rect 643 249 2093 259
rect 643 215 663 249
rect 697 215 741 249
rect 775 215 819 249
rect 853 215 897 249
rect 931 215 975 249
rect 1009 215 1043 249
rect 1077 215 1121 249
rect 1155 215 1199 249
rect 1233 215 1277 249
rect 1311 215 1355 249
rect 1389 215 1423 249
rect 1457 215 1501 249
rect 1535 215 1579 249
rect 1613 215 1657 249
rect 1691 215 1735 249
rect 1769 215 1813 249
rect 1847 215 1881 249
rect 1915 215 1959 249
rect 1993 215 2093 249
rect 643 205 2093 215
rect 643 177 673 205
rect 737 177 767 205
rect 831 177 861 205
rect 925 177 955 205
rect 1019 177 1049 205
rect 1113 177 1143 205
rect 1207 177 1237 205
rect 1301 177 1331 205
rect 1395 177 1425 205
rect 1489 177 1519 205
rect 1583 177 1613 205
rect 1677 177 1707 205
rect 1771 177 1801 205
rect 1865 177 1895 205
rect 1959 177 1989 205
rect 2063 177 2093 205
rect 79 21 109 47
rect 173 21 203 47
rect 267 21 297 47
rect 361 21 391 47
rect 455 21 485 47
rect 559 21 589 47
rect 643 21 673 47
rect 737 21 767 47
rect 831 21 861 47
rect 925 21 955 47
rect 1019 21 1049 47
rect 1113 21 1143 47
rect 1207 21 1237 47
rect 1301 21 1331 47
rect 1395 21 1425 47
rect 1489 21 1519 47
rect 1583 21 1613 47
rect 1677 21 1707 47
rect 1771 21 1801 47
rect 1865 21 1895 47
rect 1959 21 1989 47
rect 2063 21 2093 47
<< polycont >>
rect 103 215 137 249
rect 181 215 215 249
rect 259 215 293 249
rect 337 215 371 249
rect 415 215 449 249
rect 483 215 517 249
rect 663 215 697 249
rect 741 215 775 249
rect 819 215 853 249
rect 897 215 931 249
rect 975 215 1009 249
rect 1043 215 1077 249
rect 1121 215 1155 249
rect 1199 215 1233 249
rect 1277 215 1311 249
rect 1355 215 1389 249
rect 1423 215 1457 249
rect 1501 215 1535 249
rect 1579 215 1613 249
rect 1657 215 1691 249
rect 1735 215 1769 249
rect 1813 215 1847 249
rect 1881 215 1915 249
rect 1959 215 1993 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2300 561
rect 35 485 69 527
rect 35 417 69 451
rect 35 349 69 383
rect 35 289 69 315
rect 103 479 179 493
rect 103 445 129 479
rect 163 445 179 479
rect 103 411 179 445
rect 103 377 129 411
rect 163 377 179 411
rect 103 343 179 377
rect 223 485 257 527
rect 223 417 257 451
rect 223 367 257 383
rect 291 479 367 493
rect 291 445 317 479
rect 351 445 367 479
rect 291 411 367 445
rect 291 377 317 411
rect 351 377 367 411
rect 103 309 129 343
rect 163 323 179 343
rect 291 343 367 377
rect 411 485 445 527
rect 411 417 445 451
rect 411 367 445 383
rect 479 479 555 493
rect 479 445 505 479
rect 539 445 555 479
rect 479 411 555 445
rect 479 377 505 411
rect 539 377 555 411
rect 291 323 317 343
rect 163 309 317 323
rect 351 323 367 343
rect 479 343 555 377
rect 599 485 633 527
rect 599 417 633 451
rect 599 367 633 383
rect 667 479 743 493
rect 667 445 693 479
rect 727 445 743 479
rect 667 411 743 445
rect 667 377 693 411
rect 727 377 743 411
rect 479 323 505 343
rect 351 309 505 323
rect 539 323 555 343
rect 667 343 743 377
rect 787 485 821 527
rect 787 417 821 451
rect 787 367 821 383
rect 855 479 931 493
rect 855 445 881 479
rect 915 445 931 479
rect 855 411 931 445
rect 855 377 881 411
rect 915 377 931 411
rect 539 309 633 323
rect 103 289 633 309
rect 667 309 693 343
rect 727 323 743 343
rect 855 343 931 377
rect 975 485 1009 527
rect 975 417 1009 451
rect 975 367 1009 383
rect 1043 479 1119 493
rect 1043 445 1069 479
rect 1103 445 1119 479
rect 1043 411 1119 445
rect 1043 377 1069 411
rect 1103 377 1119 411
rect 855 323 881 343
rect 727 309 881 323
rect 915 323 931 343
rect 1043 343 1119 377
rect 1163 485 1197 527
rect 1163 417 1197 451
rect 1163 367 1197 383
rect 1231 479 1307 493
rect 1231 445 1257 479
rect 1291 445 1307 479
rect 1231 411 1307 445
rect 1231 377 1257 411
rect 1291 377 1307 411
rect 1043 323 1069 343
rect 915 309 1069 323
rect 1103 323 1119 343
rect 1231 343 1307 377
rect 1351 485 1385 527
rect 1351 417 1385 451
rect 1351 367 1385 383
rect 1419 479 1495 493
rect 1419 445 1445 479
rect 1479 445 1495 479
rect 1419 411 1495 445
rect 1419 377 1445 411
rect 1479 377 1495 411
rect 1231 323 1257 343
rect 1103 309 1257 323
rect 1291 323 1307 343
rect 1419 343 1495 377
rect 1539 485 1573 527
rect 1539 417 1573 451
rect 1539 367 1573 383
rect 1607 479 1683 493
rect 1607 445 1633 479
rect 1667 445 1683 479
rect 1607 411 1683 445
rect 1607 377 1633 411
rect 1667 377 1683 411
rect 1419 323 1445 343
rect 1291 309 1445 323
rect 1479 323 1495 343
rect 1607 343 1683 377
rect 1727 485 1761 527
rect 1727 417 1761 451
rect 1727 367 1761 383
rect 1795 479 1871 493
rect 1795 445 1821 479
rect 1855 445 1871 479
rect 1795 411 1871 445
rect 1795 377 1821 411
rect 1855 377 1871 411
rect 1607 323 1633 343
rect 1479 309 1633 323
rect 1667 323 1683 343
rect 1795 343 1871 377
rect 1915 485 1949 527
rect 1915 417 1949 451
rect 1915 367 1949 383
rect 1983 479 2059 493
rect 1983 445 2009 479
rect 2043 445 2059 479
rect 1983 411 2059 445
rect 1983 377 2009 411
rect 2043 377 2059 411
rect 1795 323 1821 343
rect 1667 309 1821 323
rect 1855 323 1871 343
rect 1983 343 2059 377
rect 2103 485 2137 527
rect 2103 417 2137 451
rect 2103 367 2137 383
rect 1983 323 2009 343
rect 1855 309 2009 323
rect 2043 323 2059 343
rect 2172 323 2227 472
rect 2043 309 2227 323
rect 667 289 2227 309
rect 598 255 633 289
rect 17 249 547 255
rect 17 215 103 249
rect 137 215 181 249
rect 215 215 259 249
rect 293 215 337 249
rect 371 215 415 249
rect 449 215 483 249
rect 517 215 547 249
rect 598 249 2035 255
rect 598 215 663 249
rect 697 215 741 249
rect 775 215 819 249
rect 853 215 897 249
rect 931 215 975 249
rect 1009 215 1043 249
rect 1077 215 1121 249
rect 1155 215 1199 249
rect 1233 215 1277 249
rect 1311 215 1355 249
rect 1389 215 1423 249
rect 1457 215 1501 249
rect 1535 215 1579 249
rect 1613 215 1657 249
rect 1691 215 1735 249
rect 1769 215 1813 249
rect 1847 215 1881 249
rect 1915 215 1959 249
rect 1993 215 2035 249
rect 598 181 633 215
rect 2127 181 2227 289
rect 35 165 69 181
rect 35 97 69 131
rect 35 17 69 63
rect 103 165 633 181
rect 103 131 129 165
rect 163 147 317 165
rect 163 131 179 147
rect 103 97 179 131
rect 291 131 317 147
rect 351 147 505 165
rect 351 131 367 147
rect 103 63 129 97
rect 163 63 179 97
rect 103 52 179 63
rect 223 97 257 113
rect 223 17 257 63
rect 291 97 367 131
rect 479 131 505 147
rect 539 147 633 165
rect 667 165 2227 181
rect 539 131 555 147
rect 291 63 317 97
rect 351 63 367 97
rect 291 52 367 63
rect 411 97 445 113
rect 411 17 445 63
rect 479 97 555 131
rect 667 131 693 165
rect 727 147 881 165
rect 727 131 743 147
rect 479 63 505 97
rect 539 63 555 97
rect 479 52 555 63
rect 599 97 633 113
rect 599 17 633 63
rect 667 97 743 131
rect 855 131 881 147
rect 915 147 1069 165
rect 915 131 931 147
rect 667 63 693 97
rect 727 63 743 97
rect 667 52 743 63
rect 787 97 821 113
rect 667 51 727 52
rect 787 17 821 63
rect 855 97 931 131
rect 1043 131 1069 147
rect 1103 147 1257 165
rect 1103 131 1119 147
rect 855 63 881 97
rect 915 63 931 97
rect 855 52 931 63
rect 975 97 1009 113
rect 881 51 915 52
rect 975 17 1009 63
rect 1043 97 1119 131
rect 1231 131 1257 147
rect 1291 147 1445 165
rect 1291 131 1307 147
rect 1043 63 1069 97
rect 1103 63 1119 97
rect 1043 52 1119 63
rect 1163 97 1197 113
rect 1069 51 1103 52
rect 1163 17 1197 63
rect 1231 97 1307 131
rect 1419 131 1445 147
rect 1479 147 1633 165
rect 1479 131 1495 147
rect 1231 63 1257 97
rect 1291 63 1307 97
rect 1231 52 1307 63
rect 1351 97 1385 113
rect 1351 17 1385 63
rect 1419 97 1495 131
rect 1607 131 1633 147
rect 1667 147 1821 165
rect 1667 131 1683 147
rect 1419 63 1445 97
rect 1479 63 1495 97
rect 1419 52 1495 63
rect 1539 97 1573 113
rect 1539 17 1573 63
rect 1607 97 1683 131
rect 1795 131 1821 147
rect 1855 147 2009 165
rect 1855 131 1871 147
rect 1607 63 1633 97
rect 1667 63 1683 97
rect 1607 52 1683 63
rect 1727 97 1761 113
rect 1727 17 1761 63
rect 1795 97 1871 131
rect 1983 131 2009 147
rect 2043 147 2227 165
rect 2043 131 2059 147
rect 1795 63 1821 97
rect 1855 63 1871 97
rect 1795 52 1871 63
rect 1915 97 1949 113
rect 1915 17 1949 63
rect 1983 97 2059 131
rect 1983 63 2009 97
rect 2043 63 2059 97
rect 1983 52 2059 63
rect 2103 97 2137 113
rect 2172 73 2227 147
rect 2103 17 2137 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2300 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
<< metal1 >>
rect 0 561 2300 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2300 561
rect 0 496 2300 527
rect 0 17 2300 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2300 17
rect 0 -48 2300 -17
<< labels >>
flabel corelocali s 399 221 433 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 307 221 341 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 2193 238 2193 238 0 FreeSans 200 0 0 0 X
port 6 nsew
flabel corelocali s 2104 306 2104 306 0 FreeSans 200 0 0 0 X
port 6 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew
rlabel comment s 0 0 0 0 4 buf_16
<< properties >>
string FIXED_BBOX 0 0 2300 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1656102
string GDS_START 1639570
<< end >>
