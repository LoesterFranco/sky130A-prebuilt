magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 327 307 596 349
rect 121 199 215 265
rect 489 165 596 307
rect 335 123 596 165
rect 640 125 709 349
rect 335 99 373 123
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 18 451 85 527
rect 218 455 284 527
rect 411 455 487 527
rect 599 455 675 527
rect 33 383 788 417
rect 33 265 67 383
rect 103 300 283 349
rect 249 297 283 300
rect 249 271 284 297
rect 33 199 85 265
rect 249 199 435 271
rect 249 161 291 199
rect 18 123 291 161
rect 18 51 85 123
rect 745 99 788 383
rect 211 17 277 89
rect 407 17 483 89
rect 599 17 675 89
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
rlabel locali s 640 125 709 349 6 A_N
port 1 nsew signal input
rlabel locali s 121 199 215 265 6 B
port 2 nsew signal input
rlabel locali s 489 165 596 307 6 X
port 3 nsew signal output
rlabel locali s 335 123 596 165 6 X
port 3 nsew signal output
rlabel locali s 335 99 373 123 6 X
port 3 nsew signal output
rlabel locali s 327 307 596 349 6 X
port 3 nsew signal output
rlabel metal1 s 0 -48 828 48 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 496 828 592 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1512614
string GDS_START 1506764
<< end >>
