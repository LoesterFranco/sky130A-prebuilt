magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 28 -17 62 17
<< scnmos >>
rect 87 47 117 131
rect 173 47 273 131
rect 431 93 531 177
rect 612 47 642 177
<< pmoshvt >>
rect 81 413 117 497
rect 173 413 273 497
rect 431 341 531 425
rect 606 297 642 497
<< ndiff >>
rect 379 152 431 177
rect 27 119 87 131
rect 27 85 35 119
rect 69 85 87 119
rect 27 47 87 85
rect 117 93 173 131
rect 117 59 129 93
rect 163 59 173 93
rect 117 47 173 59
rect 273 93 325 131
rect 379 118 387 152
rect 421 118 431 152
rect 379 93 431 118
rect 531 105 612 177
rect 531 93 554 105
rect 273 59 283 93
rect 317 59 325 93
rect 273 47 325 59
rect 546 71 554 93
rect 588 71 612 105
rect 546 47 612 71
rect 642 161 696 177
rect 642 127 654 161
rect 688 127 696 161
rect 642 93 696 127
rect 642 59 654 93
rect 688 59 696 93
rect 642 47 696 59
<< pdiff >>
rect 27 459 81 497
rect 27 425 35 459
rect 69 425 81 459
rect 27 413 81 425
rect 117 485 173 497
rect 117 451 129 485
rect 163 451 173 485
rect 117 413 173 451
rect 273 485 325 497
rect 273 451 283 485
rect 317 451 325 485
rect 273 413 325 451
rect 546 485 606 497
rect 546 451 554 485
rect 588 451 606 485
rect 546 425 606 451
rect 379 400 431 425
rect 379 366 387 400
rect 421 366 431 400
rect 379 341 431 366
rect 531 417 606 425
rect 531 383 554 417
rect 588 383 606 417
rect 531 341 606 383
rect 546 297 606 341
rect 642 485 696 497
rect 642 451 654 485
rect 688 451 696 485
rect 642 417 696 451
rect 642 383 654 417
rect 688 383 696 417
rect 642 349 696 383
rect 642 315 654 349
rect 688 315 696 349
rect 642 297 696 315
<< ndiffc >>
rect 35 85 69 119
rect 129 59 163 93
rect 387 118 421 152
rect 283 59 317 93
rect 554 71 588 105
rect 654 127 688 161
rect 654 59 688 93
<< pdiffc >>
rect 35 425 69 459
rect 129 451 163 485
rect 283 451 317 485
rect 554 451 588 485
rect 387 366 421 400
rect 554 383 588 417
rect 654 451 688 485
rect 654 383 688 417
rect 654 315 688 349
<< poly >>
rect 81 497 117 523
rect 173 497 273 523
rect 431 425 531 523
rect 606 497 642 523
rect 81 265 117 413
rect 173 265 273 413
rect 431 265 531 341
rect 606 265 642 297
rect 35 249 117 265
rect 35 215 45 249
rect 79 215 117 249
rect 35 199 117 215
rect 159 249 281 265
rect 159 215 169 249
rect 203 215 237 249
rect 271 215 281 249
rect 159 199 281 215
rect 367 249 531 265
rect 367 215 377 249
rect 411 215 445 249
rect 479 215 531 249
rect 367 199 531 215
rect 573 249 642 265
rect 573 215 589 249
rect 623 215 642 249
rect 573 199 642 215
rect 87 131 117 199
rect 173 131 273 199
rect 431 177 531 199
rect 612 177 642 199
rect 87 21 117 47
rect 173 21 273 47
rect 431 21 531 93
rect 612 21 642 47
<< polycont >>
rect 45 215 79 249
rect 169 215 203 249
rect 237 215 271 249
rect 377 215 411 249
rect 445 215 479 249
rect 589 215 623 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 17 459 76 493
rect 17 425 35 459
rect 69 425 76 459
rect 121 485 171 527
rect 121 451 129 485
rect 163 451 171 485
rect 121 435 171 451
rect 261 485 348 493
rect 261 451 283 485
rect 317 451 348 485
rect 261 435 348 451
rect 17 401 76 425
rect 17 357 189 401
rect 17 249 121 323
rect 17 215 45 249
rect 79 215 121 249
rect 17 211 121 215
rect 155 265 189 357
rect 155 249 280 265
rect 155 215 169 249
rect 203 215 237 249
rect 271 215 280 249
rect 155 199 280 215
rect 314 255 348 435
rect 538 485 604 527
rect 538 451 554 485
rect 588 451 604 485
rect 538 417 604 451
rect 382 400 426 416
rect 382 366 387 400
rect 421 366 426 400
rect 538 383 554 417
rect 588 383 604 417
rect 638 485 719 493
rect 638 451 654 485
rect 688 451 719 485
rect 638 417 719 451
rect 638 383 654 417
rect 688 383 719 417
rect 382 349 426 366
rect 638 349 719 383
rect 382 315 604 349
rect 562 265 604 315
rect 638 315 654 349
rect 688 315 719 349
rect 638 299 719 315
rect 314 249 495 255
rect 314 215 377 249
rect 411 215 445 249
rect 479 215 495 249
rect 562 249 631 265
rect 562 215 589 249
rect 623 215 631 249
rect 155 177 189 199
rect 19 143 189 177
rect 19 119 76 143
rect 19 85 35 119
rect 69 85 76 119
rect 314 109 348 215
rect 562 199 631 215
rect 562 181 604 199
rect 19 51 76 85
rect 120 93 163 109
rect 120 59 129 93
rect 120 17 163 59
rect 261 93 348 109
rect 382 152 604 181
rect 665 165 719 299
rect 382 118 387 152
rect 421 147 604 152
rect 638 161 719 165
rect 421 118 428 147
rect 382 102 428 118
rect 638 127 654 161
rect 688 127 719 161
rect 538 105 604 113
rect 261 59 283 93
rect 317 59 348 93
rect 261 51 348 59
rect 538 71 554 105
rect 588 71 604 105
rect 538 17 604 71
rect 638 93 719 127
rect 638 59 654 93
rect 688 59 719 93
rect 638 51 719 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel corelocali s 28 289 62 323 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 673 425 707 459 0 FreeSans 200 0 0 0 X
port 6 nsew
flabel corelocali s 673 357 707 391 0 FreeSans 200 0 0 0 X
port 6 nsew
flabel corelocali s 673 85 707 119 0 FreeSans 200 0 0 0 X
port 6 nsew
flabel corelocali s 28 221 62 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 673 153 707 187 0 FreeSans 200 0 0 0 X
port 6 nsew
flabel corelocali s 673 221 707 255 0 FreeSans 200 0 0 0 X
port 6 nsew
flabel corelocali s 673 289 707 323 0 FreeSans 200 0 0 0 X
port 6 nsew
flabel metal1 s 28 527 62 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew
flabel metal1 s 28 -17 62 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel nwell s 28 527 62 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew
flabel pwell s 28 -17 62 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew
rlabel comment s 0 0 0 0 4 dlygate4sd3_1
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3305392
string GDS_START 3299196
<< end >>
