magic
tech sky130A
magscale 1 2
timestamp 1599588238
<< locali >>
rect 21 236 155 323
rect 503 339 569 356
rect 257 273 569 339
rect 503 270 569 273
rect 673 364 751 596
rect 717 230 751 364
rect 505 196 751 230
rect 505 83 594 196
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 65 388 131 649
rect 189 424 305 596
rect 351 492 417 596
rect 451 530 539 649
rect 573 492 639 596
rect 351 458 639 492
rect 189 390 639 424
rect 189 208 223 390
rect 605 330 639 390
rect 605 264 683 330
rect 35 17 155 198
rect 189 142 328 208
rect 364 17 430 239
rect 642 17 708 149
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel locali s 21 236 155 323 6 A
port 1 nsew signal input
rlabel locali s 503 339 569 356 6 B
port 2 nsew signal input
rlabel locali s 503 270 569 273 6 B
port 2 nsew signal input
rlabel locali s 257 273 569 339 6 B
port 2 nsew signal input
rlabel locali s 717 230 751 364 6 X
port 3 nsew signal output
rlabel locali s 673 364 751 596 6 X
port 3 nsew signal output
rlabel locali s 505 196 751 230 6 X
port 3 nsew signal output
rlabel locali s 505 83 594 196 6 X
port 3 nsew signal output
rlabel metal1 s 0 -49 768 49 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 617 768 715 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 653686
string GDS_START 647426
<< end >>
