magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 920 561
rect 19 331 69 493
rect 187 331 253 425
rect 355 331 432 425
rect 19 297 432 331
rect 559 365 593 527
rect 727 365 761 527
rect 30 215 156 255
rect 214 215 340 255
rect 374 169 432 297
rect 489 215 620 255
rect 678 215 900 255
rect 103 17 169 102
rect 271 135 609 169
rect 711 17 777 102
rect 0 -17 920 17
<< obsli1 >>
rect 103 459 525 493
rect 103 365 153 459
rect 287 365 321 459
rect 475 331 525 459
rect 627 331 693 493
rect 795 331 861 493
rect 475 297 861 331
rect 19 136 237 170
rect 19 51 69 136
rect 203 101 237 136
rect 643 136 875 170
rect 643 101 677 136
rect 203 51 421 101
rect 459 51 677 101
rect 811 51 875 136
<< metal1 >>
rect 0 496 920 592
rect 0 -48 920 48
<< labels >>
rlabel locali s 489 215 620 255 6 A1
port 1 nsew signal input
rlabel locali s 678 215 900 255 6 A2
port 2 nsew signal input
rlabel locali s 214 215 340 255 6 B1
port 3 nsew signal input
rlabel locali s 30 215 156 255 6 B2
port 4 nsew signal input
rlabel locali s 374 169 432 297 6 Y
port 5 nsew signal output
rlabel locali s 355 331 432 425 6 Y
port 5 nsew signal output
rlabel locali s 271 135 609 169 6 Y
port 5 nsew signal output
rlabel locali s 187 331 253 425 6 Y
port 5 nsew signal output
rlabel locali s 19 331 69 493 6 Y
port 5 nsew signal output
rlabel locali s 19 297 432 331 6 Y
port 5 nsew signal output
rlabel locali s 711 17 777 102 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 103 17 169 102 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 920 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 920 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 727 365 761 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 559 365 593 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 920 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 920 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 920 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 4165480
string GDS_START 4156994
<< end >>
