magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 3206 704
rect 2536 312 2852 332
<< pwell >>
rect 0 0 3168 49
<< scnmos >>
rect 89 119 119 203
rect 167 119 197 203
rect 269 119 299 203
rect 341 119 371 203
rect 481 119 511 203
rect 679 98 709 246
rect 847 98 877 246
rect 1062 96 1092 180
rect 1162 96 1192 180
rect 1257 125 1287 209
rect 1388 125 1418 235
rect 1539 119 1569 229
rect 1625 119 1655 229
rect 1850 119 1880 229
rect 1922 119 1952 229
rect 2031 74 2061 158
rect 2139 74 2169 158
rect 2241 74 2271 222
rect 2327 74 2357 222
rect 2435 74 2465 222
rect 2634 138 2664 222
rect 2729 74 2759 222
rect 2938 74 2968 184
rect 3054 74 3084 222
<< pmoshvt >>
rect 86 464 116 592
rect 188 464 218 592
rect 272 464 302 592
rect 362 464 392 592
rect 564 464 594 592
rect 766 368 796 592
rect 856 368 886 592
rect 1078 419 1108 547
rect 1191 419 1221 503
rect 1275 419 1305 503
rect 1442 379 1472 547
rect 1550 379 1580 547
rect 1634 379 1664 547
rect 1736 379 1766 547
rect 1848 420 1878 588
rect 1956 504 1986 588
rect 2040 504 2070 588
rect 2244 392 2274 592
rect 2354 392 2384 592
rect 2432 392 2462 592
rect 2628 348 2658 476
rect 2731 348 2761 572
rect 2952 424 2982 592
rect 3054 368 3084 592
<< ndiff >>
rect 32 170 89 203
rect 32 136 44 170
rect 78 136 89 170
rect 32 119 89 136
rect 119 119 167 203
rect 197 178 269 203
rect 197 144 224 178
rect 258 144 269 178
rect 197 119 269 144
rect 299 119 341 203
rect 371 176 481 203
rect 371 142 382 176
rect 416 142 481 176
rect 371 119 481 142
rect 511 180 568 203
rect 511 146 522 180
rect 556 146 568 180
rect 511 119 568 146
rect 622 177 679 246
rect 622 143 634 177
rect 668 143 679 177
rect 622 98 679 143
rect 709 98 847 246
rect 877 234 945 246
rect 877 200 893 234
rect 927 200 945 234
rect 877 98 945 200
rect 774 82 832 98
rect 774 48 786 82
rect 820 48 832 82
rect 1338 209 1388 235
rect 1207 180 1257 209
rect 1005 146 1062 180
rect 1005 112 1017 146
rect 1051 112 1062 146
rect 1005 96 1062 112
rect 1092 148 1162 180
rect 1092 114 1117 148
rect 1151 114 1162 148
rect 1092 96 1162 114
rect 1192 125 1257 180
rect 1287 125 1388 209
rect 1418 229 1468 235
rect 1418 125 1539 229
rect 1192 96 1242 125
rect 1302 112 1373 125
rect 1302 78 1320 112
rect 1354 78 1373 112
rect 1433 119 1539 125
rect 1569 172 1625 229
rect 1569 138 1580 172
rect 1614 138 1625 172
rect 1569 119 1625 138
rect 1655 119 1739 229
rect 1793 186 1850 229
rect 1793 152 1805 186
rect 1839 152 1850 186
rect 1793 119 1850 152
rect 1880 119 1922 229
rect 1952 193 2009 229
rect 1952 159 1963 193
rect 1997 159 2009 193
rect 1952 158 2009 159
rect 2184 186 2241 222
rect 2184 158 2196 186
rect 1952 119 2031 158
rect 1433 112 1524 119
rect 1302 66 1373 78
rect 1433 78 1461 112
rect 1495 78 1524 112
rect 1670 112 1739 119
rect 1433 66 1524 78
rect 1670 78 1687 112
rect 1721 78 1739 112
rect 1670 66 1739 78
rect 1981 74 2031 119
rect 2061 74 2139 158
rect 2169 152 2196 158
rect 2230 152 2241 186
rect 2169 118 2241 152
rect 2169 84 2196 118
rect 2230 84 2241 118
rect 2169 74 2241 84
rect 2271 202 2327 222
rect 2271 168 2282 202
rect 2316 168 2327 202
rect 2271 118 2327 168
rect 2271 84 2282 118
rect 2316 84 2327 118
rect 2271 74 2327 84
rect 2357 177 2435 222
rect 2357 143 2390 177
rect 2424 143 2435 177
rect 2357 74 2435 143
rect 2465 186 2523 222
rect 2465 152 2477 186
rect 2511 152 2523 186
rect 2465 118 2523 152
rect 2577 185 2634 222
rect 2577 151 2589 185
rect 2623 151 2634 185
rect 2577 138 2634 151
rect 2664 184 2729 222
rect 2664 150 2679 184
rect 2713 150 2729 184
rect 2664 138 2729 150
rect 2465 84 2477 118
rect 2511 84 2523 118
rect 2465 74 2523 84
rect 2679 74 2729 138
rect 2759 194 2816 222
rect 2759 160 2770 194
rect 2804 160 2816 194
rect 2983 188 3054 222
rect 2983 184 2995 188
rect 2759 120 2816 160
rect 2759 86 2770 120
rect 2804 86 2816 120
rect 2759 74 2816 86
rect 2881 146 2938 184
rect 2881 112 2893 146
rect 2927 112 2938 146
rect 2881 74 2938 112
rect 2968 154 2995 184
rect 3029 154 3054 188
rect 2968 116 3054 154
rect 2968 82 2995 116
rect 3029 82 3054 116
rect 2968 74 3054 82
rect 3084 210 3141 222
rect 3084 176 3095 210
rect 3129 176 3141 210
rect 3084 120 3141 176
rect 3084 86 3095 120
rect 3129 86 3141 120
rect 3084 74 3141 86
rect 774 36 832 48
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 511 86 546
rect 27 477 39 511
rect 73 477 86 511
rect 27 464 86 477
rect 116 571 188 592
rect 116 537 139 571
rect 173 537 188 571
rect 116 464 188 537
rect 218 464 272 592
rect 302 520 362 592
rect 302 486 315 520
rect 349 486 362 520
rect 302 464 362 486
rect 392 567 451 592
rect 392 533 405 567
rect 439 533 451 567
rect 392 464 451 533
rect 505 567 564 592
rect 505 533 517 567
rect 551 533 564 567
rect 505 464 564 533
rect 594 580 653 592
rect 594 546 607 580
rect 641 546 653 580
rect 594 510 653 546
rect 594 476 607 510
rect 641 476 653 510
rect 594 464 653 476
rect 707 580 766 592
rect 707 546 719 580
rect 753 546 766 580
rect 707 499 766 546
rect 707 465 719 499
rect 753 465 766 499
rect 707 418 766 465
rect 707 384 719 418
rect 753 384 766 418
rect 707 368 766 384
rect 796 580 856 592
rect 796 546 809 580
rect 843 546 856 580
rect 796 486 856 546
rect 796 452 809 486
rect 843 452 856 486
rect 796 368 856 452
rect 886 580 945 592
rect 886 546 899 580
rect 933 546 945 580
rect 886 499 945 546
rect 886 465 899 499
rect 933 465 945 499
rect 886 418 945 465
rect 886 384 899 418
rect 933 384 945 418
rect 886 368 945 384
rect 1019 535 1078 547
rect 1019 501 1031 535
rect 1065 501 1078 535
rect 1019 465 1078 501
rect 1019 431 1031 465
rect 1065 431 1078 465
rect 1019 419 1078 431
rect 1108 503 1161 547
rect 2091 592 2226 594
rect 2091 588 2244 592
rect 1795 547 1848 588
rect 1323 533 1442 547
rect 1323 503 1335 533
rect 1108 491 1191 503
rect 1108 457 1137 491
rect 1171 457 1191 491
rect 1108 419 1191 457
rect 1221 419 1275 503
rect 1305 499 1335 503
rect 1369 499 1442 533
rect 1305 465 1442 499
rect 1305 431 1335 465
rect 1369 431 1442 465
rect 1305 419 1442 431
rect 1389 379 1442 419
rect 1472 531 1550 547
rect 1472 497 1503 531
rect 1537 497 1550 531
rect 1472 425 1550 497
rect 1472 391 1503 425
rect 1537 391 1550 425
rect 1472 379 1550 391
rect 1580 379 1634 547
rect 1664 535 1736 547
rect 1664 501 1683 535
rect 1717 501 1736 535
rect 1664 379 1736 501
rect 1766 420 1848 547
rect 1878 547 1956 588
rect 1878 513 1891 547
rect 1925 513 1956 547
rect 1878 504 1956 513
rect 1986 504 2040 588
rect 2070 582 2244 588
rect 2070 548 2103 582
rect 2137 548 2180 582
rect 2214 548 2244 582
rect 2070 504 2244 548
rect 1878 462 1938 504
rect 1878 428 1891 462
rect 1925 428 1938 462
rect 1878 420 1938 428
rect 1766 379 1819 420
rect 2191 392 2244 504
rect 2274 580 2354 592
rect 2274 546 2307 580
rect 2341 546 2354 580
rect 2274 512 2354 546
rect 2274 478 2307 512
rect 2341 478 2354 512
rect 2274 444 2354 478
rect 2274 410 2307 444
rect 2341 410 2354 444
rect 2274 392 2354 410
rect 2384 392 2432 592
rect 2462 546 2518 592
rect 2893 580 2952 592
rect 2462 512 2475 546
rect 2509 512 2518 546
rect 2462 392 2518 512
rect 2676 546 2731 572
rect 2676 512 2684 546
rect 2718 512 2731 546
rect 2676 476 2731 512
rect 2572 394 2628 476
rect 2572 360 2581 394
rect 2615 360 2628 394
rect 2572 348 2628 360
rect 2658 348 2731 476
rect 2761 560 2816 572
rect 2761 526 2774 560
rect 2808 526 2816 560
rect 2761 477 2816 526
rect 2761 443 2774 477
rect 2808 443 2816 477
rect 2761 394 2816 443
rect 2893 546 2905 580
rect 2939 546 2952 580
rect 2893 470 2952 546
rect 2893 436 2905 470
rect 2939 436 2952 470
rect 2893 424 2952 436
rect 2982 580 3054 592
rect 2982 546 3006 580
rect 3040 546 3054 580
rect 2982 473 3054 546
rect 2982 439 3006 473
rect 3040 439 3054 473
rect 2982 424 3054 439
rect 2761 360 2774 394
rect 2808 360 2816 394
rect 2761 348 2816 360
rect 3001 368 3054 424
rect 3084 580 3141 592
rect 3084 546 3097 580
rect 3131 546 3141 580
rect 3084 497 3141 546
rect 3084 463 3097 497
rect 3131 463 3141 497
rect 3084 414 3141 463
rect 3084 380 3097 414
rect 3131 380 3141 414
rect 3084 368 3141 380
<< ndiffc >>
rect 44 136 78 170
rect 224 144 258 178
rect 382 142 416 176
rect 522 146 556 180
rect 634 143 668 177
rect 893 200 927 234
rect 786 48 820 82
rect 1017 112 1051 146
rect 1117 114 1151 148
rect 1320 78 1354 112
rect 1580 138 1614 172
rect 1805 152 1839 186
rect 1963 159 1997 193
rect 1461 78 1495 112
rect 1687 78 1721 112
rect 2196 152 2230 186
rect 2196 84 2230 118
rect 2282 168 2316 202
rect 2282 84 2316 118
rect 2390 143 2424 177
rect 2477 152 2511 186
rect 2589 151 2623 185
rect 2679 150 2713 184
rect 2477 84 2511 118
rect 2770 160 2804 194
rect 2770 86 2804 120
rect 2893 112 2927 146
rect 2995 154 3029 188
rect 2995 82 3029 116
rect 3095 176 3129 210
rect 3095 86 3129 120
<< pdiffc >>
rect 39 546 73 580
rect 39 477 73 511
rect 139 537 173 571
rect 315 486 349 520
rect 405 533 439 567
rect 517 533 551 567
rect 607 546 641 580
rect 607 476 641 510
rect 719 546 753 580
rect 719 465 753 499
rect 719 384 753 418
rect 809 546 843 580
rect 809 452 843 486
rect 899 546 933 580
rect 899 465 933 499
rect 899 384 933 418
rect 1031 501 1065 535
rect 1031 431 1065 465
rect 1137 457 1171 491
rect 1335 499 1369 533
rect 1335 431 1369 465
rect 1503 497 1537 531
rect 1503 391 1537 425
rect 1683 501 1717 535
rect 1891 513 1925 547
rect 2103 548 2137 582
rect 2180 548 2214 582
rect 1891 428 1925 462
rect 2307 546 2341 580
rect 2307 478 2341 512
rect 2307 410 2341 444
rect 2475 512 2509 546
rect 2684 512 2718 546
rect 2581 360 2615 394
rect 2774 526 2808 560
rect 2774 443 2808 477
rect 2905 546 2939 580
rect 2905 436 2939 470
rect 3006 546 3040 580
rect 3006 439 3040 473
rect 2774 360 2808 394
rect 3097 546 3131 580
rect 3097 463 3131 497
rect 3097 380 3131 414
<< poly >>
rect 86 592 116 618
rect 188 592 218 618
rect 272 592 302 618
rect 362 592 392 618
rect 564 592 594 618
rect 766 592 796 618
rect 856 592 886 618
rect 960 615 1881 645
rect 86 449 116 464
rect 188 449 218 464
rect 272 449 302 464
rect 362 449 392 464
rect 564 449 594 464
rect 83 427 119 449
rect 44 411 119 427
rect 185 419 221 449
rect 44 377 60 411
rect 94 377 119 411
rect 44 343 119 377
rect 161 403 227 419
rect 161 369 177 403
rect 211 369 227 403
rect 161 353 227 369
rect 269 371 305 449
rect 359 419 519 449
rect 403 416 519 419
rect 403 382 469 416
rect 503 382 519 416
rect 269 355 355 371
rect 44 309 60 343
rect 94 309 119 343
rect 44 275 119 309
rect 44 241 60 275
rect 94 241 119 275
rect 44 225 119 241
rect 89 203 119 225
rect 167 203 197 353
rect 269 321 305 355
rect 339 321 355 355
rect 269 305 355 321
rect 403 366 519 382
rect 269 203 299 305
rect 403 263 433 366
rect 561 291 597 449
rect 766 353 796 368
rect 856 353 886 368
rect 763 334 799 353
rect 853 334 889 353
rect 341 233 433 263
rect 481 261 597 291
rect 679 318 799 334
rect 679 284 702 318
rect 736 304 799 318
rect 847 318 913 334
rect 736 284 793 304
rect 679 268 793 284
rect 847 284 863 318
rect 897 298 913 318
rect 960 298 990 615
rect 1078 547 1108 573
rect 1188 518 1224 615
rect 1845 603 1881 615
rect 1848 588 1878 603
rect 1956 588 1986 614
rect 2040 588 2070 614
rect 2244 592 2274 618
rect 2354 592 2384 618
rect 2432 592 2462 618
rect 1442 547 1472 573
rect 1550 547 1580 573
rect 1634 547 1664 573
rect 1736 547 1766 573
rect 1191 503 1221 518
rect 1275 503 1305 529
rect 1078 404 1108 419
rect 1075 351 1111 404
rect 1191 393 1221 419
rect 1275 404 1305 419
rect 1075 339 1105 351
rect 897 284 990 298
rect 847 268 990 284
rect 1032 323 1105 339
rect 1032 289 1048 323
rect 1082 303 1105 323
rect 1082 289 1192 303
rect 1272 297 1308 404
rect 1956 489 1986 504
rect 2040 489 2070 504
rect 1953 436 1989 489
rect 2037 472 2073 489
rect 2037 456 2169 472
rect 2037 442 2109 456
rect 1848 405 1878 420
rect 1845 388 1881 405
rect 1442 364 1472 379
rect 1550 364 1580 379
rect 1634 364 1664 379
rect 1736 364 1766 379
rect 1845 372 1917 388
rect 1439 340 1475 364
rect 1388 324 1475 340
rect 1032 273 1192 289
rect 341 203 371 233
rect 481 203 511 261
rect 679 246 709 268
rect 847 246 877 268
rect 89 93 119 119
rect 167 51 197 119
rect 269 93 299 119
rect 341 93 371 119
rect 481 51 511 119
rect 679 72 709 98
rect 167 21 511 51
rect 847 72 877 98
rect 960 81 990 268
rect 1062 180 1092 206
rect 1162 180 1192 273
rect 1250 281 1316 297
rect 1250 247 1266 281
rect 1300 247 1316 281
rect 1250 231 1316 247
rect 1388 290 1425 324
rect 1459 290 1475 324
rect 1547 317 1583 364
rect 1631 317 1667 364
rect 1733 333 1769 364
rect 1845 338 1867 372
rect 1901 338 1917 372
rect 1733 317 1803 333
rect 1845 322 1917 338
rect 1388 274 1475 290
rect 1517 301 1583 317
rect 1388 235 1418 274
rect 1517 267 1533 301
rect 1567 267 1583 301
rect 1517 251 1583 267
rect 1625 301 1691 317
rect 1625 267 1641 301
rect 1675 267 1691 301
rect 1625 251 1691 267
rect 1733 283 1753 317
rect 1787 283 1803 317
rect 1733 274 1803 283
rect 1959 274 1989 436
rect 2093 422 2109 442
rect 2143 422 2169 456
rect 2093 406 2169 422
rect 1257 209 1287 231
rect 1539 229 1569 251
rect 1625 229 1655 251
rect 1733 244 1880 274
rect 1850 229 1880 244
rect 1922 244 1989 274
rect 1922 229 1952 244
rect 2031 230 2097 246
rect 1257 99 1287 125
rect 1062 81 1092 96
rect 960 51 1092 81
rect 1162 51 1192 96
rect 1388 99 1418 125
rect 2031 196 2047 230
rect 2081 196 2097 230
rect 2031 180 2097 196
rect 2031 158 2061 180
rect 2139 158 2169 406
rect 2731 572 2761 598
rect 2952 592 2982 618
rect 3054 592 3084 618
rect 2628 476 2658 502
rect 2244 377 2274 392
rect 2354 377 2384 392
rect 2432 377 2462 392
rect 2241 360 2277 377
rect 2211 344 2277 360
rect 2211 310 2227 344
rect 2261 310 2277 344
rect 2351 310 2387 377
rect 2429 310 2465 377
rect 2952 409 2982 424
rect 2831 379 2985 409
rect 2628 333 2658 348
rect 2731 333 2761 348
rect 2625 310 2661 333
rect 2728 310 2764 333
rect 2211 294 2277 310
rect 2319 294 2385 310
rect 2241 222 2271 294
rect 2319 260 2335 294
rect 2369 260 2385 294
rect 2429 294 2555 310
rect 2429 280 2505 294
rect 2319 244 2385 260
rect 2435 260 2505 280
rect 2539 260 2555 294
rect 2435 244 2555 260
rect 2609 294 2675 310
rect 2609 260 2625 294
rect 2659 260 2675 294
rect 2609 244 2675 260
rect 2717 294 2783 310
rect 2717 260 2733 294
rect 2767 274 2783 294
rect 2831 274 2861 379
rect 3054 353 3084 368
rect 2767 260 2861 274
rect 2903 321 2969 337
rect 2903 287 2919 321
rect 2953 301 2969 321
rect 3051 301 3087 353
rect 2953 287 3084 301
rect 2903 271 3084 287
rect 2717 244 2861 260
rect 2327 222 2357 244
rect 2435 222 2465 244
rect 2634 222 2664 244
rect 2729 222 2759 244
rect 2831 229 2861 244
rect 1539 93 1569 119
rect 1625 93 1655 119
rect 1850 93 1880 119
rect 1922 51 1952 119
rect 2634 112 2664 138
rect 2831 199 2968 229
rect 3054 222 3084 271
rect 2938 184 2968 199
rect 1162 21 1952 51
rect 2031 48 2061 74
rect 2139 48 2169 74
rect 2241 48 2271 74
rect 2327 48 2357 74
rect 2435 48 2465 74
rect 2729 48 2759 74
rect 2938 48 2968 74
rect 3054 48 3084 74
<< polycont >>
rect 60 377 94 411
rect 177 369 211 403
rect 469 382 503 416
rect 60 309 94 343
rect 60 241 94 275
rect 305 321 339 355
rect 702 284 736 318
rect 863 284 897 318
rect 1048 289 1082 323
rect 1266 247 1300 281
rect 1425 290 1459 324
rect 1867 338 1901 372
rect 1533 267 1567 301
rect 1641 267 1675 301
rect 1753 283 1787 317
rect 2109 422 2143 456
rect 2047 196 2081 230
rect 2227 310 2261 344
rect 2335 260 2369 294
rect 2505 260 2539 294
rect 2625 260 2659 294
rect 2733 260 2767 294
rect 2919 287 2953 321
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3168 683
rect 23 580 89 596
rect 23 546 39 580
rect 73 546 89 580
rect 23 511 89 546
rect 123 571 189 649
rect 123 537 139 571
rect 173 537 189 571
rect 123 529 189 537
rect 223 581 455 615
rect 23 477 39 511
rect 73 495 89 511
rect 223 495 257 581
rect 389 567 455 581
rect 73 477 257 495
rect 23 461 257 477
rect 299 520 349 547
rect 299 486 315 520
rect 389 533 405 567
rect 439 533 455 567
rect 389 504 455 533
rect 501 567 551 649
rect 501 533 517 567
rect 501 504 551 533
rect 591 580 657 596
rect 591 546 607 580
rect 641 546 657 580
rect 591 510 657 546
rect 299 439 349 486
rect 591 476 607 510
rect 641 476 657 510
rect 591 470 657 476
rect 25 411 110 427
rect 25 377 60 411
rect 94 377 110 411
rect 25 343 110 377
rect 25 309 60 343
rect 94 309 110 343
rect 161 403 257 419
rect 299 405 421 439
rect 161 369 177 403
rect 211 369 257 403
rect 161 310 257 369
rect 291 355 353 371
rect 291 321 305 355
rect 339 321 353 355
rect 25 275 110 309
rect 291 305 353 321
rect 25 241 60 275
rect 94 241 110 275
rect 387 271 421 405
rect 455 436 657 470
rect 703 580 769 596
rect 703 546 719 580
rect 753 546 769 580
rect 703 499 769 546
rect 703 465 719 499
rect 753 465 769 499
rect 455 416 556 436
rect 455 382 469 416
rect 503 382 556 416
rect 703 418 769 465
rect 809 580 843 649
rect 809 486 843 546
rect 809 436 843 452
rect 883 580 981 596
rect 883 546 899 580
rect 933 546 981 580
rect 883 499 981 546
rect 883 465 899 499
rect 933 465 981 499
rect 703 402 719 418
rect 455 366 556 382
rect 25 225 110 241
rect 208 237 484 271
rect 28 170 94 191
rect 28 136 44 170
rect 78 136 94 170
rect 28 17 94 136
rect 208 178 274 237
rect 208 144 224 178
rect 258 144 274 178
rect 208 115 274 144
rect 366 176 416 203
rect 366 142 382 176
rect 366 17 416 142
rect 450 85 484 237
rect 522 207 556 366
rect 618 384 719 402
rect 753 402 769 418
rect 883 418 981 465
rect 753 384 849 402
rect 618 368 849 384
rect 883 384 899 418
rect 933 384 981 418
rect 883 368 981 384
rect 1015 535 1081 551
rect 1015 501 1031 535
rect 1065 501 1081 535
rect 1319 533 1385 649
rect 1015 465 1081 501
rect 1015 431 1031 465
rect 1065 431 1081 465
rect 1115 491 1225 507
rect 1115 457 1137 491
rect 1171 457 1225 491
rect 1115 441 1225 457
rect 1015 407 1081 431
rect 1015 373 1157 407
rect 522 180 572 207
rect 556 146 572 180
rect 522 119 572 146
rect 618 202 652 368
rect 815 334 849 368
rect 947 339 981 368
rect 686 318 752 334
rect 686 284 702 318
rect 736 284 752 318
rect 686 236 752 284
rect 815 318 913 334
rect 815 284 863 318
rect 897 284 913 318
rect 815 268 913 284
rect 947 323 1089 339
rect 947 289 1048 323
rect 1082 289 1089 323
rect 947 273 1089 289
rect 947 234 981 273
rect 1123 239 1157 373
rect 618 177 668 202
rect 872 200 893 234
rect 927 200 981 234
rect 1033 205 1157 239
rect 1191 365 1225 441
rect 1319 499 1335 533
rect 1369 499 1385 533
rect 1319 465 1385 499
rect 1319 431 1335 465
rect 1369 431 1385 465
rect 1319 415 1385 431
rect 1419 581 1621 615
rect 1191 331 1375 365
rect 1419 331 1453 581
rect 1487 531 1553 547
rect 1487 497 1503 531
rect 1537 497 1553 531
rect 1487 425 1553 497
rect 1587 467 1621 581
rect 1663 535 1737 649
rect 1663 501 1683 535
rect 1717 501 1737 535
rect 1771 581 2053 615
rect 1771 467 1805 581
rect 1587 433 1805 467
rect 1875 513 1891 547
rect 1925 513 1985 547
rect 1875 462 1985 513
rect 1487 391 1503 425
rect 1537 399 1553 425
rect 1875 428 1891 462
rect 1925 428 1985 462
rect 1875 422 1985 428
rect 1537 391 1803 399
rect 1487 365 1803 391
rect 618 143 634 177
rect 1033 166 1067 205
rect 1191 171 1225 331
rect 618 119 668 143
rect 702 146 1067 166
rect 702 132 1017 146
rect 702 85 736 132
rect 1001 112 1017 132
rect 1051 112 1067 146
rect 450 51 736 85
rect 770 82 836 98
rect 1001 92 1067 112
rect 1101 148 1225 171
rect 1101 114 1117 148
rect 1151 137 1225 148
rect 1259 281 1307 297
rect 1259 247 1266 281
rect 1300 247 1307 281
rect 1259 180 1307 247
rect 1341 248 1375 331
rect 1409 324 1475 331
rect 1409 290 1425 324
rect 1459 290 1475 324
rect 1737 317 1803 365
rect 1409 282 1475 290
rect 1517 301 1583 317
rect 1517 267 1533 301
rect 1567 267 1583 301
rect 1517 248 1583 267
rect 1341 214 1583 248
rect 1625 301 1703 317
rect 1625 267 1641 301
rect 1675 276 1703 301
rect 1625 242 1663 267
rect 1697 242 1703 276
rect 1625 236 1703 242
rect 1737 283 1753 317
rect 1787 283 1803 317
rect 1737 267 1803 283
rect 1851 372 1917 388
rect 1851 338 1867 372
rect 1901 338 1917 372
rect 1851 301 1917 338
rect 1951 369 1985 422
rect 2019 437 2053 581
rect 2087 582 2230 649
rect 2087 548 2103 582
rect 2137 548 2180 582
rect 2214 548 2230 582
rect 2087 532 2230 548
rect 2307 580 2357 596
rect 2341 546 2357 580
rect 2307 512 2357 546
rect 2093 478 2307 498
rect 2341 478 2357 512
rect 2459 546 2525 649
rect 2459 512 2475 546
rect 2509 512 2525 546
rect 2459 496 2525 512
rect 2668 546 2734 649
rect 2889 580 2955 596
rect 2668 512 2684 546
rect 2718 512 2734 546
rect 2668 496 2734 512
rect 2774 560 2855 578
rect 2808 526 2855 560
rect 2093 464 2357 478
rect 2093 456 2159 464
rect 2019 403 2059 437
rect 2093 422 2109 456
rect 2143 422 2159 456
rect 2307 462 2357 464
rect 2774 477 2855 526
rect 2307 444 2740 462
rect 2093 406 2159 422
rect 2025 372 2059 403
rect 2211 372 2273 430
rect 2341 428 2740 444
rect 2341 410 2443 428
rect 2307 394 2443 410
rect 1951 335 1991 369
rect 2025 360 2273 372
rect 2025 344 2277 360
rect 2025 338 2227 344
rect 1957 304 1991 335
rect 2211 310 2227 338
rect 2261 310 2277 344
rect 2211 304 2277 310
rect 1851 267 1923 301
rect 1737 180 1771 267
rect 1259 172 1771 180
rect 1259 146 1580 172
rect 1564 138 1580 146
rect 1614 146 1771 172
rect 1805 186 1855 210
rect 1839 152 1855 186
rect 1614 138 1630 146
rect 1151 114 1167 137
rect 1564 131 1630 138
rect 1101 92 1167 114
rect 770 48 786 82
rect 820 48 836 82
rect 770 17 836 48
rect 1298 78 1320 112
rect 1354 78 1377 112
rect 1298 17 1377 78
rect 1429 78 1461 112
rect 1495 96 1528 112
rect 1666 96 1687 112
rect 1495 78 1687 96
rect 1721 78 1743 112
rect 1429 62 1743 78
rect 1805 17 1855 152
rect 1889 85 1923 267
rect 1957 270 2177 304
rect 2319 294 2375 310
rect 2319 270 2335 294
rect 1957 193 1997 270
rect 2143 260 2335 270
rect 2369 260 2375 294
rect 2143 236 2375 260
rect 1957 159 1963 193
rect 1957 119 1997 159
rect 2031 230 2097 236
rect 2031 196 2047 230
rect 2081 196 2097 230
rect 2409 202 2443 394
rect 2545 360 2581 394
rect 2615 360 2631 394
rect 2545 344 2631 360
rect 2489 294 2579 344
rect 2706 310 2740 428
rect 2808 443 2855 477
rect 2774 394 2855 443
rect 2808 360 2855 394
rect 2774 344 2855 360
rect 2489 260 2505 294
rect 2539 276 2579 294
rect 2489 242 2527 260
rect 2561 242 2579 276
rect 2489 236 2579 242
rect 2613 294 2672 310
rect 2613 260 2625 294
rect 2659 260 2672 294
rect 2613 236 2672 260
rect 2706 294 2783 310
rect 2706 260 2733 294
rect 2767 260 2783 294
rect 2706 244 2783 260
rect 2545 202 2579 236
rect 2821 210 2855 344
rect 2031 85 2097 196
rect 1889 51 2097 85
rect 2180 186 2230 202
rect 2180 152 2196 186
rect 2180 118 2230 152
rect 2180 84 2196 118
rect 2180 17 2230 84
rect 2266 168 2282 202
rect 2316 168 2332 202
rect 2266 118 2332 168
rect 2374 177 2443 202
rect 2374 143 2390 177
rect 2424 143 2443 177
rect 2374 119 2443 143
rect 2477 186 2511 202
rect 2266 84 2282 118
rect 2316 85 2332 118
rect 2477 118 2511 152
rect 2545 185 2623 202
rect 2545 151 2589 185
rect 2545 134 2623 151
rect 2659 184 2718 200
rect 2659 150 2679 184
rect 2713 150 2718 184
rect 2316 84 2477 85
rect 2266 51 2511 84
rect 2659 17 2718 150
rect 2754 194 2855 210
rect 2754 160 2770 194
rect 2804 160 2855 194
rect 2754 120 2855 160
rect 2754 86 2770 120
rect 2804 86 2855 120
rect 2754 70 2855 86
rect 2889 546 2905 580
rect 2939 546 2955 580
rect 2889 470 2955 546
rect 2889 436 2905 470
rect 2939 436 2955 470
rect 2889 337 2955 436
rect 2989 580 3041 649
rect 2989 546 3006 580
rect 3040 546 3041 580
rect 2989 473 3041 546
rect 2989 439 3006 473
rect 3040 439 3041 473
rect 2989 423 3041 439
rect 3079 580 3147 596
rect 3079 546 3097 580
rect 3131 546 3147 580
rect 3079 497 3147 546
rect 3079 463 3097 497
rect 3131 463 3147 497
rect 3079 414 3147 463
rect 3079 380 3097 414
rect 3131 380 3147 414
rect 2889 321 2969 337
rect 2889 287 2919 321
rect 2953 287 2969 321
rect 2889 271 2969 287
rect 2889 146 2943 271
rect 3079 210 3147 380
rect 2889 112 2893 146
rect 2927 112 2943 146
rect 2889 70 2943 112
rect 2979 154 2995 188
rect 3029 154 3045 188
rect 2979 116 3045 154
rect 2979 82 2995 116
rect 3029 82 3045 116
rect 2979 17 3045 82
rect 3079 176 3095 210
rect 3129 176 3147 210
rect 3079 120 3147 176
rect 3079 86 3095 120
rect 3129 86 3147 120
rect 3079 70 3147 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3168 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 1663 267 1675 276
rect 1675 267 1697 276
rect 1663 242 1697 267
rect 2527 260 2539 276
rect 2539 260 2561 276
rect 2527 242 2561 260
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
<< metal1 >>
rect 0 683 3168 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3168 683
rect 0 617 3168 649
rect 1651 276 1709 282
rect 1651 242 1663 276
rect 1697 273 1709 276
rect 2515 276 2573 282
rect 2515 273 2527 276
rect 1697 245 2527 273
rect 1697 242 1709 245
rect 1651 236 1709 242
rect 2515 242 2527 245
rect 2561 242 2573 276
rect 2515 236 2573 242
rect 0 17 3168 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3168 17
rect 0 -49 3168 -17
<< labels >>
rlabel comment s 0 0 0 0 4 sdfbbp_1
flabel comment s 1201 629 1201 629 0 FreeSans 200 0 0 0 no_jumper_check
flabel pwell s 0 0 3168 49 0 FreeSans 200 0 0 0 VNB
port 8 nsew
flabel nwell s 0 617 3168 666 0 FreeSans 200 0 0 0 VPB
port 9 nsew
flabel metal1 s 0 617 3168 666 0 FreeSans 340 0 0 0 VPWR
port 10 nsew
flabel metal1 s 0 0 3168 49 0 FreeSans 340 0 0 0 VGND
port 7 nsew
flabel corelocali s 2815 390 2849 424 0 FreeSans 340 0 0 0 Q_N
port 12 nsew
flabel corelocali s 2815 464 2849 498 0 FreeSans 340 0 0 0 Q_N
port 12 nsew
flabel corelocali s 2815 538 2849 572 0 FreeSans 340 0 0 0 Q_N
port 12 nsew
flabel corelocali s 2623 242 2657 276 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 SCD
port 4 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 SCD
port 4 nsew
flabel corelocali s 3103 94 3137 128 0 FreeSans 340 0 0 0 Q
port 11 nsew
flabel corelocali s 3103 168 3137 202 0 FreeSans 340 0 0 0 Q
port 11 nsew
flabel corelocali s 3103 242 3137 276 0 FreeSans 340 0 0 0 Q
port 11 nsew
flabel corelocali s 3103 316 3137 350 0 FreeSans 340 0 0 0 Q
port 11 nsew
flabel corelocali s 3103 390 3137 424 0 FreeSans 340 0 0 0 Q
port 11 nsew
flabel corelocali s 3103 464 3137 498 0 FreeSans 340 0 0 0 Q
port 11 nsew
flabel corelocali s 3103 538 3137 572 0 FreeSans 340 0 0 0 Q
port 11 nsew
flabel corelocali s 703 242 737 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 2239 390 2273 424 0 FreeSans 340 0 0 0 SET_B
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 3168 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 74136
string GDS_START 50680
<< end >>
