magic
tech sky130A
magscale 1 2
timestamp 1604502711
<< locali >>
rect 111 313 177 483
rect 111 165 156 313
rect 111 63 177 165
rect 462 279 719 335
rect 462 201 523 279
rect 764 245 809 335
rect 558 211 809 245
rect 943 309 993 483
rect 958 165 993 309
rect 927 63 993 165
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 27 299 75 527
rect 27 17 75 177
rect 211 303 250 527
rect 284 441 444 475
rect 570 441 728 527
rect 284 249 318 441
rect 762 405 796 471
rect 843 441 909 527
rect 190 215 318 249
rect 211 17 250 177
rect 284 135 318 215
rect 352 371 893 405
rect 352 199 386 371
rect 859 265 893 371
rect 859 199 924 265
rect 859 177 893 199
rect 284 69 349 135
rect 399 127 601 161
rect 399 69 433 127
rect 467 17 533 93
rect 567 69 601 127
rect 692 143 893 177
rect 1029 299 1077 527
rect 692 69 726 143
rect 843 17 893 109
rect 1029 17 1077 177
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
rlabel locali s 764 245 809 335 6 A
port 1 nsew signal input
rlabel locali s 558 211 809 245 6 A
port 1 nsew signal input
rlabel locali s 462 279 719 335 6 B
port 2 nsew signal input
rlabel locali s 462 201 523 279 6 B
port 2 nsew signal input
rlabel locali s 958 165 993 309 6 COUT
port 3 nsew signal output
rlabel locali s 943 309 993 483 6 COUT
port 3 nsew signal output
rlabel locali s 927 63 993 165 6 COUT
port 3 nsew signal output
rlabel locali s 111 313 177 483 6 SUM
port 4 nsew signal output
rlabel locali s 111 165 156 313 6 SUM
port 4 nsew signal output
rlabel locali s 111 63 177 165 6 SUM
port 4 nsew signal output
rlabel metal1 s 0 -48 1104 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1104 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1104 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2131262
string GDS_START 2121692
<< end >>
