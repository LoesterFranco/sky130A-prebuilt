magic
tech sky130A
magscale 1 2
timestamp 1601050082
<< locali >>
rect 25 225 110 427
rect 161 225 263 359
rect 297 292 363 358
rect 697 270 779 356
rect 2789 301 2855 367
rect 3075 356 3125 596
rect 3075 310 3143 356
rect 3479 364 3541 596
rect 3075 244 3122 310
rect 3056 70 3122 244
rect 3507 210 3541 364
rect 3474 70 3541 210
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3391 683
rect 3425 649 3487 683
rect 3521 649 3583 683
rect 3617 649 3648 683
rect 23 495 73 596
rect 113 529 179 649
rect 213 581 437 615
rect 213 495 247 581
rect 23 461 247 495
rect 281 460 331 547
rect 371 460 437 581
rect 483 460 549 649
rect 297 426 331 460
rect 297 392 431 426
rect 397 258 431 392
rect 589 362 639 596
rect 685 424 735 596
rect 775 458 841 649
rect 685 390 847 424
rect 521 296 639 362
rect 297 224 554 258
rect 297 191 338 224
rect 28 17 94 191
rect 192 125 338 191
rect 436 17 486 190
rect 520 85 554 224
rect 588 119 639 296
rect 813 334 847 390
rect 881 368 957 596
rect 993 470 1043 649
rect 1077 581 1565 615
rect 1077 436 1111 581
rect 1380 580 1565 581
rect 813 268 889 334
rect 923 270 957 368
rect 1007 402 1111 436
rect 1168 442 1234 547
rect 1268 510 1334 547
rect 1380 546 1609 580
rect 1268 476 1541 510
rect 1168 408 1473 442
rect 1007 366 1073 402
rect 1299 368 1365 371
rect 1119 305 1365 368
rect 1119 270 1223 305
rect 1407 271 1473 408
rect 813 234 847 268
rect 923 236 1223 270
rect 1257 237 1473 271
rect 684 200 847 234
rect 673 132 904 166
rect 673 85 707 132
rect 520 51 707 85
rect 786 17 836 98
rect 870 85 904 132
rect 938 119 988 236
rect 1022 168 1223 202
rect 1022 85 1056 168
rect 870 51 1056 85
rect 1090 17 1144 134
rect 1189 87 1223 168
rect 1257 121 1323 237
rect 1507 203 1541 476
rect 1357 169 1541 203
rect 1575 459 1609 546
rect 1673 493 1739 649
rect 1781 459 1847 596
rect 1575 425 1847 459
rect 1893 458 1959 649
rect 1575 223 1609 425
rect 1781 424 1847 425
rect 2061 454 2127 596
rect 2246 520 2312 649
rect 2361 486 2427 596
rect 2461 520 2527 649
rect 2637 535 2687 596
rect 2856 569 3034 649
rect 2637 501 2931 535
rect 2637 486 2687 501
rect 1643 257 1724 391
rect 1781 390 1989 424
rect 2061 420 2182 454
rect 1758 350 1889 356
rect 1758 316 1855 350
rect 1923 316 1989 390
rect 2148 384 2182 420
rect 2216 452 2687 486
rect 2216 418 2282 452
rect 2316 384 2533 418
rect 2637 412 2687 452
rect 2031 316 2097 351
rect 2148 350 2350 384
rect 2499 378 2533 384
rect 2721 401 2815 467
rect 1758 290 1889 316
rect 1690 256 1724 257
rect 2031 256 2277 316
rect 1575 189 1656 223
rect 1690 222 1945 256
rect 2031 236 2097 256
rect 2311 222 2345 350
rect 2391 316 2431 350
rect 2499 344 2673 378
rect 2391 236 2465 316
rect 2499 260 2565 310
rect 2607 294 2673 344
rect 2721 267 2755 401
rect 2897 352 2931 501
rect 2965 390 3034 569
rect 3165 390 3231 649
rect 2897 286 2963 352
rect 3268 310 3340 588
rect 3379 364 3445 649
rect 3575 364 3625 649
rect 2721 260 2830 267
rect 1357 87 1423 169
rect 1189 53 1423 87
rect 1469 87 1554 135
rect 1590 121 1656 189
rect 1690 121 1777 187
rect 1690 87 1724 121
rect 1469 53 1724 87
rect 1811 17 1877 188
rect 1911 86 1945 222
rect 2188 188 2345 222
rect 2499 226 2830 260
rect 2499 188 2533 226
rect 2721 201 2830 226
rect 2897 201 2931 286
rect 2188 170 2222 188
rect 1992 120 2222 170
rect 2379 154 2533 188
rect 2567 167 2617 192
rect 2864 167 2931 201
rect 2268 120 2413 154
rect 2567 133 2898 167
rect 2268 86 2302 120
rect 1911 52 2302 86
rect 2336 17 2411 86
rect 2447 85 2531 120
rect 2567 119 2617 133
rect 2653 85 2719 99
rect 2447 51 2719 85
rect 2965 17 3022 226
rect 3268 244 3473 310
rect 3156 17 3222 226
rect 3268 108 3334 244
rect 3374 17 3440 210
rect 3576 17 3626 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3648 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 3199 649 3233 683
rect 3295 649 3329 683
rect 3391 649 3425 683
rect 3487 649 3521 683
rect 3583 649 3617 683
rect 1855 316 1889 350
rect 2431 316 2465 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
rect 3583 -17 3617 17
<< metal1 >>
rect 0 683 3648 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3391 683
rect 3425 649 3487 683
rect 3521 649 3583 683
rect 3617 649 3648 683
rect 0 617 3648 649
rect 1843 350 1901 356
rect 1843 316 1855 350
rect 1889 347 1901 350
rect 2419 350 2477 356
rect 2419 347 2431 350
rect 1889 319 2431 347
rect 1889 316 1901 319
rect 1843 310 1901 316
rect 2419 316 2431 319
rect 2465 316 2477 350
rect 2419 310 2477 316
rect 0 17 3648 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3648 17
rect 0 -49 3648 -17
<< obsm1 >>
rect 1171 273 1229 282
rect 2035 273 2093 282
rect 1171 245 2093 273
rect 1171 236 1229 245
rect 2035 236 2093 245
<< labels >>
rlabel locali s 297 292 363 358 6 D
port 1 nsew signal input
rlabel locali s 3507 210 3541 364 6 Q
port 2 nsew signal output
rlabel locali s 3479 364 3541 596 6 Q
port 2 nsew signal output
rlabel locali s 3474 70 3541 210 6 Q
port 2 nsew signal output
rlabel locali s 3075 356 3125 596 6 Q_N
port 3 nsew signal output
rlabel locali s 3075 310 3143 356 6 Q_N
port 3 nsew signal output
rlabel locali s 3075 244 3122 310 6 Q_N
port 3 nsew signal output
rlabel locali s 3056 70 3122 244 6 Q_N
port 3 nsew signal output
rlabel locali s 2789 301 2855 367 6 RESET_B
port 4 nsew signal input
rlabel locali s 25 225 110 427 6 SCD
port 5 nsew signal input
rlabel locali s 161 225 263 359 6 SCE
port 6 nsew signal input
rlabel metal1 s 2419 347 2477 356 6 SET_B
port 7 nsew signal input
rlabel metal1 s 2419 310 2477 319 6 SET_B
port 7 nsew signal input
rlabel metal1 s 1843 347 1901 356 6 SET_B
port 7 nsew signal input
rlabel metal1 s 1843 319 2477 347 6 SET_B
port 7 nsew signal input
rlabel metal1 s 1843 310 1901 319 6 SET_B
port 7 nsew signal input
rlabel locali s 697 270 779 356 6 CLK_N
port 8 nsew clock input
rlabel metal1 s 0 -49 3648 49 8 VGND
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 617 3648 715 6 VPWR
port 10 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 3648 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 50622
string GDS_START 24572
<< end >>
