magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 18 572 174 613
rect 18 538 127 572
rect 161 538 174 572
rect 18 442 174 538
<< viali >>
rect 127 538 161 572
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 192 683
rect 18 128 174 221
rect 18 94 31 128
rect 65 94 174 128
rect 18 53 174 94
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 192 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 31 94 65 128
rect 31 -17 65 17
rect 127 -17 161 17
<< metal1 >>
rect 0 683 192 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 192 683
rect 0 617 192 649
rect 112 572 176 581
rect 112 538 127 572
rect 161 538 176 572
rect 112 529 176 538
rect 16 128 80 137
rect 16 94 31 128
rect 65 94 80 128
rect 16 85 80 94
rect 0 17 192 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 192 17
rect 0 -49 192 -17
<< labels >>
rlabel metal1 s 16 85 80 137 6 VNB
port 1 nsew
rlabel viali s 127 538 161 572 6 VPB
port 2 nsew
rlabel locali s 18 442 174 613 6 VPB
port 2 nsew
rlabel metal1 s 112 529 176 581 6 VPB
port 2 nsew
rlabel metal1 s 0 -49 192 49 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 617 192 715 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE WELLTAP
string FIXED_BBOX 0 0 192 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 647370
string GDS_START 644542
<< end >>
