magic
tech sky130A
magscale 1 2
timestamp 1599588209
<< nwell >>
rect -38 332 710 704
<< pwell >>
rect 0 0 672 49
<< scpmos >>
rect 130 368 160 592
rect 230 368 260 592
rect 328 368 358 592
rect 442 368 472 592
rect 556 368 586 592
<< nmoslvt >>
rect 127 74 157 222
rect 236 74 266 222
rect 353 74 383 222
rect 439 74 469 222
rect 553 74 583 222
<< ndiff >>
rect 70 192 127 222
rect 70 158 82 192
rect 116 158 127 192
rect 70 120 127 158
rect 70 86 82 120
rect 116 86 127 120
rect 70 74 127 86
rect 157 210 236 222
rect 157 176 191 210
rect 225 176 236 210
rect 157 120 236 176
rect 157 86 191 120
rect 225 86 236 120
rect 157 74 236 86
rect 266 136 353 222
rect 266 102 291 136
rect 325 102 353 136
rect 266 74 353 102
rect 383 210 439 222
rect 383 176 394 210
rect 428 176 439 210
rect 383 120 439 176
rect 383 86 394 120
rect 428 86 439 120
rect 383 74 439 86
rect 469 136 553 222
rect 469 102 494 136
rect 528 102 553 136
rect 469 74 553 102
rect 583 210 640 222
rect 583 176 594 210
rect 628 176 640 210
rect 583 120 640 176
rect 583 86 594 120
rect 628 86 640 120
rect 583 74 640 86
<< pdiff >>
rect 27 580 130 592
rect 27 546 82 580
rect 116 546 130 580
rect 27 498 130 546
rect 27 464 74 498
rect 108 464 130 498
rect 27 414 130 464
rect 27 380 74 414
rect 108 380 130 414
rect 27 368 130 380
rect 160 580 230 592
rect 160 546 183 580
rect 217 546 230 580
rect 160 510 230 546
rect 160 476 183 510
rect 217 476 230 510
rect 160 440 230 476
rect 160 406 183 440
rect 217 406 230 440
rect 160 368 230 406
rect 260 368 328 592
rect 358 368 442 592
rect 472 368 556 592
rect 586 580 645 592
rect 586 546 599 580
rect 633 546 645 580
rect 586 510 645 546
rect 586 476 599 510
rect 633 476 645 510
rect 586 440 645 476
rect 586 406 599 440
rect 633 406 645 440
rect 586 368 645 406
<< ndiffc >>
rect 82 158 116 192
rect 82 86 116 120
rect 191 176 225 210
rect 191 86 225 120
rect 291 102 325 136
rect 394 176 428 210
rect 394 86 428 120
rect 494 102 528 136
rect 594 176 628 210
rect 594 86 628 120
<< pdiffc >>
rect 82 546 116 580
rect 74 464 108 498
rect 74 380 108 414
rect 183 546 217 580
rect 183 476 217 510
rect 183 406 217 440
rect 599 546 633 580
rect 599 476 633 510
rect 599 406 633 440
<< poly >>
rect 130 592 160 618
rect 230 592 260 618
rect 328 592 358 618
rect 442 592 472 618
rect 556 592 586 618
rect 130 353 160 368
rect 230 353 260 368
rect 328 353 358 368
rect 442 353 472 368
rect 556 353 586 368
rect 127 310 163 353
rect 227 336 263 353
rect 325 336 361 353
rect 439 336 475 353
rect 553 336 589 353
rect 21 294 163 310
rect 21 260 37 294
rect 71 260 163 294
rect 211 320 277 336
rect 211 286 227 320
rect 261 286 277 320
rect 211 270 277 286
rect 325 320 391 336
rect 325 286 341 320
rect 375 286 391 320
rect 325 270 391 286
rect 439 320 505 336
rect 439 286 455 320
rect 489 286 505 320
rect 439 270 505 286
rect 553 320 628 336
rect 553 286 578 320
rect 612 286 628 320
rect 553 270 628 286
rect 21 244 163 260
rect 127 222 157 244
rect 236 222 266 270
rect 353 222 383 270
rect 439 222 469 270
rect 553 222 583 270
rect 127 48 157 74
rect 236 48 266 74
rect 353 48 383 74
rect 439 48 469 74
rect 553 48 583 74
<< polycont >>
rect 37 260 71 294
rect 227 286 261 320
rect 341 286 375 320
rect 455 286 489 320
rect 578 286 612 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 23 580 133 649
rect 23 546 82 580
rect 116 546 133 580
rect 23 530 133 546
rect 167 580 233 596
rect 167 546 183 580
rect 217 546 233 580
rect 599 580 649 649
rect 23 498 109 530
rect 23 464 74 498
rect 108 464 109 498
rect 23 414 109 464
rect 167 510 233 546
rect 167 476 183 510
rect 217 476 233 510
rect 167 440 233 476
rect 167 424 183 440
rect 23 380 74 414
rect 108 380 109 414
rect 23 364 109 380
rect 143 406 183 424
rect 217 406 233 440
rect 143 390 233 406
rect 21 294 87 310
rect 143 304 177 390
rect 21 260 37 294
rect 71 260 87 294
rect 21 236 87 260
rect 121 270 177 304
rect 211 320 277 356
rect 211 286 227 320
rect 261 286 277 320
rect 211 270 277 286
rect 313 336 359 578
rect 409 384 459 578
rect 633 546 649 580
rect 599 510 649 546
rect 633 476 649 510
rect 599 440 649 476
rect 633 406 649 440
rect 599 390 649 406
rect 425 336 459 384
rect 313 320 391 336
rect 313 286 341 320
rect 375 286 391 320
rect 313 270 391 286
rect 425 320 505 336
rect 425 286 455 320
rect 489 286 505 320
rect 425 270 505 286
rect 562 320 647 356
rect 562 286 578 320
rect 612 286 647 320
rect 562 270 647 286
rect 121 202 155 270
rect 25 192 155 202
rect 25 158 82 192
rect 116 158 155 192
rect 25 120 155 158
rect 25 86 82 120
rect 116 86 155 120
rect 25 70 155 86
rect 191 210 644 236
rect 225 202 394 210
rect 225 176 241 202
rect 191 120 241 176
rect 378 176 394 202
rect 428 202 594 210
rect 428 176 444 202
rect 225 86 241 120
rect 191 70 241 86
rect 275 136 341 168
rect 275 102 291 136
rect 325 102 341 136
rect 275 17 341 102
rect 378 120 444 176
rect 578 176 594 202
rect 628 176 644 210
rect 378 86 394 120
rect 428 86 444 120
rect 378 70 444 86
rect 478 136 544 168
rect 478 102 494 136
rect 528 102 544 136
rect 478 17 544 102
rect 578 120 644 176
rect 578 86 594 120
rect 628 86 644 120
rect 578 70 644 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o41ai_1
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 319 390 353 424 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 319 464 353 498 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 319 538 353 572 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 415 390 449 424 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 415 464 449 498 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 415 538 449 572 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 B1
port 5 nsew
flabel corelocali s 31 94 65 128 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A4
port 4 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 672 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 745928
string GDS_START 739168
<< end >>
