magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 736 561
rect 291 443 362 527
rect 480 375 546 527
rect 580 357 632 493
rect 18 215 115 255
rect 153 215 248 257
rect 19 17 109 170
rect 204 135 248 215
rect 302 215 368 257
rect 402 215 483 255
rect 302 135 344 215
rect 598 117 632 357
rect 666 289 700 527
rect 471 17 537 113
rect 580 51 632 117
rect 666 17 700 197
rect 0 -17 736 17
<< obsli1 >>
rect 19 459 253 493
rect 19 325 85 459
rect 187 451 253 459
rect 119 407 165 425
rect 396 407 446 493
rect 119 359 446 407
rect 19 291 563 325
rect 529 181 563 291
rect 395 147 563 181
rect 395 101 429 147
rect 164 51 429 101
<< metal1 >>
rect 0 496 736 592
rect 0 -48 736 48
<< labels >>
rlabel locali s 302 215 368 257 6 A1
port 1 nsew signal input
rlabel locali s 302 135 344 215 6 A1
port 1 nsew signal input
rlabel locali s 402 215 483 255 6 A2
port 2 nsew signal input
rlabel locali s 204 135 248 215 6 B1
port 3 nsew signal input
rlabel locali s 153 215 248 257 6 B1
port 3 nsew signal input
rlabel locali s 18 215 115 255 6 B2
port 4 nsew signal input
rlabel locali s 598 117 632 357 6 X
port 5 nsew signal output
rlabel locali s 580 357 632 493 6 X
port 5 nsew signal output
rlabel locali s 580 51 632 117 6 X
port 5 nsew signal output
rlabel locali s 666 17 700 197 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 471 17 537 113 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 19 17 109 170 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 736 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 736 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 666 289 700 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 480 375 546 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 291 443 362 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 736 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 736 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 4141538
string GDS_START 4134790
<< end >>
