magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 21 236 87 310
rect 121 236 184 547
rect 134 125 184 236
rect 496 52 562 134
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 23 581 253 615
rect 23 364 73 581
rect 219 330 253 581
rect 293 364 343 649
rect 383 330 433 596
rect 219 296 433 330
rect 32 85 98 202
rect 220 228 442 262
rect 220 85 254 228
rect 32 51 254 85
rect 290 17 356 194
rect 390 70 442 228
rect 483 228 549 596
rect 583 460 649 649
rect 483 168 560 228
rect 596 17 649 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel locali s 21 236 87 310 6 A
port 1 nsew signal input
rlabel locali s 496 52 562 134 6 TE
port 2 nsew signal input
rlabel locali s 134 125 184 236 6 Z
port 3 nsew signal output
rlabel locali s 121 236 184 547 6 Z
port 3 nsew signal output
rlabel metal1 s 0 -49 672 49 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 617 672 715 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2090994
string GDS_START 2084272
<< end >>
