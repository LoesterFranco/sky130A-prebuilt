magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 31 326 82 487
rect 222 326 274 487
rect 31 292 431 326
rect 17 213 267 258
rect 304 179 431 292
rect 225 145 431 179
rect 225 56 270 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 126 360 178 527
rect 321 360 372 527
rect 112 17 181 122
rect 304 17 380 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
rlabel locali s 17 213 267 258 6 A
port 1 nsew signal input
rlabel locali s 304 179 431 292 6 Y
port 2 nsew signal output
rlabel locali s 225 145 431 179 6 Y
port 2 nsew signal output
rlabel locali s 225 56 270 145 6 Y
port 2 nsew signal output
rlabel locali s 222 326 274 487 6 Y
port 2 nsew signal output
rlabel locali s 31 326 82 487 6 Y
port 2 nsew signal output
rlabel locali s 31 292 431 326 6 Y
port 2 nsew signal output
rlabel metal1 s 0 -48 460 48 8 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 496 460 592 6 VPWR
port 4 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 460 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1801914
string GDS_START 1797560
<< end >>
