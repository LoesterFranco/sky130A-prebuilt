magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1380 561
rect 17 367 69 527
rect 17 191 68 333
rect 176 289 247 391
rect 176 265 238 289
rect 170 191 238 265
rect 474 415 602 527
rect 716 451 1098 527
rect 1206 451 1272 527
rect 103 17 169 89
rect 533 17 602 165
rect 1306 299 1363 493
rect 942 253 986 265
rect 942 191 1202 253
rect 1329 165 1363 299
rect 816 17 882 89
rect 1101 17 1272 89
rect 1306 51 1363 165
rect 0 -17 1380 17
<< obsli1 >>
rect 108 425 251 493
rect 285 425 440 493
rect 108 351 142 425
rect 102 292 142 351
rect 102 157 136 292
rect 281 323 372 391
rect 281 289 305 323
rect 339 289 372 323
rect 281 265 372 289
rect 272 241 372 265
rect 406 275 440 425
rect 636 417 680 493
rect 1132 417 1166 493
rect 636 383 1090 417
rect 636 381 680 383
rect 474 327 680 381
rect 474 315 508 327
rect 406 241 602 275
rect 17 123 238 157
rect 272 141 340 241
rect 374 187 431 207
rect 374 153 397 187
rect 374 141 431 153
rect 465 199 602 241
rect 17 51 69 123
rect 203 51 238 123
rect 465 107 499 199
rect 272 51 499 107
rect 636 51 680 327
rect 716 315 798 349
rect 832 323 992 349
rect 716 187 750 315
rect 832 289 859 323
rect 893 299 992 323
rect 1028 321 1090 383
rect 1132 355 1272 417
rect 832 255 893 289
rect 1028 287 1122 321
rect 1156 287 1272 355
rect 1238 265 1272 287
rect 784 221 893 255
rect 716 153 767 187
rect 835 157 893 221
rect 1238 199 1292 265
rect 1238 157 1272 199
rect 716 51 782 153
rect 835 123 966 157
rect 916 51 966 123
rect 1002 123 1272 157
rect 1002 51 1054 123
<< obsli1c >>
rect 305 289 339 323
rect 397 153 431 187
rect 859 289 893 323
rect 767 153 801 187
<< metal1 >>
rect 0 496 1380 592
rect 0 -48 1380 48
<< obsm1 >>
rect 293 323 351 329
rect 293 289 305 323
rect 339 320 351 323
rect 847 323 905 329
rect 847 320 859 323
rect 339 292 859 320
rect 339 289 351 292
rect 293 283 351 289
rect 847 289 859 292
rect 893 289 905 323
rect 847 283 905 289
rect 385 187 443 193
rect 385 153 397 187
rect 431 184 443 187
rect 755 187 813 193
rect 755 184 767 187
rect 431 156 767 184
rect 431 153 443 156
rect 385 147 443 153
rect 755 153 767 156
rect 801 153 813 187
rect 755 147 813 153
<< labels >>
rlabel locali s 176 289 247 391 6 GATE
port 1 nsew signal input
rlabel locali s 176 265 238 289 6 GATE
port 1 nsew signal input
rlabel locali s 170 191 238 265 6 GATE
port 1 nsew signal input
rlabel locali s 1329 165 1363 299 6 GCLK
port 2 nsew signal output
rlabel locali s 1306 299 1363 493 6 GCLK
port 2 nsew signal output
rlabel locali s 1306 51 1363 165 6 GCLK
port 2 nsew signal output
rlabel locali s 17 191 68 333 6 SCE
port 3 nsew signal input
rlabel locali s 942 253 986 265 6 CLK
port 4 nsew clock input
rlabel locali s 942 191 1202 253 6 CLK
port 4 nsew clock input
rlabel locali s 1101 17 1272 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 816 17 882 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 533 17 602 165 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 103 17 169 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 1380 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1380 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 1206 451 1272 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 716 451 1098 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 474 415 602 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 17 367 69 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 1380 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 1380 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1380 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 419710
string GDS_START 408734
<< end >>
