magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 89 47 119 177
rect 195 47 225 131
rect 288 47 318 131
rect 499 47 529 131
rect 593 47 623 131
rect 709 47 739 131
<< pmoshvt >>
rect 81 297 117 497
rect 188 369 224 453
rect 308 369 344 453
rect 491 369 527 453
rect 597 369 633 453
rect 711 369 747 453
<< ndiff >>
rect 27 161 89 177
rect 27 127 35 161
rect 69 127 89 161
rect 27 93 89 127
rect 27 59 35 93
rect 69 59 89 93
rect 27 47 89 59
rect 119 131 170 177
rect 119 122 195 131
rect 119 88 134 122
rect 168 88 195 122
rect 119 47 195 88
rect 225 47 288 131
rect 318 113 380 131
rect 318 79 338 113
rect 372 79 380 113
rect 318 47 380 79
rect 437 114 499 131
rect 437 80 445 114
rect 479 80 499 114
rect 437 47 499 80
rect 529 114 593 131
rect 529 80 539 114
rect 573 80 593 114
rect 529 47 593 80
rect 623 95 709 131
rect 623 61 646 95
rect 680 61 709 95
rect 623 47 709 61
rect 739 104 801 131
rect 739 70 759 104
rect 793 70 801 104
rect 739 47 801 70
<< pdiff >>
rect 27 477 81 497
rect 27 443 35 477
rect 69 443 81 477
rect 27 409 81 443
rect 27 375 35 409
rect 69 375 81 409
rect 27 297 81 375
rect 117 481 171 497
rect 117 447 129 481
rect 163 453 171 481
rect 362 481 474 493
rect 362 453 396 481
rect 163 447 188 453
rect 117 369 188 447
rect 224 369 308 453
rect 344 447 396 453
rect 430 453 474 481
rect 430 447 491 453
rect 344 369 491 447
rect 527 429 597 453
rect 527 395 541 429
rect 575 395 597 429
rect 527 369 597 395
rect 633 369 711 453
rect 747 429 801 453
rect 747 395 759 429
rect 793 395 801 429
rect 747 369 801 395
rect 117 297 171 369
rect 241 343 291 369
rect 241 309 249 343
rect 283 309 291 343
rect 241 297 291 309
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 134 88 168 122
rect 338 79 372 113
rect 445 80 479 114
rect 539 80 573 114
rect 646 61 680 95
rect 759 70 793 104
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 129 447 163 481
rect 396 447 430 481
rect 541 395 575 429
rect 759 395 793 429
rect 249 309 283 343
<< poly >>
rect 81 497 117 523
rect 188 453 224 479
rect 308 453 344 479
rect 491 453 527 479
rect 597 453 633 479
rect 711 453 747 479
rect 188 354 224 369
rect 81 282 117 297
rect 79 265 119 282
rect 186 265 226 354
rect 308 354 344 369
rect 491 354 527 369
rect 597 354 633 369
rect 711 354 747 369
rect 76 249 140 265
rect 76 215 86 249
rect 120 215 140 249
rect 76 199 140 215
rect 182 249 246 265
rect 182 215 192 249
rect 226 215 246 249
rect 306 220 346 354
rect 489 337 529 354
rect 388 321 529 337
rect 388 287 398 321
rect 432 287 529 321
rect 388 271 529 287
rect 182 199 246 215
rect 288 204 356 220
rect 89 177 119 199
rect 195 131 225 199
rect 288 170 298 204
rect 332 170 356 204
rect 288 154 356 170
rect 288 131 318 154
rect 499 131 529 271
rect 595 265 635 354
rect 571 249 635 265
rect 571 215 581 249
rect 615 215 635 249
rect 571 199 635 215
rect 709 265 749 354
rect 709 249 807 265
rect 709 215 758 249
rect 792 215 807 249
rect 709 199 807 215
rect 593 131 623 199
rect 709 131 739 199
rect 89 21 119 47
rect 195 21 225 47
rect 288 21 318 47
rect 499 21 529 47
rect 593 21 623 47
rect 709 21 739 47
<< polycont >>
rect 86 215 120 249
rect 192 215 226 249
rect 398 287 432 321
rect 298 170 332 204
rect 581 215 615 249
rect 758 215 792 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 17 477 69 493
rect 17 443 35 477
rect 103 481 179 527
rect 103 447 129 481
rect 163 447 179 481
rect 373 481 453 527
rect 373 447 396 481
rect 430 447 453 481
rect 17 409 69 443
rect 511 429 587 458
rect 511 411 541 429
rect 17 375 35 409
rect 17 359 69 375
rect 141 395 541 411
rect 575 395 587 429
rect 141 377 587 395
rect 17 165 52 359
rect 141 323 175 377
rect 86 289 175 323
rect 209 309 249 343
rect 283 321 432 343
rect 283 309 398 321
rect 209 299 398 309
rect 86 249 130 289
rect 377 287 398 299
rect 377 271 432 287
rect 466 299 587 377
rect 120 215 130 249
rect 164 249 264 255
rect 164 215 192 249
rect 226 215 264 249
rect 86 199 130 215
rect 298 204 343 220
rect 203 170 298 181
rect 332 170 343 204
rect 17 161 85 165
rect 17 127 35 161
rect 69 127 85 161
rect 17 93 85 127
rect 17 59 35 93
rect 69 59 85 93
rect 17 51 85 59
rect 134 122 168 150
rect 134 17 168 88
rect 203 147 343 170
rect 203 76 260 147
rect 377 113 411 271
rect 466 249 500 299
rect 667 265 707 485
rect 741 429 811 527
rect 741 395 759 429
rect 793 395 811 429
rect 741 363 811 395
rect 461 215 500 249
rect 544 249 707 265
rect 544 215 581 249
rect 615 215 707 249
rect 741 249 811 329
rect 741 215 758 249
rect 792 215 811 249
rect 461 138 495 215
rect 312 79 338 113
rect 372 79 411 113
rect 445 114 495 138
rect 479 80 495 114
rect 445 64 495 80
rect 539 145 811 181
rect 539 114 589 145
rect 573 80 589 114
rect 539 64 589 80
rect 627 95 697 111
rect 627 61 646 95
rect 680 61 697 95
rect 733 104 811 145
rect 733 70 759 104
rect 793 70 811 104
rect 733 64 811 70
rect 627 17 697 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel corelocali s 211 221 245 255 0 FreeSans 400 0 0 0 A1_N
port 1 nsew
flabel corelocali s 30 425 64 459 0 FreeSans 400 0 0 0 X
port 9 nsew
flabel corelocali s 214 85 248 119 0 FreeSans 400 0 0 0 A2_N
port 2 nsew
flabel corelocali s 598 242 598 242 0 FreeSans 400 0 0 0 B2
port 4 nsew
flabel corelocali s 760 238 760 238 0 FreeSans 400 0 0 0 B1
port 3 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
rlabel comment s 0 0 0 0 4 o2bb2a_1
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 938674
string GDS_START 931946
<< end >>
