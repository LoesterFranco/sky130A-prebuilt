magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1380 561
rect 125 435 177 527
rect 653 455 719 527
rect 825 455 891 527
rect 997 455 1063 527
rect 1169 455 1235 527
rect 29 215 130 323
rect 96 199 130 215
rect 312 341 545 407
rect 312 317 572 341
rect 514 179 572 317
rect 606 296 1290 341
rect 606 213 675 296
rect 709 213 994 262
rect 1041 215 1290 296
rect 514 173 977 179
rect 255 139 977 173
rect 255 123 465 139
rect 651 135 977 139
rect 144 17 221 89
rect 255 74 293 123
rect 327 17 393 89
rect 427 51 465 123
rect 499 17 617 105
rect 1097 17 1135 113
rect 1269 17 1321 177
rect 0 -17 1380 17
<< obsli1 >>
rect 25 401 91 493
rect 232 443 619 493
rect 25 357 198 401
rect 232 359 271 443
rect 387 441 619 443
rect 579 421 619 441
rect 925 421 963 493
rect 1097 421 1133 493
rect 1269 421 1321 493
rect 164 269 198 357
rect 579 375 1321 421
rect 164 207 480 269
rect 164 159 221 207
rect 18 123 221 159
rect 1011 147 1235 181
rect 18 51 89 123
rect 1011 101 1063 147
rect 653 51 1063 101
rect 1169 51 1235 147
<< metal1 >>
rect 0 496 1380 592
rect 0 -48 1380 48
<< labels >>
rlabel locali s 709 213 994 262 6 A1
port 1 nsew signal input
rlabel locali s 1041 215 1290 296 6 A2
port 2 nsew signal input
rlabel locali s 606 296 1290 341 6 A2
port 2 nsew signal input
rlabel locali s 606 213 675 296 6 A2
port 2 nsew signal input
rlabel locali s 96 199 130 215 6 B1_N
port 3 nsew signal input
rlabel locali s 29 215 130 323 6 B1_N
port 3 nsew signal input
rlabel locali s 651 135 977 139 6 Y
port 4 nsew signal output
rlabel locali s 514 179 572 317 6 Y
port 4 nsew signal output
rlabel locali s 514 173 977 179 6 Y
port 4 nsew signal output
rlabel locali s 427 51 465 123 6 Y
port 4 nsew signal output
rlabel locali s 312 341 545 407 6 Y
port 4 nsew signal output
rlabel locali s 312 317 572 341 6 Y
port 4 nsew signal output
rlabel locali s 255 139 977 173 6 Y
port 4 nsew signal output
rlabel locali s 255 123 465 139 6 Y
port 4 nsew signal output
rlabel locali s 255 74 293 123 6 Y
port 4 nsew signal output
rlabel locali s 1269 17 1321 177 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 1097 17 1135 113 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 499 17 617 105 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 327 17 393 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 144 17 221 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 1380 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1380 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 1169 455 1235 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 997 455 1063 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 825 455 891 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 653 455 719 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 125 435 177 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 1380 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 1380 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1380 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 4091804
string GDS_START 4082372
<< end >>
