magic
tech sky130A
magscale 1 2
timestamp 1604502729
<< locali >>
rect 119 424 185 596
rect 299 424 365 596
rect 591 424 657 547
rect 119 390 657 424
rect 25 270 110 356
rect 144 236 178 390
rect 217 270 403 356
rect 487 330 647 356
rect 487 264 689 330
rect 737 264 939 330
rect 873 236 939 264
rect 112 119 178 236
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 29 390 79 649
rect 225 458 259 649
rect 405 458 455 649
rect 501 581 731 615
rect 501 458 551 581
rect 697 398 731 581
rect 771 432 837 649
rect 871 398 937 596
rect 697 364 937 398
rect 26 85 76 236
rect 212 146 278 236
rect 312 230 378 236
rect 312 196 832 230
rect 312 180 378 196
rect 212 85 466 146
rect 26 51 466 85
rect 512 17 578 159
rect 614 70 648 196
rect 684 17 750 159
rect 787 70 832 196
rect 866 17 937 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
rlabel locali s 873 236 939 264 6 A1
port 1 nsew signal input
rlabel locali s 737 264 939 330 6 A1
port 1 nsew signal input
rlabel locali s 487 330 647 356 6 A2
port 2 nsew signal input
rlabel locali s 487 264 689 330 6 A2
port 2 nsew signal input
rlabel locali s 217 270 403 356 6 B1
port 3 nsew signal input
rlabel locali s 25 270 110 356 6 C1
port 4 nsew signal input
rlabel locali s 591 424 657 547 6 Y
port 5 nsew signal output
rlabel locali s 299 424 365 596 6 Y
port 5 nsew signal output
rlabel locali s 144 236 178 390 6 Y
port 5 nsew signal output
rlabel locali s 119 424 185 596 6 Y
port 5 nsew signal output
rlabel locali s 119 390 657 424 6 Y
port 5 nsew signal output
rlabel locali s 112 119 178 236 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -49 960 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 960 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1089940
string GDS_START 1080758
<< end >>
