magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 17 289 419 323
rect 17 215 125 289
rect 171 215 289 255
rect 343 215 419 289
rect 1165 391 1215 493
rect 1353 391 1403 493
rect 1165 357 1403 391
rect 1353 331 1403 357
rect 723 289 1093 323
rect 723 215 799 289
rect 833 215 977 255
rect 1011 215 1093 289
rect 1353 283 1542 331
rect 1481 181 1542 283
rect 1147 145 1542 181
rect 1147 55 1223 145
rect 1335 55 1411 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 28 359 69 527
rect 121 459 359 493
rect 121 357 171 459
rect 309 425 359 459
rect 403 425 453 527
rect 215 391 265 425
rect 497 393 555 493
rect 599 427 745 527
rect 883 427 933 527
rect 789 393 839 425
rect 977 393 1027 493
rect 497 391 573 393
rect 215 357 573 391
rect 453 321 573 357
rect 453 287 539 321
rect 453 283 573 287
rect 651 357 1027 393
rect 1071 359 1121 527
rect 1259 433 1309 527
rect 1447 365 1497 527
rect 453 215 539 283
rect 651 249 689 357
rect 573 215 689 249
rect 1133 289 1145 323
rect 1179 289 1201 323
rect 1133 249 1201 289
rect 1133 215 1417 249
rect 19 147 445 181
rect 19 145 273 147
rect 19 51 85 145
rect 129 17 163 111
rect 197 51 273 145
rect 317 17 351 111
rect 385 95 445 147
rect 479 163 539 215
rect 651 181 689 215
rect 479 129 555 163
rect 651 145 941 181
rect 865 129 941 145
rect 385 51 649 95
rect 703 17 737 111
rect 985 95 1035 179
rect 771 61 1035 95
rect 1079 17 1113 179
rect 1267 17 1301 111
rect 1455 17 1489 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 539 287 573 321
rect 1145 289 1179 323
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
<< metal1 >>
rect 0 561 1564 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 0 496 1564 527
rect 0 17 1564 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
rect 0 -48 1564 -17
<< obsm1 >>
rect 527 321 595 327
rect 527 287 539 321
rect 573 320 595 321
rect 1133 323 1192 329
rect 1133 320 1145 323
rect 573 292 1145 320
rect 573 287 595 292
rect 527 277 595 287
rect 1133 289 1145 292
rect 1179 289 1192 323
rect 1133 279 1192 289
<< labels >>
rlabel locali s 1011 215 1093 289 6 A1_N
port 1 nsew signal input
rlabel locali s 723 289 1093 323 6 A1_N
port 1 nsew signal input
rlabel locali s 723 215 799 289 6 A1_N
port 1 nsew signal input
rlabel locali s 833 215 977 255 6 A2_N
port 2 nsew signal input
rlabel locali s 343 215 419 289 6 B1
port 3 nsew signal input
rlabel locali s 17 289 419 323 6 B1
port 3 nsew signal input
rlabel locali s 17 215 125 289 6 B1
port 3 nsew signal input
rlabel locali s 171 215 289 255 6 B2
port 4 nsew signal input
rlabel locali s 1481 181 1542 283 6 X
port 5 nsew signal output
rlabel locali s 1353 391 1403 493 6 X
port 5 nsew signal output
rlabel locali s 1353 331 1403 357 6 X
port 5 nsew signal output
rlabel locali s 1353 283 1542 331 6 X
port 5 nsew signal output
rlabel locali s 1335 55 1411 145 6 X
port 5 nsew signal output
rlabel locali s 1165 391 1215 493 6 X
port 5 nsew signal output
rlabel locali s 1165 357 1403 391 6 X
port 5 nsew signal output
rlabel locali s 1147 145 1542 181 6 X
port 5 nsew signal output
rlabel locali s 1147 55 1223 145 6 X
port 5 nsew signal output
rlabel metal1 s 0 -48 1564 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 1564 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1564 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 924254
string GDS_START 912514
<< end >>
