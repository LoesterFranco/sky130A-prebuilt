magic
tech sky130A
magscale 1 2
timestamp 1599588238
<< locali >>
rect 306 492 356 596
rect 610 492 644 547
rect 306 458 644 492
rect 92 270 167 356
rect 306 236 373 458
rect 450 390 743 424
rect 450 270 516 390
rect 564 270 647 356
rect 697 330 743 390
rect 697 264 811 330
rect 323 123 373 236
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 23 390 128 572
rect 23 236 57 390
rect 201 364 267 649
rect 396 530 470 649
rect 504 581 751 615
rect 504 526 570 581
rect 684 458 751 581
rect 206 236 272 310
rect 791 364 841 649
rect 23 202 272 236
rect 23 70 73 202
rect 109 17 175 168
rect 221 85 287 168
rect 407 230 649 236
rect 407 202 837 230
rect 407 85 473 202
rect 615 196 837 202
rect 221 51 473 85
rect 507 17 573 168
rect 615 70 649 196
rect 685 17 751 162
rect 787 70 837 196
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel locali s 697 330 743 390 6 A1
port 1 nsew signal input
rlabel locali s 697 264 811 330 6 A1
port 1 nsew signal input
rlabel locali s 450 390 743 424 6 A1
port 1 nsew signal input
rlabel locali s 450 270 516 390 6 A1
port 1 nsew signal input
rlabel locali s 564 270 647 356 6 A2
port 2 nsew signal input
rlabel locali s 92 270 167 356 6 B1_N
port 3 nsew signal input
rlabel locali s 610 492 644 547 6 Y
port 4 nsew signal output
rlabel locali s 323 123 373 236 6 Y
port 4 nsew signal output
rlabel locali s 306 492 356 596 6 Y
port 4 nsew signal output
rlabel locali s 306 458 644 492 6 Y
port 4 nsew signal output
rlabel locali s 306 236 373 458 6 Y
port 4 nsew signal output
rlabel metal1 s 0 -49 864 49 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 617 864 715 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1426168
string GDS_START 1418580
<< end >>
