magic
tech sky130A
magscale 1 2
timestamp 1604502701
<< nwell >>
rect -38 332 710 704
<< pwell >>
rect 0 0 672 49
<< scpmos >>
rect 87 368 117 592
rect 177 368 207 592
rect 371 392 401 592
rect 461 392 491 592
rect 551 392 581 592
<< nmoslvt >>
rect 120 74 150 222
rect 206 74 236 222
rect 368 74 398 222
rect 454 74 484 222
rect 548 74 578 222
<< ndiff >>
rect 67 210 120 222
rect 67 176 75 210
rect 109 176 120 210
rect 67 120 120 176
rect 67 86 75 120
rect 109 86 120 120
rect 67 74 120 86
rect 150 194 206 222
rect 150 160 161 194
rect 195 160 206 194
rect 150 120 206 160
rect 150 86 161 120
rect 195 86 206 120
rect 150 74 206 86
rect 236 118 368 222
rect 236 84 247 118
rect 281 84 323 118
rect 357 84 368 118
rect 236 74 368 84
rect 398 202 454 222
rect 398 168 409 202
rect 443 168 454 202
rect 398 116 454 168
rect 398 82 409 116
rect 443 82 454 116
rect 398 74 454 82
rect 484 74 548 222
rect 578 202 635 222
rect 578 168 589 202
rect 623 168 635 202
rect 578 120 635 168
rect 578 86 589 120
rect 623 86 635 120
rect 578 74 635 86
<< pdiff >>
rect 32 580 87 592
rect 32 546 40 580
rect 74 546 87 580
rect 32 497 87 546
rect 32 463 40 497
rect 74 463 87 497
rect 32 414 87 463
rect 32 380 40 414
rect 74 380 87 414
rect 32 368 87 380
rect 117 580 177 592
rect 117 546 130 580
rect 164 546 177 580
rect 117 497 177 546
rect 117 463 130 497
rect 164 463 177 497
rect 117 414 177 463
rect 117 380 130 414
rect 164 380 177 414
rect 117 368 177 380
rect 207 580 262 592
rect 207 546 220 580
rect 254 546 262 580
rect 207 511 262 546
rect 207 477 220 511
rect 254 477 262 511
rect 207 443 262 477
rect 207 409 220 443
rect 254 409 262 443
rect 207 368 262 409
rect 316 580 371 592
rect 316 546 324 580
rect 358 546 371 580
rect 316 509 371 546
rect 316 475 324 509
rect 358 475 371 509
rect 316 438 371 475
rect 316 404 324 438
rect 358 404 371 438
rect 316 392 371 404
rect 401 580 461 592
rect 401 546 414 580
rect 448 546 461 580
rect 401 509 461 546
rect 401 475 414 509
rect 448 475 461 509
rect 401 438 461 475
rect 401 404 414 438
rect 448 404 461 438
rect 401 392 461 404
rect 491 584 551 592
rect 491 550 504 584
rect 538 550 551 584
rect 491 516 551 550
rect 491 482 504 516
rect 538 482 551 516
rect 491 448 551 482
rect 491 414 504 448
rect 538 414 551 448
rect 491 392 551 414
rect 581 580 636 592
rect 581 546 594 580
rect 628 546 636 580
rect 581 509 636 546
rect 581 475 594 509
rect 628 475 636 509
rect 581 438 636 475
rect 581 404 594 438
rect 628 404 636 438
rect 581 392 636 404
<< ndiffc >>
rect 75 176 109 210
rect 75 86 109 120
rect 161 160 195 194
rect 161 86 195 120
rect 247 84 281 118
rect 323 84 357 118
rect 409 168 443 202
rect 409 82 443 116
rect 589 168 623 202
rect 589 86 623 120
<< pdiffc >>
rect 40 546 74 580
rect 40 463 74 497
rect 40 380 74 414
rect 130 546 164 580
rect 130 463 164 497
rect 130 380 164 414
rect 220 546 254 580
rect 220 477 254 511
rect 220 409 254 443
rect 324 546 358 580
rect 324 475 358 509
rect 324 404 358 438
rect 414 546 448 580
rect 414 475 448 509
rect 414 404 448 438
rect 504 550 538 584
rect 504 482 538 516
rect 504 414 538 448
rect 594 546 628 580
rect 594 475 628 509
rect 594 404 628 438
<< poly >>
rect 87 592 117 618
rect 177 592 207 618
rect 371 592 401 618
rect 461 592 491 618
rect 551 592 581 618
rect 371 377 401 392
rect 461 377 491 392
rect 551 377 581 392
rect 87 353 117 368
rect 177 353 207 368
rect 368 358 401 377
rect 84 310 120 353
rect 174 310 210 353
rect 368 310 398 358
rect 458 310 494 377
rect 551 358 584 377
rect 554 310 584 358
rect 84 294 279 310
rect 84 260 229 294
rect 263 260 279 294
rect 84 244 279 260
rect 332 294 398 310
rect 332 260 348 294
rect 382 260 398 294
rect 332 244 398 260
rect 440 294 506 310
rect 440 260 456 294
rect 490 260 506 294
rect 440 244 506 260
rect 548 294 651 310
rect 548 260 601 294
rect 635 260 651 294
rect 548 244 651 260
rect 120 222 150 244
rect 206 222 236 244
rect 368 222 398 244
rect 454 222 484 244
rect 548 222 578 244
rect 120 48 150 74
rect 206 48 236 74
rect 368 48 398 74
rect 454 48 484 74
rect 548 48 578 74
<< polycont >>
rect 229 260 263 294
rect 348 260 382 294
rect 456 260 490 294
rect 601 260 635 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 24 580 74 649
rect 24 546 40 580
rect 24 497 74 546
rect 24 463 40 497
rect 24 414 74 463
rect 24 380 40 414
rect 24 364 74 380
rect 114 580 170 596
rect 114 546 130 580
rect 164 546 170 580
rect 114 497 170 546
rect 114 463 130 497
rect 164 463 170 497
rect 114 414 170 463
rect 114 380 130 414
rect 164 380 170 414
rect 204 580 270 649
rect 204 546 220 580
rect 254 546 270 580
rect 204 511 270 546
rect 204 477 220 511
rect 254 477 270 511
rect 204 443 270 477
rect 204 409 220 443
rect 254 409 270 443
rect 308 580 358 596
rect 308 546 324 580
rect 308 509 358 546
rect 308 475 324 509
rect 308 438 358 475
rect 114 378 170 380
rect 308 404 324 438
rect 114 310 180 378
rect 308 375 358 404
rect 59 210 109 226
rect 59 176 75 210
rect 59 120 109 176
rect 59 86 75 120
rect 59 17 109 86
rect 145 210 180 310
rect 214 341 358 375
rect 398 580 448 596
rect 398 546 414 580
rect 398 509 448 546
rect 398 475 414 509
rect 398 438 448 475
rect 398 404 414 438
rect 488 584 554 649
rect 488 550 504 584
rect 538 550 554 584
rect 488 516 554 550
rect 488 482 504 516
rect 538 482 554 516
rect 488 448 554 482
rect 488 414 504 448
rect 538 414 554 448
rect 488 412 554 414
rect 594 580 644 596
rect 628 546 644 580
rect 594 509 644 546
rect 628 475 644 509
rect 594 438 644 475
rect 398 378 448 404
rect 628 404 644 438
rect 594 378 644 404
rect 398 344 644 378
rect 214 294 279 341
rect 214 260 229 294
rect 263 260 279 294
rect 214 244 279 260
rect 145 194 211 210
rect 145 160 161 194
rect 195 160 211 194
rect 245 202 279 244
rect 313 294 398 307
rect 313 260 348 294
rect 382 260 398 294
rect 313 236 398 260
rect 440 294 551 310
rect 440 260 456 294
rect 490 260 551 294
rect 440 236 551 260
rect 585 294 651 310
rect 585 260 601 294
rect 635 260 651 294
rect 585 236 651 260
rect 245 168 409 202
rect 443 168 459 202
rect 145 120 211 160
rect 145 86 161 120
rect 195 86 211 120
rect 145 70 211 86
rect 245 118 359 134
rect 245 84 247 118
rect 281 84 323 118
rect 357 84 359 118
rect 245 17 359 84
rect 393 116 459 168
rect 393 82 409 116
rect 443 82 459 116
rect 393 70 459 82
rect 573 168 589 202
rect 623 168 639 202
rect 573 120 639 168
rect 573 86 589 120
rect 623 86 639 120
rect 573 17 639 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a21o_2
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 319 242 353 276 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 607 242 641 276 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 511 242 545 276 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 127 390 161 424 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 127 464 161 498 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 127 538 161 572 0 FreeSans 340 0 0 0 X
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 672 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 4078452
string GDS_START 4071510
<< end >>
