magic
tech sky130A
magscale 1 2
timestamp 1599588209
<< nwell >>
rect -38 332 422 704
<< pwell >>
rect 0 0 384 49
<< scpmos >>
rect 84 368 114 592
rect 168 368 198 592
rect 270 368 300 592
<< nmoslvt >>
rect 84 74 114 222
rect 170 74 200 222
rect 270 74 300 222
<< ndiff >>
rect 27 186 84 222
rect 27 152 38 186
rect 72 152 84 186
rect 27 118 84 152
rect 27 84 39 118
rect 73 84 84 118
rect 27 74 84 84
rect 114 210 170 222
rect 114 176 125 210
rect 159 176 170 210
rect 114 123 170 176
rect 114 89 125 123
rect 159 89 170 123
rect 114 74 170 89
rect 200 123 270 222
rect 200 89 211 123
rect 245 89 270 123
rect 200 74 270 89
rect 300 210 357 222
rect 300 176 311 210
rect 345 176 357 210
rect 300 120 357 176
rect 300 86 311 120
rect 345 86 357 120
rect 300 74 357 86
<< pdiff >>
rect 27 580 84 592
rect 27 546 37 580
rect 71 546 84 580
rect 27 508 84 546
rect 27 474 37 508
rect 71 474 84 508
rect 27 440 84 474
rect 27 406 37 440
rect 71 406 84 440
rect 27 368 84 406
rect 114 368 168 592
rect 198 368 270 592
rect 300 580 357 592
rect 300 546 313 580
rect 347 546 357 580
rect 300 510 357 546
rect 300 476 313 510
rect 347 476 357 510
rect 300 440 357 476
rect 300 406 313 440
rect 347 406 357 440
rect 300 368 357 406
<< ndiffc >>
rect 38 152 72 186
rect 39 84 73 118
rect 125 176 159 210
rect 125 89 159 123
rect 211 89 245 123
rect 311 176 345 210
rect 311 86 345 120
<< pdiffc >>
rect 37 546 71 580
rect 37 474 71 508
rect 37 406 71 440
rect 313 546 347 580
rect 313 476 347 510
rect 313 406 347 440
<< poly >>
rect 84 592 114 618
rect 168 592 198 618
rect 270 592 300 618
rect 84 353 114 368
rect 168 353 198 368
rect 270 353 300 368
rect 81 310 117 353
rect 165 326 201 353
rect 267 326 303 353
rect 21 294 117 310
rect 21 260 37 294
rect 71 260 117 294
rect 159 310 225 326
rect 159 276 175 310
rect 209 276 225 310
rect 159 260 225 276
rect 267 310 363 326
rect 267 276 313 310
rect 347 276 363 310
rect 267 260 363 276
rect 21 244 117 260
rect 84 222 114 244
rect 170 222 200 260
rect 270 222 300 260
rect 84 48 114 74
rect 170 48 200 74
rect 270 48 300 74
<< polycont >>
rect 37 260 71 294
rect 175 276 209 310
rect 313 276 347 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 384 683
rect 21 580 87 649
rect 21 546 37 580
rect 71 546 87 580
rect 21 508 87 546
rect 21 474 37 508
rect 71 474 87 508
rect 21 465 87 474
rect 121 580 363 596
rect 121 546 313 580
rect 347 546 363 580
rect 121 510 363 546
rect 121 476 313 510
rect 347 476 363 510
rect 21 440 71 465
rect 21 406 37 440
rect 121 440 363 476
rect 121 424 313 440
rect 21 390 71 406
rect 106 406 313 424
rect 347 406 363 440
rect 106 390 363 406
rect 21 294 72 356
rect 21 260 37 294
rect 71 260 72 294
rect 21 236 72 260
rect 106 226 140 390
rect 174 310 263 356
rect 174 276 175 310
rect 209 276 263 310
rect 174 260 263 276
rect 297 310 363 356
rect 297 276 313 310
rect 347 276 363 310
rect 297 260 363 276
rect 106 210 361 226
rect 23 186 72 202
rect 23 152 38 186
rect 106 176 125 210
rect 159 176 311 210
rect 345 176 361 210
rect 23 142 72 152
rect 23 118 89 142
rect 23 84 39 118
rect 73 84 89 118
rect 23 17 89 84
rect 123 123 161 176
rect 123 89 125 123
rect 159 89 161 123
rect 123 73 161 89
rect 195 123 261 142
rect 195 89 211 123
rect 245 89 261 123
rect 195 17 261 89
rect 295 120 361 176
rect 295 86 311 120
rect 345 86 361 120
rect 295 70 361 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 384 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
<< metal1 >>
rect 0 683 384 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 384 683
rect 0 617 384 649
rect 0 17 384 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 384 17
rect 0 -49 384 -17
<< labels >>
rlabel comment s 0 0 0 0 4 nor3_1
flabel pwell s 0 0 384 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 0 617 384 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 384 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 384 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 127 464 161 498 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 223 464 257 498 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 319 464 353 498 0 FreeSans 340 0 0 0 Y
port 8 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 384 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1579262
string GDS_START 1574480
<< end >>
