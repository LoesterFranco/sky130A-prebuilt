magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 192 236 257 350
rect 984 270 1050 356
rect 1375 236 1441 337
rect 1751 80 1801 596
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 17 452 120 596
rect 154 452 220 649
rect 274 581 779 615
rect 17 260 51 452
rect 274 418 340 581
rect 745 551 779 581
rect 85 388 340 418
rect 386 513 711 547
rect 386 388 452 513
rect 85 384 325 388
rect 85 294 150 384
rect 17 166 89 260
rect 291 200 325 384
rect 486 286 552 479
rect 593 375 643 479
rect 359 252 552 286
rect 359 166 393 252
rect 518 218 552 252
rect 17 132 393 166
rect 17 130 89 132
rect 125 17 239 98
rect 427 92 477 218
rect 518 126 570 218
rect 604 92 643 375
rect 427 58 643 92
rect 677 85 711 513
rect 745 381 879 551
rect 745 287 811 347
rect 745 153 779 287
rect 845 253 879 381
rect 813 187 879 253
rect 916 226 950 596
rect 990 390 1040 649
rect 1205 581 1521 615
rect 1081 398 1171 568
rect 1081 390 1125 398
rect 1084 272 1125 390
rect 1205 364 1239 581
rect 1161 306 1239 364
rect 1273 310 1341 547
rect 1375 405 1441 547
rect 1487 505 1521 581
rect 1487 439 1597 505
rect 1375 371 1529 405
rect 1084 238 1273 272
rect 916 153 961 226
rect 745 119 961 153
rect 995 170 1205 204
rect 995 85 1029 170
rect 677 51 1029 85
rect 1063 17 1113 136
rect 1155 85 1205 170
rect 1239 153 1273 238
rect 1307 187 1341 310
rect 1377 153 1461 185
rect 1239 119 1461 153
rect 1495 85 1529 371
rect 1155 51 1529 85
rect 1563 172 1597 439
rect 1645 390 1711 649
rect 1651 270 1717 356
rect 1563 80 1613 172
rect 1649 17 1715 236
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
<< metal1 >>
rect 0 683 1824 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 0 617 1824 649
rect 0 17 1824 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
rect 0 -49 1824 -17
<< obsm1 >>
rect 595 347 653 356
rect 1075 347 1133 356
rect 595 319 1133 347
rect 595 310 653 319
rect 1075 310 1133 319
rect 1267 347 1325 356
rect 1651 347 1709 356
rect 1267 319 1709 347
rect 1267 310 1325 319
rect 1651 310 1709 319
<< labels >>
rlabel locali s 192 236 257 350 6 A
port 1 nsew signal input
rlabel locali s 984 270 1050 356 6 B
port 2 nsew signal input
rlabel locali s 1375 236 1441 337 6 C
port 3 nsew signal input
rlabel locali s 1751 80 1801 596 6 X
port 4 nsew signal output
rlabel metal1 s 0 -49 1824 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 617 1824 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1824 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 585532
string GDS_START 571620
<< end >>
