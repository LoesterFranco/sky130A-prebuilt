magic
tech sky130A
magscale 1 2
timestamp 1604502710
<< nwell >>
rect -38 332 1286 704
<< pwell >>
rect 0 0 1248 49
<< scpmos >>
rect 83 368 119 592
rect 193 368 229 592
rect 283 368 319 592
rect 373 368 409 592
rect 463 368 499 592
rect 652 424 688 592
rect 742 424 778 592
rect 859 392 895 592
rect 949 392 985 592
rect 1039 392 1075 592
rect 1129 392 1165 592
<< nmoslvt >>
rect 90 74 120 222
rect 193 74 223 222
rect 281 74 311 222
rect 367 74 397 222
rect 453 74 483 222
rect 675 94 705 222
rect 761 94 791 222
rect 861 125 891 253
rect 961 125 991 253
rect 1047 125 1077 253
rect 1133 125 1163 253
<< ndiff >>
rect 811 222 861 253
rect 33 202 90 222
rect 33 168 45 202
rect 79 168 90 202
rect 33 120 90 168
rect 33 86 45 120
rect 79 86 90 120
rect 33 74 90 86
rect 120 202 193 222
rect 120 168 145 202
rect 179 168 193 202
rect 120 116 193 168
rect 120 82 145 116
rect 179 82 193 116
rect 120 74 193 82
rect 223 208 281 222
rect 223 174 234 208
rect 268 174 281 208
rect 223 120 281 174
rect 223 86 234 120
rect 268 86 281 120
rect 223 74 281 86
rect 311 130 367 222
rect 311 96 322 130
rect 356 96 367 130
rect 311 74 367 96
rect 397 208 453 222
rect 397 174 408 208
rect 442 174 453 208
rect 397 120 453 174
rect 397 86 408 120
rect 442 86 453 120
rect 397 74 453 86
rect 483 208 540 222
rect 483 174 494 208
rect 528 174 540 208
rect 483 120 540 174
rect 483 86 494 120
rect 528 86 540 120
rect 618 188 675 222
rect 618 154 630 188
rect 664 154 675 188
rect 618 94 675 154
rect 705 140 761 222
rect 705 106 716 140
rect 750 106 761 140
rect 705 94 761 106
rect 791 190 861 222
rect 791 156 816 190
rect 850 156 861 190
rect 791 125 861 156
rect 891 171 961 253
rect 891 137 916 171
rect 950 137 961 171
rect 891 125 961 137
rect 991 240 1047 253
rect 991 206 1002 240
rect 1036 206 1047 240
rect 991 171 1047 206
rect 991 137 1002 171
rect 1036 137 1047 171
rect 991 125 1047 137
rect 1077 171 1133 253
rect 1077 137 1088 171
rect 1122 137 1133 171
rect 1077 125 1133 137
rect 1163 240 1221 253
rect 1163 206 1174 240
rect 1208 206 1221 240
rect 1163 171 1221 206
rect 1163 137 1174 171
rect 1208 137 1221 171
rect 1163 125 1221 137
rect 791 94 841 125
rect 483 74 540 86
<< pdiff >>
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 497 83 546
rect 27 463 39 497
rect 73 463 83 497
rect 27 414 83 463
rect 27 380 39 414
rect 73 380 83 414
rect 27 368 83 380
rect 119 580 193 592
rect 119 546 144 580
rect 178 546 193 580
rect 119 368 193 546
rect 229 421 283 592
rect 229 387 239 421
rect 273 387 283 421
rect 229 368 283 387
rect 319 580 373 592
rect 319 546 329 580
rect 363 546 373 580
rect 319 368 373 546
rect 409 421 463 592
rect 409 387 419 421
rect 453 387 463 421
rect 409 368 463 387
rect 499 580 652 592
rect 499 546 509 580
rect 543 546 591 580
rect 625 546 652 580
rect 499 424 652 546
rect 688 580 742 592
rect 688 546 698 580
rect 732 546 742 580
rect 688 476 742 546
rect 688 442 698 476
rect 732 442 742 476
rect 688 424 742 442
rect 778 544 859 592
rect 778 510 805 544
rect 839 510 859 544
rect 778 424 859 510
rect 499 368 549 424
rect 809 392 859 424
rect 895 544 949 592
rect 895 510 905 544
rect 939 510 949 544
rect 895 392 949 510
rect 985 531 1039 592
rect 985 497 995 531
rect 1029 497 1039 531
rect 985 440 1039 497
rect 985 406 995 440
rect 1029 406 1039 440
rect 985 392 1039 406
rect 1075 580 1129 592
rect 1075 546 1085 580
rect 1119 546 1129 580
rect 1075 510 1129 546
rect 1075 476 1085 510
rect 1119 476 1129 510
rect 1075 440 1129 476
rect 1075 406 1085 440
rect 1119 406 1129 440
rect 1075 392 1129 406
rect 1165 580 1221 592
rect 1165 546 1175 580
rect 1209 546 1221 580
rect 1165 510 1221 546
rect 1165 476 1175 510
rect 1209 476 1221 510
rect 1165 440 1221 476
rect 1165 406 1175 440
rect 1209 406 1221 440
rect 1165 392 1221 406
<< ndiffc >>
rect 45 168 79 202
rect 45 86 79 120
rect 145 168 179 202
rect 145 82 179 116
rect 234 174 268 208
rect 234 86 268 120
rect 322 96 356 130
rect 408 174 442 208
rect 408 86 442 120
rect 494 174 528 208
rect 494 86 528 120
rect 630 154 664 188
rect 716 106 750 140
rect 816 156 850 190
rect 916 137 950 171
rect 1002 206 1036 240
rect 1002 137 1036 171
rect 1088 137 1122 171
rect 1174 206 1208 240
rect 1174 137 1208 171
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 144 546 178 580
rect 239 387 273 421
rect 329 546 363 580
rect 419 387 453 421
rect 509 546 543 580
rect 591 546 625 580
rect 698 546 732 580
rect 698 442 732 476
rect 805 510 839 544
rect 905 510 939 544
rect 995 497 1029 531
rect 995 406 1029 440
rect 1085 546 1119 580
rect 1085 476 1119 510
rect 1085 406 1119 440
rect 1175 546 1209 580
rect 1175 476 1209 510
rect 1175 406 1209 440
<< poly >>
rect 83 592 119 618
rect 193 592 229 618
rect 283 592 319 618
rect 373 592 409 618
rect 463 592 499 618
rect 652 592 688 618
rect 742 592 778 618
rect 859 592 895 618
rect 949 592 985 618
rect 1039 592 1075 618
rect 1129 592 1165 618
rect 652 392 688 424
rect 742 392 778 424
rect 632 376 778 392
rect 83 310 119 368
rect 193 310 229 368
rect 283 324 319 368
rect 373 324 409 368
rect 463 324 499 368
rect 632 342 648 376
rect 682 356 778 376
rect 859 356 895 392
rect 949 356 985 392
rect 1039 356 1075 392
rect 682 342 791 356
rect 632 326 791 342
rect 281 310 499 324
rect 83 294 151 310
rect 83 260 101 294
rect 135 260 151 294
rect 83 244 151 260
rect 193 308 499 310
rect 193 274 313 308
rect 347 274 381 308
rect 415 274 449 308
rect 483 274 499 308
rect 193 258 499 274
rect 90 222 120 244
rect 193 222 223 258
rect 281 222 311 258
rect 367 222 397 258
rect 453 222 483 258
rect 675 222 705 326
rect 761 222 791 326
rect 835 340 901 356
rect 835 306 851 340
rect 885 306 901 340
rect 835 290 901 306
rect 949 340 1075 356
rect 949 306 985 340
rect 1019 320 1075 340
rect 1019 306 1077 320
rect 949 290 1077 306
rect 861 253 891 290
rect 961 253 991 290
rect 1047 253 1077 290
rect 1129 268 1165 392
rect 1133 253 1163 268
rect 90 48 120 74
rect 193 48 223 74
rect 281 48 311 74
rect 367 48 397 74
rect 453 48 483 74
rect 675 68 705 94
rect 761 68 791 94
rect 861 51 891 125
rect 961 99 991 125
rect 1047 99 1077 125
rect 1133 51 1163 125
rect 861 21 1163 51
<< polycont >>
rect 648 342 682 376
rect 101 260 135 294
rect 313 274 347 308
rect 381 274 415 308
rect 449 274 483 308
rect 851 306 885 340
rect 985 306 1019 340
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 17 580 89 596
rect 17 546 39 580
rect 73 546 89 580
rect 123 580 199 649
rect 123 546 144 580
rect 178 546 199 580
rect 313 580 379 649
rect 313 546 329 580
rect 363 546 379 580
rect 493 580 641 649
rect 493 546 509 580
rect 543 546 591 580
rect 625 546 641 580
rect 698 580 748 596
rect 732 546 748 580
rect 17 512 89 546
rect 17 497 664 512
rect 17 463 39 497
rect 73 478 664 497
rect 73 463 89 478
rect 17 414 89 463
rect 17 380 39 414
rect 73 380 89 414
rect 17 364 89 380
rect 217 421 469 444
rect 217 387 239 421
rect 273 387 419 421
rect 453 387 469 421
rect 217 364 469 387
rect 630 392 664 478
rect 698 476 748 546
rect 789 544 855 649
rect 789 510 805 544
rect 839 510 855 544
rect 789 494 855 510
rect 889 581 1135 615
rect 889 544 955 581
rect 1069 580 1135 581
rect 889 510 905 544
rect 939 510 955 544
rect 889 494 955 510
rect 995 531 1029 547
rect 732 460 748 476
rect 995 460 1029 497
rect 732 442 1029 460
rect 698 440 1029 442
rect 698 426 995 440
rect 732 406 995 426
rect 630 376 698 392
rect 17 202 51 364
rect 217 310 263 364
rect 630 342 648 376
rect 682 342 698 376
rect 630 326 698 342
rect 732 390 1029 406
rect 1069 546 1085 580
rect 1119 546 1135 580
rect 1069 510 1135 546
rect 1069 476 1085 510
rect 1119 476 1135 510
rect 1069 440 1135 476
rect 1069 406 1085 440
rect 1119 406 1135 440
rect 1069 390 1135 406
rect 1175 580 1225 649
rect 1209 546 1225 580
rect 1175 510 1225 546
rect 1209 476 1225 510
rect 1175 440 1225 476
rect 1209 406 1225 440
rect 1175 390 1225 406
rect 85 294 167 310
rect 85 260 101 294
rect 135 260 167 294
rect 85 236 167 260
rect 229 224 263 310
rect 297 308 596 324
rect 297 274 313 308
rect 347 274 381 308
rect 415 274 449 308
rect 483 292 596 308
rect 732 292 766 390
rect 483 274 766 292
rect 835 340 935 356
rect 835 306 851 340
rect 885 306 935 340
rect 835 290 935 306
rect 969 340 1223 356
rect 969 306 985 340
rect 1019 306 1223 340
rect 969 290 1223 306
rect 297 258 766 274
rect 229 208 442 224
rect 17 168 45 202
rect 79 168 95 202
rect 17 120 95 168
rect 17 86 45 120
rect 79 86 95 120
rect 17 70 95 86
rect 129 168 145 202
rect 179 168 195 202
rect 129 116 195 168
rect 129 82 145 116
rect 179 82 195 116
rect 129 17 195 82
rect 229 174 234 208
rect 268 190 408 208
rect 229 120 268 174
rect 392 174 408 190
rect 229 86 234 120
rect 229 70 268 86
rect 306 130 356 156
rect 306 96 322 130
rect 306 17 356 96
rect 392 120 442 174
rect 392 86 408 120
rect 392 70 442 86
rect 478 208 528 224
rect 478 174 494 208
rect 478 120 528 174
rect 478 86 494 120
rect 478 17 528 86
rect 562 85 596 258
rect 800 240 1225 256
rect 800 224 1002 240
rect 630 222 1002 224
rect 630 190 866 222
rect 630 188 664 190
rect 800 156 816 190
rect 850 156 866 190
rect 986 206 1002 222
rect 1036 222 1174 240
rect 630 119 664 154
rect 700 140 766 156
rect 700 106 716 140
rect 750 106 766 140
rect 800 121 866 156
rect 900 171 950 188
rect 900 137 916 171
rect 700 85 766 106
rect 562 51 766 85
rect 900 17 950 137
rect 986 171 1036 206
rect 1158 206 1174 222
rect 1208 206 1225 240
rect 986 137 1002 171
rect 986 121 1036 137
rect 1072 171 1122 188
rect 1072 137 1088 171
rect 1072 17 1122 137
rect 1158 171 1225 206
rect 1158 137 1174 171
rect 1208 137 1225 171
rect 1158 121 1225 137
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
<< metal1 >>
rect 0 683 1248 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 0 617 1248 649
rect 0 17 1248 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
rect 0 -49 1248 -17
<< labels >>
flabel pwell s 0 0 1248 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 1248 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
rlabel comment s 0 0 0 0 4 o21ba_4
flabel metal1 s 0 617 1248 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 1248 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 1183 316 1217 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 127 242 161 276 0 FreeSans 340 0 0 0 B1_N
port 3 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 223 390 257 424 0 FreeSans 340 0 0 0 X
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 1248 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1101342
string GDS_START 1091676
<< end >>
