magic
tech sky130A
magscale 1 2
timestamp 1599588209
<< nwell >>
rect -38 332 1670 704
rect 925 316 1139 332
<< pwell >>
rect 0 0 1632 49
<< scpmos >>
rect 120 424 150 592
rect 220 424 250 592
rect 432 392 462 560
rect 541 392 571 592
rect 625 392 655 592
rect 775 392 805 476
rect 872 392 902 476
rect 1017 352 1047 576
rect 1216 368 1246 592
rect 1317 424 1347 592
rect 1516 368 1546 592
<< nmoslvt >>
rect 84 120 114 230
rect 202 82 232 230
rect 429 80 459 228
rect 545 79 575 207
rect 623 79 653 207
rect 822 123 852 207
rect 900 123 930 207
rect 1014 74 1044 222
rect 1219 74 1249 222
rect 1321 112 1351 222
rect 1519 74 1549 222
<< ndiff >>
rect 27 184 84 230
rect 27 150 39 184
rect 73 150 84 184
rect 27 120 84 150
rect 114 120 202 230
rect 129 82 202 120
rect 232 218 289 230
rect 232 184 243 218
rect 277 184 289 218
rect 232 82 289 184
rect 343 218 429 228
rect 343 184 369 218
rect 403 184 429 218
rect 129 48 141 82
rect 175 48 187 82
rect 343 80 429 184
rect 459 207 509 228
rect 964 207 1014 222
rect 459 82 545 207
rect 459 80 484 82
rect 129 36 187 48
rect 474 48 484 80
rect 518 79 545 82
rect 575 79 623 207
rect 653 195 822 207
rect 653 161 684 195
rect 718 161 777 195
rect 811 161 822 195
rect 653 123 822 161
rect 852 123 900 207
rect 930 192 1014 207
rect 930 158 957 192
rect 991 158 1014 192
rect 930 124 1014 158
rect 930 123 957 124
rect 653 79 703 123
rect 518 48 530 79
rect 474 36 530 48
rect 945 90 957 123
rect 991 90 1014 124
rect 945 74 1014 90
rect 1044 192 1103 222
rect 1044 158 1057 192
rect 1091 158 1103 192
rect 1044 124 1103 158
rect 1044 90 1057 124
rect 1091 90 1103 124
rect 1044 74 1103 90
rect 1162 204 1219 222
rect 1162 170 1174 204
rect 1208 170 1219 204
rect 1162 120 1219 170
rect 1162 86 1174 120
rect 1208 86 1219 120
rect 1162 74 1219 86
rect 1249 195 1321 222
rect 1249 161 1269 195
rect 1303 161 1321 195
rect 1249 112 1321 161
rect 1351 184 1408 222
rect 1351 150 1362 184
rect 1396 150 1408 184
rect 1351 112 1408 150
rect 1462 210 1519 222
rect 1462 176 1474 210
rect 1508 176 1519 210
rect 1462 120 1519 176
rect 1249 74 1299 112
rect 1462 86 1474 120
rect 1508 86 1519 120
rect 1462 74 1519 86
rect 1549 210 1605 222
rect 1549 176 1560 210
rect 1594 176 1605 210
rect 1549 120 1605 176
rect 1549 86 1560 120
rect 1594 86 1605 120
rect 1549 74 1605 86
<< pdiff >>
rect 50 580 120 592
rect 50 546 59 580
rect 93 546 120 580
rect 50 470 120 546
rect 50 436 59 470
rect 93 436 120 470
rect 50 424 120 436
rect 150 580 220 592
rect 150 546 163 580
rect 197 546 220 580
rect 150 498 220 546
rect 150 464 163 498
rect 197 464 220 498
rect 150 424 220 464
rect 250 580 309 592
rect 250 546 263 580
rect 297 546 309 580
rect 480 580 541 592
rect 480 560 492 580
rect 250 498 309 546
rect 250 464 263 498
rect 297 464 309 498
rect 250 424 309 464
rect 373 441 432 560
rect 373 407 385 441
rect 419 407 432 441
rect 373 392 432 407
rect 462 546 492 560
rect 526 546 541 580
rect 462 392 541 546
rect 571 392 625 592
rect 655 476 708 592
rect 1160 580 1216 592
rect 958 564 1017 576
rect 958 530 970 564
rect 1004 530 1017 564
rect 958 476 1017 530
rect 655 444 775 476
rect 655 410 689 444
rect 723 410 775 444
rect 655 392 775 410
rect 805 392 872 476
rect 902 452 1017 476
rect 902 418 933 452
rect 967 418 1017 452
rect 902 392 1017 418
rect 961 352 1017 392
rect 1047 564 1103 576
rect 1047 530 1060 564
rect 1094 530 1103 564
rect 1047 481 1103 530
rect 1047 447 1060 481
rect 1094 447 1103 481
rect 1047 398 1103 447
rect 1047 364 1060 398
rect 1094 364 1103 398
rect 1160 546 1169 580
rect 1203 546 1216 580
rect 1160 497 1216 546
rect 1160 463 1169 497
rect 1203 463 1216 497
rect 1160 414 1216 463
rect 1160 380 1169 414
rect 1203 380 1216 414
rect 1160 368 1216 380
rect 1246 580 1317 592
rect 1246 546 1260 580
rect 1294 546 1317 580
rect 1246 470 1317 546
rect 1246 436 1260 470
rect 1294 436 1317 470
rect 1246 424 1317 436
rect 1347 580 1406 592
rect 1347 546 1361 580
rect 1395 546 1406 580
rect 1347 470 1406 546
rect 1347 436 1361 470
rect 1395 436 1406 470
rect 1347 424 1406 436
rect 1460 580 1516 592
rect 1460 546 1469 580
rect 1503 546 1516 580
rect 1460 497 1516 546
rect 1460 463 1469 497
rect 1503 463 1516 497
rect 1246 368 1299 424
rect 1460 414 1516 463
rect 1047 352 1103 364
rect 1460 380 1469 414
rect 1503 380 1516 414
rect 1460 368 1516 380
rect 1546 580 1605 592
rect 1546 546 1559 580
rect 1593 546 1605 580
rect 1546 497 1605 546
rect 1546 463 1559 497
rect 1593 463 1605 497
rect 1546 414 1605 463
rect 1546 380 1559 414
rect 1593 380 1605 414
rect 1546 368 1605 380
<< ndiffc >>
rect 39 150 73 184
rect 243 184 277 218
rect 369 184 403 218
rect 141 48 175 82
rect 484 48 518 82
rect 684 161 718 195
rect 777 161 811 195
rect 957 158 991 192
rect 957 90 991 124
rect 1057 158 1091 192
rect 1057 90 1091 124
rect 1174 170 1208 204
rect 1174 86 1208 120
rect 1269 161 1303 195
rect 1362 150 1396 184
rect 1474 176 1508 210
rect 1474 86 1508 120
rect 1560 176 1594 210
rect 1560 86 1594 120
<< pdiffc >>
rect 59 546 93 580
rect 59 436 93 470
rect 163 546 197 580
rect 163 464 197 498
rect 263 546 297 580
rect 263 464 297 498
rect 385 407 419 441
rect 492 546 526 580
rect 970 530 1004 564
rect 689 410 723 444
rect 933 418 967 452
rect 1060 530 1094 564
rect 1060 447 1094 481
rect 1060 364 1094 398
rect 1169 546 1203 580
rect 1169 463 1203 497
rect 1169 380 1203 414
rect 1260 546 1294 580
rect 1260 436 1294 470
rect 1361 546 1395 580
rect 1361 436 1395 470
rect 1469 546 1503 580
rect 1469 463 1503 497
rect 1469 380 1503 414
rect 1559 546 1593 580
rect 1559 463 1593 497
rect 1559 380 1593 414
<< poly >>
rect 120 592 150 618
rect 220 592 250 618
rect 541 592 571 618
rect 625 592 655 618
rect 432 560 462 586
rect 120 409 150 424
rect 220 409 250 424
rect 117 386 153 409
rect 217 392 253 409
rect 1017 576 1047 602
rect 1216 592 1246 618
rect 1317 592 1347 618
rect 1516 592 1546 618
rect 775 476 805 502
rect 872 476 902 502
rect 84 370 153 386
rect 84 336 103 370
rect 137 336 153 370
rect 84 302 153 336
rect 201 376 267 392
rect 432 377 462 392
rect 541 377 571 392
rect 625 377 655 392
rect 775 377 805 392
rect 872 377 902 392
rect 201 342 217 376
rect 251 342 267 376
rect 201 326 267 342
rect 84 268 103 302
rect 137 268 153 302
rect 84 252 153 268
rect 84 230 114 252
rect 202 230 232 326
rect 315 300 381 316
rect 315 266 331 300
rect 365 280 381 300
rect 429 280 465 377
rect 538 316 574 377
rect 622 360 658 377
rect 772 360 808 377
rect 869 360 905 377
rect 617 344 683 360
rect 365 266 465 280
rect 315 250 465 266
rect 507 300 575 316
rect 507 266 523 300
rect 557 266 575 300
rect 617 310 633 344
rect 667 310 683 344
rect 617 294 683 310
rect 744 344 821 360
rect 744 310 771 344
rect 805 310 821 344
rect 744 294 821 310
rect 863 344 930 360
rect 1317 409 1347 424
rect 1216 353 1246 368
rect 863 310 879 344
rect 913 310 930 344
rect 1017 337 1047 352
rect 1014 310 1050 337
rect 1213 320 1249 353
rect 1314 320 1350 409
rect 1516 353 1546 368
rect 1513 326 1549 353
rect 863 294 930 310
rect 507 250 575 266
rect 744 252 774 294
rect 84 94 114 120
rect 429 228 459 250
rect 202 56 232 82
rect 545 207 575 250
rect 623 222 774 252
rect 623 207 653 222
rect 822 207 852 233
rect 900 207 930 294
rect 978 294 1050 310
rect 978 260 994 294
rect 1028 260 1050 294
rect 978 244 1050 260
rect 1092 304 1350 320
rect 1092 270 1108 304
rect 1142 270 1350 304
rect 1092 267 1350 270
rect 1434 310 1549 326
rect 1434 276 1450 310
rect 1484 276 1549 310
rect 1092 254 1351 267
rect 1434 260 1549 276
rect 1014 222 1044 244
rect 1219 237 1351 254
rect 1219 222 1249 237
rect 1321 222 1351 237
rect 1519 222 1549 260
rect 429 54 459 80
rect 822 101 852 123
rect 786 85 852 101
rect 900 97 930 123
rect 545 53 575 79
rect 623 53 653 79
rect 786 51 802 85
rect 836 51 852 85
rect 1321 86 1351 112
rect 786 35 852 51
rect 1014 48 1044 74
rect 1219 48 1249 74
rect 1519 48 1549 74
<< polycont >>
rect 103 336 137 370
rect 217 342 251 376
rect 103 268 137 302
rect 331 266 365 300
rect 523 266 557 300
rect 633 310 667 344
rect 771 310 805 344
rect 879 310 913 344
rect 994 260 1028 294
rect 1108 270 1142 304
rect 1450 276 1484 310
rect 802 51 836 85
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 19 580 109 596
rect 19 546 59 580
rect 93 546 109 580
rect 19 470 109 546
rect 19 436 59 470
rect 93 436 109 470
rect 147 580 213 649
rect 147 546 163 580
rect 197 546 213 580
rect 147 498 213 546
rect 147 464 163 498
rect 197 464 213 498
rect 247 580 313 596
rect 247 546 263 580
rect 297 546 313 580
rect 476 580 542 649
rect 476 546 492 580
rect 526 546 542 580
rect 896 564 1004 649
rect 1153 580 1226 596
rect 247 512 313 546
rect 896 530 970 564
rect 247 498 829 512
rect 247 464 263 498
rect 297 478 829 498
rect 297 464 335 478
rect 19 420 109 436
rect 19 218 53 420
rect 87 370 167 386
rect 87 336 103 370
rect 137 336 167 370
rect 201 376 267 430
rect 201 342 217 376
rect 251 342 267 376
rect 201 338 267 342
rect 87 302 167 336
rect 301 304 335 464
rect 369 441 582 444
rect 369 407 385 441
rect 419 407 582 441
rect 652 410 689 444
rect 723 410 761 444
rect 369 376 582 407
rect 415 344 668 376
rect 415 342 633 344
rect 87 268 103 302
rect 137 268 167 302
rect 87 252 167 268
rect 227 300 381 304
rect 227 266 331 300
rect 365 266 381 300
rect 227 252 381 266
rect 227 218 293 252
rect 415 218 449 342
rect 607 310 633 342
rect 667 310 668 344
rect 19 184 89 218
rect 227 184 243 218
rect 277 184 293 218
rect 339 184 369 218
rect 403 184 449 218
rect 507 300 573 302
rect 507 266 523 300
rect 557 266 573 300
rect 19 150 39 184
rect 73 150 89 184
rect 507 150 573 266
rect 19 116 573 150
rect 607 294 668 310
rect 607 101 641 294
rect 702 260 736 410
rect 795 360 829 478
rect 896 452 1004 530
rect 896 418 933 452
rect 967 418 1004 452
rect 896 412 1004 418
rect 1044 564 1112 580
rect 1044 530 1060 564
rect 1094 530 1112 564
rect 1044 481 1112 530
rect 1044 447 1060 481
rect 1094 447 1112 481
rect 1044 398 1112 447
rect 1044 378 1060 398
rect 770 344 829 360
rect 770 310 771 344
rect 805 310 829 344
rect 770 294 829 310
rect 863 364 1060 378
rect 1094 364 1112 398
rect 1153 546 1169 580
rect 1203 546 1226 580
rect 1153 497 1226 546
rect 1153 463 1169 497
rect 1203 463 1226 497
rect 1153 414 1226 463
rect 1260 580 1310 649
rect 1294 546 1310 580
rect 1260 470 1310 546
rect 1294 436 1310 470
rect 1260 420 1310 436
rect 1344 580 1413 596
rect 1344 546 1361 580
rect 1395 546 1413 580
rect 1344 470 1413 546
rect 1344 436 1361 470
rect 1395 436 1413 470
rect 1153 380 1169 414
rect 1203 380 1226 414
rect 1153 364 1226 380
rect 863 344 1112 364
rect 863 310 879 344
rect 913 310 929 344
rect 1078 320 1112 344
rect 863 294 929 310
rect 978 294 1044 310
rect 978 260 994 294
rect 1028 260 1044 294
rect 702 226 1044 260
rect 1078 304 1158 320
rect 1078 270 1108 304
rect 1142 270 1158 304
rect 1078 254 1158 270
rect 702 211 827 226
rect 675 195 827 211
rect 675 161 684 195
rect 718 161 777 195
rect 811 161 827 195
rect 1078 192 1112 254
rect 1192 220 1226 364
rect 1344 326 1413 436
rect 1453 580 1503 649
rect 1453 546 1469 580
rect 1453 497 1503 546
rect 1453 463 1469 497
rect 1453 414 1503 463
rect 1453 380 1469 414
rect 1453 364 1503 380
rect 1543 580 1610 596
rect 1543 546 1559 580
rect 1593 546 1610 580
rect 1543 497 1610 546
rect 1543 463 1559 497
rect 1593 463 1610 497
rect 1543 414 1610 463
rect 1543 380 1559 414
rect 1593 380 1610 414
rect 1344 310 1500 326
rect 1344 276 1450 310
rect 1484 276 1500 310
rect 1344 260 1500 276
rect 675 145 827 161
rect 941 158 957 192
rect 991 158 1007 192
rect 941 124 1007 158
rect 607 85 852 101
rect 125 48 141 82
rect 175 48 191 82
rect 125 17 191 48
rect 468 48 484 82
rect 518 48 535 82
rect 607 51 802 85
rect 836 51 852 85
rect 941 90 957 124
rect 991 90 1007 124
rect 468 17 535 48
rect 941 17 1007 90
rect 1041 158 1057 192
rect 1091 158 1112 192
rect 1041 124 1112 158
rect 1041 90 1057 124
rect 1091 90 1112 124
rect 1041 70 1112 90
rect 1158 204 1226 220
rect 1158 170 1174 204
rect 1208 170 1226 204
rect 1158 120 1226 170
rect 1158 86 1174 120
rect 1208 86 1226 120
rect 1158 70 1226 86
rect 1260 195 1310 226
rect 1260 161 1269 195
rect 1303 161 1310 195
rect 1260 17 1310 161
rect 1344 184 1412 260
rect 1344 150 1362 184
rect 1396 150 1412 184
rect 1344 108 1412 150
rect 1458 210 1508 226
rect 1458 176 1474 210
rect 1458 120 1508 176
rect 1458 86 1474 120
rect 1458 17 1508 86
rect 1543 210 1610 380
rect 1543 176 1560 210
rect 1594 176 1610 210
rect 1543 120 1610 176
rect 1543 86 1560 120
rect 1594 86 1610 120
rect 1543 70 1610 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dlxbn_1
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nwell s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 1 nsew
flabel corelocali s 1567 94 1601 128 0 FreeSans 340 0 0 0 Q_N
port 8 nsew
flabel corelocali s 1567 168 1601 202 0 FreeSans 340 0 0 0 Q_N
port 8 nsew
flabel corelocali s 1567 242 1601 276 0 FreeSans 340 0 0 0 Q_N
port 8 nsew
flabel corelocali s 1567 316 1601 350 0 FreeSans 340 0 0 0 Q_N
port 8 nsew
flabel corelocali s 1567 390 1601 424 0 FreeSans 340 0 0 0 Q_N
port 8 nsew
flabel corelocali s 1567 464 1601 498 0 FreeSans 340 0 0 0 Q_N
port 8 nsew
flabel corelocali s 1567 538 1601 572 0 FreeSans 340 0 0 0 Q_N
port 8 nsew
flabel corelocali s 1183 94 1217 128 0 FreeSans 340 0 0 0 Q
port 7 nsew
flabel corelocali s 1183 168 1217 202 0 FreeSans 340 0 0 0 Q
port 7 nsew
flabel corelocali s 223 390 257 424 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 1632 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 2201714
string GDS_START 2188728
<< end >>
