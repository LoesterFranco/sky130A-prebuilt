magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1472 561
rect 115 367 165 527
rect 283 367 333 527
rect 451 367 501 527
rect 619 367 669 527
rect 787 323 837 425
rect 955 323 1005 425
rect 1123 323 1173 425
rect 1291 323 1341 425
rect 787 289 1455 323
rect 72 215 706 255
rect 760 215 1308 255
rect 1342 181 1455 289
rect 18 17 73 181
rect 107 145 1455 181
rect 107 51 173 145
rect 207 17 241 111
rect 275 51 341 145
rect 375 17 409 111
rect 443 51 509 145
rect 543 17 577 111
rect 611 51 677 145
rect 711 17 745 111
rect 779 51 845 145
rect 879 17 913 111
rect 947 51 1013 145
rect 1047 17 1081 111
rect 1115 51 1181 145
rect 1215 17 1249 111
rect 1283 51 1349 145
rect 1383 17 1441 111
rect 0 -17 1472 17
<< obsli1 >>
rect 18 333 81 493
rect 199 333 249 493
rect 367 333 417 493
rect 535 333 585 493
rect 703 459 1425 493
rect 703 333 753 459
rect 18 291 753 333
rect 871 357 921 459
rect 1039 357 1089 459
rect 1207 357 1257 459
rect 1375 357 1425 459
<< metal1 >>
rect 0 496 1472 592
rect 0 -48 1472 48
<< labels >>
rlabel locali s 72 215 706 255 6 A
port 1 nsew signal input
rlabel locali s 760 215 1308 255 6 B
port 2 nsew signal input
rlabel locali s 1342 181 1455 289 6 Y
port 3 nsew signal output
rlabel locali s 1291 323 1341 425 6 Y
port 3 nsew signal output
rlabel locali s 1283 51 1349 145 6 Y
port 3 nsew signal output
rlabel locali s 1123 323 1173 425 6 Y
port 3 nsew signal output
rlabel locali s 1115 51 1181 145 6 Y
port 3 nsew signal output
rlabel locali s 955 323 1005 425 6 Y
port 3 nsew signal output
rlabel locali s 947 51 1013 145 6 Y
port 3 nsew signal output
rlabel locali s 787 323 837 425 6 Y
port 3 nsew signal output
rlabel locali s 787 289 1455 323 6 Y
port 3 nsew signal output
rlabel locali s 779 51 845 145 6 Y
port 3 nsew signal output
rlabel locali s 611 51 677 145 6 Y
port 3 nsew signal output
rlabel locali s 443 51 509 145 6 Y
port 3 nsew signal output
rlabel locali s 275 51 341 145 6 Y
port 3 nsew signal output
rlabel locali s 107 145 1455 181 6 Y
port 3 nsew signal output
rlabel locali s 107 51 173 145 6 Y
port 3 nsew signal output
rlabel locali s 1383 17 1441 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 1215 17 1249 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 1047 17 1081 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 879 17 913 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 711 17 745 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 543 17 577 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 375 17 409 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 207 17 241 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 18 17 73 181 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 1472 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1472 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 619 367 669 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 451 367 501 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 283 367 333 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 115 367 165 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 1472 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 1472 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1472 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1949518
string GDS_START 1938120
<< end >>
