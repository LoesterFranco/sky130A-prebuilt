magic
tech sky130A
magscale 1 2
timestamp 1601050056
<< nwell >>
rect -38 332 518 704
<< pwell >>
rect 0 0 480 49
<< scpmos >>
rect 83 368 119 536
rect 217 368 253 592
rect 317 368 353 592
<< nmoslvt >>
rect 84 112 114 222
rect 239 74 269 222
rect 317 74 347 222
<< ndiff >>
rect 27 184 84 222
rect 27 150 39 184
rect 73 150 84 184
rect 27 112 84 150
rect 114 158 239 222
rect 114 124 126 158
rect 160 124 194 158
rect 228 124 239 158
rect 114 112 239 124
rect 129 74 239 112
rect 269 74 317 222
rect 347 210 433 222
rect 347 176 371 210
rect 405 176 433 210
rect 347 120 433 176
rect 347 86 371 120
rect 405 86 433 120
rect 347 74 433 86
<< pdiff >>
rect 134 576 217 592
rect 134 542 147 576
rect 181 542 217 576
rect 134 536 217 542
rect 27 524 83 536
rect 27 490 39 524
rect 73 490 83 524
rect 27 440 83 490
rect 27 406 39 440
rect 73 406 83 440
rect 27 368 83 406
rect 119 508 217 536
rect 119 474 147 508
rect 181 474 217 508
rect 119 368 217 474
rect 253 580 317 592
rect 253 546 263 580
rect 297 546 317 580
rect 253 508 317 546
rect 253 474 263 508
rect 297 474 317 508
rect 253 368 317 474
rect 353 580 410 592
rect 353 546 363 580
rect 397 546 410 580
rect 353 368 410 546
<< ndiffc >>
rect 39 150 73 184
rect 126 124 160 158
rect 194 124 228 158
rect 371 176 405 210
rect 371 86 405 120
<< pdiffc >>
rect 147 542 181 576
rect 39 490 73 524
rect 39 406 73 440
rect 147 474 181 508
rect 263 546 297 580
rect 263 474 297 508
rect 363 546 397 580
<< poly >>
rect 217 592 253 618
rect 317 592 353 618
rect 83 536 119 562
rect 83 326 119 368
rect 217 336 253 368
rect 21 310 155 326
rect 21 276 37 310
rect 71 276 105 310
rect 139 276 155 310
rect 21 260 155 276
rect 203 320 269 336
rect 203 286 219 320
rect 253 286 269 320
rect 203 270 269 286
rect 84 222 114 260
rect 239 222 269 270
rect 317 326 353 368
rect 317 310 383 326
rect 317 276 333 310
rect 367 276 383 310
rect 317 260 383 276
rect 317 222 347 260
rect 84 86 114 112
rect 239 48 269 74
rect 317 48 347 74
<< polycont >>
rect 37 276 71 310
rect 105 276 139 310
rect 219 286 253 320
rect 333 276 367 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 130 576 183 649
rect 130 542 147 576
rect 181 542 183 576
rect 23 524 89 540
rect 23 490 39 524
rect 73 490 89 524
rect 23 440 89 490
rect 130 508 183 542
rect 130 474 147 508
rect 181 474 183 508
rect 130 458 183 474
rect 217 580 313 596
rect 217 546 263 580
rect 297 546 313 580
rect 217 508 313 546
rect 347 580 414 649
rect 347 546 363 580
rect 397 546 414 580
rect 347 530 414 546
rect 217 474 263 508
rect 297 492 313 508
rect 297 474 451 492
rect 217 458 451 474
rect 23 406 39 440
rect 73 424 89 440
rect 73 406 337 424
rect 23 390 337 406
rect 21 310 167 356
rect 21 276 37 310
rect 71 276 105 310
rect 139 276 167 310
rect 21 260 167 276
rect 203 320 269 356
rect 203 286 219 320
rect 253 286 269 320
rect 203 270 269 286
rect 303 326 337 390
rect 303 310 383 326
rect 303 276 333 310
rect 367 276 383 310
rect 303 260 383 276
rect 303 226 337 260
rect 417 226 451 458
rect 23 192 337 226
rect 371 210 451 226
rect 23 184 76 192
rect 23 150 39 184
rect 73 150 76 184
rect 405 176 451 210
rect 23 108 76 150
rect 110 124 126 158
rect 160 124 194 158
rect 228 124 244 158
rect 110 17 244 124
rect 371 120 451 176
rect 405 86 451 120
rect 371 70 451 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< metal1 >>
rect 0 683 480 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 0 617 480 649
rect 0 17 480 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
rect 0 -49 480 -17
<< labels >>
flabel pwell s 0 0 480 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 0 617 480 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
rlabel comment s 0 0 0 0 4 nand2b_1
flabel metal1 s 0 617 480 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 480 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 223 464 257 498 0 FreeSans 340 0 0 0 Y
port 7 nsew
flabel corelocali s 223 538 257 572 0 FreeSans 340 0 0 0 Y
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 480 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 2008040
string GDS_START 2003424
<< end >>
