magic
tech sky130A
magscale 1 2
timestamp 1601050088
<< locali >>
rect 85 196 161 398
rect 303 222 369 288
rect 690 236 756 310
rect 2415 310 2481 596
rect 2415 226 2469 310
rect 2403 70 2469 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2592 683
rect 17 470 87 596
rect 189 504 239 649
rect 273 581 443 615
rect 273 470 307 581
rect 17 436 307 470
rect 17 162 51 436
rect 195 356 261 402
rect 341 356 375 547
rect 409 424 443 581
rect 477 458 527 649
rect 734 530 800 649
rect 1004 530 1054 649
rect 1199 538 1249 596
rect 620 496 695 524
rect 1088 504 1249 538
rect 1283 504 1355 596
rect 1482 550 1548 649
rect 1701 550 1767 649
rect 1088 496 1122 504
rect 620 462 1122 496
rect 620 424 695 462
rect 409 390 654 424
rect 195 322 477 356
rect 195 188 261 322
rect 411 277 477 322
rect 511 209 586 356
rect 17 68 106 162
rect 195 154 364 188
rect 620 175 654 390
rect 790 294 980 428
rect 1026 330 1060 462
rect 1165 428 1249 460
rect 1094 394 1249 428
rect 1094 364 1199 394
rect 1026 296 1131 330
rect 790 202 824 294
rect 204 17 270 120
rect 314 83 364 154
rect 400 17 466 175
rect 558 83 654 175
rect 688 17 722 202
rect 758 70 824 202
rect 867 17 917 226
rect 953 85 1019 226
rect 1065 119 1131 296
rect 1165 85 1199 364
rect 1283 360 1317 504
rect 1389 482 1960 516
rect 1389 466 1423 482
rect 1351 400 1423 466
rect 1589 414 1688 448
rect 1540 360 1606 366
rect 1233 326 1606 360
rect 1233 153 1267 326
rect 1540 323 1606 326
rect 1654 321 1688 414
rect 1926 345 1960 482
rect 1994 419 2044 600
rect 2169 505 2277 649
rect 2311 464 2377 590
rect 2133 419 2377 464
rect 1994 385 2081 419
rect 2047 351 2189 385
rect 1426 289 1492 292
rect 1654 289 1788 321
rect 1301 221 1392 262
rect 1426 255 1788 289
rect 1822 275 1892 310
rect 1926 309 2013 345
rect 2055 275 2121 317
rect 1301 187 1552 221
rect 1233 119 1324 153
rect 1358 85 1392 187
rect 953 51 1392 85
rect 1434 17 1484 153
rect 1518 85 1552 187
rect 1586 119 1620 255
rect 1822 241 2121 275
rect 2155 267 2189 351
rect 2329 310 2377 419
rect 2521 364 2571 649
rect 1822 221 1856 241
rect 1654 187 1856 221
rect 2155 201 2301 267
rect 1654 85 1688 187
rect 1890 167 2189 201
rect 1518 51 1688 85
rect 1722 17 1772 153
rect 1890 70 1956 167
rect 2335 162 2369 310
rect 2070 17 2262 133
rect 2298 67 2369 162
rect 2503 17 2569 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2592 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
<< metal1 >>
rect 0 683 2592 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2592 683
rect 0 617 2592 649
rect 0 17 2592 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2592 17
rect 0 -49 2592 -17
<< obsm1 >>
rect 499 347 557 356
rect 2323 347 2381 356
rect 499 319 2381 347
rect 499 310 557 319
rect 2323 310 2381 319
<< labels >>
rlabel locali s 85 196 161 398 6 D
port 1 nsew signal input
rlabel locali s 303 222 369 288 6 DE
port 2 nsew signal input
rlabel locali s 2415 310 2481 596 6 Q
port 3 nsew signal output
rlabel locali s 2415 226 2469 310 6 Q
port 3 nsew signal output
rlabel locali s 2403 70 2469 226 6 Q
port 3 nsew signal output
rlabel locali s 690 236 756 310 6 CLK
port 4 nsew clock input
rlabel metal1 s 0 -49 2592 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 617 2592 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2592 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 2310562
string GDS_START 2292598
<< end >>
