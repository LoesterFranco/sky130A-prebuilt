magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 1190 704
<< pwell >>
rect 0 0 1152 49
<< scnmos >>
rect 97 74 127 222
rect 183 74 213 222
rect 269 74 299 222
rect 369 74 399 222
rect 567 74 597 222
rect 667 74 697 222
rect 753 74 783 222
rect 843 74 873 222
rect 929 74 959 222
rect 1029 74 1059 222
<< pmoshvt >>
rect 94 368 124 592
rect 184 368 214 592
rect 284 368 314 592
rect 374 368 404 592
rect 464 368 494 592
rect 554 368 584 592
rect 756 368 786 592
rect 846 368 876 592
rect 936 368 966 592
rect 1036 368 1066 592
<< ndiff >>
rect 40 202 97 222
rect 40 168 52 202
rect 86 168 97 202
rect 40 120 97 168
rect 40 86 52 120
rect 86 86 97 120
rect 40 74 97 86
rect 127 189 183 222
rect 127 155 138 189
rect 172 155 183 189
rect 127 74 183 155
rect 213 210 269 222
rect 213 176 224 210
rect 258 176 269 210
rect 213 120 269 176
rect 213 86 224 120
rect 258 86 269 120
rect 213 74 269 86
rect 299 127 369 222
rect 299 93 310 127
rect 344 93 369 127
rect 299 74 369 93
rect 399 189 456 222
rect 399 155 410 189
rect 444 155 456 189
rect 399 74 456 155
rect 510 189 567 222
rect 510 155 522 189
rect 556 155 567 189
rect 510 74 567 155
rect 597 144 667 222
rect 597 110 622 144
rect 656 110 667 144
rect 597 74 667 110
rect 697 210 753 222
rect 697 176 708 210
rect 742 176 753 210
rect 697 120 753 176
rect 697 86 708 120
rect 742 86 753 120
rect 697 74 753 86
rect 783 136 843 222
rect 783 102 794 136
rect 828 102 843 136
rect 783 74 843 102
rect 873 210 929 222
rect 873 176 884 210
rect 918 176 929 210
rect 873 120 929 176
rect 873 86 884 120
rect 918 86 929 120
rect 873 74 929 86
rect 959 136 1029 222
rect 959 102 984 136
rect 1018 102 1029 136
rect 959 74 1029 102
rect 1059 210 1116 222
rect 1059 176 1070 210
rect 1104 176 1116 210
rect 1059 120 1116 176
rect 1059 86 1070 120
rect 1104 86 1116 120
rect 1059 74 1116 86
<< pdiff >>
rect 35 580 94 592
rect 35 546 47 580
rect 81 546 94 580
rect 35 497 94 546
rect 35 463 47 497
rect 81 463 94 497
rect 35 414 94 463
rect 35 380 47 414
rect 81 380 94 414
rect 35 368 94 380
rect 124 580 184 592
rect 124 546 137 580
rect 171 546 184 580
rect 124 497 184 546
rect 124 463 137 497
rect 171 463 184 497
rect 124 414 184 463
rect 124 380 137 414
rect 171 380 184 414
rect 124 368 184 380
rect 214 580 284 592
rect 214 546 237 580
rect 271 546 284 580
rect 214 478 284 546
rect 214 444 237 478
rect 271 444 284 478
rect 214 368 284 444
rect 314 580 374 592
rect 314 546 327 580
rect 361 546 374 580
rect 314 497 374 546
rect 314 463 327 497
rect 361 463 374 497
rect 314 414 374 463
rect 314 380 327 414
rect 361 380 374 414
rect 314 368 374 380
rect 404 580 464 592
rect 404 546 417 580
rect 451 546 464 580
rect 404 508 464 546
rect 404 474 417 508
rect 451 474 464 508
rect 404 368 464 474
rect 494 580 554 592
rect 494 546 507 580
rect 541 546 554 580
rect 494 510 554 546
rect 494 476 507 510
rect 541 476 554 510
rect 494 440 554 476
rect 494 406 507 440
rect 541 406 554 440
rect 494 368 554 406
rect 584 580 643 592
rect 584 546 597 580
rect 631 546 643 580
rect 584 508 643 546
rect 584 474 597 508
rect 631 474 643 508
rect 584 368 643 474
rect 697 580 756 592
rect 697 546 709 580
rect 743 546 756 580
rect 697 508 756 546
rect 697 474 709 508
rect 743 474 756 508
rect 697 368 756 474
rect 786 531 846 592
rect 786 497 799 531
rect 833 497 846 531
rect 786 440 846 497
rect 786 406 799 440
rect 833 406 846 440
rect 786 368 846 406
rect 876 580 936 592
rect 876 546 889 580
rect 923 546 936 580
rect 876 510 936 546
rect 876 476 889 510
rect 923 476 936 510
rect 876 440 936 476
rect 876 406 889 440
rect 923 406 936 440
rect 876 368 936 406
rect 966 580 1036 592
rect 966 546 979 580
rect 1013 546 1036 580
rect 966 508 1036 546
rect 966 474 979 508
rect 1013 474 1036 508
rect 966 368 1036 474
rect 1066 580 1125 592
rect 1066 546 1079 580
rect 1113 546 1125 580
rect 1066 510 1125 546
rect 1066 476 1079 510
rect 1113 476 1125 510
rect 1066 440 1125 476
rect 1066 406 1079 440
rect 1113 406 1125 440
rect 1066 368 1125 406
<< ndiffc >>
rect 52 168 86 202
rect 52 86 86 120
rect 138 155 172 189
rect 224 176 258 210
rect 224 86 258 120
rect 310 93 344 127
rect 410 155 444 189
rect 522 155 556 189
rect 622 110 656 144
rect 708 176 742 210
rect 708 86 742 120
rect 794 102 828 136
rect 884 176 918 210
rect 884 86 918 120
rect 984 102 1018 136
rect 1070 176 1104 210
rect 1070 86 1104 120
<< pdiffc >>
rect 47 546 81 580
rect 47 463 81 497
rect 47 380 81 414
rect 137 546 171 580
rect 137 463 171 497
rect 137 380 171 414
rect 237 546 271 580
rect 237 444 271 478
rect 327 546 361 580
rect 327 463 361 497
rect 327 380 361 414
rect 417 546 451 580
rect 417 474 451 508
rect 507 546 541 580
rect 507 476 541 510
rect 507 406 541 440
rect 597 546 631 580
rect 597 474 631 508
rect 709 546 743 580
rect 709 474 743 508
rect 799 497 833 531
rect 799 406 833 440
rect 889 546 923 580
rect 889 476 923 510
rect 889 406 923 440
rect 979 546 1013 580
rect 979 474 1013 508
rect 1079 546 1113 580
rect 1079 476 1113 510
rect 1079 406 1113 440
<< poly >>
rect 94 592 124 618
rect 184 592 214 618
rect 284 592 314 618
rect 374 592 404 618
rect 464 592 494 618
rect 554 592 584 618
rect 756 592 786 618
rect 846 592 876 618
rect 936 592 966 618
rect 1036 592 1066 618
rect 94 353 124 368
rect 184 353 214 368
rect 284 353 314 368
rect 374 353 404 368
rect 464 353 494 368
rect 554 353 584 368
rect 756 353 786 368
rect 846 353 876 368
rect 936 353 966 368
rect 1036 353 1066 368
rect 91 310 127 353
rect 181 310 217 353
rect 281 326 317 353
rect 371 326 407 353
rect 21 294 217 310
rect 21 260 37 294
rect 71 260 217 294
rect 21 244 217 260
rect 269 310 407 326
rect 269 276 285 310
rect 319 276 353 310
rect 387 276 407 310
rect 461 336 497 353
rect 551 336 587 353
rect 753 336 789 353
rect 843 336 879 353
rect 461 320 697 336
rect 461 306 573 320
rect 269 260 407 276
rect 557 286 573 306
rect 607 286 641 320
rect 675 286 697 320
rect 557 270 697 286
rect 97 222 127 244
rect 183 222 213 244
rect 269 222 299 260
rect 369 222 399 260
rect 567 222 597 270
rect 667 222 697 270
rect 753 320 879 336
rect 753 286 809 320
rect 843 286 879 320
rect 933 333 969 353
rect 1033 336 1069 353
rect 1017 333 1083 336
rect 933 320 1083 333
rect 933 300 1033 320
rect 753 270 879 286
rect 929 286 1033 300
rect 1067 286 1083 320
rect 929 270 1083 286
rect 753 222 783 270
rect 843 222 873 270
rect 929 222 959 270
rect 1029 222 1059 270
rect 97 48 127 74
rect 183 48 213 74
rect 269 48 299 74
rect 369 48 399 74
rect 567 48 597 74
rect 667 48 697 74
rect 753 48 783 74
rect 843 48 873 74
rect 929 48 959 74
rect 1029 48 1059 74
<< polycont >>
rect 37 260 71 294
rect 285 276 319 310
rect 353 276 387 310
rect 573 286 607 320
rect 641 286 675 320
rect 809 286 843 320
rect 1033 286 1067 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 31 580 81 649
rect 31 546 47 580
rect 31 497 81 546
rect 31 463 47 497
rect 31 414 81 463
rect 31 380 47 414
rect 31 364 81 380
rect 121 580 187 596
rect 121 546 137 580
rect 171 546 187 580
rect 121 497 187 546
rect 121 463 137 497
rect 171 463 187 497
rect 121 414 187 463
rect 221 580 271 649
rect 221 546 237 580
rect 221 478 271 546
rect 221 444 237 478
rect 221 428 271 444
rect 311 580 377 596
rect 311 546 327 580
rect 361 546 377 580
rect 311 497 377 546
rect 311 463 327 497
rect 361 463 377 497
rect 121 380 137 414
rect 171 394 187 414
rect 311 424 377 463
rect 417 580 451 649
rect 417 508 451 546
rect 417 458 451 474
rect 491 580 557 596
rect 491 546 507 580
rect 541 546 557 580
rect 491 510 557 546
rect 491 476 507 510
rect 541 476 557 510
rect 491 440 557 476
rect 597 580 647 649
rect 631 546 647 580
rect 597 508 647 546
rect 631 474 647 508
rect 597 458 647 474
rect 693 581 923 615
rect 693 580 743 581
rect 693 546 709 580
rect 889 580 923 581
rect 693 508 743 546
rect 693 474 709 508
rect 693 458 743 474
rect 783 531 849 547
rect 783 497 799 531
rect 833 497 849 531
rect 491 424 507 440
rect 311 414 507 424
rect 311 394 327 414
rect 171 380 327 394
rect 361 406 507 414
rect 541 424 557 440
rect 783 440 849 497
rect 783 424 799 440
rect 541 406 799 424
rect 833 406 849 440
rect 361 390 849 406
rect 889 510 923 546
rect 889 440 923 476
rect 963 580 1029 649
rect 963 546 979 580
rect 1013 546 1029 580
rect 963 508 1029 546
rect 963 474 979 508
rect 1013 474 1029 508
rect 963 458 1029 474
rect 1063 580 1129 596
rect 1063 546 1079 580
rect 1113 546 1129 580
rect 1063 510 1129 546
rect 1063 476 1079 510
rect 1113 476 1129 510
rect 1063 440 1129 476
rect 1063 424 1079 440
rect 923 406 1079 424
rect 1113 406 1129 440
rect 889 390 1129 406
rect 361 380 377 390
rect 121 360 377 380
rect 21 294 87 310
rect 21 260 37 294
rect 71 260 87 294
rect 21 236 87 260
rect 121 236 187 360
rect 269 310 403 326
rect 269 276 285 310
rect 319 276 353 310
rect 387 276 403 310
rect 269 260 403 276
rect 505 320 743 356
rect 505 286 573 320
rect 607 286 641 320
rect 675 286 743 320
rect 505 270 743 286
rect 793 320 935 356
rect 793 286 809 320
rect 843 286 935 320
rect 793 270 935 286
rect 985 320 1127 356
rect 985 286 1033 320
rect 1067 286 1127 320
rect 985 270 1127 286
rect 313 236 359 260
rect 138 226 187 236
rect 36 168 52 202
rect 86 168 102 202
rect 36 120 102 168
rect 36 86 52 120
rect 86 86 102 120
rect 138 189 188 226
rect 172 155 188 189
rect 138 119 188 155
rect 224 210 258 226
rect 394 202 460 226
rect 258 189 460 202
rect 258 176 410 189
rect 224 168 410 176
rect 224 120 258 168
rect 394 155 410 168
rect 444 155 460 189
rect 36 85 102 86
rect 224 85 258 86
rect 36 51 258 85
rect 294 127 360 134
rect 294 93 310 127
rect 344 93 360 127
rect 394 119 460 155
rect 506 210 1120 236
rect 506 202 708 210
rect 506 189 572 202
rect 506 155 522 189
rect 556 155 572 189
rect 742 202 884 210
rect 506 119 572 155
rect 606 144 672 168
rect 294 85 360 93
rect 606 110 622 144
rect 656 110 672 144
rect 606 85 672 110
rect 294 51 672 85
rect 708 120 742 176
rect 918 202 1070 210
rect 918 176 934 202
rect 708 70 742 86
rect 778 136 844 168
rect 778 102 794 136
rect 828 102 844 136
rect 778 17 844 102
rect 884 120 934 176
rect 1104 176 1120 210
rect 918 86 934 120
rect 884 70 934 86
rect 968 136 1034 168
rect 968 102 984 136
rect 1018 102 1034 136
rect 968 17 1034 102
rect 1070 120 1120 176
rect 1104 86 1120 120
rect 1070 70 1120 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o2111ai_2
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 D1
port 5 nsew
flabel corelocali s 319 242 353 276 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 127 242 161 276 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 127 390 161 424 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 127 464 161 498 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 127 538 161 572 0 FreeSans 340 0 0 0 Y
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 1152 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1330000
string GDS_START 1319084
<< end >>
