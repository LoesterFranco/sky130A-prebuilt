magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 122 391 172 493
rect 508 391 558 425
rect 900 391 950 425
rect 122 357 950 391
rect 122 289 180 357
rect 17 215 87 255
rect 131 173 180 289
rect 224 289 712 323
rect 224 215 437 289
rect 471 215 602 255
rect 636 215 712 289
rect 746 289 1053 323
rect 746 215 822 289
rect 1019 255 1053 289
rect 856 215 975 255
rect 1019 215 1167 255
rect 104 129 180 173
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 28 291 78 527
rect 216 425 370 527
rect 414 459 652 493
rect 414 425 464 459
rect 602 425 652 459
rect 696 425 762 527
rect 806 459 1044 493
rect 806 425 856 459
rect 994 357 1044 459
rect 20 95 70 179
rect 1097 291 1138 527
rect 224 129 660 181
rect 704 147 1146 181
rect 224 95 274 129
rect 704 95 770 147
rect 882 145 1146 147
rect 20 51 274 95
rect 312 51 770 95
rect 814 17 848 111
rect 882 51 958 145
rect 1002 17 1036 111
rect 1070 51 1146 145
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
rlabel locali s 1019 255 1053 289 6 A1
port 1 nsew signal input
rlabel locali s 1019 215 1167 255 6 A1
port 1 nsew signal input
rlabel locali s 746 289 1053 323 6 A1
port 1 nsew signal input
rlabel locali s 746 215 822 289 6 A1
port 1 nsew signal input
rlabel locali s 856 215 975 255 6 A2
port 2 nsew signal input
rlabel locali s 636 215 712 289 6 B1
port 3 nsew signal input
rlabel locali s 224 289 712 323 6 B1
port 3 nsew signal input
rlabel locali s 224 215 437 289 6 B1
port 3 nsew signal input
rlabel locali s 471 215 602 255 6 B2
port 4 nsew signal input
rlabel locali s 17 215 87 255 6 C1
port 5 nsew signal input
rlabel locali s 900 391 950 425 6 Y
port 6 nsew signal output
rlabel locali s 508 391 558 425 6 Y
port 6 nsew signal output
rlabel locali s 131 173 180 289 6 Y
port 6 nsew signal output
rlabel locali s 122 391 172 493 6 Y
port 6 nsew signal output
rlabel locali s 122 357 950 391 6 Y
port 6 nsew signal output
rlabel locali s 122 289 180 357 6 Y
port 6 nsew signal output
rlabel locali s 104 129 180 173 6 Y
port 6 nsew signal output
rlabel metal1 s 0 -48 1196 48 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 496 1196 592 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 829230
string GDS_START 820084
<< end >>
