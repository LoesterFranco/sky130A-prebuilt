magic
tech sky130A
magscale 1 2
timestamp 1601050056
<< nwell >>
rect -38 332 1670 704
<< pwell >>
rect 0 0 1632 49
<< scpmos >>
rect 87 424 123 592
rect 197 424 233 592
rect 425 392 461 560
rect 558 392 594 592
rect 642 392 678 592
rect 756 508 792 592
rect 840 508 876 592
rect 1026 424 1062 592
rect 1127 424 1163 592
rect 1228 368 1264 592
rect 1333 368 1369 592
rect 1423 368 1459 592
rect 1513 368 1549 592
<< nmoslvt >>
rect 84 115 114 225
rect 202 114 232 262
rect 456 74 486 222
rect 628 79 658 207
rect 706 79 736 207
rect 865 123 895 207
rect 937 123 967 207
rect 1039 79 1069 207
rect 1125 79 1155 207
rect 1228 74 1258 222
rect 1332 74 1362 222
rect 1418 74 1448 222
rect 1513 74 1543 222
<< ndiff >>
rect 152 225 202 262
rect 27 185 84 225
rect 27 151 39 185
rect 73 151 84 185
rect 27 115 84 151
rect 114 115 202 225
rect 129 114 202 115
rect 232 250 289 262
rect 232 216 243 250
rect 277 216 289 250
rect 232 114 289 216
rect 399 189 456 222
rect 399 155 411 189
rect 445 155 456 189
rect 129 82 187 114
rect 129 48 141 82
rect 175 48 187 82
rect 399 74 456 155
rect 486 207 536 222
rect 1178 207 1228 222
rect 486 194 628 207
rect 486 160 579 194
rect 613 160 628 194
rect 486 125 628 160
rect 486 91 579 125
rect 613 91 628 125
rect 486 79 628 91
rect 658 79 706 207
rect 736 195 865 207
rect 736 161 747 195
rect 781 161 820 195
rect 854 161 865 195
rect 736 123 865 161
rect 895 123 937 207
rect 967 182 1039 207
rect 967 148 978 182
rect 1012 148 1039 182
rect 967 123 1039 148
rect 736 79 786 123
rect 486 74 536 79
rect 989 79 1039 123
rect 1069 195 1125 207
rect 1069 161 1080 195
rect 1114 161 1125 195
rect 1069 125 1125 161
rect 1069 91 1080 125
rect 1114 91 1125 125
rect 1069 79 1125 91
rect 1155 135 1228 207
rect 1155 101 1166 135
rect 1200 101 1228 135
rect 1155 79 1228 101
rect 1178 74 1228 79
rect 1258 210 1332 222
rect 1258 176 1271 210
rect 1305 176 1332 210
rect 1258 120 1332 176
rect 1258 86 1271 120
rect 1305 86 1332 120
rect 1258 74 1332 86
rect 1362 141 1418 222
rect 1362 107 1373 141
rect 1407 107 1418 141
rect 1362 74 1418 107
rect 1448 210 1513 222
rect 1448 176 1459 210
rect 1493 176 1513 210
rect 1448 120 1513 176
rect 1448 86 1459 120
rect 1493 86 1513 120
rect 1448 74 1513 86
rect 1543 141 1605 222
rect 1543 107 1559 141
rect 1593 107 1605 141
rect 1543 74 1605 107
rect 129 36 187 48
<< pdiff >>
rect 31 580 87 592
rect 31 546 43 580
rect 77 546 87 580
rect 31 470 87 546
rect 31 436 43 470
rect 77 436 87 470
rect 31 424 87 436
rect 123 580 197 592
rect 123 546 143 580
rect 177 546 197 580
rect 123 508 197 546
rect 123 474 143 508
rect 177 474 197 508
rect 123 424 197 474
rect 233 580 289 592
rect 233 546 243 580
rect 277 546 289 580
rect 476 580 558 592
rect 476 560 501 580
rect 233 470 289 546
rect 233 436 243 470
rect 277 436 289 470
rect 233 424 289 436
rect 369 441 425 560
rect 369 407 381 441
rect 415 407 425 441
rect 369 392 425 407
rect 461 546 501 560
rect 535 546 558 580
rect 461 392 558 546
rect 594 392 642 592
rect 678 531 756 592
rect 678 497 688 531
rect 722 508 756 531
rect 792 508 840 592
rect 876 568 1026 592
rect 876 534 887 568
rect 921 534 979 568
rect 1013 534 1026 568
rect 876 508 1026 534
rect 722 497 734 508
rect 678 462 734 497
rect 678 428 688 462
rect 722 428 734 462
rect 678 392 734 428
rect 976 424 1026 508
rect 1062 580 1127 592
rect 1062 546 1079 580
rect 1113 546 1127 580
rect 1062 470 1127 546
rect 1062 436 1079 470
rect 1113 436 1127 470
rect 1062 424 1127 436
rect 1163 580 1228 592
rect 1163 546 1179 580
rect 1213 546 1228 580
rect 1163 482 1228 546
rect 1163 448 1179 482
rect 1213 448 1228 482
rect 1163 424 1228 448
rect 1178 368 1228 424
rect 1264 580 1333 592
rect 1264 546 1279 580
rect 1313 546 1333 580
rect 1264 497 1333 546
rect 1264 463 1279 497
rect 1313 463 1333 497
rect 1264 414 1333 463
rect 1264 380 1279 414
rect 1313 380 1333 414
rect 1264 368 1333 380
rect 1369 580 1423 592
rect 1369 546 1379 580
rect 1413 546 1423 580
rect 1369 470 1423 546
rect 1369 436 1379 470
rect 1413 436 1423 470
rect 1369 368 1423 436
rect 1459 580 1513 592
rect 1459 546 1469 580
rect 1503 546 1513 580
rect 1459 497 1513 546
rect 1459 463 1469 497
rect 1503 463 1513 497
rect 1459 414 1513 463
rect 1459 380 1469 414
rect 1503 380 1513 414
rect 1459 368 1513 380
rect 1549 580 1605 592
rect 1549 546 1559 580
rect 1593 546 1605 580
rect 1549 498 1605 546
rect 1549 464 1559 498
rect 1593 464 1605 498
rect 1549 368 1605 464
<< ndiffc >>
rect 39 151 73 185
rect 243 216 277 250
rect 411 155 445 189
rect 141 48 175 82
rect 579 160 613 194
rect 579 91 613 125
rect 747 161 781 195
rect 820 161 854 195
rect 978 148 1012 182
rect 1080 161 1114 195
rect 1080 91 1114 125
rect 1166 101 1200 135
rect 1271 176 1305 210
rect 1271 86 1305 120
rect 1373 107 1407 141
rect 1459 176 1493 210
rect 1459 86 1493 120
rect 1559 107 1593 141
<< pdiffc >>
rect 43 546 77 580
rect 43 436 77 470
rect 143 546 177 580
rect 143 474 177 508
rect 243 546 277 580
rect 243 436 277 470
rect 381 407 415 441
rect 501 546 535 580
rect 688 497 722 531
rect 887 534 921 568
rect 979 534 1013 568
rect 688 428 722 462
rect 1079 546 1113 580
rect 1079 436 1113 470
rect 1179 546 1213 580
rect 1179 448 1213 482
rect 1279 546 1313 580
rect 1279 463 1313 497
rect 1279 380 1313 414
rect 1379 546 1413 580
rect 1379 436 1413 470
rect 1469 546 1503 580
rect 1469 463 1503 497
rect 1469 380 1503 414
rect 1559 546 1593 580
rect 1559 464 1593 498
<< poly >>
rect 87 592 123 618
rect 197 592 233 618
rect 558 592 594 618
rect 642 592 678 618
rect 756 592 792 618
rect 840 592 876 618
rect 1026 592 1062 618
rect 1127 592 1163 618
rect 1228 592 1264 618
rect 1333 592 1369 618
rect 1423 592 1459 618
rect 1513 592 1549 618
rect 425 560 461 586
rect 87 326 123 424
rect 25 310 123 326
rect 25 276 41 310
rect 75 276 123 310
rect 197 366 233 424
rect 197 350 263 366
rect 425 354 461 392
rect 197 316 213 350
rect 247 316 263 350
rect 197 300 263 316
rect 311 338 461 354
rect 311 304 327 338
rect 361 304 461 338
rect 558 310 594 392
rect 642 360 678 392
rect 642 344 708 360
rect 642 310 658 344
rect 692 310 708 344
rect 25 260 123 276
rect 202 262 232 300
rect 311 270 461 304
rect 84 225 114 260
rect 84 89 114 115
rect 311 236 327 270
rect 361 267 461 270
rect 534 294 600 310
rect 642 294 708 310
rect 756 347 792 508
rect 840 461 876 508
rect 840 445 954 461
rect 840 411 894 445
rect 928 411 954 445
rect 840 395 954 411
rect 924 382 954 395
rect 924 352 967 382
rect 756 331 876 347
rect 756 297 826 331
rect 860 297 876 331
rect 361 237 486 267
rect 534 260 550 294
rect 584 260 600 294
rect 534 252 600 260
rect 756 281 876 297
rect 756 252 786 281
rect 534 244 658 252
rect 361 236 377 237
rect 311 202 377 236
rect 456 222 486 237
rect 570 222 658 244
rect 311 168 327 202
rect 361 168 377 202
rect 311 152 377 168
rect 202 88 232 114
rect 628 207 658 222
rect 706 222 786 252
rect 706 207 736 222
rect 865 207 895 233
rect 937 207 967 352
rect 1026 330 1062 424
rect 1127 330 1163 424
rect 1228 330 1264 368
rect 1333 330 1369 368
rect 1423 330 1459 368
rect 1513 330 1549 368
rect 1032 314 1157 330
rect 1032 280 1048 314
rect 1082 280 1157 314
rect 1032 264 1157 280
rect 1228 314 1549 330
rect 1228 280 1244 314
rect 1278 280 1312 314
rect 1346 280 1380 314
rect 1414 280 1448 314
rect 1482 294 1549 314
rect 1482 280 1543 294
rect 1228 264 1543 280
rect 1039 207 1069 264
rect 1125 207 1155 264
rect 1228 222 1258 264
rect 1332 222 1362 264
rect 1418 222 1448 264
rect 1513 222 1543 264
rect 865 101 895 123
rect 823 85 895 101
rect 937 97 967 123
rect 456 48 486 74
rect 628 53 658 79
rect 706 53 736 79
rect 823 51 839 85
rect 873 51 895 85
rect 1039 53 1069 79
rect 1125 53 1155 79
rect 823 35 895 51
rect 1228 48 1258 74
rect 1332 48 1362 74
rect 1418 48 1448 74
rect 1513 48 1543 74
<< polycont >>
rect 41 276 75 310
rect 213 316 247 350
rect 327 304 361 338
rect 658 310 692 344
rect 327 236 361 270
rect 894 411 928 445
rect 826 297 860 331
rect 550 260 584 294
rect 327 168 361 202
rect 1048 280 1082 314
rect 1244 280 1278 314
rect 1312 280 1346 314
rect 1380 280 1414 314
rect 1448 280 1482 314
rect 839 51 873 85
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 27 580 93 596
rect 27 546 43 580
rect 77 546 93 580
rect 27 470 93 546
rect 27 436 43 470
rect 77 436 93 470
rect 127 580 193 649
rect 127 546 143 580
rect 177 546 193 580
rect 127 508 193 546
rect 127 474 143 508
rect 177 474 193 508
rect 127 458 193 474
rect 227 580 331 596
rect 227 546 243 580
rect 277 546 331 580
rect 472 580 564 649
rect 472 546 501 580
rect 535 546 564 580
rect 598 581 844 615
rect 227 512 331 546
rect 598 512 632 581
rect 227 478 632 512
rect 672 531 776 547
rect 672 497 688 531
rect 722 497 776 531
rect 227 470 331 478
rect 27 424 93 436
rect 227 436 243 470
rect 277 436 331 470
rect 672 462 776 497
rect 27 390 159 424
rect 227 420 331 436
rect 25 310 91 356
rect 25 276 41 310
rect 75 276 91 310
rect 25 260 91 276
rect 125 226 159 390
rect 197 350 263 366
rect 197 316 213 350
rect 247 316 263 350
rect 197 300 263 316
rect 297 354 331 420
rect 365 441 445 444
rect 365 407 381 441
rect 415 407 445 441
rect 672 428 688 462
rect 722 428 776 462
rect 672 412 776 428
rect 365 388 445 407
rect 411 378 445 388
rect 297 338 377 354
rect 297 304 327 338
rect 361 304 377 338
rect 297 270 377 304
rect 297 266 327 270
rect 23 185 159 226
rect 227 250 327 266
rect 227 216 243 250
rect 277 236 327 250
rect 361 236 377 270
rect 277 216 377 236
rect 227 202 377 216
rect 227 200 327 202
rect 23 151 39 185
rect 73 166 159 185
rect 297 168 327 200
rect 361 168 377 202
rect 73 151 263 166
rect 297 152 377 168
rect 411 344 708 378
rect 411 189 461 344
rect 642 310 658 344
rect 692 310 708 344
rect 445 155 461 189
rect 23 132 263 151
rect 23 111 89 132
rect 125 82 191 98
rect 125 48 141 82
rect 175 48 191 82
rect 229 85 263 132
rect 411 119 461 155
rect 495 294 600 310
rect 642 294 708 310
rect 495 260 550 294
rect 584 260 600 294
rect 495 244 600 260
rect 495 85 529 244
rect 229 51 529 85
rect 563 194 629 210
rect 563 160 579 194
rect 613 160 629 194
rect 563 125 629 160
rect 563 91 579 125
rect 613 91 629 125
rect 125 17 191 48
rect 563 17 629 91
rect 663 101 697 294
rect 742 211 776 412
rect 810 347 844 581
rect 878 568 1029 649
rect 878 534 887 568
rect 921 534 979 568
rect 1013 534 1029 568
rect 878 518 1029 534
rect 1063 580 1129 596
rect 1063 546 1079 580
rect 1113 546 1129 580
rect 1063 470 1129 546
rect 1063 461 1079 470
rect 878 445 1079 461
rect 878 411 894 445
rect 928 436 1079 445
rect 1113 436 1129 470
rect 928 411 1129 436
rect 1163 580 1229 649
rect 1163 546 1179 580
rect 1213 546 1229 580
rect 1163 482 1229 546
rect 1163 448 1179 482
rect 1213 448 1229 482
rect 1163 432 1229 448
rect 1263 580 1329 596
rect 1263 546 1279 580
rect 1313 546 1329 580
rect 1263 497 1329 546
rect 1263 463 1279 497
rect 1313 463 1329 497
rect 878 398 1129 411
rect 1263 414 1329 463
rect 1363 580 1429 649
rect 1363 546 1379 580
rect 1413 546 1429 580
rect 1363 470 1429 546
rect 1363 436 1379 470
rect 1413 436 1429 470
rect 1363 432 1429 436
rect 1463 580 1509 596
rect 1463 546 1469 580
rect 1503 546 1509 580
rect 1463 497 1509 546
rect 1463 463 1469 497
rect 1503 463 1509 497
rect 1543 580 1609 649
rect 1543 546 1559 580
rect 1593 546 1609 580
rect 1543 498 1609 546
rect 1543 464 1559 498
rect 1593 464 1609 498
rect 878 395 1166 398
rect 1063 364 1166 395
rect 1263 380 1279 414
rect 1313 398 1329 414
rect 1463 430 1509 463
rect 1463 414 1607 430
rect 1463 398 1469 414
rect 1313 380 1469 398
rect 1503 380 1607 414
rect 1263 364 1607 380
rect 810 331 876 347
rect 810 297 826 331
rect 860 297 876 331
rect 1132 330 1166 364
rect 810 281 876 297
rect 910 314 1098 330
rect 910 280 1048 314
rect 1082 280 1098 314
rect 910 264 1098 280
rect 1132 314 1498 330
rect 1132 280 1244 314
rect 1278 280 1312 314
rect 1346 280 1380 314
rect 1414 280 1448 314
rect 1482 280 1498 314
rect 1132 264 1498 280
rect 910 211 944 264
rect 1132 230 1166 264
rect 1561 230 1607 364
rect 731 195 944 211
rect 731 161 747 195
rect 781 161 820 195
rect 854 161 944 195
rect 731 145 944 161
rect 978 182 1028 211
rect 1012 148 1028 182
rect 663 85 889 101
rect 663 51 839 85
rect 873 51 889 85
rect 978 17 1028 148
rect 1064 196 1166 230
rect 1253 210 1607 230
rect 1064 195 1114 196
rect 1064 161 1080 195
rect 1253 176 1271 210
rect 1305 196 1459 210
rect 1305 176 1323 196
rect 1064 125 1114 161
rect 1064 91 1080 125
rect 1064 75 1114 91
rect 1150 135 1216 162
rect 1150 101 1166 135
rect 1200 101 1216 135
rect 1150 17 1216 101
rect 1253 120 1323 176
rect 1493 196 1607 210
rect 1493 176 1509 196
rect 1253 86 1271 120
rect 1305 86 1323 120
rect 1253 70 1323 86
rect 1357 141 1423 162
rect 1357 107 1373 141
rect 1407 107 1423 141
rect 1357 17 1423 107
rect 1459 120 1509 176
rect 1493 86 1509 120
rect 1459 70 1509 86
rect 1543 141 1609 162
rect 1543 107 1559 141
rect 1593 107 1609 141
rect 1543 17 1609 107
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
rlabel comment s 0 0 0 0 4 dlxtn_4
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 D
port 1 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew
flabel corelocali s 1567 242 1601 276 0 FreeSans 340 0 0 0 Q
port 7 nsew
flabel corelocali s 1567 316 1601 350 0 FreeSans 340 0 0 0 Q
port 7 nsew
flabel corelocali s 1567 390 1601 424 0 FreeSans 340 0 0 0 Q
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 1632 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 2199536
string GDS_START 2187576
<< end >>
