magic
tech sky130A
magscale 1 2
timestamp 1599588238
<< locali >>
rect 25 270 114 356
rect 167 270 263 356
rect 297 270 363 356
rect 503 364 559 596
rect 525 226 559 364
rect 486 70 559 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 23 424 89 572
rect 311 458 463 649
rect 23 390 452 424
rect 418 326 452 390
rect 418 260 491 326
rect 418 236 452 260
rect 23 202 452 236
rect 23 70 73 202
rect 109 17 175 162
rect 209 91 352 202
rect 386 17 452 162
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
rlabel locali s 297 270 363 356 6 A
port 1 nsew signal input
rlabel locali s 167 270 263 356 6 B
port 2 nsew signal input
rlabel locali s 25 270 114 356 6 C
port 3 nsew signal input
rlabel locali s 525 226 559 364 6 X
port 4 nsew signal output
rlabel locali s 503 364 559 596 6 X
port 4 nsew signal output
rlabel locali s 486 70 559 226 6 X
port 4 nsew signal output
rlabel metal1 s 0 -49 576 49 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 617 576 715 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 576 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 987414
string GDS_START 982148
<< end >>
