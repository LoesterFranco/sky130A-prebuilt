magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 287 3074 582
rect -38 261 1057 287
rect 1597 261 3074 287
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 89 47 119 131
rect 183 47 213 131
rect 383 47 413 131
rect 455 47 485 131
rect 661 47 691 131
rect 749 47 779 131
rect 871 47 901 131
rect 955 47 985 131
rect 1239 119 1269 203
rect 1343 119 1373 203
rect 1415 119 1445 203
rect 1600 47 1630 119
rect 1708 47 1738 119
rect 1814 47 1844 131
rect 1953 47 1983 175
rect 2151 47 2181 131
rect 2248 47 2278 119
rect 2361 47 2391 119
rect 2456 47 2486 131
rect 2568 47 2598 177
rect 2783 47 2813 131
rect 2900 47 2930 177
<< pmoshvt >>
rect 81 363 117 491
rect 175 363 211 491
rect 373 369 409 497
rect 455 369 491 497
rect 653 369 689 497
rect 751 369 787 497
rect 863 369 899 497
rect 965 369 1001 497
rect 1221 369 1257 497
rect 1340 369 1376 497
rect 1446 369 1482 497
rect 1575 413 1611 497
rect 1676 413 1712 497
rect 1789 413 1825 497
rect 1931 347 1967 497
rect 2129 413 2165 497
rect 2230 413 2266 497
rect 2324 413 2360 497
rect 2458 413 2494 497
rect 2565 297 2601 497
rect 2785 369 2821 497
rect 2892 297 2928 497
<< ndiff >>
rect 27 119 89 131
rect 27 85 35 119
rect 69 85 89 119
rect 27 47 89 85
rect 119 93 183 131
rect 119 59 129 93
rect 163 59 183 93
rect 119 47 183 59
rect 213 119 265 131
rect 213 85 223 119
rect 257 85 265 119
rect 213 47 265 85
rect 319 100 383 131
rect 319 66 327 100
rect 361 66 383 100
rect 319 47 383 66
rect 413 47 455 131
rect 485 93 545 131
rect 485 59 503 93
rect 537 59 545 93
rect 485 47 545 59
rect 599 119 661 131
rect 599 85 607 119
rect 641 85 661 119
rect 599 47 661 85
rect 691 106 749 131
rect 691 72 703 106
rect 737 72 749 106
rect 691 47 749 72
rect 779 47 871 131
rect 901 106 955 131
rect 901 72 911 106
rect 945 72 955 106
rect 901 47 955 72
rect 985 106 1047 131
rect 985 72 1005 106
rect 1039 72 1047 106
rect 985 47 1047 72
rect 1187 167 1239 203
rect 1187 133 1195 167
rect 1229 133 1239 167
rect 1187 119 1239 133
rect 1269 165 1343 203
rect 1269 131 1289 165
rect 1323 131 1343 165
rect 1269 119 1343 131
rect 1373 119 1415 203
rect 1445 180 1558 203
rect 1445 146 1467 180
rect 1501 146 1558 180
rect 1445 119 1558 146
rect 1893 131 1953 175
rect 1764 119 1814 131
rect 1470 99 1600 119
rect 1470 65 1534 99
rect 1568 65 1600 99
rect 1470 47 1600 65
rect 1630 99 1708 119
rect 1630 65 1650 99
rect 1684 65 1708 99
rect 1630 47 1708 65
rect 1738 47 1814 119
rect 1844 101 1953 131
rect 1844 67 1865 101
rect 1899 67 1953 101
rect 1844 47 1953 67
rect 1983 163 2035 175
rect 1983 129 1993 163
rect 2027 129 2035 163
rect 1983 95 2035 129
rect 1983 61 1993 95
rect 2027 61 2035 95
rect 1983 47 2035 61
rect 2089 107 2151 131
rect 2089 73 2097 107
rect 2131 73 2151 107
rect 2089 47 2151 73
rect 2181 119 2231 131
rect 2516 164 2568 177
rect 2516 131 2524 164
rect 2406 119 2456 131
rect 2181 47 2248 119
rect 2278 104 2361 119
rect 2278 70 2301 104
rect 2335 70 2361 104
rect 2278 47 2361 70
rect 2391 47 2456 119
rect 2486 130 2524 131
rect 2558 130 2568 164
rect 2486 96 2568 130
rect 2486 62 2524 96
rect 2558 62 2568 96
rect 2486 47 2568 62
rect 2598 164 2650 177
rect 2598 130 2608 164
rect 2642 130 2650 164
rect 2838 164 2900 177
rect 2838 131 2846 164
rect 2598 96 2650 130
rect 2598 62 2608 96
rect 2642 62 2650 96
rect 2598 47 2650 62
rect 2731 94 2783 131
rect 2731 60 2739 94
rect 2773 60 2783 94
rect 2731 47 2783 60
rect 2813 130 2846 131
rect 2880 130 2900 164
rect 2813 96 2900 130
rect 2813 62 2846 96
rect 2880 62 2900 96
rect 2813 47 2900 62
rect 2930 164 2991 177
rect 2930 130 2949 164
rect 2983 130 2991 164
rect 2930 96 2991 130
rect 2930 62 2949 96
rect 2983 62 2991 96
rect 2930 47 2991 62
<< pdiff >>
rect 27 477 81 491
rect 27 443 35 477
rect 69 443 81 477
rect 27 409 81 443
rect 27 375 35 409
rect 69 375 81 409
rect 27 363 81 375
rect 117 461 175 491
rect 117 427 129 461
rect 163 427 175 461
rect 117 363 175 427
rect 211 477 265 491
rect 211 443 223 477
rect 257 443 265 477
rect 211 409 265 443
rect 211 375 223 409
rect 257 375 265 409
rect 211 363 265 375
rect 319 485 373 497
rect 319 451 327 485
rect 361 451 373 485
rect 319 415 373 451
rect 319 381 327 415
rect 361 381 373 415
rect 319 369 373 381
rect 409 369 455 497
rect 491 485 545 497
rect 491 451 503 485
rect 537 451 545 485
rect 491 417 545 451
rect 491 383 503 417
rect 537 383 545 417
rect 491 369 545 383
rect 599 485 653 497
rect 599 451 607 485
rect 641 451 653 485
rect 599 415 653 451
rect 599 381 607 415
rect 641 381 653 415
rect 599 369 653 381
rect 689 485 751 497
rect 689 451 703 485
rect 737 451 751 485
rect 689 415 751 451
rect 689 381 703 415
rect 737 381 751 415
rect 689 369 751 381
rect 787 369 863 497
rect 899 485 965 497
rect 899 451 911 485
rect 945 451 965 485
rect 899 417 965 451
rect 899 383 911 417
rect 945 383 965 417
rect 899 369 965 383
rect 1001 485 1065 497
rect 1001 451 1023 485
rect 1057 451 1065 485
rect 1001 417 1065 451
rect 1001 383 1023 417
rect 1057 383 1065 417
rect 1001 369 1065 383
rect 1166 485 1221 497
rect 1166 451 1174 485
rect 1208 451 1221 485
rect 1166 417 1221 451
rect 1166 383 1174 417
rect 1208 383 1221 417
rect 1166 369 1221 383
rect 1257 485 1340 497
rect 1257 451 1281 485
rect 1315 451 1340 485
rect 1257 369 1340 451
rect 1376 369 1446 497
rect 1482 485 1575 497
rect 1482 451 1508 485
rect 1542 451 1575 485
rect 1482 417 1575 451
rect 1482 383 1508 417
rect 1542 413 1575 417
rect 1611 472 1676 497
rect 1611 438 1626 472
rect 1660 438 1676 472
rect 1611 413 1676 438
rect 1712 413 1789 497
rect 1825 485 1931 497
rect 1825 451 1879 485
rect 1913 451 1931 485
rect 1825 417 1931 451
rect 1825 413 1879 417
rect 1542 383 1558 413
rect 1482 369 1558 383
rect 1842 383 1879 413
rect 1913 383 1931 417
rect 1842 347 1931 383
rect 1967 485 2021 497
rect 1967 451 1979 485
rect 2013 451 2021 485
rect 1967 393 2021 451
rect 2075 472 2129 497
rect 2075 438 2083 472
rect 2117 438 2129 472
rect 2075 413 2129 438
rect 2165 413 2230 497
rect 2266 469 2324 497
rect 2266 435 2278 469
rect 2312 435 2324 469
rect 2266 413 2324 435
rect 2360 413 2458 497
rect 2494 485 2565 497
rect 2494 451 2519 485
rect 2553 451 2565 485
rect 2494 417 2565 451
rect 2494 413 2519 417
rect 1967 359 1979 393
rect 2013 359 2021 393
rect 1967 347 2021 359
rect 2511 383 2519 413
rect 2553 383 2565 417
rect 2511 349 2565 383
rect 2511 315 2519 349
rect 2553 315 2565 349
rect 2511 297 2565 315
rect 2601 479 2655 497
rect 2601 445 2613 479
rect 2647 445 2655 479
rect 2601 411 2655 445
rect 2601 377 2613 411
rect 2647 377 2655 411
rect 2601 343 2655 377
rect 2729 485 2785 497
rect 2729 451 2737 485
rect 2771 451 2785 485
rect 2729 415 2785 451
rect 2729 381 2737 415
rect 2771 381 2785 415
rect 2729 369 2785 381
rect 2821 479 2892 497
rect 2821 445 2846 479
rect 2880 445 2892 479
rect 2821 411 2892 445
rect 2821 377 2846 411
rect 2880 377 2892 411
rect 2821 369 2892 377
rect 2601 309 2613 343
rect 2647 309 2655 343
rect 2601 297 2655 309
rect 2838 343 2892 369
rect 2838 309 2846 343
rect 2880 309 2892 343
rect 2838 297 2892 309
rect 2928 479 2991 497
rect 2928 445 2949 479
rect 2983 445 2991 479
rect 2928 411 2991 445
rect 2928 377 2949 411
rect 2983 377 2991 411
rect 2928 343 2991 377
rect 2928 309 2949 343
rect 2983 309 2991 343
rect 2928 297 2991 309
<< ndiffc >>
rect 35 85 69 119
rect 129 59 163 93
rect 223 85 257 119
rect 327 66 361 100
rect 503 59 537 93
rect 607 85 641 119
rect 703 72 737 106
rect 911 72 945 106
rect 1005 72 1039 106
rect 1195 133 1229 167
rect 1289 131 1323 165
rect 1467 146 1501 180
rect 1534 65 1568 99
rect 1650 65 1684 99
rect 1865 67 1899 101
rect 1993 129 2027 163
rect 1993 61 2027 95
rect 2097 73 2131 107
rect 2301 70 2335 104
rect 2524 130 2558 164
rect 2524 62 2558 96
rect 2608 130 2642 164
rect 2608 62 2642 96
rect 2739 60 2773 94
rect 2846 130 2880 164
rect 2846 62 2880 96
rect 2949 130 2983 164
rect 2949 62 2983 96
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 129 427 163 461
rect 223 443 257 477
rect 223 375 257 409
rect 327 451 361 485
rect 327 381 361 415
rect 503 451 537 485
rect 503 383 537 417
rect 607 451 641 485
rect 607 381 641 415
rect 703 451 737 485
rect 703 381 737 415
rect 911 451 945 485
rect 911 383 945 417
rect 1023 451 1057 485
rect 1023 383 1057 417
rect 1174 451 1208 485
rect 1174 383 1208 417
rect 1281 451 1315 485
rect 1508 451 1542 485
rect 1508 383 1542 417
rect 1626 438 1660 472
rect 1879 451 1913 485
rect 1879 383 1913 417
rect 1979 451 2013 485
rect 2083 438 2117 472
rect 2278 435 2312 469
rect 2519 451 2553 485
rect 1979 359 2013 393
rect 2519 383 2553 417
rect 2519 315 2553 349
rect 2613 445 2647 479
rect 2613 377 2647 411
rect 2737 451 2771 485
rect 2737 381 2771 415
rect 2846 445 2880 479
rect 2846 377 2880 411
rect 2613 309 2647 343
rect 2846 309 2880 343
rect 2949 445 2983 479
rect 2949 377 2983 411
rect 2949 309 2983 343
<< poly >>
rect 81 491 117 517
rect 175 491 211 517
rect 373 497 409 523
rect 455 497 491 523
rect 653 497 689 523
rect 751 497 787 523
rect 863 497 899 523
rect 965 497 1001 523
rect 1221 497 1257 523
rect 1340 497 1376 523
rect 1446 497 1482 523
rect 1575 497 1611 523
rect 1676 497 1712 523
rect 1789 497 1825 523
rect 1931 497 1967 523
rect 2129 497 2165 523
rect 2230 497 2266 523
rect 2324 497 2360 523
rect 2458 497 2494 523
rect 2565 497 2601 523
rect 2785 497 2821 523
rect 2892 497 2928 523
rect 1575 398 1611 413
rect 1676 398 1712 413
rect 1789 398 1825 413
rect 81 348 117 363
rect 175 348 211 363
rect 373 354 409 369
rect 455 354 491 369
rect 653 354 689 369
rect 751 354 787 369
rect 863 354 899 369
rect 965 354 1001 369
rect 1221 354 1257 369
rect 1340 354 1376 369
rect 1446 354 1482 369
rect 47 318 119 348
rect 47 265 77 318
rect 173 274 213 348
rect 371 330 411 354
rect 23 249 77 265
rect 23 215 33 249
rect 67 215 77 249
rect 129 264 213 274
rect 129 230 145 264
rect 179 230 213 264
rect 129 220 213 230
rect 23 199 77 215
rect 47 176 77 199
rect 47 146 119 176
rect 89 131 119 146
rect 183 131 213 220
rect 343 314 413 330
rect 455 324 589 354
rect 343 280 359 314
rect 393 280 413 314
rect 343 246 413 280
rect 523 321 589 324
rect 523 287 539 321
rect 573 287 589 321
rect 523 277 589 287
rect 651 322 691 354
rect 749 322 789 354
rect 861 330 901 354
rect 651 292 789 322
rect 851 314 915 330
rect 343 212 359 246
rect 393 212 413 246
rect 343 196 413 212
rect 383 131 413 196
rect 455 219 531 235
rect 455 185 471 219
rect 505 200 531 219
rect 651 200 691 292
rect 851 280 861 314
rect 895 280 915 314
rect 963 315 1003 354
rect 1219 315 1259 354
rect 1338 337 1378 354
rect 1444 337 1484 354
rect 963 305 1259 315
rect 963 285 1134 305
rect 851 264 915 280
rect 1114 271 1134 285
rect 1168 271 1259 305
rect 1314 321 1378 337
rect 1314 287 1324 321
rect 1358 287 1378 321
rect 1314 271 1378 287
rect 1420 321 1484 337
rect 1420 287 1430 321
rect 1464 287 1484 321
rect 1573 297 1613 398
rect 1674 381 1714 398
rect 1674 365 1745 381
rect 1674 331 1691 365
rect 1725 331 1745 365
rect 1674 315 1745 331
rect 1420 271 1484 287
rect 1560 287 1636 297
rect 505 185 691 200
rect 455 170 691 185
rect 455 162 531 170
rect 455 131 485 162
rect 661 131 691 170
rect 733 219 797 235
rect 733 185 743 219
rect 777 185 797 219
rect 733 169 797 185
rect 749 131 779 169
rect 871 131 901 264
rect 1114 261 1259 271
rect 1219 247 1259 261
rect 1219 218 1269 247
rect 1239 203 1269 218
rect 1343 203 1373 271
rect 1560 253 1576 287
rect 1610 273 1636 287
rect 1610 253 1738 273
rect 1560 243 1738 253
rect 1415 203 1445 229
rect 955 153 1156 183
rect 955 131 985 153
rect 1126 101 1156 153
rect 1580 191 1656 201
rect 1580 157 1596 191
rect 1630 157 1656 191
rect 1580 147 1656 157
rect 1600 119 1630 147
rect 1708 119 1738 243
rect 1787 213 1827 398
rect 2129 398 2165 413
rect 2230 398 2266 413
rect 2324 398 2360 413
rect 2458 398 2494 413
rect 1931 332 1967 347
rect 1929 309 1969 332
rect 1869 299 1969 309
rect 1869 265 1885 299
rect 1919 265 1969 299
rect 2127 275 2167 398
rect 2228 315 2268 398
rect 2322 375 2362 398
rect 2321 365 2397 375
rect 2321 331 2337 365
rect 2371 331 2397 365
rect 2321 321 2397 331
rect 1869 255 1969 265
rect 1929 220 1969 255
rect 2102 259 2167 275
rect 2102 225 2112 259
rect 2146 225 2167 259
rect 2215 299 2279 315
rect 2215 265 2225 299
rect 2259 279 2279 299
rect 2259 265 2391 279
rect 2215 249 2391 265
rect 1787 203 1871 213
rect 1787 169 1811 203
rect 1845 169 1871 203
rect 1929 190 1983 220
rect 1953 175 1983 190
rect 2102 209 2167 225
rect 2102 179 2181 209
rect 1787 159 1871 169
rect 1814 131 1844 159
rect 1126 85 1180 101
rect 1126 51 1136 85
rect 1170 51 1180 85
rect 89 21 119 47
rect 183 21 213 47
rect 383 21 413 47
rect 455 21 485 47
rect 661 21 691 47
rect 749 21 779 47
rect 871 21 901 47
rect 955 21 985 47
rect 1126 35 1180 51
rect 1239 51 1269 119
rect 1343 93 1373 119
rect 1415 51 1445 119
rect 1239 21 1445 51
rect 2151 131 2181 179
rect 2248 191 2319 207
rect 2248 157 2275 191
rect 2309 157 2319 191
rect 2248 141 2319 157
rect 2248 119 2278 141
rect 2361 119 2391 249
rect 2456 244 2496 398
rect 2785 354 2821 369
rect 2565 282 2601 297
rect 2563 244 2603 282
rect 2783 265 2823 354
rect 2892 282 2928 297
rect 2890 265 2930 282
rect 2783 249 2930 265
rect 2456 228 2741 244
rect 2456 207 2697 228
rect 2456 131 2486 207
rect 2568 177 2598 207
rect 2687 194 2697 207
rect 2731 194 2741 228
rect 2687 178 2741 194
rect 2783 215 2839 249
rect 2873 215 2930 249
rect 2783 199 2930 215
rect 2783 131 2813 199
rect 2900 177 2930 199
rect 1600 21 1630 47
rect 1708 21 1738 47
rect 1814 21 1844 47
rect 1953 21 1983 47
rect 2151 21 2181 47
rect 2248 21 2278 47
rect 2361 21 2391 47
rect 2456 21 2486 47
rect 2568 21 2598 47
rect 2783 21 2813 47
rect 2900 21 2930 47
<< polycont >>
rect 33 215 67 249
rect 145 230 179 264
rect 359 280 393 314
rect 539 287 573 321
rect 359 212 393 246
rect 471 185 505 219
rect 861 280 895 314
rect 1134 271 1168 305
rect 1324 287 1358 321
rect 1430 287 1464 321
rect 1691 331 1725 365
rect 743 185 777 219
rect 1576 253 1610 287
rect 1596 157 1630 191
rect 1885 265 1919 299
rect 2337 331 2371 365
rect 2112 225 2146 259
rect 2225 265 2259 299
rect 1811 169 1845 203
rect 1136 51 1170 85
rect 2275 157 2309 191
rect 2697 194 2731 228
rect 2839 215 2873 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3036 561
rect 35 477 69 493
rect 35 409 69 443
rect 103 461 179 527
rect 103 427 129 461
rect 163 427 179 461
rect 223 477 257 493
rect 223 409 257 443
rect 69 391 179 393
rect 69 375 137 391
rect 35 359 137 375
rect 133 357 137 359
rect 171 357 179 391
rect 19 249 89 325
rect 19 215 33 249
rect 67 215 89 249
rect 19 195 89 215
rect 133 264 179 357
rect 133 230 145 264
rect 133 161 179 230
rect 35 127 179 161
rect 223 323 257 375
rect 35 119 69 127
rect 223 119 257 289
rect 35 69 69 85
rect 103 59 129 93
rect 163 59 179 93
rect 223 69 257 85
rect 291 485 377 493
rect 291 451 327 485
rect 361 451 377 485
rect 291 415 377 451
rect 291 381 327 415
rect 361 381 377 415
rect 291 378 377 381
rect 477 485 553 527
rect 703 485 742 527
rect 477 451 503 485
rect 537 451 553 485
rect 477 417 553 451
rect 477 383 503 417
rect 537 383 553 417
rect 477 378 553 383
rect 591 451 607 485
rect 641 451 657 485
rect 591 415 657 451
rect 591 381 607 415
rect 641 381 657 415
rect 291 119 325 378
rect 591 344 657 381
rect 737 451 742 485
rect 703 415 742 451
rect 737 381 742 415
rect 703 365 742 381
rect 885 485 961 493
rect 885 451 911 485
rect 945 451 961 485
rect 885 417 961 451
rect 1007 485 1073 493
rect 1007 451 1023 485
rect 1057 451 1073 485
rect 1007 442 1073 451
rect 885 383 911 417
rect 945 404 961 417
rect 1017 417 1073 442
rect 945 383 973 404
rect 885 364 973 383
rect 359 314 431 344
rect 393 280 431 314
rect 359 246 431 280
rect 539 321 657 344
rect 573 287 657 321
rect 393 212 431 246
rect 359 153 431 212
rect 465 237 505 274
rect 539 271 657 287
rect 465 219 553 237
rect 465 185 471 219
rect 505 185 553 219
rect 465 153 553 185
rect 596 235 657 271
rect 821 314 905 330
rect 821 280 861 314
rect 895 280 905 314
rect 821 264 905 280
rect 596 219 777 235
rect 596 185 743 219
rect 596 169 777 185
rect 821 187 855 264
rect 939 230 973 364
rect 596 119 641 169
rect 821 137 855 153
rect 889 196 973 230
rect 1017 383 1023 417
rect 1057 383 1073 417
rect 1017 357 1073 383
rect 1158 485 1226 493
rect 1158 451 1174 485
rect 1208 451 1226 485
rect 1158 417 1226 451
rect 1270 485 1339 527
rect 1270 451 1281 485
rect 1315 451 1339 485
rect 1270 435 1339 451
rect 1492 485 1558 493
rect 1492 451 1508 485
rect 1542 451 1558 485
rect 1872 485 1919 527
rect 1492 430 1558 451
rect 1600 472 1838 475
rect 1600 438 1626 472
rect 1660 438 1838 472
rect 1600 435 1838 438
rect 1158 383 1174 417
rect 1208 401 1226 417
rect 1508 417 1558 430
rect 1208 383 1474 401
rect 1158 367 1474 383
rect 325 100 377 103
rect 325 85 327 100
rect 103 17 179 59
rect 291 66 327 85
rect 361 66 377 100
rect 291 51 377 66
rect 477 93 553 103
rect 477 59 503 93
rect 537 59 553 93
rect 477 17 553 59
rect 596 85 607 119
rect 596 51 641 85
rect 677 106 753 122
rect 677 72 703 106
rect 737 72 753 106
rect 677 17 753 72
rect 889 119 953 196
rect 1017 165 1051 357
rect 1121 305 1177 323
rect 1121 271 1134 305
rect 1168 271 1177 305
rect 1121 221 1177 271
rect 1211 187 1245 367
rect 1289 321 1390 333
rect 1289 287 1324 321
rect 1358 287 1390 321
rect 1289 221 1390 287
rect 1424 321 1474 367
rect 1424 287 1430 321
rect 1464 287 1474 321
rect 1424 271 1474 287
rect 1542 383 1558 417
rect 1508 373 1558 383
rect 1657 391 1760 401
rect 1508 237 1542 373
rect 1657 357 1669 391
rect 1703 365 1760 391
rect 889 85 907 119
rect 941 106 953 119
rect 889 72 911 85
rect 945 72 953 106
rect 889 51 953 72
rect 999 129 1051 165
rect 1179 167 1245 187
rect 1179 133 1195 167
rect 1229 133 1245 167
rect 999 119 1039 129
rect 999 85 1003 119
rect 1037 106 1039 119
rect 1179 103 1245 133
rect 999 72 1005 85
rect 999 51 1039 72
rect 1073 85 1245 103
rect 1073 51 1136 85
rect 1170 51 1245 85
rect 1289 165 1339 181
rect 1323 131 1339 165
rect 1289 17 1339 131
rect 1460 180 1542 237
rect 1576 323 1623 344
rect 1576 289 1582 323
rect 1616 289 1623 323
rect 1576 287 1623 289
rect 1610 253 1623 287
rect 1576 225 1623 253
rect 1657 191 1691 357
rect 1725 331 1760 365
rect 1794 315 1838 435
rect 1872 451 1879 485
rect 1913 451 1919 485
rect 1872 417 1919 451
rect 1872 383 1879 417
rect 1913 383 1919 417
rect 1872 367 1919 383
rect 1953 485 2029 493
rect 1953 451 1979 485
rect 2013 451 2029 485
rect 1953 393 2029 451
rect 2071 472 2129 527
rect 2071 438 2083 472
rect 2117 438 2129 472
rect 2519 485 2553 527
rect 2071 421 2129 438
rect 2252 469 2475 471
rect 2252 435 2278 469
rect 2312 435 2475 469
rect 2252 433 2475 435
rect 1953 359 1979 393
rect 2013 359 2029 393
rect 1794 299 1919 315
rect 1794 297 1885 299
rect 1460 146 1467 180
rect 1501 146 1542 180
rect 1580 157 1596 191
rect 1630 157 1691 191
rect 1580 147 1691 157
rect 1739 265 1885 297
rect 1739 263 1919 265
rect 1460 119 1542 146
rect 1460 85 1463 119
rect 1497 113 1542 119
rect 1739 113 1773 263
rect 1885 249 1919 263
rect 1953 275 2029 359
rect 2225 391 2273 393
rect 2225 357 2232 391
rect 2266 357 2273 391
rect 2225 299 2273 357
rect 1953 259 2146 275
rect 1953 225 2112 259
rect 2259 265 2273 299
rect 2225 249 2273 265
rect 2307 365 2381 399
rect 2307 331 2337 365
rect 2371 331 2381 365
rect 2307 323 2381 331
rect 2307 289 2326 323
rect 2360 289 2381 323
rect 1811 213 1861 219
rect 1953 213 2146 225
rect 1811 209 2146 213
rect 1811 203 2044 209
rect 2307 207 2381 289
rect 1845 169 2044 203
rect 1811 163 2044 169
rect 1811 153 1993 163
rect 1497 99 1584 113
rect 1497 85 1534 99
rect 1460 65 1534 85
rect 1568 65 1584 99
rect 1460 51 1584 65
rect 1628 99 1773 113
rect 1953 129 1993 153
rect 2027 129 2044 163
rect 2275 191 2381 207
rect 2309 157 2381 191
rect 2275 141 2381 157
rect 2425 255 2475 433
rect 2519 417 2553 451
rect 2519 349 2553 383
rect 2519 299 2553 315
rect 2592 479 2663 493
rect 2592 445 2613 479
rect 2647 445 2663 479
rect 2592 411 2663 445
rect 2592 377 2613 411
rect 2647 377 2663 411
rect 2592 343 2663 377
rect 2592 309 2613 343
rect 2647 309 2663 343
rect 2425 221 2433 255
rect 2467 221 2475 255
rect 1628 65 1650 99
rect 1684 65 1773 99
rect 1628 51 1773 65
rect 1836 101 1915 112
rect 1836 67 1865 101
rect 1899 67 1915 101
rect 1836 17 1915 67
rect 1953 95 2044 129
rect 1953 61 1993 95
rect 2027 61 2044 95
rect 1953 51 2044 61
rect 2090 107 2145 123
rect 2425 107 2475 221
rect 2090 73 2097 107
rect 2131 73 2145 107
rect 2090 17 2145 73
rect 2282 104 2475 107
rect 2282 70 2301 104
rect 2335 70 2475 104
rect 2282 66 2475 70
rect 2509 164 2558 180
rect 2509 130 2524 164
rect 2509 96 2558 130
rect 2509 62 2524 96
rect 2509 17 2558 62
rect 2592 164 2663 309
rect 2721 485 2789 493
rect 2721 451 2737 485
rect 2771 451 2789 485
rect 2721 415 2789 451
rect 2721 381 2737 415
rect 2771 381 2789 415
rect 2721 244 2789 381
rect 2833 479 2880 527
rect 2833 445 2846 479
rect 2833 411 2880 445
rect 2833 377 2846 411
rect 2833 343 2880 377
rect 2833 309 2846 343
rect 2833 293 2880 309
rect 2931 479 3014 484
rect 2931 445 2949 479
rect 2983 445 3014 479
rect 2931 411 3014 445
rect 2931 377 2949 411
rect 2983 377 3014 411
rect 2931 343 3014 377
rect 2931 309 2949 343
rect 2983 309 3014 343
rect 2697 228 2789 244
rect 2731 194 2789 228
rect 2823 255 2889 259
rect 2823 215 2839 255
rect 2873 215 2889 255
rect 2823 214 2889 215
rect 2697 187 2789 194
rect 2697 178 2740 187
rect 2592 130 2608 164
rect 2642 130 2663 164
rect 2592 96 2663 130
rect 2592 62 2608 96
rect 2642 62 2663 96
rect 2592 51 2663 62
rect 2721 153 2740 178
rect 2774 153 2789 187
rect 2721 94 2789 153
rect 2721 60 2739 94
rect 2773 60 2789 94
rect 2721 51 2789 60
rect 2833 164 2880 180
rect 2833 130 2846 164
rect 2833 96 2880 130
rect 2833 62 2846 96
rect 2833 17 2880 62
rect 2931 164 3014 309
rect 2931 130 2949 164
rect 2983 130 3014 164
rect 2931 96 3014 130
rect 2931 62 2949 96
rect 2983 62 3014 96
rect 2931 51 3014 62
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3036 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 2881 527 2915 561
rect 2973 527 3007 561
rect 137 357 171 391
rect 223 289 257 323
rect 291 85 325 119
rect 821 153 855 187
rect 1669 365 1703 391
rect 1669 357 1691 365
rect 1691 357 1703 365
rect 907 106 941 119
rect 907 85 911 106
rect 911 85 941 106
rect 1003 106 1037 119
rect 1003 85 1005 106
rect 1005 85 1037 106
rect 1582 289 1616 323
rect 1463 85 1497 119
rect 2232 357 2266 391
rect 2326 289 2360 323
rect 2433 221 2467 255
rect 2839 249 2873 255
rect 2839 221 2873 249
rect 2740 153 2774 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
rect 2881 -17 2915 17
rect 2973 -17 3007 17
<< metal1 >>
rect 0 561 3036 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3036 561
rect 0 496 3036 527
rect 125 391 183 397
rect 125 357 137 391
rect 171 388 183 391
rect 1657 391 1725 397
rect 1657 388 1669 391
rect 171 360 1669 388
rect 171 357 183 360
rect 125 351 183 357
rect 1657 357 1669 360
rect 1703 388 1725 391
rect 2215 391 2283 397
rect 2215 388 2232 391
rect 1703 360 2232 388
rect 1703 357 1725 360
rect 1657 351 1725 357
rect 2215 357 2232 360
rect 2266 357 2283 391
rect 2215 351 2283 357
rect 201 323 269 329
rect 201 289 223 323
rect 257 320 269 323
rect 1565 323 1633 329
rect 1565 320 1582 323
rect 257 292 1582 320
rect 257 289 269 292
rect 201 283 269 289
rect 1565 289 1582 292
rect 1616 320 1633 323
rect 2309 323 2377 329
rect 2309 320 2326 323
rect 1616 292 2326 320
rect 1616 289 1633 292
rect 1565 283 1633 289
rect 2309 289 2326 292
rect 2360 289 2377 323
rect 2309 283 2377 289
rect 2421 255 2479 261
rect 2421 221 2433 255
rect 2467 252 2479 255
rect 2827 255 2885 261
rect 2827 252 2839 255
rect 2467 224 2839 252
rect 2467 221 2479 224
rect 2421 215 2479 221
rect 2827 221 2839 224
rect 2873 221 2885 255
rect 2827 215 2885 221
rect 809 187 867 193
rect 809 153 821 187
rect 855 184 867 187
rect 2728 187 2786 193
rect 2728 184 2740 187
rect 855 156 2740 184
rect 855 153 867 156
rect 809 147 867 153
rect 2728 153 2740 156
rect 2774 153 2786 187
rect 2728 147 2786 153
rect 279 119 337 125
rect 279 85 291 119
rect 325 116 337 119
rect 885 119 953 125
rect 885 116 907 119
rect 325 85 907 116
rect 941 85 953 119
rect 279 79 953 85
rect 981 119 1049 125
rect 981 85 1003 119
rect 1037 116 1049 119
rect 1441 119 1509 125
rect 1441 116 1463 119
rect 1037 85 1463 116
rect 1497 85 1509 119
rect 981 79 1509 85
rect 0 17 3036 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3036 17
rect 0 -48 3036 -17
<< labels >>
rlabel comment s 0 0 0 0 4 sedfxbp_1
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew
flabel corelocali s 1134 286 1168 320 0 FreeSans 400 0 0 0 SCE
port 5 nsew
flabel corelocali s 2961 221 2995 255 0 FreeSans 400 0 0 0 Q
port 10 nsew
flabel corelocali s 394 221 428 255 0 FreeSans 400 0 0 0 D
port 2 nsew
flabel corelocali s 503 190 503 190 0 FreeSans 400 0 0 0 DE
port 3 nsew
flabel corelocali s 1316 221 1350 255 0 FreeSans 400 0 0 0 SCD
port 4 nsew
flabel corelocali s 2603 221 2637 255 0 FreeSans 400 0 0 0 Q_N
port 11 nsew
flabel corelocali s 29 221 63 255 0 FreeSans 400 0 0 0 CLK
port 1 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel nbase s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel pwell s 296 0 296 0 0 FreeSans 400 0 0 0 VNB
port 7 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 3036 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 429640
string GDS_START 407262
<< end >>
