magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1932 561
rect 103 427 169 527
rect 291 427 357 527
rect 17 195 87 325
rect 686 451 762 527
rect 354 201 436 325
rect 866 451 932 527
rect 1184 451 1268 527
rect 103 17 169 93
rect 291 17 357 93
rect 722 147 804 213
rect 1402 389 1468 527
rect 722 17 804 105
rect 952 17 1016 109
rect 1332 201 1402 213
rect 1332 147 1468 201
rect 1338 17 1466 113
rect 1694 299 1728 527
rect 1762 323 1828 492
rect 1862 357 1915 527
rect 1762 299 1915 323
rect 1795 289 1915 299
rect 1804 179 1915 289
rect 1798 171 1915 179
rect 1795 165 1915 171
rect 1678 17 1744 165
rect 1778 153 1915 165
rect 1778 53 1827 153
rect 1861 17 1915 119
rect 0 -17 1932 17
<< obsli1 >>
rect 17 393 69 493
rect 203 409 247 493
rect 17 391 167 393
rect 17 359 121 391
rect 155 357 167 391
rect 121 161 167 357
rect 17 127 167 161
rect 201 187 247 409
rect 391 393 425 493
rect 472 450 638 484
rect 201 153 213 187
rect 17 69 69 127
rect 201 113 247 153
rect 286 359 425 393
rect 286 165 320 359
rect 470 357 489 391
rect 523 357 570 391
rect 470 315 570 357
rect 286 127 425 165
rect 470 141 514 315
rect 604 281 638 450
rect 798 417 832 475
rect 1022 433 1148 483
rect 1114 417 1148 433
rect 1308 417 1356 475
rect 672 367 942 417
rect 672 315 722 367
rect 824 281 874 313
rect 604 247 874 281
rect 604 239 688 247
rect 550 187 620 203
rect 550 153 581 187
rect 615 153 620 187
rect 550 129 620 153
rect 203 69 247 113
rect 391 61 425 127
rect 654 93 688 239
rect 908 213 942 367
rect 862 145 942 213
rect 976 391 1080 393
rect 976 357 1041 391
rect 1075 357 1080 391
rect 976 331 1080 357
rect 1114 383 1356 417
rect 976 179 1010 331
rect 1044 255 1080 295
rect 1044 221 1045 255
rect 1079 221 1080 255
rect 1114 281 1148 383
rect 1502 353 1536 475
rect 1594 383 1660 485
rect 1502 349 1576 353
rect 1182 315 1576 349
rect 1114 247 1498 281
rect 1044 213 1080 221
rect 1160 179 1230 203
rect 976 145 1230 179
rect 485 53 688 93
rect 862 59 912 145
rect 1264 95 1298 247
rect 1428 235 1498 247
rect 1538 136 1576 315
rect 1128 61 1298 95
rect 1506 70 1576 136
rect 1610 265 1660 383
rect 1610 199 1770 265
rect 1610 69 1644 199
<< obsli1c >>
rect 121 357 155 391
rect 213 153 247 187
rect 489 357 523 391
rect 581 153 615 187
rect 1041 357 1075 391
rect 1045 221 1079 255
<< metal1 >>
rect 0 496 1932 592
rect 753 184 811 193
rect 1397 184 1455 193
rect 753 156 1455 184
rect 753 147 811 156
rect 1397 147 1455 156
rect 0 -48 1932 48
<< obsm1 >>
rect 109 391 167 397
rect 109 357 121 391
rect 155 388 167 391
rect 477 391 535 397
rect 477 388 489 391
rect 155 360 489 388
rect 155 357 167 360
rect 109 351 167 357
rect 477 357 489 360
rect 523 388 535 391
rect 1029 391 1087 397
rect 1029 388 1041 391
rect 523 360 1041 388
rect 523 357 535 360
rect 477 351 535 357
rect 1029 357 1041 360
rect 1075 357 1087 391
rect 1029 351 1087 357
rect 1033 255 1091 261
rect 1033 252 1045 255
rect 584 224 1045 252
rect 584 193 627 224
rect 1033 221 1045 224
rect 1079 221 1091 255
rect 1033 215 1091 221
rect 201 187 259 193
rect 201 153 213 187
rect 247 184 259 187
rect 569 187 627 193
rect 569 184 581 187
rect 247 156 581 184
rect 247 153 259 156
rect 201 147 259 153
rect 569 153 581 156
rect 615 153 627 187
rect 569 147 627 153
<< labels >>
rlabel locali s 354 201 436 325 6 D
port 1 nsew signal input
rlabel locali s 1804 179 1915 289 6 Q
port 2 nsew signal output
rlabel locali s 1798 171 1915 179 6 Q
port 2 nsew signal output
rlabel locali s 1795 289 1915 299 6 Q
port 2 nsew signal output
rlabel locali s 1795 165 1915 171 6 Q
port 2 nsew signal output
rlabel locali s 1778 153 1915 165 6 Q
port 2 nsew signal output
rlabel locali s 1778 53 1827 153 6 Q
port 2 nsew signal output
rlabel locali s 1762 323 1828 492 6 Q
port 2 nsew signal output
rlabel locali s 1762 299 1915 323 6 Q
port 2 nsew signal output
rlabel locali s 722 147 804 213 6 SET_B
port 3 nsew signal input
rlabel locali s 1332 201 1402 213 6 SET_B
port 3 nsew signal input
rlabel locali s 1332 147 1468 201 6 SET_B
port 3 nsew signal input
rlabel metal1 s 1397 184 1455 193 6 SET_B
port 3 nsew signal input
rlabel metal1 s 1397 147 1455 156 6 SET_B
port 3 nsew signal input
rlabel metal1 s 753 184 811 193 6 SET_B
port 3 nsew signal input
rlabel metal1 s 753 156 1455 184 6 SET_B
port 3 nsew signal input
rlabel metal1 s 753 147 811 156 6 SET_B
port 3 nsew signal input
rlabel locali s 17 195 87 325 6 CLK
port 4 nsew clock input
rlabel locali s 1861 17 1915 119 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 1678 17 1744 165 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 1338 17 1466 113 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 952 17 1016 109 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 722 17 804 105 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 291 17 357 93 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 103 17 169 93 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 1932 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1932 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 1862 357 1915 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 1694 299 1728 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 1402 389 1468 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 1184 451 1268 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 866 451 932 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 686 451 762 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 291 427 357 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 103 427 169 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 1932 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 1932 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1932 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2476390
string GDS_START 2460278
<< end >>
