magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 5006 827
<< pwell >>
rect 29 1071 63 1105
rect 1225 1071 1259 1105
rect 3709 1071 3743 1105
rect 29 -17 63 17
rect 1225 -17 1259 17
rect 3709 -17 3743 17
<< scnmos >>
rect 114 957 144 1041
rect 198 957 228 1041
rect 457 918 487 1022
rect 541 918 571 1022
rect 625 918 655 1022
rect 709 918 739 1022
rect 897 911 927 1041
rect 981 911 1011 1041
rect 1085 911 1115 1041
rect 1169 911 1199 1041
rect 1285 911 1315 1041
rect 1369 911 1399 1041
rect 1473 911 1503 1041
rect 1557 911 1587 1041
rect 1745 918 1775 1022
rect 1829 918 1859 1022
rect 1913 918 1943 1022
rect 1997 918 2027 1022
rect 2256 957 2286 1041
rect 2340 957 2370 1041
rect 2598 957 2628 1041
rect 2682 957 2712 1041
rect 2941 918 2971 1022
rect 3025 918 3055 1022
rect 3109 918 3139 1022
rect 3193 918 3223 1022
rect 3381 911 3411 1041
rect 3465 911 3495 1041
rect 3569 911 3599 1041
rect 3653 911 3683 1041
rect 3769 911 3799 1041
rect 3853 911 3883 1041
rect 3957 911 3987 1041
rect 4041 911 4071 1041
rect 4229 918 4259 1022
rect 4313 918 4343 1022
rect 4397 918 4427 1022
rect 4481 918 4511 1022
rect 4740 957 4770 1041
rect 4824 957 4854 1041
rect 114 47 144 131
rect 198 47 228 131
rect 457 66 487 170
rect 541 66 571 170
rect 625 66 655 170
rect 709 66 739 170
rect 897 47 927 177
rect 981 47 1011 177
rect 1085 47 1115 177
rect 1169 47 1199 177
rect 1285 47 1315 177
rect 1369 47 1399 177
rect 1473 47 1503 177
rect 1557 47 1587 177
rect 1745 66 1775 170
rect 1829 66 1859 170
rect 1913 66 1943 170
rect 1997 66 2027 170
rect 2256 47 2286 131
rect 2340 47 2370 131
rect 2598 47 2628 131
rect 2682 47 2712 131
rect 2941 66 2971 170
rect 3025 66 3055 170
rect 3109 66 3139 170
rect 3193 66 3223 170
rect 3381 47 3411 177
rect 3465 47 3495 177
rect 3569 47 3599 177
rect 3653 47 3683 177
rect 3769 47 3799 177
rect 3853 47 3883 177
rect 3957 47 3987 177
rect 4041 47 4071 177
rect 4229 66 4259 170
rect 4313 66 4343 170
rect 4397 66 4427 170
rect 4481 66 4511 170
rect 4740 47 4770 131
rect 4824 47 4854 131
<< pmoshvt >>
rect 106 599 142 763
rect 200 599 236 763
rect 409 613 445 777
rect 503 613 539 777
rect 597 613 633 777
rect 691 613 727 777
rect 889 591 925 791
rect 983 591 1019 791
rect 1077 591 1113 791
rect 1171 591 1207 791
rect 1277 591 1313 791
rect 1371 591 1407 791
rect 1465 591 1501 791
rect 1559 591 1595 791
rect 1757 613 1793 777
rect 1851 613 1887 777
rect 1945 613 1981 777
rect 2039 613 2075 777
rect 2248 599 2284 763
rect 2342 599 2378 763
rect 2590 599 2626 763
rect 2684 599 2720 763
rect 2893 613 2929 777
rect 2987 613 3023 777
rect 3081 613 3117 777
rect 3175 613 3211 777
rect 3373 591 3409 791
rect 3467 591 3503 791
rect 3561 591 3597 791
rect 3655 591 3691 791
rect 3761 591 3797 791
rect 3855 591 3891 791
rect 3949 591 3985 791
rect 4043 591 4079 791
rect 4241 613 4277 777
rect 4335 613 4371 777
rect 4429 613 4465 777
rect 4523 613 4559 777
rect 4732 599 4768 763
rect 4826 599 4862 763
rect 106 325 142 489
rect 200 325 236 489
rect 409 311 445 475
rect 503 311 539 475
rect 597 311 633 475
rect 691 311 727 475
rect 889 297 925 497
rect 983 297 1019 497
rect 1077 297 1113 497
rect 1171 297 1207 497
rect 1277 297 1313 497
rect 1371 297 1407 497
rect 1465 297 1501 497
rect 1559 297 1595 497
rect 1757 311 1793 475
rect 1851 311 1887 475
rect 1945 311 1981 475
rect 2039 311 2075 475
rect 2248 325 2284 489
rect 2342 325 2378 489
rect 2590 325 2626 489
rect 2684 325 2720 489
rect 2893 311 2929 475
rect 2987 311 3023 475
rect 3081 311 3117 475
rect 3175 311 3211 475
rect 3373 297 3409 497
rect 3467 297 3503 497
rect 3561 297 3597 497
rect 3655 297 3691 497
rect 3761 297 3797 497
rect 3855 297 3891 497
rect 3949 297 3985 497
rect 4043 297 4079 497
rect 4241 311 4277 475
rect 4335 311 4371 475
rect 4429 311 4465 475
rect 4523 311 4559 475
rect 4732 325 4768 489
rect 4826 325 4862 489
<< ndiff >>
rect 62 1016 114 1041
rect 62 982 70 1016
rect 104 982 114 1016
rect 62 957 114 982
rect 144 1016 198 1041
rect 144 982 154 1016
rect 188 982 198 1016
rect 144 957 198 982
rect 228 1016 280 1041
rect 228 982 238 1016
rect 272 982 280 1016
rect 228 957 280 982
rect 845 1029 897 1041
rect 405 987 457 1022
rect 405 953 413 987
rect 447 953 457 987
rect 405 918 457 953
rect 487 969 541 1022
rect 487 935 497 969
rect 531 935 541 969
rect 487 918 541 935
rect 571 987 625 1022
rect 571 953 581 987
rect 615 953 625 987
rect 571 918 625 953
rect 655 969 709 1022
rect 655 935 665 969
rect 699 935 709 969
rect 655 918 709 935
rect 739 987 791 1022
rect 739 953 749 987
rect 783 953 791 987
rect 739 918 791 953
rect 845 995 853 1029
rect 887 995 897 1029
rect 845 911 897 995
rect 927 1029 981 1041
rect 927 995 937 1029
rect 971 995 981 1029
rect 927 961 981 995
rect 927 927 937 961
rect 971 927 981 961
rect 927 911 981 927
rect 1011 1029 1085 1041
rect 1011 995 1031 1029
rect 1065 995 1085 1029
rect 1011 911 1085 995
rect 1115 1029 1169 1041
rect 1115 995 1125 1029
rect 1159 995 1169 1029
rect 1115 961 1169 995
rect 1115 927 1125 961
rect 1159 927 1169 961
rect 1115 911 1169 927
rect 1199 1029 1285 1041
rect 1199 995 1225 1029
rect 1259 995 1285 1029
rect 1199 961 1285 995
rect 1199 927 1225 961
rect 1259 927 1285 961
rect 1199 911 1285 927
rect 1315 1029 1369 1041
rect 1315 995 1325 1029
rect 1359 995 1369 1029
rect 1315 961 1369 995
rect 1315 927 1325 961
rect 1359 927 1369 961
rect 1315 911 1369 927
rect 1399 1029 1473 1041
rect 1399 995 1419 1029
rect 1453 995 1473 1029
rect 1399 911 1473 995
rect 1503 1029 1557 1041
rect 1503 995 1513 1029
rect 1547 995 1557 1029
rect 1503 961 1557 995
rect 1503 927 1513 961
rect 1547 927 1557 961
rect 1503 911 1557 927
rect 1587 1029 1639 1041
rect 1587 995 1597 1029
rect 1631 995 1639 1029
rect 1587 911 1639 995
rect 1693 987 1745 1022
rect 1693 953 1701 987
rect 1735 953 1745 987
rect 1693 918 1745 953
rect 1775 969 1829 1022
rect 1775 935 1785 969
rect 1819 935 1829 969
rect 1775 918 1829 935
rect 1859 987 1913 1022
rect 1859 953 1869 987
rect 1903 953 1913 987
rect 1859 918 1913 953
rect 1943 969 1997 1022
rect 1943 935 1953 969
rect 1987 935 1997 969
rect 1943 918 1997 935
rect 2027 987 2079 1022
rect 2027 953 2037 987
rect 2071 953 2079 987
rect 2027 918 2079 953
rect 2204 1016 2256 1041
rect 2204 982 2212 1016
rect 2246 982 2256 1016
rect 2204 957 2256 982
rect 2286 1016 2340 1041
rect 2286 982 2296 1016
rect 2330 982 2340 1016
rect 2286 957 2340 982
rect 2370 1016 2422 1041
rect 2370 982 2380 1016
rect 2414 982 2422 1016
rect 2370 957 2422 982
rect 2546 1016 2598 1041
rect 2546 982 2554 1016
rect 2588 982 2598 1016
rect 2546 957 2598 982
rect 2628 1016 2682 1041
rect 2628 982 2638 1016
rect 2672 982 2682 1016
rect 2628 957 2682 982
rect 2712 1016 2764 1041
rect 2712 982 2722 1016
rect 2756 982 2764 1016
rect 2712 957 2764 982
rect 3329 1029 3381 1041
rect 2889 987 2941 1022
rect 2889 953 2897 987
rect 2931 953 2941 987
rect 2889 918 2941 953
rect 2971 969 3025 1022
rect 2971 935 2981 969
rect 3015 935 3025 969
rect 2971 918 3025 935
rect 3055 987 3109 1022
rect 3055 953 3065 987
rect 3099 953 3109 987
rect 3055 918 3109 953
rect 3139 969 3193 1022
rect 3139 935 3149 969
rect 3183 935 3193 969
rect 3139 918 3193 935
rect 3223 987 3275 1022
rect 3223 953 3233 987
rect 3267 953 3275 987
rect 3223 918 3275 953
rect 3329 995 3337 1029
rect 3371 995 3381 1029
rect 3329 911 3381 995
rect 3411 1029 3465 1041
rect 3411 995 3421 1029
rect 3455 995 3465 1029
rect 3411 961 3465 995
rect 3411 927 3421 961
rect 3455 927 3465 961
rect 3411 911 3465 927
rect 3495 1029 3569 1041
rect 3495 995 3515 1029
rect 3549 995 3569 1029
rect 3495 911 3569 995
rect 3599 1029 3653 1041
rect 3599 995 3609 1029
rect 3643 995 3653 1029
rect 3599 961 3653 995
rect 3599 927 3609 961
rect 3643 927 3653 961
rect 3599 911 3653 927
rect 3683 1029 3769 1041
rect 3683 995 3709 1029
rect 3743 995 3769 1029
rect 3683 961 3769 995
rect 3683 927 3709 961
rect 3743 927 3769 961
rect 3683 911 3769 927
rect 3799 1029 3853 1041
rect 3799 995 3809 1029
rect 3843 995 3853 1029
rect 3799 961 3853 995
rect 3799 927 3809 961
rect 3843 927 3853 961
rect 3799 911 3853 927
rect 3883 1029 3957 1041
rect 3883 995 3903 1029
rect 3937 995 3957 1029
rect 3883 911 3957 995
rect 3987 1029 4041 1041
rect 3987 995 3997 1029
rect 4031 995 4041 1029
rect 3987 961 4041 995
rect 3987 927 3997 961
rect 4031 927 4041 961
rect 3987 911 4041 927
rect 4071 1029 4123 1041
rect 4071 995 4081 1029
rect 4115 995 4123 1029
rect 4071 911 4123 995
rect 4177 987 4229 1022
rect 4177 953 4185 987
rect 4219 953 4229 987
rect 4177 918 4229 953
rect 4259 969 4313 1022
rect 4259 935 4269 969
rect 4303 935 4313 969
rect 4259 918 4313 935
rect 4343 987 4397 1022
rect 4343 953 4353 987
rect 4387 953 4397 987
rect 4343 918 4397 953
rect 4427 969 4481 1022
rect 4427 935 4437 969
rect 4471 935 4481 969
rect 4427 918 4481 935
rect 4511 987 4563 1022
rect 4511 953 4521 987
rect 4555 953 4563 987
rect 4511 918 4563 953
rect 4688 1016 4740 1041
rect 4688 982 4696 1016
rect 4730 982 4740 1016
rect 4688 957 4740 982
rect 4770 1016 4824 1041
rect 4770 982 4780 1016
rect 4814 982 4824 1016
rect 4770 957 4824 982
rect 4854 1016 4906 1041
rect 4854 982 4864 1016
rect 4898 982 4906 1016
rect 4854 957 4906 982
rect 62 106 114 131
rect 62 72 70 106
rect 104 72 114 106
rect 62 47 114 72
rect 144 106 198 131
rect 144 72 154 106
rect 188 72 198 106
rect 144 47 198 72
rect 228 106 280 131
rect 228 72 238 106
rect 272 72 280 106
rect 228 47 280 72
rect 405 135 457 170
rect 405 101 413 135
rect 447 101 457 135
rect 405 66 457 101
rect 487 153 541 170
rect 487 119 497 153
rect 531 119 541 153
rect 487 66 541 119
rect 571 135 625 170
rect 571 101 581 135
rect 615 101 625 135
rect 571 66 625 101
rect 655 153 709 170
rect 655 119 665 153
rect 699 119 709 153
rect 655 66 709 119
rect 739 135 791 170
rect 739 101 749 135
rect 783 101 791 135
rect 739 66 791 101
rect 845 93 897 177
rect 845 59 853 93
rect 887 59 897 93
rect 845 47 897 59
rect 927 161 981 177
rect 927 127 937 161
rect 971 127 981 161
rect 927 93 981 127
rect 927 59 937 93
rect 971 59 981 93
rect 927 47 981 59
rect 1011 93 1085 177
rect 1011 59 1031 93
rect 1065 59 1085 93
rect 1011 47 1085 59
rect 1115 161 1169 177
rect 1115 127 1125 161
rect 1159 127 1169 161
rect 1115 93 1169 127
rect 1115 59 1125 93
rect 1159 59 1169 93
rect 1115 47 1169 59
rect 1199 161 1285 177
rect 1199 127 1225 161
rect 1259 127 1285 161
rect 1199 93 1285 127
rect 1199 59 1225 93
rect 1259 59 1285 93
rect 1199 47 1285 59
rect 1315 161 1369 177
rect 1315 127 1325 161
rect 1359 127 1369 161
rect 1315 93 1369 127
rect 1315 59 1325 93
rect 1359 59 1369 93
rect 1315 47 1369 59
rect 1399 93 1473 177
rect 1399 59 1419 93
rect 1453 59 1473 93
rect 1399 47 1473 59
rect 1503 161 1557 177
rect 1503 127 1513 161
rect 1547 127 1557 161
rect 1503 93 1557 127
rect 1503 59 1513 93
rect 1547 59 1557 93
rect 1503 47 1557 59
rect 1587 93 1639 177
rect 1587 59 1597 93
rect 1631 59 1639 93
rect 1693 135 1745 170
rect 1693 101 1701 135
rect 1735 101 1745 135
rect 1693 66 1745 101
rect 1775 153 1829 170
rect 1775 119 1785 153
rect 1819 119 1829 153
rect 1775 66 1829 119
rect 1859 135 1913 170
rect 1859 101 1869 135
rect 1903 101 1913 135
rect 1859 66 1913 101
rect 1943 153 1997 170
rect 1943 119 1953 153
rect 1987 119 1997 153
rect 1943 66 1997 119
rect 2027 135 2079 170
rect 2027 101 2037 135
rect 2071 101 2079 135
rect 2027 66 2079 101
rect 1587 47 1639 59
rect 2204 106 2256 131
rect 2204 72 2212 106
rect 2246 72 2256 106
rect 2204 47 2256 72
rect 2286 106 2340 131
rect 2286 72 2296 106
rect 2330 72 2340 106
rect 2286 47 2340 72
rect 2370 106 2422 131
rect 2370 72 2380 106
rect 2414 72 2422 106
rect 2370 47 2422 72
rect 2546 106 2598 131
rect 2546 72 2554 106
rect 2588 72 2598 106
rect 2546 47 2598 72
rect 2628 106 2682 131
rect 2628 72 2638 106
rect 2672 72 2682 106
rect 2628 47 2682 72
rect 2712 106 2764 131
rect 2712 72 2722 106
rect 2756 72 2764 106
rect 2712 47 2764 72
rect 2889 135 2941 170
rect 2889 101 2897 135
rect 2931 101 2941 135
rect 2889 66 2941 101
rect 2971 153 3025 170
rect 2971 119 2981 153
rect 3015 119 3025 153
rect 2971 66 3025 119
rect 3055 135 3109 170
rect 3055 101 3065 135
rect 3099 101 3109 135
rect 3055 66 3109 101
rect 3139 153 3193 170
rect 3139 119 3149 153
rect 3183 119 3193 153
rect 3139 66 3193 119
rect 3223 135 3275 170
rect 3223 101 3233 135
rect 3267 101 3275 135
rect 3223 66 3275 101
rect 3329 93 3381 177
rect 3329 59 3337 93
rect 3371 59 3381 93
rect 3329 47 3381 59
rect 3411 161 3465 177
rect 3411 127 3421 161
rect 3455 127 3465 161
rect 3411 93 3465 127
rect 3411 59 3421 93
rect 3455 59 3465 93
rect 3411 47 3465 59
rect 3495 93 3569 177
rect 3495 59 3515 93
rect 3549 59 3569 93
rect 3495 47 3569 59
rect 3599 161 3653 177
rect 3599 127 3609 161
rect 3643 127 3653 161
rect 3599 93 3653 127
rect 3599 59 3609 93
rect 3643 59 3653 93
rect 3599 47 3653 59
rect 3683 161 3769 177
rect 3683 127 3709 161
rect 3743 127 3769 161
rect 3683 93 3769 127
rect 3683 59 3709 93
rect 3743 59 3769 93
rect 3683 47 3769 59
rect 3799 161 3853 177
rect 3799 127 3809 161
rect 3843 127 3853 161
rect 3799 93 3853 127
rect 3799 59 3809 93
rect 3843 59 3853 93
rect 3799 47 3853 59
rect 3883 93 3957 177
rect 3883 59 3903 93
rect 3937 59 3957 93
rect 3883 47 3957 59
rect 3987 161 4041 177
rect 3987 127 3997 161
rect 4031 127 4041 161
rect 3987 93 4041 127
rect 3987 59 3997 93
rect 4031 59 4041 93
rect 3987 47 4041 59
rect 4071 93 4123 177
rect 4071 59 4081 93
rect 4115 59 4123 93
rect 4177 135 4229 170
rect 4177 101 4185 135
rect 4219 101 4229 135
rect 4177 66 4229 101
rect 4259 153 4313 170
rect 4259 119 4269 153
rect 4303 119 4313 153
rect 4259 66 4313 119
rect 4343 135 4397 170
rect 4343 101 4353 135
rect 4387 101 4397 135
rect 4343 66 4397 101
rect 4427 153 4481 170
rect 4427 119 4437 153
rect 4471 119 4481 153
rect 4427 66 4481 119
rect 4511 135 4563 170
rect 4511 101 4521 135
rect 4555 101 4563 135
rect 4511 66 4563 101
rect 4071 47 4123 59
rect 4688 106 4740 131
rect 4688 72 4696 106
rect 4730 72 4740 106
rect 4688 47 4740 72
rect 4770 106 4824 131
rect 4770 72 4780 106
rect 4814 72 4824 106
rect 4770 47 4824 72
rect 4854 106 4906 131
rect 4854 72 4864 106
rect 4898 72 4906 106
rect 4854 47 4906 72
<< pdiff >>
rect 52 751 106 763
rect 52 717 60 751
rect 94 717 106 751
rect 52 645 106 717
rect 52 611 60 645
rect 94 611 106 645
rect 52 599 106 611
rect 142 751 200 763
rect 142 717 154 751
rect 188 717 200 751
rect 142 645 200 717
rect 142 611 154 645
rect 188 611 200 645
rect 142 599 200 611
rect 236 751 290 763
rect 236 717 248 751
rect 282 717 290 751
rect 236 645 290 717
rect 236 611 248 645
rect 282 611 290 645
rect 355 759 409 777
rect 355 725 363 759
rect 397 725 409 759
rect 355 659 409 725
rect 355 625 363 659
rect 397 625 409 659
rect 355 613 409 625
rect 445 765 503 777
rect 445 731 457 765
rect 491 731 503 765
rect 445 659 503 731
rect 445 625 457 659
rect 491 625 503 659
rect 445 613 503 625
rect 539 765 597 777
rect 539 731 551 765
rect 585 731 597 765
rect 539 659 597 731
rect 539 625 551 659
rect 585 625 597 659
rect 539 613 597 625
rect 633 765 691 777
rect 633 731 645 765
rect 679 731 691 765
rect 633 659 691 731
rect 633 625 645 659
rect 679 625 691 659
rect 633 613 691 625
rect 727 765 781 777
rect 727 731 739 765
rect 773 731 781 765
rect 727 659 781 731
rect 727 625 739 659
rect 773 625 781 659
rect 727 613 781 625
rect 835 705 889 791
rect 835 671 843 705
rect 877 671 889 705
rect 835 637 889 671
rect 236 599 290 611
rect 835 603 843 637
rect 877 603 889 637
rect 835 591 889 603
rect 925 773 983 791
rect 925 739 937 773
rect 971 739 983 773
rect 925 705 983 739
rect 925 671 937 705
rect 971 671 983 705
rect 925 637 983 671
rect 925 603 937 637
rect 971 603 983 637
rect 925 591 983 603
rect 1019 705 1077 791
rect 1019 671 1031 705
rect 1065 671 1077 705
rect 1019 637 1077 671
rect 1019 603 1031 637
rect 1065 603 1077 637
rect 1019 591 1077 603
rect 1113 773 1171 791
rect 1113 739 1125 773
rect 1159 739 1171 773
rect 1113 705 1171 739
rect 1113 671 1125 705
rect 1159 671 1171 705
rect 1113 637 1171 671
rect 1113 603 1125 637
rect 1159 603 1171 637
rect 1113 591 1171 603
rect 1207 773 1277 791
rect 1207 739 1225 773
rect 1259 739 1277 773
rect 1207 705 1277 739
rect 1207 671 1225 705
rect 1259 671 1277 705
rect 1207 637 1277 671
rect 1207 603 1225 637
rect 1259 603 1277 637
rect 1207 591 1277 603
rect 1313 773 1371 791
rect 1313 739 1325 773
rect 1359 739 1371 773
rect 1313 705 1371 739
rect 1313 671 1325 705
rect 1359 671 1371 705
rect 1313 637 1371 671
rect 1313 603 1325 637
rect 1359 603 1371 637
rect 1313 591 1371 603
rect 1407 705 1465 791
rect 1407 671 1419 705
rect 1453 671 1465 705
rect 1407 637 1465 671
rect 1407 603 1419 637
rect 1453 603 1465 637
rect 1407 591 1465 603
rect 1501 773 1559 791
rect 1501 739 1513 773
rect 1547 739 1559 773
rect 1501 705 1559 739
rect 1501 671 1513 705
rect 1547 671 1559 705
rect 1501 637 1559 671
rect 1501 603 1513 637
rect 1547 603 1559 637
rect 1501 591 1559 603
rect 1595 705 1649 791
rect 1595 671 1607 705
rect 1641 671 1649 705
rect 1595 637 1649 671
rect 1595 603 1607 637
rect 1641 603 1649 637
rect 1703 765 1757 777
rect 1703 731 1711 765
rect 1745 731 1757 765
rect 1703 659 1757 731
rect 1703 625 1711 659
rect 1745 625 1757 659
rect 1703 613 1757 625
rect 1793 765 1851 777
rect 1793 731 1805 765
rect 1839 731 1851 765
rect 1793 659 1851 731
rect 1793 625 1805 659
rect 1839 625 1851 659
rect 1793 613 1851 625
rect 1887 765 1945 777
rect 1887 731 1899 765
rect 1933 731 1945 765
rect 1887 659 1945 731
rect 1887 625 1899 659
rect 1933 625 1945 659
rect 1887 613 1945 625
rect 1981 765 2039 777
rect 1981 731 1993 765
rect 2027 731 2039 765
rect 1981 659 2039 731
rect 1981 625 1993 659
rect 2027 625 2039 659
rect 1981 613 2039 625
rect 2075 759 2129 777
rect 2075 725 2087 759
rect 2121 725 2129 759
rect 2075 659 2129 725
rect 2075 625 2087 659
rect 2121 625 2129 659
rect 2075 613 2129 625
rect 2194 751 2248 763
rect 2194 717 2202 751
rect 2236 717 2248 751
rect 2194 645 2248 717
rect 1595 591 1649 603
rect 2194 611 2202 645
rect 2236 611 2248 645
rect 2194 599 2248 611
rect 2284 751 2342 763
rect 2284 717 2296 751
rect 2330 717 2342 751
rect 2284 645 2342 717
rect 2284 611 2296 645
rect 2330 611 2342 645
rect 2284 599 2342 611
rect 2378 751 2432 763
rect 2378 717 2390 751
rect 2424 717 2432 751
rect 2378 645 2432 717
rect 2378 611 2390 645
rect 2424 611 2432 645
rect 2378 599 2432 611
rect 2536 751 2590 763
rect 2536 717 2544 751
rect 2578 717 2590 751
rect 2536 645 2590 717
rect 2536 611 2544 645
rect 2578 611 2590 645
rect 2536 599 2590 611
rect 2626 751 2684 763
rect 2626 717 2638 751
rect 2672 717 2684 751
rect 2626 645 2684 717
rect 2626 611 2638 645
rect 2672 611 2684 645
rect 2626 599 2684 611
rect 2720 751 2774 763
rect 2720 717 2732 751
rect 2766 717 2774 751
rect 2720 645 2774 717
rect 2720 611 2732 645
rect 2766 611 2774 645
rect 2839 759 2893 777
rect 2839 725 2847 759
rect 2881 725 2893 759
rect 2839 659 2893 725
rect 2839 625 2847 659
rect 2881 625 2893 659
rect 2839 613 2893 625
rect 2929 765 2987 777
rect 2929 731 2941 765
rect 2975 731 2987 765
rect 2929 659 2987 731
rect 2929 625 2941 659
rect 2975 625 2987 659
rect 2929 613 2987 625
rect 3023 765 3081 777
rect 3023 731 3035 765
rect 3069 731 3081 765
rect 3023 659 3081 731
rect 3023 625 3035 659
rect 3069 625 3081 659
rect 3023 613 3081 625
rect 3117 765 3175 777
rect 3117 731 3129 765
rect 3163 731 3175 765
rect 3117 659 3175 731
rect 3117 625 3129 659
rect 3163 625 3175 659
rect 3117 613 3175 625
rect 3211 765 3265 777
rect 3211 731 3223 765
rect 3257 731 3265 765
rect 3211 659 3265 731
rect 3211 625 3223 659
rect 3257 625 3265 659
rect 3211 613 3265 625
rect 3319 705 3373 791
rect 3319 671 3327 705
rect 3361 671 3373 705
rect 3319 637 3373 671
rect 2720 599 2774 611
rect 3319 603 3327 637
rect 3361 603 3373 637
rect 3319 591 3373 603
rect 3409 773 3467 791
rect 3409 739 3421 773
rect 3455 739 3467 773
rect 3409 705 3467 739
rect 3409 671 3421 705
rect 3455 671 3467 705
rect 3409 637 3467 671
rect 3409 603 3421 637
rect 3455 603 3467 637
rect 3409 591 3467 603
rect 3503 705 3561 791
rect 3503 671 3515 705
rect 3549 671 3561 705
rect 3503 637 3561 671
rect 3503 603 3515 637
rect 3549 603 3561 637
rect 3503 591 3561 603
rect 3597 773 3655 791
rect 3597 739 3609 773
rect 3643 739 3655 773
rect 3597 705 3655 739
rect 3597 671 3609 705
rect 3643 671 3655 705
rect 3597 637 3655 671
rect 3597 603 3609 637
rect 3643 603 3655 637
rect 3597 591 3655 603
rect 3691 773 3761 791
rect 3691 739 3709 773
rect 3743 739 3761 773
rect 3691 705 3761 739
rect 3691 671 3709 705
rect 3743 671 3761 705
rect 3691 637 3761 671
rect 3691 603 3709 637
rect 3743 603 3761 637
rect 3691 591 3761 603
rect 3797 773 3855 791
rect 3797 739 3809 773
rect 3843 739 3855 773
rect 3797 705 3855 739
rect 3797 671 3809 705
rect 3843 671 3855 705
rect 3797 637 3855 671
rect 3797 603 3809 637
rect 3843 603 3855 637
rect 3797 591 3855 603
rect 3891 705 3949 791
rect 3891 671 3903 705
rect 3937 671 3949 705
rect 3891 637 3949 671
rect 3891 603 3903 637
rect 3937 603 3949 637
rect 3891 591 3949 603
rect 3985 773 4043 791
rect 3985 739 3997 773
rect 4031 739 4043 773
rect 3985 705 4043 739
rect 3985 671 3997 705
rect 4031 671 4043 705
rect 3985 637 4043 671
rect 3985 603 3997 637
rect 4031 603 4043 637
rect 3985 591 4043 603
rect 4079 705 4133 791
rect 4079 671 4091 705
rect 4125 671 4133 705
rect 4079 637 4133 671
rect 4079 603 4091 637
rect 4125 603 4133 637
rect 4187 765 4241 777
rect 4187 731 4195 765
rect 4229 731 4241 765
rect 4187 659 4241 731
rect 4187 625 4195 659
rect 4229 625 4241 659
rect 4187 613 4241 625
rect 4277 765 4335 777
rect 4277 731 4289 765
rect 4323 731 4335 765
rect 4277 659 4335 731
rect 4277 625 4289 659
rect 4323 625 4335 659
rect 4277 613 4335 625
rect 4371 765 4429 777
rect 4371 731 4383 765
rect 4417 731 4429 765
rect 4371 659 4429 731
rect 4371 625 4383 659
rect 4417 625 4429 659
rect 4371 613 4429 625
rect 4465 765 4523 777
rect 4465 731 4477 765
rect 4511 731 4523 765
rect 4465 659 4523 731
rect 4465 625 4477 659
rect 4511 625 4523 659
rect 4465 613 4523 625
rect 4559 759 4613 777
rect 4559 725 4571 759
rect 4605 725 4613 759
rect 4559 659 4613 725
rect 4559 625 4571 659
rect 4605 625 4613 659
rect 4559 613 4613 625
rect 4678 751 4732 763
rect 4678 717 4686 751
rect 4720 717 4732 751
rect 4678 645 4732 717
rect 4079 591 4133 603
rect 4678 611 4686 645
rect 4720 611 4732 645
rect 4678 599 4732 611
rect 4768 751 4826 763
rect 4768 717 4780 751
rect 4814 717 4826 751
rect 4768 645 4826 717
rect 4768 611 4780 645
rect 4814 611 4826 645
rect 4768 599 4826 611
rect 4862 751 4916 763
rect 4862 717 4874 751
rect 4908 717 4916 751
rect 4862 645 4916 717
rect 4862 611 4874 645
rect 4908 611 4916 645
rect 4862 599 4916 611
rect 52 477 106 489
rect 52 443 60 477
rect 94 443 106 477
rect 52 371 106 443
rect 52 337 60 371
rect 94 337 106 371
rect 52 325 106 337
rect 142 477 200 489
rect 142 443 154 477
rect 188 443 200 477
rect 142 371 200 443
rect 142 337 154 371
rect 188 337 200 371
rect 142 325 200 337
rect 236 477 290 489
rect 236 443 248 477
rect 282 443 290 477
rect 835 485 889 497
rect 236 371 290 443
rect 236 337 248 371
rect 282 337 290 371
rect 236 325 290 337
rect 355 463 409 475
rect 355 429 363 463
rect 397 429 409 463
rect 355 363 409 429
rect 355 329 363 363
rect 397 329 409 363
rect 355 311 409 329
rect 445 463 503 475
rect 445 429 457 463
rect 491 429 503 463
rect 445 357 503 429
rect 445 323 457 357
rect 491 323 503 357
rect 445 311 503 323
rect 539 463 597 475
rect 539 429 551 463
rect 585 429 597 463
rect 539 357 597 429
rect 539 323 551 357
rect 585 323 597 357
rect 539 311 597 323
rect 633 463 691 475
rect 633 429 645 463
rect 679 429 691 463
rect 633 357 691 429
rect 633 323 645 357
rect 679 323 691 357
rect 633 311 691 323
rect 727 463 781 475
rect 727 429 739 463
rect 773 429 781 463
rect 727 357 781 429
rect 727 323 739 357
rect 773 323 781 357
rect 727 311 781 323
rect 835 451 843 485
rect 877 451 889 485
rect 835 417 889 451
rect 835 383 843 417
rect 877 383 889 417
rect 835 297 889 383
rect 925 485 983 497
rect 925 451 937 485
rect 971 451 983 485
rect 925 417 983 451
rect 925 383 937 417
rect 971 383 983 417
rect 925 349 983 383
rect 925 315 937 349
rect 971 315 983 349
rect 925 297 983 315
rect 1019 485 1077 497
rect 1019 451 1031 485
rect 1065 451 1077 485
rect 1019 417 1077 451
rect 1019 383 1031 417
rect 1065 383 1077 417
rect 1019 297 1077 383
rect 1113 485 1171 497
rect 1113 451 1125 485
rect 1159 451 1171 485
rect 1113 417 1171 451
rect 1113 383 1125 417
rect 1159 383 1171 417
rect 1113 349 1171 383
rect 1113 315 1125 349
rect 1159 315 1171 349
rect 1113 297 1171 315
rect 1207 485 1277 497
rect 1207 451 1225 485
rect 1259 451 1277 485
rect 1207 417 1277 451
rect 1207 383 1225 417
rect 1259 383 1277 417
rect 1207 349 1277 383
rect 1207 315 1225 349
rect 1259 315 1277 349
rect 1207 297 1277 315
rect 1313 485 1371 497
rect 1313 451 1325 485
rect 1359 451 1371 485
rect 1313 417 1371 451
rect 1313 383 1325 417
rect 1359 383 1371 417
rect 1313 349 1371 383
rect 1313 315 1325 349
rect 1359 315 1371 349
rect 1313 297 1371 315
rect 1407 485 1465 497
rect 1407 451 1419 485
rect 1453 451 1465 485
rect 1407 417 1465 451
rect 1407 383 1419 417
rect 1453 383 1465 417
rect 1407 297 1465 383
rect 1501 485 1559 497
rect 1501 451 1513 485
rect 1547 451 1559 485
rect 1501 417 1559 451
rect 1501 383 1513 417
rect 1547 383 1559 417
rect 1501 349 1559 383
rect 1501 315 1513 349
rect 1547 315 1559 349
rect 1501 297 1559 315
rect 1595 485 1649 497
rect 1595 451 1607 485
rect 1641 451 1649 485
rect 2194 477 2248 489
rect 1595 417 1649 451
rect 1595 383 1607 417
rect 1641 383 1649 417
rect 1595 297 1649 383
rect 1703 463 1757 475
rect 1703 429 1711 463
rect 1745 429 1757 463
rect 1703 357 1757 429
rect 1703 323 1711 357
rect 1745 323 1757 357
rect 1703 311 1757 323
rect 1793 463 1851 475
rect 1793 429 1805 463
rect 1839 429 1851 463
rect 1793 357 1851 429
rect 1793 323 1805 357
rect 1839 323 1851 357
rect 1793 311 1851 323
rect 1887 463 1945 475
rect 1887 429 1899 463
rect 1933 429 1945 463
rect 1887 357 1945 429
rect 1887 323 1899 357
rect 1933 323 1945 357
rect 1887 311 1945 323
rect 1981 463 2039 475
rect 1981 429 1993 463
rect 2027 429 2039 463
rect 1981 357 2039 429
rect 1981 323 1993 357
rect 2027 323 2039 357
rect 1981 311 2039 323
rect 2075 463 2129 475
rect 2075 429 2087 463
rect 2121 429 2129 463
rect 2075 363 2129 429
rect 2075 329 2087 363
rect 2121 329 2129 363
rect 2075 311 2129 329
rect 2194 443 2202 477
rect 2236 443 2248 477
rect 2194 371 2248 443
rect 2194 337 2202 371
rect 2236 337 2248 371
rect 2194 325 2248 337
rect 2284 477 2342 489
rect 2284 443 2296 477
rect 2330 443 2342 477
rect 2284 371 2342 443
rect 2284 337 2296 371
rect 2330 337 2342 371
rect 2284 325 2342 337
rect 2378 477 2432 489
rect 2378 443 2390 477
rect 2424 443 2432 477
rect 2378 371 2432 443
rect 2378 337 2390 371
rect 2424 337 2432 371
rect 2378 325 2432 337
rect 2536 477 2590 489
rect 2536 443 2544 477
rect 2578 443 2590 477
rect 2536 371 2590 443
rect 2536 337 2544 371
rect 2578 337 2590 371
rect 2536 325 2590 337
rect 2626 477 2684 489
rect 2626 443 2638 477
rect 2672 443 2684 477
rect 2626 371 2684 443
rect 2626 337 2638 371
rect 2672 337 2684 371
rect 2626 325 2684 337
rect 2720 477 2774 489
rect 2720 443 2732 477
rect 2766 443 2774 477
rect 3319 485 3373 497
rect 2720 371 2774 443
rect 2720 337 2732 371
rect 2766 337 2774 371
rect 2720 325 2774 337
rect 2839 463 2893 475
rect 2839 429 2847 463
rect 2881 429 2893 463
rect 2839 363 2893 429
rect 2839 329 2847 363
rect 2881 329 2893 363
rect 2839 311 2893 329
rect 2929 463 2987 475
rect 2929 429 2941 463
rect 2975 429 2987 463
rect 2929 357 2987 429
rect 2929 323 2941 357
rect 2975 323 2987 357
rect 2929 311 2987 323
rect 3023 463 3081 475
rect 3023 429 3035 463
rect 3069 429 3081 463
rect 3023 357 3081 429
rect 3023 323 3035 357
rect 3069 323 3081 357
rect 3023 311 3081 323
rect 3117 463 3175 475
rect 3117 429 3129 463
rect 3163 429 3175 463
rect 3117 357 3175 429
rect 3117 323 3129 357
rect 3163 323 3175 357
rect 3117 311 3175 323
rect 3211 463 3265 475
rect 3211 429 3223 463
rect 3257 429 3265 463
rect 3211 357 3265 429
rect 3211 323 3223 357
rect 3257 323 3265 357
rect 3211 311 3265 323
rect 3319 451 3327 485
rect 3361 451 3373 485
rect 3319 417 3373 451
rect 3319 383 3327 417
rect 3361 383 3373 417
rect 3319 297 3373 383
rect 3409 485 3467 497
rect 3409 451 3421 485
rect 3455 451 3467 485
rect 3409 417 3467 451
rect 3409 383 3421 417
rect 3455 383 3467 417
rect 3409 349 3467 383
rect 3409 315 3421 349
rect 3455 315 3467 349
rect 3409 297 3467 315
rect 3503 485 3561 497
rect 3503 451 3515 485
rect 3549 451 3561 485
rect 3503 417 3561 451
rect 3503 383 3515 417
rect 3549 383 3561 417
rect 3503 297 3561 383
rect 3597 485 3655 497
rect 3597 451 3609 485
rect 3643 451 3655 485
rect 3597 417 3655 451
rect 3597 383 3609 417
rect 3643 383 3655 417
rect 3597 349 3655 383
rect 3597 315 3609 349
rect 3643 315 3655 349
rect 3597 297 3655 315
rect 3691 485 3761 497
rect 3691 451 3709 485
rect 3743 451 3761 485
rect 3691 417 3761 451
rect 3691 383 3709 417
rect 3743 383 3761 417
rect 3691 349 3761 383
rect 3691 315 3709 349
rect 3743 315 3761 349
rect 3691 297 3761 315
rect 3797 485 3855 497
rect 3797 451 3809 485
rect 3843 451 3855 485
rect 3797 417 3855 451
rect 3797 383 3809 417
rect 3843 383 3855 417
rect 3797 349 3855 383
rect 3797 315 3809 349
rect 3843 315 3855 349
rect 3797 297 3855 315
rect 3891 485 3949 497
rect 3891 451 3903 485
rect 3937 451 3949 485
rect 3891 417 3949 451
rect 3891 383 3903 417
rect 3937 383 3949 417
rect 3891 297 3949 383
rect 3985 485 4043 497
rect 3985 451 3997 485
rect 4031 451 4043 485
rect 3985 417 4043 451
rect 3985 383 3997 417
rect 4031 383 4043 417
rect 3985 349 4043 383
rect 3985 315 3997 349
rect 4031 315 4043 349
rect 3985 297 4043 315
rect 4079 485 4133 497
rect 4079 451 4091 485
rect 4125 451 4133 485
rect 4678 477 4732 489
rect 4079 417 4133 451
rect 4079 383 4091 417
rect 4125 383 4133 417
rect 4079 297 4133 383
rect 4187 463 4241 475
rect 4187 429 4195 463
rect 4229 429 4241 463
rect 4187 357 4241 429
rect 4187 323 4195 357
rect 4229 323 4241 357
rect 4187 311 4241 323
rect 4277 463 4335 475
rect 4277 429 4289 463
rect 4323 429 4335 463
rect 4277 357 4335 429
rect 4277 323 4289 357
rect 4323 323 4335 357
rect 4277 311 4335 323
rect 4371 463 4429 475
rect 4371 429 4383 463
rect 4417 429 4429 463
rect 4371 357 4429 429
rect 4371 323 4383 357
rect 4417 323 4429 357
rect 4371 311 4429 323
rect 4465 463 4523 475
rect 4465 429 4477 463
rect 4511 429 4523 463
rect 4465 357 4523 429
rect 4465 323 4477 357
rect 4511 323 4523 357
rect 4465 311 4523 323
rect 4559 463 4613 475
rect 4559 429 4571 463
rect 4605 429 4613 463
rect 4559 363 4613 429
rect 4559 329 4571 363
rect 4605 329 4613 363
rect 4559 311 4613 329
rect 4678 443 4686 477
rect 4720 443 4732 477
rect 4678 371 4732 443
rect 4678 337 4686 371
rect 4720 337 4732 371
rect 4678 325 4732 337
rect 4768 477 4826 489
rect 4768 443 4780 477
rect 4814 443 4826 477
rect 4768 371 4826 443
rect 4768 337 4780 371
rect 4814 337 4826 371
rect 4768 325 4826 337
rect 4862 477 4916 489
rect 4862 443 4874 477
rect 4908 443 4916 477
rect 4862 371 4916 443
rect 4862 337 4874 371
rect 4908 337 4916 371
rect 4862 325 4916 337
<< ndiffc >>
rect 70 982 104 1016
rect 154 982 188 1016
rect 238 982 272 1016
rect 413 953 447 987
rect 497 935 531 969
rect 581 953 615 987
rect 665 935 699 969
rect 749 953 783 987
rect 853 995 887 1029
rect 937 995 971 1029
rect 937 927 971 961
rect 1031 995 1065 1029
rect 1125 995 1159 1029
rect 1125 927 1159 961
rect 1225 995 1259 1029
rect 1225 927 1259 961
rect 1325 995 1359 1029
rect 1325 927 1359 961
rect 1419 995 1453 1029
rect 1513 995 1547 1029
rect 1513 927 1547 961
rect 1597 995 1631 1029
rect 1701 953 1735 987
rect 1785 935 1819 969
rect 1869 953 1903 987
rect 1953 935 1987 969
rect 2037 953 2071 987
rect 2212 982 2246 1016
rect 2296 982 2330 1016
rect 2380 982 2414 1016
rect 2554 982 2588 1016
rect 2638 982 2672 1016
rect 2722 982 2756 1016
rect 2897 953 2931 987
rect 2981 935 3015 969
rect 3065 953 3099 987
rect 3149 935 3183 969
rect 3233 953 3267 987
rect 3337 995 3371 1029
rect 3421 995 3455 1029
rect 3421 927 3455 961
rect 3515 995 3549 1029
rect 3609 995 3643 1029
rect 3609 927 3643 961
rect 3709 995 3743 1029
rect 3709 927 3743 961
rect 3809 995 3843 1029
rect 3809 927 3843 961
rect 3903 995 3937 1029
rect 3997 995 4031 1029
rect 3997 927 4031 961
rect 4081 995 4115 1029
rect 4185 953 4219 987
rect 4269 935 4303 969
rect 4353 953 4387 987
rect 4437 935 4471 969
rect 4521 953 4555 987
rect 4696 982 4730 1016
rect 4780 982 4814 1016
rect 4864 982 4898 1016
rect 70 72 104 106
rect 154 72 188 106
rect 238 72 272 106
rect 413 101 447 135
rect 497 119 531 153
rect 581 101 615 135
rect 665 119 699 153
rect 749 101 783 135
rect 853 59 887 93
rect 937 127 971 161
rect 937 59 971 93
rect 1031 59 1065 93
rect 1125 127 1159 161
rect 1125 59 1159 93
rect 1225 127 1259 161
rect 1225 59 1259 93
rect 1325 127 1359 161
rect 1325 59 1359 93
rect 1419 59 1453 93
rect 1513 127 1547 161
rect 1513 59 1547 93
rect 1597 59 1631 93
rect 1701 101 1735 135
rect 1785 119 1819 153
rect 1869 101 1903 135
rect 1953 119 1987 153
rect 2037 101 2071 135
rect 2212 72 2246 106
rect 2296 72 2330 106
rect 2380 72 2414 106
rect 2554 72 2588 106
rect 2638 72 2672 106
rect 2722 72 2756 106
rect 2897 101 2931 135
rect 2981 119 3015 153
rect 3065 101 3099 135
rect 3149 119 3183 153
rect 3233 101 3267 135
rect 3337 59 3371 93
rect 3421 127 3455 161
rect 3421 59 3455 93
rect 3515 59 3549 93
rect 3609 127 3643 161
rect 3609 59 3643 93
rect 3709 127 3743 161
rect 3709 59 3743 93
rect 3809 127 3843 161
rect 3809 59 3843 93
rect 3903 59 3937 93
rect 3997 127 4031 161
rect 3997 59 4031 93
rect 4081 59 4115 93
rect 4185 101 4219 135
rect 4269 119 4303 153
rect 4353 101 4387 135
rect 4437 119 4471 153
rect 4521 101 4555 135
rect 4696 72 4730 106
rect 4780 72 4814 106
rect 4864 72 4898 106
<< pdiffc >>
rect 60 717 94 751
rect 60 611 94 645
rect 154 717 188 751
rect 154 611 188 645
rect 248 717 282 751
rect 248 611 282 645
rect 363 725 397 759
rect 363 625 397 659
rect 457 731 491 765
rect 457 625 491 659
rect 551 731 585 765
rect 551 625 585 659
rect 645 731 679 765
rect 645 625 679 659
rect 739 731 773 765
rect 739 625 773 659
rect 843 671 877 705
rect 843 603 877 637
rect 937 739 971 773
rect 937 671 971 705
rect 937 603 971 637
rect 1031 671 1065 705
rect 1031 603 1065 637
rect 1125 739 1159 773
rect 1125 671 1159 705
rect 1125 603 1159 637
rect 1225 739 1259 773
rect 1225 671 1259 705
rect 1225 603 1259 637
rect 1325 739 1359 773
rect 1325 671 1359 705
rect 1325 603 1359 637
rect 1419 671 1453 705
rect 1419 603 1453 637
rect 1513 739 1547 773
rect 1513 671 1547 705
rect 1513 603 1547 637
rect 1607 671 1641 705
rect 1607 603 1641 637
rect 1711 731 1745 765
rect 1711 625 1745 659
rect 1805 731 1839 765
rect 1805 625 1839 659
rect 1899 731 1933 765
rect 1899 625 1933 659
rect 1993 731 2027 765
rect 1993 625 2027 659
rect 2087 725 2121 759
rect 2087 625 2121 659
rect 2202 717 2236 751
rect 2202 611 2236 645
rect 2296 717 2330 751
rect 2296 611 2330 645
rect 2390 717 2424 751
rect 2390 611 2424 645
rect 2544 717 2578 751
rect 2544 611 2578 645
rect 2638 717 2672 751
rect 2638 611 2672 645
rect 2732 717 2766 751
rect 2732 611 2766 645
rect 2847 725 2881 759
rect 2847 625 2881 659
rect 2941 731 2975 765
rect 2941 625 2975 659
rect 3035 731 3069 765
rect 3035 625 3069 659
rect 3129 731 3163 765
rect 3129 625 3163 659
rect 3223 731 3257 765
rect 3223 625 3257 659
rect 3327 671 3361 705
rect 3327 603 3361 637
rect 3421 739 3455 773
rect 3421 671 3455 705
rect 3421 603 3455 637
rect 3515 671 3549 705
rect 3515 603 3549 637
rect 3609 739 3643 773
rect 3609 671 3643 705
rect 3609 603 3643 637
rect 3709 739 3743 773
rect 3709 671 3743 705
rect 3709 603 3743 637
rect 3809 739 3843 773
rect 3809 671 3843 705
rect 3809 603 3843 637
rect 3903 671 3937 705
rect 3903 603 3937 637
rect 3997 739 4031 773
rect 3997 671 4031 705
rect 3997 603 4031 637
rect 4091 671 4125 705
rect 4091 603 4125 637
rect 4195 731 4229 765
rect 4195 625 4229 659
rect 4289 731 4323 765
rect 4289 625 4323 659
rect 4383 731 4417 765
rect 4383 625 4417 659
rect 4477 731 4511 765
rect 4477 625 4511 659
rect 4571 725 4605 759
rect 4571 625 4605 659
rect 4686 717 4720 751
rect 4686 611 4720 645
rect 4780 717 4814 751
rect 4780 611 4814 645
rect 4874 717 4908 751
rect 4874 611 4908 645
rect 60 443 94 477
rect 60 337 94 371
rect 154 443 188 477
rect 154 337 188 371
rect 248 443 282 477
rect 248 337 282 371
rect 363 429 397 463
rect 363 329 397 363
rect 457 429 491 463
rect 457 323 491 357
rect 551 429 585 463
rect 551 323 585 357
rect 645 429 679 463
rect 645 323 679 357
rect 739 429 773 463
rect 739 323 773 357
rect 843 451 877 485
rect 843 383 877 417
rect 937 451 971 485
rect 937 383 971 417
rect 937 315 971 349
rect 1031 451 1065 485
rect 1031 383 1065 417
rect 1125 451 1159 485
rect 1125 383 1159 417
rect 1125 315 1159 349
rect 1225 451 1259 485
rect 1225 383 1259 417
rect 1225 315 1259 349
rect 1325 451 1359 485
rect 1325 383 1359 417
rect 1325 315 1359 349
rect 1419 451 1453 485
rect 1419 383 1453 417
rect 1513 451 1547 485
rect 1513 383 1547 417
rect 1513 315 1547 349
rect 1607 451 1641 485
rect 1607 383 1641 417
rect 1711 429 1745 463
rect 1711 323 1745 357
rect 1805 429 1839 463
rect 1805 323 1839 357
rect 1899 429 1933 463
rect 1899 323 1933 357
rect 1993 429 2027 463
rect 1993 323 2027 357
rect 2087 429 2121 463
rect 2087 329 2121 363
rect 2202 443 2236 477
rect 2202 337 2236 371
rect 2296 443 2330 477
rect 2296 337 2330 371
rect 2390 443 2424 477
rect 2390 337 2424 371
rect 2544 443 2578 477
rect 2544 337 2578 371
rect 2638 443 2672 477
rect 2638 337 2672 371
rect 2732 443 2766 477
rect 2732 337 2766 371
rect 2847 429 2881 463
rect 2847 329 2881 363
rect 2941 429 2975 463
rect 2941 323 2975 357
rect 3035 429 3069 463
rect 3035 323 3069 357
rect 3129 429 3163 463
rect 3129 323 3163 357
rect 3223 429 3257 463
rect 3223 323 3257 357
rect 3327 451 3361 485
rect 3327 383 3361 417
rect 3421 451 3455 485
rect 3421 383 3455 417
rect 3421 315 3455 349
rect 3515 451 3549 485
rect 3515 383 3549 417
rect 3609 451 3643 485
rect 3609 383 3643 417
rect 3609 315 3643 349
rect 3709 451 3743 485
rect 3709 383 3743 417
rect 3709 315 3743 349
rect 3809 451 3843 485
rect 3809 383 3843 417
rect 3809 315 3843 349
rect 3903 451 3937 485
rect 3903 383 3937 417
rect 3997 451 4031 485
rect 3997 383 4031 417
rect 3997 315 4031 349
rect 4091 451 4125 485
rect 4091 383 4125 417
rect 4195 429 4229 463
rect 4195 323 4229 357
rect 4289 429 4323 463
rect 4289 323 4323 357
rect 4383 429 4417 463
rect 4383 323 4417 357
rect 4477 429 4511 463
rect 4477 323 4511 357
rect 4571 429 4605 463
rect 4571 329 4605 363
rect 4686 443 4720 477
rect 4686 337 4720 371
rect 4780 443 4814 477
rect 4780 337 4814 371
rect 4874 443 4908 477
rect 4874 337 4908 371
<< poly >>
rect 114 1041 144 1067
rect 198 1041 228 1067
rect 305 1037 739 1067
rect 897 1041 927 1067
rect 981 1041 1011 1069
rect 1085 1041 1115 1067
rect 1169 1041 1199 1069
rect 1285 1041 1315 1069
rect 1369 1041 1399 1067
rect 1473 1041 1503 1069
rect 1557 1041 1587 1067
rect 114 941 144 957
rect 198 941 228 957
rect 305 941 335 1037
rect 457 1022 487 1037
rect 541 1022 571 1037
rect 625 1022 655 1037
rect 709 1022 739 1037
rect 114 911 335 941
rect 114 889 144 911
rect 21 873 144 889
rect 21 839 31 873
rect 65 839 99 873
rect 133 839 144 873
rect 21 823 144 839
rect 104 778 144 823
rect 198 778 238 911
rect 457 892 487 918
rect 541 892 571 918
rect 625 892 655 918
rect 709 892 739 918
rect 1745 1037 2179 1067
rect 2256 1041 2286 1067
rect 2340 1041 2370 1067
rect 2598 1041 2628 1067
rect 2682 1041 2712 1067
rect 1745 1022 1775 1037
rect 1829 1022 1859 1037
rect 1913 1022 1943 1037
rect 1997 1022 2027 1037
rect 2149 941 2179 1037
rect 2789 1037 3223 1067
rect 3381 1041 3411 1067
rect 3465 1041 3495 1069
rect 3569 1041 3599 1067
rect 3653 1041 3683 1069
rect 3769 1041 3799 1069
rect 3853 1041 3883 1067
rect 3957 1041 3987 1069
rect 4041 1041 4071 1067
rect 2256 941 2286 957
rect 2340 941 2370 957
rect 897 883 927 911
rect 981 883 1011 911
rect 1085 883 1115 911
rect 1169 883 1199 911
rect 1285 883 1315 911
rect 1369 883 1399 911
rect 1473 883 1503 911
rect 1557 883 1587 911
rect 1745 892 1775 918
rect 1829 892 1859 918
rect 1913 892 1943 918
rect 1997 892 2027 918
rect 2149 911 2370 941
rect 887 873 1209 883
rect 280 859 414 869
rect 280 825 296 859
rect 330 825 364 859
rect 398 825 414 859
rect 887 839 947 873
rect 981 839 1015 873
rect 1049 839 1083 873
rect 1117 839 1151 873
rect 1185 839 1209 873
rect 887 829 1209 839
rect 1275 873 1597 883
rect 1275 839 1299 873
rect 1333 839 1367 873
rect 1401 839 1435 873
rect 1469 839 1503 873
rect 1537 839 1597 873
rect 1275 829 1597 839
rect 2070 859 2204 869
rect 280 823 414 825
rect 280 815 729 823
rect 363 793 729 815
rect 106 763 142 778
rect 200 763 236 778
rect 409 777 445 793
rect 503 777 539 793
rect 597 777 633 793
rect 691 777 727 793
rect 889 791 925 829
rect 983 791 1019 829
rect 1077 791 1113 829
rect 1171 791 1207 829
rect 1277 791 1313 829
rect 1371 791 1407 829
rect 1465 791 1501 829
rect 1559 791 1595 829
rect 2070 825 2086 859
rect 2120 825 2154 859
rect 2188 825 2204 859
rect 2070 823 2204 825
rect 1755 815 2204 823
rect 1755 793 2121 815
rect 106 565 142 599
rect 200 565 236 599
rect 409 565 445 613
rect 503 565 539 613
rect 597 565 633 613
rect 691 565 727 613
rect 1757 777 1793 793
rect 1851 777 1887 793
rect 1945 777 1981 793
rect 2039 777 2075 793
rect 2246 778 2286 911
rect 2340 889 2370 911
rect 2598 941 2628 957
rect 2682 941 2712 957
rect 2789 941 2819 1037
rect 2941 1022 2971 1037
rect 3025 1022 3055 1037
rect 3109 1022 3139 1037
rect 3193 1022 3223 1037
rect 2598 911 2819 941
rect 2598 889 2628 911
rect 2340 873 2463 889
rect 2340 839 2351 873
rect 2385 839 2419 873
rect 2453 839 2463 873
rect 2340 823 2463 839
rect 2505 873 2628 889
rect 2505 839 2515 873
rect 2549 839 2583 873
rect 2617 839 2628 873
rect 2505 823 2628 839
rect 2340 778 2380 823
rect 2588 778 2628 823
rect 2682 778 2722 911
rect 2941 892 2971 918
rect 3025 892 3055 918
rect 3109 892 3139 918
rect 3193 892 3223 918
rect 4229 1037 4663 1067
rect 4740 1041 4770 1067
rect 4824 1041 4854 1067
rect 4229 1022 4259 1037
rect 4313 1022 4343 1037
rect 4397 1022 4427 1037
rect 4481 1022 4511 1037
rect 4633 941 4663 1037
rect 4740 941 4770 957
rect 4824 941 4854 957
rect 3381 883 3411 911
rect 3465 883 3495 911
rect 3569 883 3599 911
rect 3653 883 3683 911
rect 3769 883 3799 911
rect 3853 883 3883 911
rect 3957 883 3987 911
rect 4041 883 4071 911
rect 4229 892 4259 918
rect 4313 892 4343 918
rect 4397 892 4427 918
rect 4481 892 4511 918
rect 4633 911 4854 941
rect 3371 873 3693 883
rect 2764 859 2898 869
rect 2764 825 2780 859
rect 2814 825 2848 859
rect 2882 825 2898 859
rect 3371 839 3431 873
rect 3465 839 3499 873
rect 3533 839 3567 873
rect 3601 839 3635 873
rect 3669 839 3693 873
rect 3371 829 3693 839
rect 3759 873 4081 883
rect 3759 839 3783 873
rect 3817 839 3851 873
rect 3885 839 3919 873
rect 3953 839 3987 873
rect 4021 839 4081 873
rect 3759 829 4081 839
rect 4554 859 4688 869
rect 2764 823 2898 825
rect 2764 815 3213 823
rect 2847 793 3213 815
rect 2248 763 2284 778
rect 2342 763 2378 778
rect 2590 763 2626 778
rect 2684 763 2720 778
rect 2893 777 2929 793
rect 2987 777 3023 793
rect 3081 777 3117 793
rect 3175 777 3211 793
rect 3373 791 3409 829
rect 3467 791 3503 829
rect 3561 791 3597 829
rect 3655 791 3691 829
rect 3761 791 3797 829
rect 3855 791 3891 829
rect 3949 791 3985 829
rect 4043 791 4079 829
rect 4554 825 4570 859
rect 4604 825 4638 859
rect 4672 825 4688 859
rect 4554 823 4688 825
rect 4239 815 4688 823
rect 4239 793 4605 815
rect 889 565 925 591
rect 983 565 1019 591
rect 1077 565 1113 591
rect 1171 565 1207 591
rect 1277 565 1313 591
rect 1371 565 1407 591
rect 1465 565 1501 591
rect 1559 565 1595 591
rect 1757 565 1793 613
rect 1851 565 1887 613
rect 1945 565 1981 613
rect 2039 565 2075 613
rect 2248 565 2284 599
rect 2342 565 2378 599
rect 2590 565 2626 599
rect 2684 565 2720 599
rect 2893 565 2929 613
rect 2987 565 3023 613
rect 3081 565 3117 613
rect 3175 565 3211 613
rect 4241 777 4277 793
rect 4335 777 4371 793
rect 4429 777 4465 793
rect 4523 777 4559 793
rect 4730 778 4770 911
rect 4824 889 4854 911
rect 4824 873 4947 889
rect 4824 839 4835 873
rect 4869 839 4903 873
rect 4937 839 4947 873
rect 4824 823 4947 839
rect 4824 778 4864 823
rect 4732 763 4768 778
rect 4826 763 4862 778
rect 3373 565 3409 591
rect 3467 565 3503 591
rect 3561 565 3597 591
rect 3655 565 3691 591
rect 3761 565 3797 591
rect 3855 565 3891 591
rect 3949 565 3985 591
rect 4043 565 4079 591
rect 4241 565 4277 613
rect 4335 565 4371 613
rect 4429 565 4465 613
rect 4523 565 4559 613
rect 4732 565 4768 599
rect 4826 565 4862 599
rect 106 489 142 523
rect 200 489 236 523
rect 409 475 445 523
rect 503 475 539 523
rect 597 475 633 523
rect 691 475 727 523
rect 889 497 925 523
rect 983 497 1019 523
rect 1077 497 1113 523
rect 1171 497 1207 523
rect 1277 497 1313 523
rect 1371 497 1407 523
rect 1465 497 1501 523
rect 1559 497 1595 523
rect 106 310 142 325
rect 200 310 236 325
rect 104 265 144 310
rect 21 249 144 265
rect 21 215 31 249
rect 65 215 99 249
rect 133 215 144 249
rect 21 199 144 215
rect 114 177 144 199
rect 198 177 238 310
rect 409 295 445 311
rect 503 295 539 311
rect 597 295 633 311
rect 691 295 727 311
rect 1757 475 1793 523
rect 1851 475 1887 523
rect 1945 475 1981 523
rect 2039 475 2075 523
rect 2248 489 2284 523
rect 2342 489 2378 523
rect 2590 489 2626 523
rect 2684 489 2720 523
rect 2893 475 2929 523
rect 2987 475 3023 523
rect 3081 475 3117 523
rect 3175 475 3211 523
rect 3373 497 3409 523
rect 3467 497 3503 523
rect 3561 497 3597 523
rect 3655 497 3691 523
rect 3761 497 3797 523
rect 3855 497 3891 523
rect 3949 497 3985 523
rect 4043 497 4079 523
rect 363 273 729 295
rect 280 265 729 273
rect 280 263 414 265
rect 280 229 296 263
rect 330 229 364 263
rect 398 229 414 263
rect 889 259 925 297
rect 983 259 1019 297
rect 1077 259 1113 297
rect 1171 259 1207 297
rect 1277 259 1313 297
rect 1371 259 1407 297
rect 1465 259 1501 297
rect 1559 259 1595 297
rect 1757 295 1793 311
rect 1851 295 1887 311
rect 1945 295 1981 311
rect 2039 295 2075 311
rect 2248 310 2284 325
rect 2342 310 2378 325
rect 2590 310 2626 325
rect 2684 310 2720 325
rect 1755 273 2121 295
rect 1755 265 2204 273
rect 2070 263 2204 265
rect 280 219 414 229
rect 887 249 1209 259
rect 887 215 947 249
rect 981 215 1015 249
rect 1049 215 1083 249
rect 1117 215 1151 249
rect 1185 215 1209 249
rect 887 205 1209 215
rect 1275 249 1597 259
rect 1275 215 1299 249
rect 1333 215 1367 249
rect 1401 215 1435 249
rect 1469 215 1503 249
rect 1537 215 1597 249
rect 2070 229 2086 263
rect 2120 229 2154 263
rect 2188 229 2204 263
rect 2070 219 2204 229
rect 1275 205 1597 215
rect 114 147 335 177
rect 457 170 487 196
rect 541 170 571 196
rect 625 170 655 196
rect 709 170 739 196
rect 897 177 927 205
rect 981 177 1011 205
rect 1085 177 1115 205
rect 1169 177 1199 205
rect 1285 177 1315 205
rect 1369 177 1399 205
rect 1473 177 1503 205
rect 1557 177 1587 205
rect 114 131 144 147
rect 198 131 228 147
rect 305 51 335 147
rect 457 51 487 66
rect 541 51 571 66
rect 625 51 655 66
rect 709 51 739 66
rect 114 21 144 47
rect 198 21 228 47
rect 305 21 739 51
rect 1745 170 1775 196
rect 1829 170 1859 196
rect 1913 170 1943 196
rect 1997 170 2027 196
rect 2246 177 2286 310
rect 2340 265 2380 310
rect 2588 265 2628 310
rect 2340 249 2463 265
rect 2340 215 2351 249
rect 2385 215 2419 249
rect 2453 215 2463 249
rect 2340 199 2463 215
rect 2505 249 2628 265
rect 2505 215 2515 249
rect 2549 215 2583 249
rect 2617 215 2628 249
rect 2505 199 2628 215
rect 2340 177 2370 199
rect 2149 147 2370 177
rect 1745 51 1775 66
rect 1829 51 1859 66
rect 1913 51 1943 66
rect 1997 51 2027 66
rect 2149 51 2179 147
rect 2256 131 2286 147
rect 2340 131 2370 147
rect 2598 177 2628 199
rect 2682 177 2722 310
rect 2893 295 2929 311
rect 2987 295 3023 311
rect 3081 295 3117 311
rect 3175 295 3211 311
rect 4241 475 4277 523
rect 4335 475 4371 523
rect 4429 475 4465 523
rect 4523 475 4559 523
rect 4732 489 4768 523
rect 4826 489 4862 523
rect 2847 273 3213 295
rect 2764 265 3213 273
rect 2764 263 2898 265
rect 2764 229 2780 263
rect 2814 229 2848 263
rect 2882 229 2898 263
rect 3373 259 3409 297
rect 3467 259 3503 297
rect 3561 259 3597 297
rect 3655 259 3691 297
rect 3761 259 3797 297
rect 3855 259 3891 297
rect 3949 259 3985 297
rect 4043 259 4079 297
rect 4241 295 4277 311
rect 4335 295 4371 311
rect 4429 295 4465 311
rect 4523 295 4559 311
rect 4732 310 4768 325
rect 4826 310 4862 325
rect 4239 273 4605 295
rect 4239 265 4688 273
rect 4554 263 4688 265
rect 2764 219 2898 229
rect 3371 249 3693 259
rect 3371 215 3431 249
rect 3465 215 3499 249
rect 3533 215 3567 249
rect 3601 215 3635 249
rect 3669 215 3693 249
rect 3371 205 3693 215
rect 3759 249 4081 259
rect 3759 215 3783 249
rect 3817 215 3851 249
rect 3885 215 3919 249
rect 3953 215 3987 249
rect 4021 215 4081 249
rect 4554 229 4570 263
rect 4604 229 4638 263
rect 4672 229 4688 263
rect 4554 219 4688 229
rect 3759 205 4081 215
rect 2598 147 2819 177
rect 2941 170 2971 196
rect 3025 170 3055 196
rect 3109 170 3139 196
rect 3193 170 3223 196
rect 3381 177 3411 205
rect 3465 177 3495 205
rect 3569 177 3599 205
rect 3653 177 3683 205
rect 3769 177 3799 205
rect 3853 177 3883 205
rect 3957 177 3987 205
rect 4041 177 4071 205
rect 2598 131 2628 147
rect 2682 131 2712 147
rect 897 21 927 47
rect 981 19 1011 47
rect 1085 21 1115 47
rect 1169 19 1199 47
rect 1285 19 1315 47
rect 1369 21 1399 47
rect 1473 19 1503 47
rect 1557 21 1587 47
rect 1745 21 2179 51
rect 2789 51 2819 147
rect 2941 51 2971 66
rect 3025 51 3055 66
rect 3109 51 3139 66
rect 3193 51 3223 66
rect 2256 21 2286 47
rect 2340 21 2370 47
rect 2598 21 2628 47
rect 2682 21 2712 47
rect 2789 21 3223 51
rect 4229 170 4259 196
rect 4313 170 4343 196
rect 4397 170 4427 196
rect 4481 170 4511 196
rect 4730 177 4770 310
rect 4824 265 4864 310
rect 4824 249 4947 265
rect 4824 215 4835 249
rect 4869 215 4903 249
rect 4937 215 4947 249
rect 4824 199 4947 215
rect 4824 177 4854 199
rect 4633 147 4854 177
rect 4229 51 4259 66
rect 4313 51 4343 66
rect 4397 51 4427 66
rect 4481 51 4511 66
rect 4633 51 4663 147
rect 4740 131 4770 147
rect 4824 131 4854 147
rect 3381 21 3411 47
rect 3465 19 3495 47
rect 3569 21 3599 47
rect 3653 19 3683 47
rect 3769 19 3799 47
rect 3853 21 3883 47
rect 3957 19 3987 47
rect 4041 21 4071 47
rect 4229 21 4663 51
rect 4740 21 4770 47
rect 4824 21 4854 47
<< polycont >>
rect 31 839 65 873
rect 99 839 133 873
rect 296 825 330 859
rect 364 825 398 859
rect 947 839 981 873
rect 1015 839 1049 873
rect 1083 839 1117 873
rect 1151 839 1185 873
rect 1299 839 1333 873
rect 1367 839 1401 873
rect 1435 839 1469 873
rect 1503 839 1537 873
rect 2086 825 2120 859
rect 2154 825 2188 859
rect 2351 839 2385 873
rect 2419 839 2453 873
rect 2515 839 2549 873
rect 2583 839 2617 873
rect 2780 825 2814 859
rect 2848 825 2882 859
rect 3431 839 3465 873
rect 3499 839 3533 873
rect 3567 839 3601 873
rect 3635 839 3669 873
rect 3783 839 3817 873
rect 3851 839 3885 873
rect 3919 839 3953 873
rect 3987 839 4021 873
rect 4570 825 4604 859
rect 4638 825 4672 859
rect 4835 839 4869 873
rect 4903 839 4937 873
rect 31 215 65 249
rect 99 215 133 249
rect 296 229 330 263
rect 364 229 398 263
rect 947 215 981 249
rect 1015 215 1049 249
rect 1083 215 1117 249
rect 1151 215 1185 249
rect 1299 215 1333 249
rect 1367 215 1401 249
rect 1435 215 1469 249
rect 1503 215 1537 249
rect 2086 229 2120 263
rect 2154 229 2188 263
rect 2351 215 2385 249
rect 2419 215 2453 249
rect 2515 215 2549 249
rect 2583 215 2617 249
rect 2780 229 2814 263
rect 2848 229 2882 263
rect 3431 215 3465 249
rect 3499 215 3533 249
rect 3567 215 3601 249
rect 3635 215 3669 249
rect 3783 215 3817 249
rect 3851 215 3885 249
rect 3919 215 3953 249
rect 3987 215 4021 249
rect 4570 229 4604 263
rect 4638 229 4672 263
rect 4835 215 4869 249
rect 4903 215 4937 249
<< locali >>
rect 0 1071 29 1105
rect 63 1071 121 1105
rect 155 1071 213 1105
rect 247 1071 305 1105
rect 339 1071 397 1105
rect 431 1071 489 1105
rect 523 1071 581 1105
rect 615 1071 673 1105
rect 707 1071 765 1105
rect 799 1071 857 1105
rect 891 1071 949 1105
rect 983 1071 1041 1105
rect 1075 1071 1133 1105
rect 1167 1071 1225 1105
rect 1259 1071 1317 1105
rect 1351 1071 1409 1105
rect 1443 1071 1501 1105
rect 1535 1071 1593 1105
rect 1627 1071 1685 1105
rect 1719 1071 1777 1105
rect 1811 1071 1869 1105
rect 1903 1071 1961 1105
rect 1995 1071 2053 1105
rect 2087 1071 2145 1105
rect 2179 1071 2237 1105
rect 2271 1071 2329 1105
rect 2363 1071 2421 1105
rect 2455 1071 2513 1105
rect 2547 1071 2605 1105
rect 2639 1071 2697 1105
rect 2731 1071 2789 1105
rect 2823 1071 2881 1105
rect 2915 1071 2973 1105
rect 3007 1071 3065 1105
rect 3099 1071 3157 1105
rect 3191 1071 3249 1105
rect 3283 1071 3341 1105
rect 3375 1071 3433 1105
rect 3467 1071 3525 1105
rect 3559 1071 3617 1105
rect 3651 1071 3709 1105
rect 3743 1071 3801 1105
rect 3835 1071 3893 1105
rect 3927 1071 3985 1105
rect 4019 1071 4077 1105
rect 4111 1071 4169 1105
rect 4203 1071 4261 1105
rect 4295 1071 4353 1105
rect 4387 1071 4445 1105
rect 4479 1071 4537 1105
rect 4571 1071 4629 1105
rect 4663 1071 4721 1105
rect 4755 1071 4813 1105
rect 4847 1071 4905 1105
rect 4939 1071 4968 1105
rect 54 1016 112 1071
rect 54 982 70 1016
rect 104 982 112 1016
rect 54 966 112 982
rect 154 1016 204 1032
rect 188 982 204 1016
rect 154 923 204 982
rect 238 1016 296 1071
rect 272 982 296 1016
rect 238 966 296 982
rect 397 1003 803 1037
rect 397 987 447 1003
rect 397 953 413 987
rect 581 987 615 1003
rect 397 934 447 953
rect 481 935 497 969
rect 531 935 547 969
rect 17 873 136 889
rect 17 839 31 873
rect 65 839 99 873
rect 133 839 136 873
rect 17 823 136 839
rect 170 875 204 923
rect 481 875 547 935
rect 749 987 803 1003
rect 581 934 615 953
rect 649 935 665 969
rect 699 935 715 969
rect 649 911 715 935
rect 783 953 803 987
rect 837 1029 887 1071
rect 837 995 853 1029
rect 837 979 887 995
rect 921 1029 987 1037
rect 921 995 937 1029
rect 971 995 987 1029
rect 749 945 803 953
rect 921 961 987 995
rect 1021 1029 1075 1071
rect 1021 995 1031 1029
rect 1065 995 1075 1029
rect 1021 979 1075 995
rect 1109 1029 1175 1037
rect 1109 995 1125 1029
rect 1159 995 1175 1029
rect 921 945 937 961
rect 749 927 937 945
rect 971 945 987 961
rect 1109 961 1175 995
rect 1109 945 1125 961
rect 971 927 1125 945
rect 1159 927 1175 961
rect 749 911 1175 927
rect 1209 1029 1275 1071
rect 1209 995 1225 1029
rect 1259 995 1275 1029
rect 1209 961 1275 995
rect 1209 927 1225 961
rect 1259 927 1275 961
rect 1209 911 1275 927
rect 1309 1029 1375 1037
rect 1309 995 1325 1029
rect 1359 995 1375 1029
rect 1309 961 1375 995
rect 1409 1029 1463 1071
rect 1409 995 1419 1029
rect 1453 995 1463 1029
rect 1409 979 1463 995
rect 1497 1029 1563 1037
rect 1497 995 1513 1029
rect 1547 995 1563 1029
rect 1309 927 1325 961
rect 1359 945 1375 961
rect 1497 961 1563 995
rect 1597 1029 1647 1071
rect 1631 995 1647 1029
rect 1597 979 1647 995
rect 1681 1003 2087 1037
rect 1681 987 1735 1003
rect 1497 945 1513 961
rect 1359 927 1513 945
rect 1547 945 1563 961
rect 1681 953 1701 987
rect 1869 987 1903 1003
rect 1681 945 1735 953
rect 1547 927 1735 945
rect 1309 911 1735 927
rect 1769 935 1785 969
rect 1819 935 1835 969
rect 1769 911 1835 935
rect 2037 987 2087 1003
rect 1869 934 1903 953
rect 1937 935 1953 969
rect 1987 935 2003 969
rect 649 875 695 911
rect 170 859 407 875
rect 170 825 296 859
rect 330 825 364 859
rect 398 825 407 859
rect 170 809 407 825
rect 441 815 695 875
rect 931 873 1209 877
rect 931 839 947 873
rect 981 839 1015 873
rect 1049 839 1083 873
rect 1117 839 1151 873
rect 1185 839 1209 873
rect 931 823 1209 839
rect 1275 873 1553 877
rect 1275 839 1299 873
rect 1333 839 1367 873
rect 1401 839 1435 873
rect 1469 839 1503 873
rect 1537 839 1553 873
rect 1275 823 1553 839
rect 1789 875 1835 911
rect 1937 875 2003 935
rect 2071 953 2087 987
rect 2188 1016 2246 1071
rect 2188 982 2212 1016
rect 2188 966 2246 982
rect 2280 1016 2330 1032
rect 2280 982 2296 1016
rect 2037 934 2087 953
rect 2280 923 2330 982
rect 2372 1016 2430 1071
rect 2372 982 2380 1016
rect 2414 982 2430 1016
rect 2372 966 2430 982
rect 2538 1016 2596 1071
rect 2538 982 2554 1016
rect 2588 982 2596 1016
rect 2538 966 2596 982
rect 2638 1016 2688 1032
rect 2672 982 2688 1016
rect 2638 923 2688 982
rect 2722 1016 2780 1071
rect 2756 982 2780 1016
rect 2722 966 2780 982
rect 2881 1003 3287 1037
rect 2881 987 2931 1003
rect 2881 953 2897 987
rect 3065 987 3099 1003
rect 2881 934 2931 953
rect 2965 935 2981 969
rect 3015 935 3031 969
rect 2280 875 2314 923
rect 170 767 204 809
rect 44 751 104 767
rect 44 717 60 751
rect 94 717 104 751
rect 44 645 104 717
rect 44 611 60 645
rect 94 611 104 645
rect 44 561 104 611
rect 138 751 204 767
rect 138 717 154 751
rect 188 717 204 751
rect 138 645 204 717
rect 138 611 154 645
rect 188 611 204 645
rect 138 595 204 611
rect 243 751 298 767
rect 243 717 248 751
rect 282 717 298 751
rect 243 645 298 717
rect 243 611 248 645
rect 282 611 298 645
rect 243 561 298 611
rect 347 759 407 775
rect 347 725 363 759
rect 397 725 407 759
rect 347 660 407 725
rect 347 626 361 660
rect 395 659 407 660
rect 347 625 363 626
rect 397 625 407 659
rect 347 595 407 625
rect 441 765 507 815
rect 441 697 457 765
rect 491 697 507 765
rect 441 659 507 697
rect 441 625 457 659
rect 491 625 507 659
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 407 561
rect 44 477 104 527
rect 44 443 60 477
rect 94 443 104 477
rect 44 371 104 443
rect 44 337 60 371
rect 94 337 104 371
rect 44 321 104 337
rect 138 477 204 493
rect 138 443 154 477
rect 188 443 204 477
rect 138 371 204 443
rect 138 337 154 371
rect 188 337 204 371
rect 138 321 204 337
rect 243 477 298 527
rect 243 443 248 477
rect 282 443 298 477
rect 243 371 298 443
rect 243 337 248 371
rect 282 337 298 371
rect 243 321 298 337
rect 347 463 407 493
rect 347 462 363 463
rect 347 428 361 462
rect 397 429 407 463
rect 395 428 407 429
rect 347 363 407 428
rect 347 329 363 363
rect 397 329 407 363
rect 170 279 204 321
rect 347 313 407 329
rect 441 463 507 625
rect 541 765 595 781
rect 541 731 551 765
rect 585 731 595 765
rect 541 660 595 731
rect 541 625 551 660
rect 585 625 595 660
rect 541 595 595 625
rect 629 765 695 815
rect 1789 815 2043 875
rect 629 697 645 765
rect 679 697 695 765
rect 629 659 695 697
rect 629 625 645 659
rect 679 625 695 659
rect 441 429 457 463
rect 491 429 507 463
rect 441 391 507 429
rect 441 323 457 391
rect 491 323 507 391
rect 17 249 136 265
rect 17 215 31 249
rect 65 215 99 249
rect 133 215 136 249
rect 17 199 136 215
rect 170 263 407 279
rect 170 229 296 263
rect 330 229 364 263
rect 398 229 407 263
rect 170 213 407 229
rect 441 273 507 323
rect 541 463 595 493
rect 541 428 551 463
rect 585 428 595 463
rect 541 357 595 428
rect 541 323 551 357
rect 585 323 595 357
rect 541 307 595 323
rect 629 463 695 625
rect 729 773 1175 789
rect 729 765 937 773
rect 729 731 739 765
rect 773 755 937 765
rect 773 731 789 755
rect 729 660 789 731
rect 921 739 937 755
rect 971 755 1125 773
rect 971 739 987 755
rect 729 659 741 660
rect 729 625 739 659
rect 775 626 789 660
rect 773 625 789 626
rect 729 595 789 625
rect 833 705 887 721
rect 833 671 843 705
rect 877 671 887 705
rect 833 637 887 671
rect 833 603 843 637
rect 877 603 887 637
rect 833 561 887 603
rect 921 705 987 739
rect 1109 739 1125 755
rect 1159 739 1175 773
rect 921 671 937 705
rect 971 671 987 705
rect 921 660 987 671
rect 921 603 937 660
rect 971 603 987 660
rect 921 595 987 603
rect 1021 705 1075 721
rect 1021 671 1031 705
rect 1065 671 1075 705
rect 1021 637 1075 671
rect 1021 603 1031 637
rect 1065 603 1075 637
rect 1021 561 1075 603
rect 1109 705 1175 739
rect 1109 671 1125 705
rect 1159 671 1175 705
rect 1109 660 1175 671
rect 1109 603 1125 660
rect 1159 603 1175 660
rect 1109 595 1175 603
rect 1209 773 1275 789
rect 1209 739 1225 773
rect 1259 739 1275 773
rect 1209 705 1275 739
rect 1209 671 1225 705
rect 1259 671 1275 705
rect 1209 637 1275 671
rect 1209 603 1225 637
rect 1259 603 1275 637
rect 1209 561 1275 603
rect 1309 773 1755 789
rect 1309 739 1325 773
rect 1359 755 1513 773
rect 1359 739 1375 755
rect 1309 705 1375 739
rect 1497 739 1513 755
rect 1547 765 1755 773
rect 1547 755 1711 765
rect 1547 739 1563 755
rect 1309 671 1325 705
rect 1359 671 1375 705
rect 1309 660 1375 671
rect 1309 603 1325 660
rect 1359 603 1375 660
rect 1309 595 1375 603
rect 1409 705 1463 721
rect 1409 671 1419 705
rect 1453 671 1463 705
rect 1409 637 1463 671
rect 1409 603 1419 637
rect 1453 603 1463 637
rect 1409 561 1463 603
rect 1497 705 1563 739
rect 1695 731 1711 755
rect 1745 731 1755 765
rect 1497 671 1513 705
rect 1547 671 1563 705
rect 1497 660 1563 671
rect 1497 603 1513 660
rect 1547 603 1563 660
rect 1497 595 1563 603
rect 1597 705 1651 721
rect 1597 671 1607 705
rect 1641 671 1651 705
rect 1597 637 1651 671
rect 1597 603 1607 637
rect 1641 603 1651 637
rect 1597 561 1651 603
rect 1695 660 1755 731
rect 1695 626 1709 660
rect 1743 659 1755 660
rect 1695 625 1711 626
rect 1745 625 1755 659
rect 1695 595 1755 625
rect 1789 765 1855 815
rect 1789 697 1805 765
rect 1839 697 1855 765
rect 1789 659 1855 697
rect 1789 625 1805 659
rect 1839 625 1855 659
rect 729 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1755 561
rect 629 429 645 463
rect 679 429 695 463
rect 629 391 695 429
rect 629 323 645 391
rect 679 323 695 391
rect 629 273 695 323
rect 729 463 789 493
rect 729 429 739 463
rect 773 462 789 463
rect 729 428 741 429
rect 775 428 789 462
rect 729 357 789 428
rect 833 485 887 527
rect 833 451 843 485
rect 877 451 887 485
rect 833 417 887 451
rect 833 383 843 417
rect 877 383 887 417
rect 833 367 887 383
rect 921 485 987 493
rect 921 428 937 485
rect 971 428 987 485
rect 921 417 987 428
rect 921 383 937 417
rect 971 383 987 417
rect 729 323 739 357
rect 773 333 789 357
rect 921 349 987 383
rect 1021 485 1075 527
rect 1021 451 1031 485
rect 1065 451 1075 485
rect 1021 417 1075 451
rect 1021 383 1031 417
rect 1065 383 1075 417
rect 1021 367 1075 383
rect 1109 485 1175 493
rect 1109 428 1125 485
rect 1159 428 1175 485
rect 1109 417 1175 428
rect 1109 383 1125 417
rect 1159 383 1175 417
rect 921 333 937 349
rect 773 323 937 333
rect 729 315 937 323
rect 971 333 987 349
rect 1109 349 1175 383
rect 1109 333 1125 349
rect 971 315 1125 333
rect 1159 315 1175 349
rect 729 299 1175 315
rect 1209 485 1275 527
rect 1209 451 1225 485
rect 1259 451 1275 485
rect 1209 417 1275 451
rect 1209 383 1225 417
rect 1259 383 1275 417
rect 1209 349 1275 383
rect 1209 315 1225 349
rect 1259 315 1275 349
rect 1209 299 1275 315
rect 1309 485 1375 493
rect 1309 428 1325 485
rect 1359 428 1375 485
rect 1309 417 1375 428
rect 1309 383 1325 417
rect 1359 383 1375 417
rect 1309 349 1375 383
rect 1409 485 1463 527
rect 1409 451 1419 485
rect 1453 451 1463 485
rect 1409 417 1463 451
rect 1409 383 1419 417
rect 1453 383 1463 417
rect 1409 367 1463 383
rect 1497 485 1563 493
rect 1497 428 1513 485
rect 1547 428 1563 485
rect 1497 417 1563 428
rect 1497 383 1513 417
rect 1547 383 1563 417
rect 1309 315 1325 349
rect 1359 333 1375 349
rect 1497 349 1563 383
rect 1597 485 1651 527
rect 1597 451 1607 485
rect 1641 451 1651 485
rect 1597 417 1651 451
rect 1597 383 1607 417
rect 1641 383 1651 417
rect 1597 367 1651 383
rect 1695 463 1755 493
rect 1695 462 1711 463
rect 1695 428 1709 462
rect 1745 429 1755 463
rect 1743 428 1755 429
rect 1497 333 1513 349
rect 1359 315 1513 333
rect 1547 333 1563 349
rect 1695 357 1755 428
rect 1695 333 1711 357
rect 1547 323 1711 333
rect 1745 323 1755 357
rect 1547 315 1755 323
rect 1309 299 1755 315
rect 1789 463 1855 625
rect 1889 765 1943 781
rect 1889 731 1899 765
rect 1933 731 1943 765
rect 1889 660 1943 731
rect 1889 625 1899 660
rect 1933 625 1943 660
rect 1889 595 1943 625
rect 1977 765 2043 815
rect 2077 859 2314 875
rect 2077 825 2086 859
rect 2120 825 2154 859
rect 2188 825 2314 859
rect 2077 809 2314 825
rect 2348 873 2467 889
rect 2348 839 2351 873
rect 2385 839 2419 873
rect 2453 839 2467 873
rect 2348 823 2467 839
rect 2501 873 2620 889
rect 2501 839 2515 873
rect 2549 839 2583 873
rect 2617 839 2620 873
rect 2501 823 2620 839
rect 2654 875 2688 923
rect 2965 875 3031 935
rect 3233 987 3287 1003
rect 3065 934 3099 953
rect 3133 935 3149 969
rect 3183 935 3199 969
rect 3133 911 3199 935
rect 3267 953 3287 987
rect 3321 1029 3371 1071
rect 3321 995 3337 1029
rect 3321 979 3371 995
rect 3405 1029 3471 1037
rect 3405 995 3421 1029
rect 3455 995 3471 1029
rect 3233 945 3287 953
rect 3405 961 3471 995
rect 3505 1029 3559 1071
rect 3505 995 3515 1029
rect 3549 995 3559 1029
rect 3505 979 3559 995
rect 3593 1029 3659 1037
rect 3593 995 3609 1029
rect 3643 995 3659 1029
rect 3405 945 3421 961
rect 3233 927 3421 945
rect 3455 945 3471 961
rect 3593 961 3659 995
rect 3593 945 3609 961
rect 3455 927 3609 945
rect 3643 927 3659 961
rect 3233 911 3659 927
rect 3693 1029 3759 1071
rect 3693 995 3709 1029
rect 3743 995 3759 1029
rect 3693 961 3759 995
rect 3693 927 3709 961
rect 3743 927 3759 961
rect 3693 911 3759 927
rect 3793 1029 3859 1037
rect 3793 995 3809 1029
rect 3843 995 3859 1029
rect 3793 961 3859 995
rect 3893 1029 3947 1071
rect 3893 995 3903 1029
rect 3937 995 3947 1029
rect 3893 979 3947 995
rect 3981 1029 4047 1037
rect 3981 995 3997 1029
rect 4031 995 4047 1029
rect 3793 927 3809 961
rect 3843 945 3859 961
rect 3981 961 4047 995
rect 4081 1029 4131 1071
rect 4115 995 4131 1029
rect 4081 979 4131 995
rect 4165 1003 4571 1037
rect 4165 987 4219 1003
rect 3981 945 3997 961
rect 3843 927 3997 945
rect 4031 945 4047 961
rect 4165 953 4185 987
rect 4353 987 4387 1003
rect 4165 945 4219 953
rect 4031 927 4219 945
rect 3793 911 4219 927
rect 4253 935 4269 969
rect 4303 935 4319 969
rect 4253 911 4319 935
rect 4521 987 4571 1003
rect 4353 934 4387 953
rect 4421 935 4437 969
rect 4471 935 4487 969
rect 3133 875 3179 911
rect 2654 859 2891 875
rect 2654 825 2780 859
rect 2814 825 2848 859
rect 2882 825 2891 859
rect 1977 697 1993 765
rect 2027 697 2043 765
rect 1977 659 2043 697
rect 1977 625 1993 659
rect 2027 625 2043 659
rect 1789 429 1805 463
rect 1839 429 1855 463
rect 1789 391 1855 429
rect 1789 323 1805 391
rect 1839 323 1855 391
rect 441 213 695 273
rect 1789 273 1855 323
rect 1889 463 1943 493
rect 1889 428 1899 463
rect 1933 428 1943 463
rect 1889 357 1943 428
rect 1889 323 1899 357
rect 1933 323 1943 357
rect 1889 307 1943 323
rect 1977 463 2043 625
rect 2077 759 2137 775
rect 2280 767 2314 809
rect 2654 809 2891 825
rect 2925 815 3179 875
rect 3415 873 3693 877
rect 3415 839 3431 873
rect 3465 839 3499 873
rect 3533 839 3567 873
rect 3601 839 3635 873
rect 3669 839 3693 873
rect 3415 823 3693 839
rect 3759 873 4037 877
rect 3759 839 3783 873
rect 3817 839 3851 873
rect 3885 839 3919 873
rect 3953 839 3987 873
rect 4021 839 4037 873
rect 3759 823 4037 839
rect 4273 875 4319 911
rect 4421 875 4487 935
rect 4555 953 4571 987
rect 4672 1016 4730 1071
rect 4672 982 4696 1016
rect 4672 966 4730 982
rect 4764 1016 4814 1032
rect 4764 982 4780 1016
rect 4521 934 4571 953
rect 4764 923 4814 982
rect 4856 1016 4914 1071
rect 4856 982 4864 1016
rect 4898 982 4914 1016
rect 4856 966 4914 982
rect 4764 875 4798 923
rect 2654 767 2688 809
rect 2077 725 2087 759
rect 2121 725 2137 759
rect 2077 660 2137 725
rect 2077 659 2089 660
rect 2077 625 2087 659
rect 2123 626 2137 660
rect 2121 625 2137 626
rect 2077 595 2137 625
rect 2186 751 2241 767
rect 2186 717 2202 751
rect 2236 717 2241 751
rect 2186 645 2241 717
rect 2186 611 2202 645
rect 2236 611 2241 645
rect 2186 561 2241 611
rect 2280 751 2346 767
rect 2280 717 2296 751
rect 2330 717 2346 751
rect 2280 645 2346 717
rect 2280 611 2296 645
rect 2330 611 2346 645
rect 2280 595 2346 611
rect 2380 751 2440 767
rect 2380 717 2390 751
rect 2424 717 2440 751
rect 2380 645 2440 717
rect 2380 611 2390 645
rect 2424 611 2440 645
rect 2380 561 2440 611
rect 2528 751 2588 767
rect 2528 717 2544 751
rect 2578 717 2588 751
rect 2528 645 2588 717
rect 2528 611 2544 645
rect 2578 611 2588 645
rect 2528 561 2588 611
rect 2622 751 2688 767
rect 2622 717 2638 751
rect 2672 717 2688 751
rect 2622 645 2688 717
rect 2622 611 2638 645
rect 2672 611 2688 645
rect 2622 595 2688 611
rect 2727 751 2782 767
rect 2727 717 2732 751
rect 2766 717 2782 751
rect 2727 645 2782 717
rect 2727 611 2732 645
rect 2766 611 2782 645
rect 2727 561 2782 611
rect 2831 759 2891 775
rect 2831 725 2847 759
rect 2881 725 2891 759
rect 2831 660 2891 725
rect 2831 626 2845 660
rect 2879 659 2891 660
rect 2831 625 2847 626
rect 2881 625 2891 659
rect 2831 595 2891 625
rect 2925 765 2991 815
rect 2925 697 2941 765
rect 2975 697 2991 765
rect 2925 659 2991 697
rect 2925 625 2941 659
rect 2975 625 2991 659
rect 2077 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2891 561
rect 1977 429 1993 463
rect 2027 429 2043 463
rect 1977 391 2043 429
rect 1977 323 1993 391
rect 2027 323 2043 391
rect 1977 273 2043 323
rect 2077 463 2137 493
rect 2077 429 2087 463
rect 2121 462 2137 463
rect 2077 428 2089 429
rect 2123 428 2137 462
rect 2077 363 2137 428
rect 2077 329 2087 363
rect 2121 329 2137 363
rect 2077 313 2137 329
rect 2186 477 2241 527
rect 2186 443 2202 477
rect 2236 443 2241 477
rect 2186 371 2241 443
rect 2186 337 2202 371
rect 2236 337 2241 371
rect 2186 321 2241 337
rect 2280 477 2346 493
rect 2280 443 2296 477
rect 2330 443 2346 477
rect 2280 371 2346 443
rect 2280 337 2296 371
rect 2330 337 2346 371
rect 2280 321 2346 337
rect 2380 477 2440 527
rect 2380 443 2390 477
rect 2424 443 2440 477
rect 2380 371 2440 443
rect 2380 337 2390 371
rect 2424 337 2440 371
rect 2380 321 2440 337
rect 2528 477 2588 527
rect 2528 443 2544 477
rect 2578 443 2588 477
rect 2528 371 2588 443
rect 2528 337 2544 371
rect 2578 337 2588 371
rect 2528 321 2588 337
rect 2622 477 2688 493
rect 2622 443 2638 477
rect 2672 443 2688 477
rect 2622 371 2688 443
rect 2622 337 2638 371
rect 2672 337 2688 371
rect 2622 321 2688 337
rect 2727 477 2782 527
rect 2727 443 2732 477
rect 2766 443 2782 477
rect 2727 371 2782 443
rect 2727 337 2732 371
rect 2766 337 2782 371
rect 2727 321 2782 337
rect 2831 463 2891 493
rect 2831 462 2847 463
rect 2831 428 2845 462
rect 2881 429 2891 463
rect 2879 428 2891 429
rect 2831 363 2891 428
rect 2831 329 2847 363
rect 2881 329 2891 363
rect 2280 279 2314 321
rect 170 165 204 213
rect 54 106 112 122
rect 54 72 70 106
rect 104 72 112 106
rect 54 17 112 72
rect 154 106 204 165
rect 397 135 447 154
rect 188 72 204 106
rect 154 56 204 72
rect 238 106 296 122
rect 272 72 296 106
rect 238 17 296 72
rect 397 101 413 135
rect 481 153 547 213
rect 649 177 695 213
rect 931 249 1209 265
rect 931 215 947 249
rect 981 215 1015 249
rect 1049 215 1083 249
rect 1117 215 1151 249
rect 1185 215 1209 249
rect 931 211 1209 215
rect 1275 249 1553 265
rect 1275 215 1299 249
rect 1333 215 1367 249
rect 1401 215 1435 249
rect 1469 215 1503 249
rect 1537 215 1553 249
rect 1275 211 1553 215
rect 1789 213 2043 273
rect 2077 263 2314 279
rect 2654 279 2688 321
rect 2831 313 2891 329
rect 2925 463 2991 625
rect 3025 765 3079 781
rect 3025 731 3035 765
rect 3069 731 3079 765
rect 3025 660 3079 731
rect 3025 625 3035 660
rect 3069 625 3079 660
rect 3025 595 3079 625
rect 3113 765 3179 815
rect 4273 815 4527 875
rect 3113 697 3129 765
rect 3163 697 3179 765
rect 3113 659 3179 697
rect 3113 625 3129 659
rect 3163 625 3179 659
rect 2925 429 2941 463
rect 2975 429 2991 463
rect 2925 391 2991 429
rect 2925 323 2941 391
rect 2975 323 2991 391
rect 2077 229 2086 263
rect 2120 229 2154 263
rect 2188 229 2314 263
rect 2077 213 2314 229
rect 1789 177 1835 213
rect 481 119 497 153
rect 531 119 547 153
rect 581 135 615 154
rect 397 85 447 101
rect 649 153 715 177
rect 649 119 665 153
rect 699 119 715 153
rect 749 161 1175 177
rect 749 143 937 161
rect 749 135 803 143
rect 581 85 615 101
rect 783 101 803 135
rect 921 127 937 143
rect 971 143 1125 161
rect 971 127 987 143
rect 749 85 803 101
rect 397 51 803 85
rect 837 93 887 109
rect 837 59 853 93
rect 837 17 887 59
rect 921 93 987 127
rect 1109 127 1125 143
rect 1159 127 1175 161
rect 921 59 937 93
rect 971 59 987 93
rect 921 51 987 59
rect 1021 93 1075 109
rect 1021 59 1031 93
rect 1065 59 1075 93
rect 1021 17 1075 59
rect 1109 93 1175 127
rect 1109 59 1125 93
rect 1159 59 1175 93
rect 1109 51 1175 59
rect 1209 161 1275 177
rect 1209 127 1225 161
rect 1259 127 1275 161
rect 1209 93 1275 127
rect 1209 59 1225 93
rect 1259 59 1275 93
rect 1209 17 1275 59
rect 1309 161 1735 177
rect 1309 127 1325 161
rect 1359 143 1513 161
rect 1359 127 1375 143
rect 1309 93 1375 127
rect 1497 127 1513 143
rect 1547 143 1735 161
rect 1547 127 1563 143
rect 1309 59 1325 93
rect 1359 59 1375 93
rect 1309 51 1375 59
rect 1409 93 1463 109
rect 1409 59 1419 93
rect 1453 59 1463 93
rect 1409 17 1463 59
rect 1497 93 1563 127
rect 1681 135 1735 143
rect 1497 59 1513 93
rect 1547 59 1563 93
rect 1497 51 1563 59
rect 1597 93 1647 109
rect 1631 59 1647 93
rect 1597 17 1647 59
rect 1681 101 1701 135
rect 1769 153 1835 177
rect 1769 119 1785 153
rect 1819 119 1835 153
rect 1869 135 1903 154
rect 1681 85 1735 101
rect 1937 153 2003 213
rect 2280 165 2314 213
rect 2348 249 2467 265
rect 2348 215 2351 249
rect 2385 215 2419 249
rect 2453 215 2467 249
rect 2348 199 2467 215
rect 2501 249 2620 265
rect 2501 215 2515 249
rect 2549 215 2583 249
rect 2617 215 2620 249
rect 2501 199 2620 215
rect 2654 263 2891 279
rect 2654 229 2780 263
rect 2814 229 2848 263
rect 2882 229 2891 263
rect 2654 213 2891 229
rect 2925 273 2991 323
rect 3025 463 3079 493
rect 3025 428 3035 463
rect 3069 428 3079 463
rect 3025 357 3079 428
rect 3025 323 3035 357
rect 3069 323 3079 357
rect 3025 307 3079 323
rect 3113 463 3179 625
rect 3213 773 3659 789
rect 3213 765 3421 773
rect 3213 731 3223 765
rect 3257 755 3421 765
rect 3257 731 3273 755
rect 3213 660 3273 731
rect 3405 739 3421 755
rect 3455 755 3609 773
rect 3455 739 3471 755
rect 3213 659 3225 660
rect 3213 625 3223 659
rect 3259 626 3273 660
rect 3257 625 3273 626
rect 3213 595 3273 625
rect 3317 705 3371 721
rect 3317 671 3327 705
rect 3361 671 3371 705
rect 3317 637 3371 671
rect 3317 603 3327 637
rect 3361 603 3371 637
rect 3317 561 3371 603
rect 3405 705 3471 739
rect 3593 739 3609 755
rect 3643 739 3659 773
rect 3405 671 3421 705
rect 3455 671 3471 705
rect 3405 660 3471 671
rect 3405 603 3421 660
rect 3455 603 3471 660
rect 3405 595 3471 603
rect 3505 705 3559 721
rect 3505 671 3515 705
rect 3549 671 3559 705
rect 3505 637 3559 671
rect 3505 603 3515 637
rect 3549 603 3559 637
rect 3505 561 3559 603
rect 3593 705 3659 739
rect 3593 671 3609 705
rect 3643 671 3659 705
rect 3593 660 3659 671
rect 3593 603 3609 660
rect 3643 603 3659 660
rect 3593 595 3659 603
rect 3693 773 3759 789
rect 3693 739 3709 773
rect 3743 739 3759 773
rect 3693 705 3759 739
rect 3693 671 3709 705
rect 3743 671 3759 705
rect 3693 637 3759 671
rect 3693 603 3709 637
rect 3743 603 3759 637
rect 3693 561 3759 603
rect 3793 773 4239 789
rect 3793 739 3809 773
rect 3843 755 3997 773
rect 3843 739 3859 755
rect 3793 705 3859 739
rect 3981 739 3997 755
rect 4031 765 4239 773
rect 4031 755 4195 765
rect 4031 739 4047 755
rect 3793 671 3809 705
rect 3843 671 3859 705
rect 3793 660 3859 671
rect 3793 603 3809 660
rect 3843 603 3859 660
rect 3793 595 3859 603
rect 3893 705 3947 721
rect 3893 671 3903 705
rect 3937 671 3947 705
rect 3893 637 3947 671
rect 3893 603 3903 637
rect 3937 603 3947 637
rect 3893 561 3947 603
rect 3981 705 4047 739
rect 4179 731 4195 755
rect 4229 731 4239 765
rect 3981 671 3997 705
rect 4031 671 4047 705
rect 3981 660 4047 671
rect 3981 603 3997 660
rect 4031 603 4047 660
rect 3981 595 4047 603
rect 4081 705 4135 721
rect 4081 671 4091 705
rect 4125 671 4135 705
rect 4081 637 4135 671
rect 4081 603 4091 637
rect 4125 603 4135 637
rect 4081 561 4135 603
rect 4179 660 4239 731
rect 4179 626 4193 660
rect 4227 659 4239 660
rect 4179 625 4195 626
rect 4229 625 4239 659
rect 4179 595 4239 625
rect 4273 765 4339 815
rect 4273 697 4289 765
rect 4323 697 4339 765
rect 4273 659 4339 697
rect 4273 625 4289 659
rect 4323 625 4339 659
rect 3213 527 3249 561
rect 3283 527 3341 561
rect 3375 527 3433 561
rect 3467 527 3525 561
rect 3559 527 3617 561
rect 3651 527 3709 561
rect 3743 527 3801 561
rect 3835 527 3893 561
rect 3927 527 3985 561
rect 4019 527 4077 561
rect 4111 527 4169 561
rect 4203 527 4239 561
rect 3113 429 3129 463
rect 3163 429 3179 463
rect 3113 391 3179 429
rect 3113 323 3129 391
rect 3163 323 3179 391
rect 3113 273 3179 323
rect 3213 463 3273 493
rect 3213 429 3223 463
rect 3257 462 3273 463
rect 3213 428 3225 429
rect 3259 428 3273 462
rect 3213 357 3273 428
rect 3317 485 3371 527
rect 3317 451 3327 485
rect 3361 451 3371 485
rect 3317 417 3371 451
rect 3317 383 3327 417
rect 3361 383 3371 417
rect 3317 367 3371 383
rect 3405 485 3471 493
rect 3405 428 3421 485
rect 3455 428 3471 485
rect 3405 417 3471 428
rect 3405 383 3421 417
rect 3455 383 3471 417
rect 3213 323 3223 357
rect 3257 333 3273 357
rect 3405 349 3471 383
rect 3505 485 3559 527
rect 3505 451 3515 485
rect 3549 451 3559 485
rect 3505 417 3559 451
rect 3505 383 3515 417
rect 3549 383 3559 417
rect 3505 367 3559 383
rect 3593 485 3659 493
rect 3593 428 3609 485
rect 3643 428 3659 485
rect 3593 417 3659 428
rect 3593 383 3609 417
rect 3643 383 3659 417
rect 3405 333 3421 349
rect 3257 323 3421 333
rect 3213 315 3421 323
rect 3455 333 3471 349
rect 3593 349 3659 383
rect 3593 333 3609 349
rect 3455 315 3609 333
rect 3643 315 3659 349
rect 3213 299 3659 315
rect 3693 485 3759 527
rect 3693 451 3709 485
rect 3743 451 3759 485
rect 3693 417 3759 451
rect 3693 383 3709 417
rect 3743 383 3759 417
rect 3693 349 3759 383
rect 3693 315 3709 349
rect 3743 315 3759 349
rect 3693 299 3759 315
rect 3793 485 3859 493
rect 3793 428 3809 485
rect 3843 428 3859 485
rect 3793 417 3859 428
rect 3793 383 3809 417
rect 3843 383 3859 417
rect 3793 349 3859 383
rect 3893 485 3947 527
rect 3893 451 3903 485
rect 3937 451 3947 485
rect 3893 417 3947 451
rect 3893 383 3903 417
rect 3937 383 3947 417
rect 3893 367 3947 383
rect 3981 485 4047 493
rect 3981 428 3997 485
rect 4031 428 4047 485
rect 3981 417 4047 428
rect 3981 383 3997 417
rect 4031 383 4047 417
rect 3793 315 3809 349
rect 3843 333 3859 349
rect 3981 349 4047 383
rect 4081 485 4135 527
rect 4081 451 4091 485
rect 4125 451 4135 485
rect 4081 417 4135 451
rect 4081 383 4091 417
rect 4125 383 4135 417
rect 4081 367 4135 383
rect 4179 463 4239 493
rect 4179 462 4195 463
rect 4179 428 4193 462
rect 4229 429 4239 463
rect 4227 428 4239 429
rect 3981 333 3997 349
rect 3843 315 3997 333
rect 4031 333 4047 349
rect 4179 357 4239 428
rect 4179 333 4195 357
rect 4031 323 4195 333
rect 4229 323 4239 357
rect 4031 315 4239 323
rect 3793 299 4239 315
rect 4273 463 4339 625
rect 4373 765 4427 781
rect 4373 731 4383 765
rect 4417 731 4427 765
rect 4373 660 4427 731
rect 4373 625 4383 660
rect 4417 625 4427 660
rect 4373 595 4427 625
rect 4461 765 4527 815
rect 4561 859 4798 875
rect 4561 825 4570 859
rect 4604 825 4638 859
rect 4672 825 4798 859
rect 4561 809 4798 825
rect 4832 873 4951 889
rect 4832 839 4835 873
rect 4869 839 4903 873
rect 4937 839 4951 873
rect 4832 823 4951 839
rect 4461 697 4477 765
rect 4511 697 4527 765
rect 4461 659 4527 697
rect 4461 625 4477 659
rect 4511 625 4527 659
rect 4273 429 4289 463
rect 4323 429 4339 463
rect 4273 391 4339 429
rect 4273 323 4289 391
rect 4323 323 4339 391
rect 2925 213 3179 273
rect 4273 273 4339 323
rect 4373 463 4427 493
rect 4373 428 4383 463
rect 4417 428 4427 463
rect 4373 357 4427 428
rect 4373 323 4383 357
rect 4417 323 4427 357
rect 4373 307 4427 323
rect 4461 463 4527 625
rect 4561 759 4621 775
rect 4764 767 4798 809
rect 4561 725 4571 759
rect 4605 725 4621 759
rect 4561 660 4621 725
rect 4561 659 4573 660
rect 4561 625 4571 659
rect 4607 626 4621 660
rect 4605 625 4621 626
rect 4561 595 4621 625
rect 4670 751 4725 767
rect 4670 717 4686 751
rect 4720 717 4725 751
rect 4670 645 4725 717
rect 4670 611 4686 645
rect 4720 611 4725 645
rect 4670 561 4725 611
rect 4764 751 4830 767
rect 4764 717 4780 751
rect 4814 717 4830 751
rect 4764 645 4830 717
rect 4764 611 4780 645
rect 4814 611 4830 645
rect 4764 595 4830 611
rect 4864 751 4924 767
rect 4864 717 4874 751
rect 4908 717 4924 751
rect 4864 645 4924 717
rect 4864 611 4874 645
rect 4908 611 4924 645
rect 4864 561 4924 611
rect 4561 527 4629 561
rect 4663 527 4721 561
rect 4755 527 4813 561
rect 4847 527 4905 561
rect 4939 527 4968 561
rect 4461 429 4477 463
rect 4511 429 4527 463
rect 4461 391 4527 429
rect 4461 323 4477 391
rect 4511 323 4527 391
rect 4461 273 4527 323
rect 4561 463 4621 493
rect 4561 429 4571 463
rect 4605 462 4621 463
rect 4561 428 4573 429
rect 4607 428 4621 462
rect 4561 363 4621 428
rect 4561 329 4571 363
rect 4605 329 4621 363
rect 4561 313 4621 329
rect 4670 477 4725 527
rect 4670 443 4686 477
rect 4720 443 4725 477
rect 4670 371 4725 443
rect 4670 337 4686 371
rect 4720 337 4725 371
rect 4670 321 4725 337
rect 4764 477 4830 493
rect 4764 443 4780 477
rect 4814 443 4830 477
rect 4764 371 4830 443
rect 4764 337 4780 371
rect 4814 337 4830 371
rect 4764 321 4830 337
rect 4864 477 4924 527
rect 4864 443 4874 477
rect 4908 443 4924 477
rect 4864 371 4924 443
rect 4864 337 4874 371
rect 4908 337 4924 371
rect 4864 321 4924 337
rect 4764 279 4798 321
rect 2654 165 2688 213
rect 1937 119 1953 153
rect 1987 119 2003 153
rect 2037 135 2087 154
rect 1869 85 1903 101
rect 2071 101 2087 135
rect 2037 85 2087 101
rect 1681 51 2087 85
rect 2188 106 2246 122
rect 2188 72 2212 106
rect 2188 17 2246 72
rect 2280 106 2330 165
rect 2280 72 2296 106
rect 2280 56 2330 72
rect 2372 106 2430 122
rect 2372 72 2380 106
rect 2414 72 2430 106
rect 2372 17 2430 72
rect 2538 106 2596 122
rect 2538 72 2554 106
rect 2588 72 2596 106
rect 2538 17 2596 72
rect 2638 106 2688 165
rect 2881 135 2931 154
rect 2672 72 2688 106
rect 2638 56 2688 72
rect 2722 106 2780 122
rect 2756 72 2780 106
rect 2722 17 2780 72
rect 2881 101 2897 135
rect 2965 153 3031 213
rect 3133 177 3179 213
rect 3415 249 3693 265
rect 3415 215 3431 249
rect 3465 215 3499 249
rect 3533 215 3567 249
rect 3601 215 3635 249
rect 3669 215 3693 249
rect 3415 211 3693 215
rect 3759 249 4037 265
rect 3759 215 3783 249
rect 3817 215 3851 249
rect 3885 215 3919 249
rect 3953 215 3987 249
rect 4021 215 4037 249
rect 3759 211 4037 215
rect 4273 213 4527 273
rect 4561 263 4798 279
rect 4561 229 4570 263
rect 4604 229 4638 263
rect 4672 229 4798 263
rect 4561 213 4798 229
rect 4273 177 4319 213
rect 2965 119 2981 153
rect 3015 119 3031 153
rect 3065 135 3099 154
rect 2881 85 2931 101
rect 3133 153 3199 177
rect 3133 119 3149 153
rect 3183 119 3199 153
rect 3233 161 3659 177
rect 3233 143 3421 161
rect 3233 135 3287 143
rect 3065 85 3099 101
rect 3267 101 3287 135
rect 3405 127 3421 143
rect 3455 143 3609 161
rect 3455 127 3471 143
rect 3233 85 3287 101
rect 2881 51 3287 85
rect 3321 93 3371 109
rect 3321 59 3337 93
rect 3321 17 3371 59
rect 3405 93 3471 127
rect 3593 127 3609 143
rect 3643 127 3659 161
rect 3405 59 3421 93
rect 3455 59 3471 93
rect 3405 51 3471 59
rect 3505 93 3559 109
rect 3505 59 3515 93
rect 3549 59 3559 93
rect 3505 17 3559 59
rect 3593 93 3659 127
rect 3593 59 3609 93
rect 3643 59 3659 93
rect 3593 51 3659 59
rect 3693 161 3759 177
rect 3693 127 3709 161
rect 3743 127 3759 161
rect 3693 93 3759 127
rect 3693 59 3709 93
rect 3743 59 3759 93
rect 3693 17 3759 59
rect 3793 161 4219 177
rect 3793 127 3809 161
rect 3843 143 3997 161
rect 3843 127 3859 143
rect 3793 93 3859 127
rect 3981 127 3997 143
rect 4031 143 4219 161
rect 4031 127 4047 143
rect 3793 59 3809 93
rect 3843 59 3859 93
rect 3793 51 3859 59
rect 3893 93 3947 109
rect 3893 59 3903 93
rect 3937 59 3947 93
rect 3893 17 3947 59
rect 3981 93 4047 127
rect 4165 135 4219 143
rect 3981 59 3997 93
rect 4031 59 4047 93
rect 3981 51 4047 59
rect 4081 93 4131 109
rect 4115 59 4131 93
rect 4081 17 4131 59
rect 4165 101 4185 135
rect 4253 153 4319 177
rect 4253 119 4269 153
rect 4303 119 4319 153
rect 4353 135 4387 154
rect 4165 85 4219 101
rect 4421 153 4487 213
rect 4764 165 4798 213
rect 4832 249 4951 265
rect 4832 215 4835 249
rect 4869 215 4903 249
rect 4937 215 4951 249
rect 4832 199 4951 215
rect 4421 119 4437 153
rect 4471 119 4487 153
rect 4521 135 4571 154
rect 4353 85 4387 101
rect 4555 101 4571 135
rect 4521 85 4571 101
rect 4165 51 4571 85
rect 4672 106 4730 122
rect 4672 72 4696 106
rect 4672 17 4730 72
rect 4764 106 4814 165
rect 4764 72 4780 106
rect 4764 56 4814 72
rect 4856 106 4914 122
rect 4856 72 4864 106
rect 4898 72 4914 106
rect 4856 17 4914 72
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3341 17
rect 3375 -17 3433 17
rect 3467 -17 3525 17
rect 3559 -17 3617 17
rect 3651 -17 3709 17
rect 3743 -17 3801 17
rect 3835 -17 3893 17
rect 3927 -17 3985 17
rect 4019 -17 4077 17
rect 4111 -17 4169 17
rect 4203 -17 4261 17
rect 4295 -17 4353 17
rect 4387 -17 4445 17
rect 4479 -17 4537 17
rect 4571 -17 4629 17
rect 4663 -17 4721 17
rect 4755 -17 4813 17
rect 4847 -17 4905 17
rect 4939 -17 4968 17
<< viali >>
rect 29 1071 63 1105
rect 121 1071 155 1105
rect 213 1071 247 1105
rect 305 1071 339 1105
rect 397 1071 431 1105
rect 489 1071 523 1105
rect 581 1071 615 1105
rect 673 1071 707 1105
rect 765 1071 799 1105
rect 857 1071 891 1105
rect 949 1071 983 1105
rect 1041 1071 1075 1105
rect 1133 1071 1167 1105
rect 1225 1071 1259 1105
rect 1317 1071 1351 1105
rect 1409 1071 1443 1105
rect 1501 1071 1535 1105
rect 1593 1071 1627 1105
rect 1685 1071 1719 1105
rect 1777 1071 1811 1105
rect 1869 1071 1903 1105
rect 1961 1071 1995 1105
rect 2053 1071 2087 1105
rect 2145 1071 2179 1105
rect 2237 1071 2271 1105
rect 2329 1071 2363 1105
rect 2421 1071 2455 1105
rect 2513 1071 2547 1105
rect 2605 1071 2639 1105
rect 2697 1071 2731 1105
rect 2789 1071 2823 1105
rect 2881 1071 2915 1105
rect 2973 1071 3007 1105
rect 3065 1071 3099 1105
rect 3157 1071 3191 1105
rect 3249 1071 3283 1105
rect 3341 1071 3375 1105
rect 3433 1071 3467 1105
rect 3525 1071 3559 1105
rect 3617 1071 3651 1105
rect 3709 1071 3743 1105
rect 3801 1071 3835 1105
rect 3893 1071 3927 1105
rect 3985 1071 4019 1105
rect 4077 1071 4111 1105
rect 4169 1071 4203 1105
rect 4261 1071 4295 1105
rect 4353 1071 4387 1105
rect 4445 1071 4479 1105
rect 4537 1071 4571 1105
rect 4629 1071 4663 1105
rect 4721 1071 4755 1105
rect 4813 1071 4847 1105
rect 4905 1071 4939 1105
rect 361 659 395 660
rect 361 626 363 659
rect 363 626 395 659
rect 457 697 491 731
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 361 429 363 462
rect 363 429 395 462
rect 361 428 395 429
rect 551 659 585 660
rect 551 626 585 659
rect 645 697 679 731
rect 457 357 491 391
rect 551 429 585 462
rect 551 428 585 429
rect 741 659 775 660
rect 741 626 773 659
rect 773 626 775 659
rect 937 637 971 660
rect 937 626 971 637
rect 1125 637 1159 660
rect 1125 626 1159 637
rect 1325 637 1359 660
rect 1325 626 1359 637
rect 1513 637 1547 660
rect 1513 626 1547 637
rect 1709 659 1743 660
rect 1709 626 1711 659
rect 1711 626 1743 659
rect 1805 697 1839 731
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 645 357 679 391
rect 741 429 773 462
rect 773 429 775 462
rect 741 428 775 429
rect 937 451 971 462
rect 937 428 971 451
rect 1125 451 1159 462
rect 1125 428 1159 451
rect 1325 451 1359 462
rect 1325 428 1359 451
rect 1513 451 1547 462
rect 1513 428 1547 451
rect 1709 429 1711 462
rect 1711 429 1743 462
rect 1709 428 1743 429
rect 1899 659 1933 660
rect 1899 626 1933 659
rect 1993 697 2027 731
rect 1805 357 1839 391
rect 1899 429 1933 462
rect 1899 428 1933 429
rect 2089 659 2123 660
rect 2089 626 2121 659
rect 2121 626 2123 659
rect 2845 659 2879 660
rect 2845 626 2847 659
rect 2847 626 2879 659
rect 2941 697 2975 731
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 1993 357 2027 391
rect 2089 429 2121 462
rect 2121 429 2123 462
rect 2089 428 2123 429
rect 2845 429 2847 462
rect 2847 429 2879 462
rect 2845 428 2879 429
rect 3035 659 3069 660
rect 3035 626 3069 659
rect 3129 697 3163 731
rect 2941 357 2975 391
rect 3035 429 3069 462
rect 3035 428 3069 429
rect 3225 659 3259 660
rect 3225 626 3257 659
rect 3257 626 3259 659
rect 3421 637 3455 660
rect 3421 626 3455 637
rect 3609 637 3643 660
rect 3609 626 3643 637
rect 3809 637 3843 660
rect 3809 626 3843 637
rect 3997 637 4031 660
rect 3997 626 4031 637
rect 4193 659 4227 660
rect 4193 626 4195 659
rect 4195 626 4227 659
rect 4289 697 4323 731
rect 3249 527 3283 561
rect 3341 527 3375 561
rect 3433 527 3467 561
rect 3525 527 3559 561
rect 3617 527 3651 561
rect 3709 527 3743 561
rect 3801 527 3835 561
rect 3893 527 3927 561
rect 3985 527 4019 561
rect 4077 527 4111 561
rect 4169 527 4203 561
rect 3129 357 3163 391
rect 3225 429 3257 462
rect 3257 429 3259 462
rect 3225 428 3259 429
rect 3421 451 3455 462
rect 3421 428 3455 451
rect 3609 451 3643 462
rect 3609 428 3643 451
rect 3809 451 3843 462
rect 3809 428 3843 451
rect 3997 451 4031 462
rect 3997 428 4031 451
rect 4193 429 4195 462
rect 4195 429 4227 462
rect 4193 428 4227 429
rect 4383 659 4417 660
rect 4383 626 4417 659
rect 4477 697 4511 731
rect 4289 357 4323 391
rect 4383 429 4417 462
rect 4383 428 4417 429
rect 4573 659 4607 660
rect 4573 626 4605 659
rect 4605 626 4607 659
rect 4629 527 4663 561
rect 4721 527 4755 561
rect 4813 527 4847 561
rect 4905 527 4939 561
rect 4477 357 4511 391
rect 4573 429 4605 462
rect 4605 429 4607 462
rect 4573 428 4607 429
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
rect 2881 -17 2915 17
rect 2973 -17 3007 17
rect 3065 -17 3099 17
rect 3157 -17 3191 17
rect 3249 -17 3283 17
rect 3341 -17 3375 17
rect 3433 -17 3467 17
rect 3525 -17 3559 17
rect 3617 -17 3651 17
rect 3709 -17 3743 17
rect 3801 -17 3835 17
rect 3893 -17 3927 17
rect 3985 -17 4019 17
rect 4077 -17 4111 17
rect 4169 -17 4203 17
rect 4261 -17 4295 17
rect 4353 -17 4387 17
rect 4445 -17 4479 17
rect 4537 -17 4571 17
rect 4629 -17 4663 17
rect 4721 -17 4755 17
rect 4813 -17 4847 17
rect 4905 -17 4939 17
<< metal1 >>
rect 0 1105 4968 1136
rect 0 1071 29 1105
rect 63 1071 121 1105
rect 155 1071 213 1105
rect 247 1071 305 1105
rect 339 1071 397 1105
rect 431 1071 489 1105
rect 523 1071 581 1105
rect 615 1071 673 1105
rect 707 1071 765 1105
rect 799 1071 857 1105
rect 891 1071 949 1105
rect 983 1071 1041 1105
rect 1075 1071 1133 1105
rect 1167 1071 1225 1105
rect 1259 1071 1317 1105
rect 1351 1071 1409 1105
rect 1443 1071 1501 1105
rect 1535 1071 1593 1105
rect 1627 1071 1685 1105
rect 1719 1071 1777 1105
rect 1811 1071 1869 1105
rect 1903 1071 1961 1105
rect 1995 1071 2053 1105
rect 2087 1071 2145 1105
rect 2179 1071 2237 1105
rect 2271 1071 2329 1105
rect 2363 1071 2421 1105
rect 2455 1071 2513 1105
rect 2547 1071 2605 1105
rect 2639 1071 2697 1105
rect 2731 1071 2789 1105
rect 2823 1071 2881 1105
rect 2915 1071 2973 1105
rect 3007 1071 3065 1105
rect 3099 1071 3157 1105
rect 3191 1071 3249 1105
rect 3283 1071 3341 1105
rect 3375 1071 3433 1105
rect 3467 1071 3525 1105
rect 3559 1071 3617 1105
rect 3651 1071 3709 1105
rect 3743 1071 3801 1105
rect 3835 1071 3893 1105
rect 3927 1071 3985 1105
rect 4019 1071 4077 1105
rect 4111 1071 4169 1105
rect 4203 1071 4261 1105
rect 4295 1071 4353 1105
rect 4387 1071 4445 1105
rect 4479 1071 4537 1105
rect 4571 1071 4629 1105
rect 4663 1071 4721 1105
rect 4755 1071 4813 1105
rect 4847 1071 4905 1105
rect 4939 1071 4968 1105
rect 0 1040 4968 1071
rect 445 731 503 737
rect 445 697 457 731
rect 491 728 503 731
rect 633 731 691 737
rect 633 728 645 731
rect 491 700 645 728
rect 491 697 503 700
rect 445 691 503 697
rect 633 697 645 700
rect 679 728 691 731
rect 1793 731 1851 737
rect 1793 728 1805 731
rect 679 700 1805 728
rect 679 697 691 700
rect 633 691 691 697
rect 1793 697 1805 700
rect 1839 728 1851 731
rect 1981 731 2039 737
rect 1981 728 1993 731
rect 1839 700 1993 728
rect 1839 697 1851 700
rect 1793 691 1851 697
rect 1981 697 1993 700
rect 2027 728 2039 731
rect 2929 731 2987 737
rect 2929 728 2941 731
rect 2027 700 2941 728
rect 2027 697 2039 700
rect 1981 691 2039 697
rect 2929 697 2941 700
rect 2975 728 2987 731
rect 3117 731 3175 737
rect 3117 728 3129 731
rect 2975 700 3129 728
rect 2975 697 2987 700
rect 2929 691 2987 697
rect 3117 697 3129 700
rect 3163 728 3175 731
rect 4277 731 4335 737
rect 4277 728 4289 731
rect 3163 700 4289 728
rect 3163 697 3175 700
rect 3117 691 3175 697
rect 4277 697 4289 700
rect 4323 728 4335 731
rect 4465 731 4523 737
rect 4465 728 4477 731
rect 4323 700 4477 728
rect 4323 697 4335 700
rect 4277 691 4335 697
rect 4465 697 4477 700
rect 4511 697 4523 731
rect 4465 691 4523 697
rect 349 660 407 666
rect 349 626 361 660
rect 395 657 407 660
rect 539 660 597 666
rect 539 657 551 660
rect 395 629 551 657
rect 395 626 407 629
rect 349 620 407 626
rect 539 626 551 629
rect 585 657 597 660
rect 729 660 787 666
rect 729 657 741 660
rect 585 629 741 657
rect 585 626 597 629
rect 539 620 597 626
rect 729 626 741 629
rect 775 657 787 660
rect 925 660 983 666
rect 925 657 937 660
rect 775 629 937 657
rect 775 626 787 629
rect 729 620 787 626
rect 925 626 937 629
rect 971 657 983 660
rect 1113 660 1171 666
rect 1113 657 1125 660
rect 971 629 1125 657
rect 971 626 983 629
rect 925 620 983 626
rect 1113 626 1125 629
rect 1159 626 1171 660
rect 1113 620 1171 626
rect 1313 660 1371 666
rect 1313 626 1325 660
rect 1359 657 1371 660
rect 1501 660 1559 666
rect 1501 657 1513 660
rect 1359 629 1513 657
rect 1359 626 1371 629
rect 1313 620 1371 626
rect 1501 626 1513 629
rect 1547 657 1559 660
rect 1697 660 1755 666
rect 1697 657 1709 660
rect 1547 629 1709 657
rect 1547 626 1559 629
rect 1501 620 1559 626
rect 1697 626 1709 629
rect 1743 657 1755 660
rect 1887 660 1945 666
rect 1887 657 1899 660
rect 1743 629 1899 657
rect 1743 626 1755 629
rect 1697 620 1755 626
rect 1887 626 1899 629
rect 1933 657 1945 660
rect 2077 660 2135 666
rect 2077 657 2089 660
rect 1933 629 2089 657
rect 1933 626 1945 629
rect 1887 620 1945 626
rect 2077 626 2089 629
rect 2123 626 2135 660
rect 2077 620 2135 626
rect 2833 660 2891 666
rect 2833 626 2845 660
rect 2879 657 2891 660
rect 3023 660 3081 666
rect 3023 657 3035 660
rect 2879 629 3035 657
rect 2879 626 2891 629
rect 2833 620 2891 626
rect 3023 626 3035 629
rect 3069 657 3081 660
rect 3213 660 3271 666
rect 3213 657 3225 660
rect 3069 629 3225 657
rect 3069 626 3081 629
rect 3023 620 3081 626
rect 3213 626 3225 629
rect 3259 657 3271 660
rect 3409 660 3467 666
rect 3409 657 3421 660
rect 3259 629 3421 657
rect 3259 626 3271 629
rect 3213 620 3271 626
rect 3409 626 3421 629
rect 3455 657 3467 660
rect 3597 660 3655 666
rect 3597 657 3609 660
rect 3455 629 3609 657
rect 3455 626 3467 629
rect 3409 620 3467 626
rect 3597 626 3609 629
rect 3643 626 3655 660
rect 3597 620 3655 626
rect 3797 660 3855 666
rect 3797 626 3809 660
rect 3843 657 3855 660
rect 3985 660 4043 666
rect 3985 657 3997 660
rect 3843 629 3997 657
rect 3843 626 3855 629
rect 3797 620 3855 626
rect 3985 626 3997 629
rect 4031 657 4043 660
rect 4181 660 4239 666
rect 4181 657 4193 660
rect 4031 629 4193 657
rect 4031 626 4043 629
rect 3985 620 4043 626
rect 4181 626 4193 629
rect 4227 657 4239 660
rect 4371 660 4429 666
rect 4371 657 4383 660
rect 4227 629 4383 657
rect 4227 626 4239 629
rect 4181 620 4239 626
rect 4371 626 4383 629
rect 4417 657 4429 660
rect 4561 660 4619 666
rect 4561 657 4573 660
rect 4417 629 4573 657
rect 4417 626 4429 629
rect 4371 620 4429 626
rect 4561 626 4573 629
rect 4607 626 4619 660
rect 4561 620 4619 626
rect 0 561 4968 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 3249 561
rect 3283 527 3341 561
rect 3375 527 3433 561
rect 3467 527 3525 561
rect 3559 527 3617 561
rect 3651 527 3709 561
rect 3743 527 3801 561
rect 3835 527 3893 561
rect 3927 527 3985 561
rect 4019 527 4077 561
rect 4111 527 4169 561
rect 4203 527 4629 561
rect 4663 527 4721 561
rect 4755 527 4813 561
rect 4847 527 4905 561
rect 4939 527 4968 561
rect 0 496 4968 527
rect 349 462 407 468
rect 349 428 361 462
rect 395 459 407 462
rect 539 462 597 468
rect 539 459 551 462
rect 395 431 551 459
rect 395 428 407 431
rect 349 422 407 428
rect 539 428 551 431
rect 585 459 597 462
rect 729 462 787 468
rect 729 459 741 462
rect 585 431 741 459
rect 585 428 597 431
rect 539 422 597 428
rect 729 428 741 431
rect 775 459 787 462
rect 925 462 983 468
rect 925 459 937 462
rect 775 431 937 459
rect 775 428 787 431
rect 729 422 787 428
rect 925 428 937 431
rect 971 459 983 462
rect 1113 462 1171 468
rect 1113 459 1125 462
rect 971 431 1125 459
rect 971 428 983 431
rect 925 422 983 428
rect 1113 428 1125 431
rect 1159 428 1171 462
rect 1113 422 1171 428
rect 1313 462 1371 468
rect 1313 428 1325 462
rect 1359 459 1371 462
rect 1501 462 1559 468
rect 1501 459 1513 462
rect 1359 431 1513 459
rect 1359 428 1371 431
rect 1313 422 1371 428
rect 1501 428 1513 431
rect 1547 459 1559 462
rect 1697 462 1755 468
rect 1697 459 1709 462
rect 1547 431 1709 459
rect 1547 428 1559 431
rect 1501 422 1559 428
rect 1697 428 1709 431
rect 1743 459 1755 462
rect 1887 462 1945 468
rect 1887 459 1899 462
rect 1743 431 1899 459
rect 1743 428 1755 431
rect 1697 422 1755 428
rect 1887 428 1899 431
rect 1933 459 1945 462
rect 2077 462 2135 468
rect 2077 459 2089 462
rect 1933 431 2089 459
rect 1933 428 1945 431
rect 1887 422 1945 428
rect 2077 428 2089 431
rect 2123 428 2135 462
rect 2077 422 2135 428
rect 2833 462 2891 468
rect 2833 428 2845 462
rect 2879 459 2891 462
rect 3023 462 3081 468
rect 3023 459 3035 462
rect 2879 431 3035 459
rect 2879 428 2891 431
rect 2833 422 2891 428
rect 3023 428 3035 431
rect 3069 459 3081 462
rect 3213 462 3271 468
rect 3213 459 3225 462
rect 3069 431 3225 459
rect 3069 428 3081 431
rect 3023 422 3081 428
rect 3213 428 3225 431
rect 3259 459 3271 462
rect 3409 462 3467 468
rect 3409 459 3421 462
rect 3259 431 3421 459
rect 3259 428 3271 431
rect 3213 422 3271 428
rect 3409 428 3421 431
rect 3455 459 3467 462
rect 3597 462 3655 468
rect 3597 459 3609 462
rect 3455 431 3609 459
rect 3455 428 3467 431
rect 3409 422 3467 428
rect 3597 428 3609 431
rect 3643 428 3655 462
rect 3597 422 3655 428
rect 3797 462 3855 468
rect 3797 428 3809 462
rect 3843 459 3855 462
rect 3985 462 4043 468
rect 3985 459 3997 462
rect 3843 431 3997 459
rect 3843 428 3855 431
rect 3797 422 3855 428
rect 3985 428 3997 431
rect 4031 459 4043 462
rect 4181 462 4239 468
rect 4181 459 4193 462
rect 4031 431 4193 459
rect 4031 428 4043 431
rect 3985 422 4043 428
rect 4181 428 4193 431
rect 4227 459 4239 462
rect 4371 462 4429 468
rect 4371 459 4383 462
rect 4227 431 4383 459
rect 4227 428 4239 431
rect 4181 422 4239 428
rect 4371 428 4383 431
rect 4417 459 4429 462
rect 4561 462 4619 468
rect 4561 459 4573 462
rect 4417 431 4573 459
rect 4417 428 4429 431
rect 4371 422 4429 428
rect 4561 428 4573 431
rect 4607 428 4619 462
rect 4561 422 4619 428
rect 445 391 503 397
rect 445 357 457 391
rect 491 388 503 391
rect 633 391 691 397
rect 633 388 645 391
rect 491 360 645 388
rect 491 357 503 360
rect 445 351 503 357
rect 633 357 645 360
rect 679 388 691 391
rect 1793 391 1851 397
rect 1793 388 1805 391
rect 679 360 1805 388
rect 679 357 691 360
rect 633 351 691 357
rect 1793 357 1805 360
rect 1839 388 1851 391
rect 1981 391 2039 397
rect 1981 388 1993 391
rect 1839 360 1993 388
rect 1839 357 1851 360
rect 1793 351 1851 357
rect 1981 357 1993 360
rect 2027 388 2039 391
rect 2929 391 2987 397
rect 2929 388 2941 391
rect 2027 360 2941 388
rect 2027 357 2039 360
rect 1981 351 2039 357
rect 2929 357 2941 360
rect 2975 388 2987 391
rect 3117 391 3175 397
rect 3117 388 3129 391
rect 2975 360 3129 388
rect 2975 357 2987 360
rect 2929 351 2987 357
rect 3117 357 3129 360
rect 3163 388 3175 391
rect 4277 391 4335 397
rect 4277 388 4289 391
rect 3163 360 4289 388
rect 3163 357 3175 360
rect 3117 351 3175 357
rect 4277 357 4289 360
rect 4323 388 4335 391
rect 4465 391 4523 397
rect 4465 388 4477 391
rect 4323 360 4477 388
rect 4323 357 4335 360
rect 4277 351 4335 357
rect 4465 357 4477 360
rect 4511 357 4523 391
rect 4465 351 4523 357
rect 0 17 4968 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3341 17
rect 3375 -17 3433 17
rect 3467 -17 3525 17
rect 3559 -17 3617 17
rect 3651 -17 3709 17
rect 3743 -17 3801 17
rect 3835 -17 3893 17
rect 3927 -17 3985 17
rect 4019 -17 4077 17
rect 4111 -17 4169 17
rect 4203 -17 4261 17
rect 4295 -17 4353 17
rect 4387 -17 4445 17
rect 4479 -17 4537 17
rect 4571 -17 4629 17
rect 4663 -17 4721 17
rect 4755 -17 4813 17
rect 4847 -17 4905 17
rect 4939 -17 4968 17
rect 0 -48 4968 -17
<< labels >>
rlabel comment s 0 0 0 0 4 muxb8to1_4
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 17 nsew
flabel metal1 s 469 697 503 731 0 FreeSans 200 0 0 0 Z
port 21 nsew
flabel metal1 s 29 1071 63 1105 0 FreeSans 200 0 0 0 VGND
port 17 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 20 nsew
flabel metal1 s 469 357 503 391 0 FreeSans 200 0 0 0 Z
port 21 nsew
flabel metal1 s 3709 527 3743 561 0 FreeSans 200 0 0 0 VPWR
port 20 nsew
flabel metal1 s 3709 1071 3743 1105 0 FreeSans 200 0 0 0 VGND
port 17 nsew
flabel metal1 s 3726 544 3726 544 0 FreeSans 200 180 0 0 VPWR
port 20 nsew
flabel metal1 s 3726 1088 3726 1088 0 FreeSans 200 180 0 0 VGND
port 17 nsew
flabel metal1 s 3726 544 3726 544 0 FreeSans 200 180 0 0 VPWR
port 20 nsew
flabel metal1 s 3709 -17 3743 17 0 FreeSans 200 180 0 0 VGND
port 17 nsew
flabel metal1 s 3726 544 3726 544 0 FreeSans 200 0 0 0 VPWR
port 20 nsew
flabel metal1 s 3726 0 3726 0 0 FreeSans 200 0 0 0 VGND
port 17 nsew
flabel metal1 s 1225 527 1259 561 0 FreeSans 200 180 0 0 VPWR
port 20 nsew
flabel metal1 s 1225 1071 1259 1105 0 FreeSans 200 180 0 0 VGND
port 17 nsew
flabel metal1 s 1242 544 1242 544 0 FreeSans 200 180 0 0 VPWR
port 20 nsew
flabel metal1 s 1225 -17 1259 17 0 FreeSans 200 180 0 0 VGND
port 17 nsew
flabel metal1 s 1242 544 1242 544 0 FreeSans 200 0 0 0 VPWR
port 20 nsew
flabel metal1 s 1242 0 1242 0 0 FreeSans 200 0 0 0 VGND
port 17 nsew
flabel metal1 s 1242 544 1242 544 0 FreeSans 200 0 0 0 VPWR
port 20 nsew
flabel metal1 s 1242 1088 1242 1088 0 FreeSans 200 0 0 0 VGND
port 17 nsew
flabel pwell s 29 1071 63 1105 0 FreeSans 200 0 0 0 VNB
port 18 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 18 nsew
flabel pwell s 3709 1071 3743 1105 0 FreeSans 200 0 0 0 VNB
port 18 nsew
flabel pwell s 3726 1088 3726 1088 0 FreeSans 200 180 0 0 VNB
port 18 nsew
flabel pwell s 3709 -17 3743 17 0 FreeSans 200 180 0 0 VNB
port 18 nsew
flabel pwell s 3726 0 3726 0 0 FreeSans 200 0 0 0 VNB
port 18 nsew
flabel pwell s 1225 1071 1259 1105 0 FreeSans 200 180 0 0 VNB
port 18 nsew
flabel pwell s 1225 -17 1259 17 0 FreeSans 200 180 0 0 VNB
port 18 nsew
flabel pwell s 1242 0 1242 0 0 FreeSans 200 0 0 0 VNB
port 18 nsew
flabel pwell s 1242 1088 1242 1088 0 FreeSans 200 0 0 0 VNB
port 18 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 19 nsew
flabel nbase s 3709 527 3743 561 0 FreeSans 200 0 0 0 VPB
port 19 nsew
flabel nbase s 3726 544 3726 544 0 FreeSans 200 180 0 0 VPB
port 19 nsew
flabel nbase s 3726 544 3726 544 0 FreeSans 200 180 0 0 VPB
port 19 nsew
flabel nbase s 3726 544 3726 544 0 FreeSans 200 0 0 0 VPB
port 19 nsew
flabel nbase s 1225 527 1259 561 0 FreeSans 200 180 0 0 VPB
port 19 nsew
flabel nbase s 1242 544 1242 544 0 FreeSans 200 180 0 0 VPB
port 19 nsew
flabel nbase s 1242 544 1242 544 0 FreeSans 200 0 0 0 VPB
port 19 nsew
flabel nbase s 1242 544 1242 544 0 FreeSans 200 0 0 0 VPB
port 19 nsew
flabel corelocali s 4905 221 4939 255 0 FreeSans 200 0 0 0 S[6]
port 10 nsew
flabel corelocali s 1317 833 1351 867 0 FreeSans 200 0 0 0 D[3]
port 5 nsew
flabel corelocali s 1133 221 1167 255 0 FreeSans 200 0 0 0 D[0]
port 8 nsew
flabel corelocali s 3617 221 3651 255 0 FreeSans 200 0 0 0 D[4]
port 4 nsew
flabel corelocali s 3617 833 3651 867 0 FreeSans 200 0 0 0 D[5]
port 3 nsew
flabel corelocali s 1317 221 1351 255 0 FreeSans 200 0 0 0 D[2]
port 6 nsew
flabel corelocali s 1133 833 1167 867 0 FreeSans 200 0 0 0 D[1]
port 7 nsew
flabel corelocali s 3801 221 3835 255 0 FreeSans 200 0 0 0 D[6]
port 2 nsew
flabel corelocali s 2421 221 2455 255 0 FreeSans 200 0 0 0 S[2]
port 14 nsew
flabel corelocali s 2421 833 2455 867 0 FreeSans 200 0 0 0 S[3]
port 13 nsew
flabel corelocali s 4905 833 4939 867 0 FreeSans 200 0 0 0 S[7]
port 9 nsew
flabel corelocali s 29 221 63 255 0 FreeSans 200 0 0 0 S[0]
port 16 nsew
flabel corelocali s 29 833 63 867 0 FreeSans 200 0 0 0 S[1]
port 15 nsew
flabel corelocali s 2513 221 2547 255 0 FreeSans 200 0 0 0 S[4]
port 12 nsew
flabel corelocali s 2513 833 2547 867 0 FreeSans 200 0 0 0 S[5]
port 11 nsew
flabel corelocali s 3801 833 3835 867 0 FreeSans 200 0 0 0 D[7]
port 1 nsew
<< properties >>
string FIXED_BBOX -2 0 4966 1088
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2964294
string GDS_START 2893498
<< end >>
