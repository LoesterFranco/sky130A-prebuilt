magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 103 427 179 527
rect 18 195 88 325
rect 103 17 179 93
rect 311 427 377 527
rect 746 451 822 527
rect 374 201 466 325
rect 936 451 1012 527
rect 1294 451 1388 527
rect 311 17 377 93
rect 1542 389 1608 527
rect 782 17 874 105
rect 1028 17 1106 109
rect 1464 17 1606 113
rect 1840 299 1874 527
rect 1908 323 2003 492
rect 2037 357 2090 527
rect 1908 299 2097 323
rect 1950 165 2097 299
rect 1814 17 1890 165
rect 1937 149 2097 165
rect 1937 53 2003 149
rect 2037 17 2090 115
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
<< obsli1 >>
rect 35 393 69 493
rect 35 359 178 393
rect 132 161 178 359
rect 35 127 178 161
rect 35 69 69 127
rect 223 69 268 493
rect 421 393 455 493
rect 502 450 688 484
rect 306 359 455 393
rect 306 165 340 359
rect 500 315 620 391
rect 306 127 455 165
rect 500 141 554 315
rect 654 281 688 450
rect 868 417 902 475
rect 1112 433 1258 483
rect 1214 417 1258 433
rect 1428 417 1476 475
rect 722 367 1022 417
rect 722 315 782 367
rect 894 281 954 313
rect 654 247 954 281
rect 654 246 748 247
rect 590 129 670 203
rect 421 61 455 127
rect 704 93 748 246
rect 988 213 1022 367
rect 782 187 902 213
rect 782 153 856 187
rect 890 153 902 187
rect 782 147 902 153
rect 958 145 1022 213
rect 1066 331 1180 393
rect 1214 383 1476 417
rect 1066 179 1100 331
rect 1144 213 1180 295
rect 1214 281 1258 383
rect 1642 353 1676 475
rect 1730 383 1796 485
rect 1642 349 1710 353
rect 1292 315 1710 349
rect 1214 247 1634 281
rect 1274 179 1350 203
rect 1066 145 1350 179
rect 525 53 748 93
rect 958 59 992 145
rect 1384 95 1418 247
rect 1558 235 1634 247
rect 1452 201 1528 213
rect 1452 187 1556 201
rect 1452 153 1501 187
rect 1535 153 1556 187
rect 1452 147 1556 153
rect 1668 136 1710 315
rect 1238 61 1418 95
rect 1642 70 1710 136
rect 1746 265 1796 383
rect 1746 199 1916 265
rect 1746 69 1780 199
<< obsli1c >>
rect 856 153 890 187
rect 1501 153 1535 187
<< metal1 >>
rect 0 561 2116 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 0 496 2116 527
rect 844 187 902 193
rect 844 153 856 187
rect 890 184 902 187
rect 1489 187 1547 193
rect 1489 184 1501 187
rect 890 156 1501 184
rect 890 153 902 156
rect 844 147 902 153
rect 1489 153 1501 156
rect 1535 153 1547 187
rect 1489 147 1547 153
rect 0 17 2116 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
rect 0 -48 2116 -17
<< obsm1 >>
rect 121 360 1187 388
rect 121 342 179 360
rect 517 342 575 360
rect 1129 342 1187 360
rect 1133 252 1191 262
rect 634 224 1191 252
rect 634 184 677 224
rect 1133 216 1191 224
rect 221 156 677 184
rect 221 138 279 156
rect 619 138 677 156
<< labels >>
rlabel locali s 18 195 88 325 6 CLK
port 1 nsew signal input
rlabel locali s 374 201 466 325 6 D
port 2 nsew signal input
rlabel locali s 1950 165 2097 299 6 Q
port 3 nsew signal output
rlabel locali s 1937 149 2097 165 6 Q
port 3 nsew signal output
rlabel locali s 1937 53 2003 149 6 Q
port 3 nsew signal output
rlabel locali s 1908 323 2003 492 6 Q
port 3 nsew signal output
rlabel locali s 1908 299 2097 323 6 Q
port 3 nsew signal output
rlabel metal1 s 1489 184 1547 193 6 SET_B
port 4 nsew signal input
rlabel metal1 s 1489 147 1547 156 6 SET_B
port 4 nsew signal input
rlabel metal1 s 844 184 902 193 6 SET_B
port 4 nsew signal input
rlabel metal1 s 844 156 1547 184 6 SET_B
port 4 nsew signal input
rlabel metal1 s 844 147 902 156 6 SET_B
port 4 nsew signal input
rlabel viali s 2053 -17 2087 17 8 VGND
port 5 nsew ground bidirectional
rlabel viali s 1961 -17 1995 17 8 VGND
port 5 nsew ground bidirectional
rlabel viali s 1869 -17 1903 17 8 VGND
port 5 nsew ground bidirectional
rlabel viali s 1777 -17 1811 17 8 VGND
port 5 nsew ground bidirectional
rlabel viali s 1685 -17 1719 17 8 VGND
port 5 nsew ground bidirectional
rlabel viali s 1593 -17 1627 17 8 VGND
port 5 nsew ground bidirectional
rlabel viali s 1501 -17 1535 17 8 VGND
port 5 nsew ground bidirectional
rlabel viali s 1409 -17 1443 17 8 VGND
port 5 nsew ground bidirectional
rlabel viali s 1317 -17 1351 17 8 VGND
port 5 nsew ground bidirectional
rlabel viali s 1225 -17 1259 17 8 VGND
port 5 nsew ground bidirectional
rlabel viali s 1133 -17 1167 17 8 VGND
port 5 nsew ground bidirectional
rlabel viali s 1041 -17 1075 17 8 VGND
port 5 nsew ground bidirectional
rlabel viali s 949 -17 983 17 8 VGND
port 5 nsew ground bidirectional
rlabel viali s 857 -17 891 17 8 VGND
port 5 nsew ground bidirectional
rlabel viali s 765 -17 799 17 8 VGND
port 5 nsew ground bidirectional
rlabel viali s 673 -17 707 17 8 VGND
port 5 nsew ground bidirectional
rlabel viali s 581 -17 615 17 8 VGND
port 5 nsew ground bidirectional
rlabel viali s 489 -17 523 17 8 VGND
port 5 nsew ground bidirectional
rlabel viali s 397 -17 431 17 8 VGND
port 5 nsew ground bidirectional
rlabel viali s 305 -17 339 17 8 VGND
port 5 nsew ground bidirectional
rlabel viali s 213 -17 247 17 8 VGND
port 5 nsew ground bidirectional
rlabel viali s 121 -17 155 17 8 VGND
port 5 nsew ground bidirectional
rlabel viali s 29 -17 63 17 8 VGND
port 5 nsew ground bidirectional
rlabel locali s 2037 17 2090 115 6 VGND
port 5 nsew ground bidirectional
rlabel locali s 1814 17 1890 165 6 VGND
port 5 nsew ground bidirectional
rlabel locali s 1464 17 1606 113 6 VGND
port 5 nsew ground bidirectional
rlabel locali s 1028 17 1106 109 6 VGND
port 5 nsew ground bidirectional
rlabel locali s 782 17 874 105 6 VGND
port 5 nsew ground bidirectional
rlabel locali s 311 17 377 93 6 VGND
port 5 nsew ground bidirectional
rlabel locali s 103 17 179 93 6 VGND
port 5 nsew ground bidirectional
rlabel locali s 0 -17 2116 17 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 -48 2116 48 8 VGND
port 5 nsew ground bidirectional
rlabel viali s 2053 527 2087 561 6 VPWR
port 6 nsew power bidirectional
rlabel viali s 1961 527 1995 561 6 VPWR
port 6 nsew power bidirectional
rlabel viali s 1869 527 1903 561 6 VPWR
port 6 nsew power bidirectional
rlabel viali s 1777 527 1811 561 6 VPWR
port 6 nsew power bidirectional
rlabel viali s 1685 527 1719 561 6 VPWR
port 6 nsew power bidirectional
rlabel viali s 1593 527 1627 561 6 VPWR
port 6 nsew power bidirectional
rlabel viali s 1501 527 1535 561 6 VPWR
port 6 nsew power bidirectional
rlabel viali s 1409 527 1443 561 6 VPWR
port 6 nsew power bidirectional
rlabel viali s 1317 527 1351 561 6 VPWR
port 6 nsew power bidirectional
rlabel viali s 1225 527 1259 561 6 VPWR
port 6 nsew power bidirectional
rlabel viali s 1133 527 1167 561 6 VPWR
port 6 nsew power bidirectional
rlabel viali s 1041 527 1075 561 6 VPWR
port 6 nsew power bidirectional
rlabel viali s 949 527 983 561 6 VPWR
port 6 nsew power bidirectional
rlabel viali s 857 527 891 561 6 VPWR
port 6 nsew power bidirectional
rlabel viali s 765 527 799 561 6 VPWR
port 6 nsew power bidirectional
rlabel viali s 673 527 707 561 6 VPWR
port 6 nsew power bidirectional
rlabel viali s 581 527 615 561 6 VPWR
port 6 nsew power bidirectional
rlabel viali s 489 527 523 561 6 VPWR
port 6 nsew power bidirectional
rlabel viali s 397 527 431 561 6 VPWR
port 6 nsew power bidirectional
rlabel viali s 305 527 339 561 6 VPWR
port 6 nsew power bidirectional
rlabel viali s 213 527 247 561 6 VPWR
port 6 nsew power bidirectional
rlabel viali s 121 527 155 561 6 VPWR
port 6 nsew power bidirectional
rlabel viali s 29 527 63 561 6 VPWR
port 6 nsew power bidirectional
rlabel locali s 2037 357 2090 527 6 VPWR
port 6 nsew power bidirectional
rlabel locali s 1840 299 1874 527 6 VPWR
port 6 nsew power bidirectional
rlabel locali s 1542 389 1608 527 6 VPWR
port 6 nsew power bidirectional
rlabel locali s 1294 451 1388 527 6 VPWR
port 6 nsew power bidirectional
rlabel locali s 936 451 1012 527 6 VPWR
port 6 nsew power bidirectional
rlabel locali s 746 451 822 527 6 VPWR
port 6 nsew power bidirectional
rlabel locali s 311 427 377 527 6 VPWR
port 6 nsew power bidirectional
rlabel locali s 103 427 179 527 6 VPWR
port 6 nsew power bidirectional
rlabel locali s 0 527 2116 561 6 VPWR
port 6 nsew power bidirectional
rlabel metal1 s 0 496 2116 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2116 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1909744
string GDS_START 1893024
<< end >>
