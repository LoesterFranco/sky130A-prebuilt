magic
tech sky130A
magscale 1 2
timestamp 1599588218
<< nwell >>
rect -38 332 1190 704
<< pwell >>
rect 0 0 1152 49
<< scpmos >>
rect 121 368 157 592
rect 211 368 247 592
rect 301 368 337 592
rect 391 368 427 592
rect 585 368 621 592
rect 675 368 711 592
rect 765 368 801 592
rect 855 368 891 592
rect 945 368 981 592
rect 1035 368 1071 592
<< nmoslvt >>
rect 193 74 223 222
rect 301 74 331 222
rect 409 74 439 222
rect 775 74 805 222
rect 861 74 891 222
rect 947 74 977 222
rect 1035 74 1065 222
<< ndiff >>
rect 136 152 193 222
rect 136 118 148 152
rect 182 118 193 152
rect 136 74 193 118
rect 223 210 301 222
rect 223 176 248 210
rect 282 176 301 210
rect 223 120 301 176
rect 223 86 248 120
rect 282 86 301 120
rect 223 74 301 86
rect 331 152 409 222
rect 331 118 349 152
rect 383 118 409 152
rect 331 74 409 118
rect 439 210 492 222
rect 439 176 450 210
rect 484 176 492 210
rect 439 120 492 176
rect 439 86 450 120
rect 484 86 492 120
rect 439 74 492 86
rect 722 120 775 222
rect 722 86 730 120
rect 764 86 775 120
rect 722 74 775 86
rect 805 207 861 222
rect 805 173 816 207
rect 850 173 861 207
rect 805 74 861 173
rect 891 210 947 222
rect 891 176 902 210
rect 936 176 947 210
rect 891 120 947 176
rect 891 86 902 120
rect 936 86 947 120
rect 891 74 947 86
rect 977 152 1035 222
rect 977 118 989 152
rect 1023 118 1035 152
rect 977 74 1035 118
rect 1065 210 1118 222
rect 1065 176 1076 210
rect 1110 176 1118 210
rect 1065 120 1118 176
rect 1065 86 1076 120
rect 1110 86 1118 120
rect 1065 74 1118 86
<< pdiff >>
rect 69 580 121 592
rect 69 546 77 580
rect 111 546 121 580
rect 69 508 121 546
rect 69 474 77 508
rect 111 474 121 508
rect 69 368 121 474
rect 157 531 211 592
rect 157 497 167 531
rect 201 497 211 531
rect 157 440 211 497
rect 157 406 167 440
rect 201 406 211 440
rect 157 368 211 406
rect 247 580 301 592
rect 247 546 257 580
rect 291 546 301 580
rect 247 510 301 546
rect 247 476 257 510
rect 291 476 301 510
rect 247 440 301 476
rect 247 406 257 440
rect 291 406 301 440
rect 247 368 301 406
rect 337 531 391 592
rect 337 497 347 531
rect 381 497 391 531
rect 337 440 391 497
rect 337 406 347 440
rect 381 406 391 440
rect 337 368 391 406
rect 427 580 479 592
rect 427 546 437 580
rect 471 546 479 580
rect 427 508 479 546
rect 427 474 437 508
rect 471 474 479 508
rect 427 368 479 474
rect 533 580 585 592
rect 533 546 541 580
rect 575 546 585 580
rect 533 508 585 546
rect 533 474 541 508
rect 575 474 585 508
rect 533 368 585 474
rect 621 531 675 592
rect 621 497 631 531
rect 665 497 675 531
rect 621 414 675 497
rect 621 380 631 414
rect 665 380 675 414
rect 621 368 675 380
rect 711 580 765 592
rect 711 546 721 580
rect 755 546 765 580
rect 711 506 765 546
rect 711 472 721 506
rect 755 472 765 506
rect 711 424 765 472
rect 711 390 721 424
rect 755 390 765 424
rect 711 368 765 390
rect 801 580 855 592
rect 801 546 811 580
rect 845 546 855 580
rect 801 508 855 546
rect 801 474 811 508
rect 845 474 855 508
rect 801 368 855 474
rect 891 580 945 592
rect 891 546 901 580
rect 935 546 945 580
rect 891 506 945 546
rect 891 472 901 506
rect 935 472 945 506
rect 891 424 945 472
rect 891 390 901 424
rect 935 390 945 424
rect 891 368 945 390
rect 981 580 1035 592
rect 981 546 991 580
rect 1025 546 1035 580
rect 981 498 1035 546
rect 981 464 991 498
rect 1025 464 1035 498
rect 981 368 1035 464
rect 1071 580 1123 592
rect 1071 546 1081 580
rect 1115 546 1123 580
rect 1071 497 1123 546
rect 1071 463 1081 497
rect 1115 463 1123 497
rect 1071 414 1123 463
rect 1071 380 1081 414
rect 1115 380 1123 414
rect 1071 368 1123 380
<< ndiffc >>
rect 148 118 182 152
rect 248 176 282 210
rect 248 86 282 120
rect 349 118 383 152
rect 450 176 484 210
rect 450 86 484 120
rect 730 86 764 120
rect 816 173 850 207
rect 902 176 936 210
rect 902 86 936 120
rect 989 118 1023 152
rect 1076 176 1110 210
rect 1076 86 1110 120
<< pdiffc >>
rect 77 546 111 580
rect 77 474 111 508
rect 167 497 201 531
rect 167 406 201 440
rect 257 546 291 580
rect 257 476 291 510
rect 257 406 291 440
rect 347 497 381 531
rect 347 406 381 440
rect 437 546 471 580
rect 437 474 471 508
rect 541 546 575 580
rect 541 474 575 508
rect 631 497 665 531
rect 631 380 665 414
rect 721 546 755 580
rect 721 472 755 506
rect 721 390 755 424
rect 811 546 845 580
rect 811 474 845 508
rect 901 546 935 580
rect 901 472 935 506
rect 901 390 935 424
rect 991 546 1025 580
rect 991 464 1025 498
rect 1081 546 1115 580
rect 1081 463 1115 497
rect 1081 380 1115 414
<< poly >>
rect 121 592 157 618
rect 211 592 247 618
rect 301 592 337 618
rect 391 592 427 618
rect 585 592 621 618
rect 675 592 711 618
rect 765 592 801 618
rect 855 592 891 618
rect 945 592 981 618
rect 1035 592 1071 618
rect 121 336 157 368
rect 211 336 247 368
rect 301 345 337 368
rect 391 345 427 368
rect 121 320 259 336
rect 121 286 209 320
rect 243 286 259 320
rect 121 270 259 286
rect 301 320 427 345
rect 301 286 317 320
rect 351 315 427 320
rect 351 286 367 315
rect 301 270 367 286
rect 585 310 621 368
rect 675 310 711 368
rect 585 294 711 310
rect 193 222 223 270
rect 301 222 331 270
rect 585 267 661 294
rect 409 260 661 267
rect 695 260 711 294
rect 765 336 801 368
rect 855 336 891 368
rect 765 320 891 336
rect 765 286 809 320
rect 843 286 891 320
rect 765 270 891 286
rect 945 336 981 368
rect 1035 336 1071 368
rect 945 320 1071 336
rect 945 286 986 320
rect 1020 300 1071 320
rect 1020 286 1065 300
rect 945 270 1065 286
rect 409 237 711 260
rect 409 222 439 237
rect 775 222 805 270
rect 861 222 891 270
rect 947 222 977 270
rect 1035 222 1065 270
rect 193 48 223 74
rect 301 48 331 74
rect 409 48 439 74
rect 775 48 805 74
rect 861 48 891 74
rect 947 48 977 74
rect 1035 48 1065 74
<< polycont >>
rect 209 286 243 320
rect 317 286 351 320
rect 661 260 695 294
rect 809 286 843 320
rect 986 286 1020 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 61 581 487 615
rect 61 580 111 581
rect 61 546 77 580
rect 257 580 291 581
rect 61 508 111 546
rect 61 474 77 508
rect 61 458 111 474
rect 151 531 217 547
rect 151 497 167 531
rect 201 497 217 531
rect 151 440 217 497
rect 151 424 167 440
rect 25 406 167 424
rect 201 406 217 440
rect 25 390 217 406
rect 437 580 487 581
rect 257 510 291 546
rect 257 440 291 476
rect 257 390 291 406
rect 331 531 397 547
rect 331 497 347 531
rect 381 497 397 531
rect 331 440 397 497
rect 471 546 487 580
rect 437 508 487 546
rect 471 474 487 508
rect 437 458 487 474
rect 525 581 771 615
rect 525 580 581 581
rect 525 546 541 580
rect 575 546 581 580
rect 705 580 771 581
rect 525 508 581 546
rect 525 474 541 508
rect 575 474 581 508
rect 525 458 581 474
rect 615 531 665 547
rect 615 497 631 531
rect 331 406 347 440
rect 381 424 397 440
rect 615 424 665 497
rect 381 414 665 424
rect 381 406 631 414
rect 331 390 631 406
rect 25 236 71 390
rect 615 380 631 390
rect 705 546 721 580
rect 755 546 771 580
rect 705 506 771 546
rect 705 472 721 506
rect 755 472 771 506
rect 705 424 771 472
rect 811 580 845 649
rect 811 508 845 546
rect 811 458 845 474
rect 885 580 935 596
rect 885 546 901 580
rect 885 506 935 546
rect 885 472 901 506
rect 885 424 935 472
rect 975 580 1041 649
rect 975 546 991 580
rect 1025 546 1041 580
rect 975 498 1041 546
rect 975 464 991 498
rect 1025 464 1041 498
rect 975 458 1041 464
rect 1081 580 1131 596
rect 1115 546 1131 580
rect 1081 497 1131 546
rect 1115 463 1131 497
rect 1081 424 1131 463
rect 705 390 721 424
rect 755 390 901 424
rect 935 414 1131 424
rect 935 390 1081 414
rect 615 364 665 380
rect 1115 380 1131 414
rect 1081 364 1131 380
rect 121 320 263 356
rect 121 286 209 320
rect 243 286 263 320
rect 121 270 263 286
rect 301 320 551 356
rect 301 286 317 320
rect 351 286 551 320
rect 793 320 935 356
rect 301 270 551 286
rect 601 294 743 310
rect 601 260 661 294
rect 695 260 743 294
rect 793 286 809 320
rect 843 286 935 320
rect 793 270 935 286
rect 970 320 1036 356
rect 970 286 986 320
rect 1020 286 1036 320
rect 970 270 1036 286
rect 601 236 743 260
rect 25 210 500 236
rect 25 202 248 210
rect 232 176 248 202
rect 282 202 450 210
rect 282 176 298 202
rect 132 152 198 168
rect 132 118 148 152
rect 182 118 198 152
rect 132 17 198 118
rect 232 120 298 176
rect 434 176 450 202
rect 484 195 500 210
rect 800 207 866 226
rect 800 195 816 207
rect 484 176 816 195
rect 434 173 816 176
rect 850 173 866 207
rect 232 86 248 120
rect 282 86 298 120
rect 232 70 298 86
rect 332 152 400 168
rect 332 118 349 152
rect 383 118 400 152
rect 332 17 400 118
rect 434 154 866 173
rect 902 210 1126 236
rect 936 202 1076 210
rect 434 120 500 154
rect 902 120 936 176
rect 1110 176 1126 210
rect 434 86 450 120
rect 484 86 500 120
rect 434 70 500 86
rect 714 86 730 120
rect 764 86 902 120
rect 714 70 936 86
rect 972 152 1040 168
rect 972 118 989 152
rect 1023 118 1040 152
rect 972 17 1040 118
rect 1076 120 1126 176
rect 1110 86 1126 120
rect 1076 70 1126 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
rlabel comment s 0 0 0 0 4 a2111oi_2
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 D1
port 5 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 D1
port 5 nsew
flabel corelocali s 607 242 641 276 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 703 242 737 276 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 1152 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3862148
string GDS_START 3852556
<< end >>
