magic
tech sky130A
magscale 1 2
timestamp 1599588238
<< locali >>
rect 120 424 186 596
rect 300 424 366 596
rect 120 390 455 424
rect 25 270 360 356
rect 409 236 455 390
rect 123 202 455 236
rect 123 70 173 202
rect 321 70 355 202
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 30 390 80 649
rect 226 458 260 649
rect 406 458 456 649
rect 23 17 89 226
rect 209 17 275 168
rect 391 17 457 168
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< metal1 >>
rect 0 683 480 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 0 617 480 649
rect 0 17 480 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
rect 0 -49 480 -17
<< labels >>
rlabel locali s 25 270 360 356 6 A
port 1 nsew signal input
rlabel locali s 409 236 455 390 6 Y
port 2 nsew signal output
rlabel locali s 321 70 355 202 6 Y
port 2 nsew signal output
rlabel locali s 300 424 366 596 6 Y
port 2 nsew signal output
rlabel locali s 123 202 455 236 6 Y
port 2 nsew signal output
rlabel locali s 123 70 173 202 6 Y
port 2 nsew signal output
rlabel locali s 120 424 186 596 6 Y
port 2 nsew signal output
rlabel locali s 120 390 455 424 6 Y
port 2 nsew signal output
rlabel metal1 s 0 -49 480 49 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 617 480 715 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 480 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2405640
string GDS_START 2400486
<< end >>
