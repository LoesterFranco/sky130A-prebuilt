magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 828 561
rect 103 439 169 527
rect 311 451 445 527
rect 568 439 634 527
rect 27 148 67 326
rect 19 17 85 93
rect 305 84 349 349
rect 392 84 455 339
rect 489 129 555 323
rect 668 349 709 493
rect 743 383 810 527
rect 668 307 811 349
rect 685 165 811 307
rect 652 128 811 165
rect 552 17 618 93
rect 652 51 709 128
rect 743 17 810 93
rect 0 -17 828 17
<< obsli1 >>
rect 35 400 69 493
rect 203 417 237 493
rect 488 417 522 493
rect 35 366 161 400
rect 127 265 161 366
rect 203 393 522 417
rect 203 383 633 393
rect 203 332 263 383
rect 488 359 633 383
rect 127 199 195 265
rect 127 117 161 199
rect 229 117 263 332
rect 119 51 161 117
rect 219 51 263 117
rect 599 265 633 359
rect 599 199 651 265
<< metal1 >>
rect 0 496 828 592
rect 0 -48 828 48
<< labels >>
rlabel locali s 27 148 67 326 6 A_N
port 1 nsew signal input
rlabel locali s 305 84 349 349 6 B
port 2 nsew signal input
rlabel locali s 392 84 455 339 6 C
port 3 nsew signal input
rlabel locali s 489 129 555 323 6 D
port 4 nsew signal input
rlabel locali s 685 165 811 307 6 X
port 5 nsew signal output
rlabel locali s 668 349 709 493 6 X
port 5 nsew signal output
rlabel locali s 668 307 811 349 6 X
port 5 nsew signal output
rlabel locali s 652 128 811 165 6 X
port 5 nsew signal output
rlabel locali s 652 51 709 128 6 X
port 5 nsew signal output
rlabel locali s 743 17 810 93 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 552 17 618 93 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 19 17 85 93 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 828 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 828 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 743 383 810 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 568 439 634 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 311 451 445 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 103 439 169 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 828 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 828 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3851210
string GDS_START 3842998
<< end >>
