magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 636 325 678 425
rect 489 257 587 325
rect 636 291 799 325
rect 27 215 203 257
rect 247 215 455 257
rect 489 215 662 257
rect 696 181 799 291
rect 107 145 799 181
rect 107 51 183 145
rect 295 51 371 145
rect 610 51 686 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 30 325 81 493
rect 125 359 175 527
rect 219 325 269 493
rect 313 459 772 493
rect 313 359 363 459
rect 407 325 455 425
rect 542 359 584 459
rect 722 359 772 459
rect 30 291 455 325
rect 18 17 73 181
rect 227 17 261 111
rect 415 17 576 111
rect 730 17 788 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
rlabel locali s 27 215 203 257 6 A
port 1 nsew signal input
rlabel locali s 247 215 455 257 6 B
port 2 nsew signal input
rlabel locali s 489 257 587 325 6 C
port 3 nsew signal input
rlabel locali s 489 215 662 257 6 C
port 3 nsew signal input
rlabel locali s 696 181 799 291 6 Y
port 4 nsew signal output
rlabel locali s 636 325 678 425 6 Y
port 4 nsew signal output
rlabel locali s 636 291 799 325 6 Y
port 4 nsew signal output
rlabel locali s 610 51 686 145 6 Y
port 4 nsew signal output
rlabel locali s 295 51 371 145 6 Y
port 4 nsew signal output
rlabel locali s 107 145 799 181 6 Y
port 4 nsew signal output
rlabel locali s 107 51 183 145 6 Y
port 4 nsew signal output
rlabel metal1 s 0 -48 828 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 828 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2441178
string GDS_START 2434278
<< end >>
