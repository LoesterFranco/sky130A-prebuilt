magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 17 341 73 493
rect 380 436 501 493
rect 380 341 493 436
rect 17 299 493 341
rect 571 323 625 481
rect 17 199 93 265
rect 135 165 169 299
rect 527 289 625 323
rect 203 199 319 265
rect 363 199 465 265
rect 527 249 579 289
rect 501 215 579 249
rect 613 215 715 255
rect 17 129 169 165
rect 17 73 69 129
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 120 375 316 527
rect 663 291 715 527
rect 489 165 715 173
rect 250 139 715 165
rect 250 129 512 139
rect 103 61 413 95
rect 457 56 512 129
rect 569 17 603 105
rect 637 56 715 139
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel locali s 613 215 715 255 6 A1
port 1 nsew signal input
rlabel locali s 571 323 625 481 6 A2
port 2 nsew signal input
rlabel locali s 527 289 625 323 6 A2
port 2 nsew signal input
rlabel locali s 527 249 579 289 6 A2
port 2 nsew signal input
rlabel locali s 501 215 579 249 6 A2
port 2 nsew signal input
rlabel locali s 203 199 319 265 6 B1
port 3 nsew signal input
rlabel locali s 363 199 465 265 6 B2
port 4 nsew signal input
rlabel locali s 17 199 93 265 6 C1
port 5 nsew signal input
rlabel locali s 380 436 501 493 6 Y
port 6 nsew signal output
rlabel locali s 380 341 493 436 6 Y
port 6 nsew signal output
rlabel locali s 135 165 169 299 6 Y
port 6 nsew signal output
rlabel locali s 17 341 73 493 6 Y
port 6 nsew signal output
rlabel locali s 17 299 493 341 6 Y
port 6 nsew signal output
rlabel locali s 17 129 169 165 6 Y
port 6 nsew signal output
rlabel locali s 17 73 69 129 6 Y
port 6 nsew signal output
rlabel metal1 s 0 -48 736 48 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 496 736 592 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 835850
string GDS_START 829290
<< end >>
