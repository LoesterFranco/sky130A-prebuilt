magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 203 340 241 493
rect 395 340 431 493
rect 18 306 431 340
rect 18 161 70 306
rect 547 215 697 323
rect 752 299 1176 341
rect 752 198 823 299
rect 884 199 1014 265
rect 1082 199 1176 299
rect 18 127 373 161
rect 129 123 373 127
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 83 374 159 527
rect 275 374 351 527
rect 467 451 547 527
rect 591 421 639 493
rect 703 455 769 527
rect 899 421 975 489
rect 591 417 975 421
rect 465 375 975 417
rect 1091 387 1173 527
rect 465 366 639 375
rect 465 267 513 366
rect 104 199 513 267
rect 463 174 513 199
rect 463 131 677 174
rect 711 123 1167 157
rect 711 97 777 123
rect 19 17 85 93
rect 211 17 277 89
rect 403 17 469 93
rect 517 51 777 97
rect 811 17 879 89
rect 995 17 1071 89
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
rlabel locali s 1082 199 1176 299 6 A1
port 1 nsew signal input
rlabel locali s 752 299 1176 341 6 A1
port 1 nsew signal input
rlabel locali s 752 198 823 299 6 A1
port 1 nsew signal input
rlabel locali s 884 199 1014 265 6 A2
port 2 nsew signal input
rlabel locali s 547 215 697 323 6 B1
port 3 nsew signal input
rlabel locali s 395 340 431 493 6 X
port 4 nsew signal output
rlabel locali s 203 340 241 493 6 X
port 4 nsew signal output
rlabel locali s 129 123 373 127 6 X
port 4 nsew signal output
rlabel locali s 18 306 431 340 6 X
port 4 nsew signal output
rlabel locali s 18 161 70 306 6 X
port 4 nsew signal output
rlabel locali s 18 127 373 161 6 X
port 4 nsew signal output
rlabel metal1 s 0 -48 1196 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 1196 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1022888
string GDS_START 1014548
<< end >>
