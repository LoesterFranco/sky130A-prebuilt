magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 552 561
rect 19 53 71 491
rect 105 381 173 527
rect 379 385 445 527
rect 203 203 296 265
rect 332 203 437 265
rect 123 17 257 91
rect 391 75 437 203
rect 473 199 533 265
rect 473 17 531 163
rect 0 -17 552 17
<< obsli1 >>
rect 209 345 263 491
rect 109 301 263 345
rect 299 349 345 491
rect 479 349 531 491
rect 299 301 531 349
rect 109 167 167 301
rect 109 127 355 167
rect 293 53 355 127
<< metal1 >>
rect 0 496 552 592
rect 0 -48 552 48
<< labels >>
rlabel locali s 391 75 437 203 6 A1
port 1 nsew signal input
rlabel locali s 332 203 437 265 6 A1
port 1 nsew signal input
rlabel locali s 473 199 533 265 6 A2
port 2 nsew signal input
rlabel locali s 203 203 296 265 6 B1
port 3 nsew signal input
rlabel locali s 19 53 71 491 6 X
port 4 nsew signal output
rlabel locali s 473 17 531 163 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 123 17 257 91 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 552 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 552 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 379 385 445 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 105 381 173 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 552 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 552 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 552 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 4082314
string GDS_START 4076324
<< end >>
