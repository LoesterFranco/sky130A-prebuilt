magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 19 337 74 491
rect 19 299 146 337
rect 19 135 67 265
rect 101 165 146 299
rect 180 199 259 265
rect 305 199 364 265
rect 101 129 177 165
rect 132 53 177 129
rect 213 75 259 199
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 108 405 184 491
rect 228 439 267 527
rect 303 405 379 491
rect 108 371 379 405
rect 180 305 379 371
rect 22 17 88 95
rect 319 17 379 163
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
rlabel locali s 213 75 259 199 6 A1
port 1 nsew signal input
rlabel locali s 180 199 259 265 6 A1
port 1 nsew signal input
rlabel locali s 305 199 364 265 6 A2
port 2 nsew signal input
rlabel locali s 19 135 67 265 6 B1
port 3 nsew signal input
rlabel locali s 132 53 177 129 6 Y
port 4 nsew signal output
rlabel locali s 101 165 146 299 6 Y
port 4 nsew signal output
rlabel locali s 101 129 177 165 6 Y
port 4 nsew signal output
rlabel locali s 19 337 74 491 6 Y
port 4 nsew signal output
rlabel locali s 19 299 146 337 6 Y
port 4 nsew signal output
rlabel metal1 s 0 -48 460 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 460 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 460 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1199586
string GDS_START 1194660
<< end >>
