magic
tech sky130A
magscale 1 2
timestamp 1599588238
<< locali >>
rect 21 260 75 356
rect 186 290 257 356
rect 1255 364 1327 596
rect 1087 270 1153 356
rect 1293 168 1327 364
rect 1220 70 1327 168
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 23 512 89 596
rect 123 546 189 649
rect 466 546 541 649
rect 581 581 809 615
rect 23 478 539 512
rect 23 420 143 478
rect 109 226 143 420
rect 230 394 325 444
rect 359 404 434 444
rect 291 356 325 394
rect 291 290 366 356
rect 291 226 325 290
rect 400 256 434 404
rect 505 360 539 478
rect 581 428 615 581
rect 649 481 707 547
rect 581 394 639 428
rect 505 294 571 360
rect 605 290 639 394
rect 673 379 707 481
rect 743 413 809 581
rect 887 530 1015 649
rect 1049 476 1115 596
rect 861 413 1115 476
rect 1019 390 1115 413
rect 1149 390 1215 649
rect 673 345 985 379
rect 605 256 665 290
rect 44 108 143 226
rect 177 17 211 226
rect 247 188 325 226
rect 359 222 665 256
rect 247 154 604 188
rect 699 185 733 345
rect 247 70 325 154
rect 459 17 536 120
rect 570 85 604 154
rect 638 119 733 185
rect 767 245 819 311
rect 933 294 985 345
rect 767 85 801 245
rect 1019 236 1053 390
rect 1195 236 1259 310
rect 954 202 1259 236
rect 570 51 801 85
rect 842 17 908 162
rect 954 70 1020 202
rect 1118 17 1184 168
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
<< metal1 >>
rect 0 683 1344 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 0 617 1344 649
rect 0 17 1344 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
rect 0 -49 1344 -17
<< labels >>
rlabel locali s 21 260 75 356 6 D
port 1 nsew signal input
rlabel locali s 1293 168 1327 364 6 Q
port 2 nsew signal output
rlabel locali s 1255 364 1327 596 6 Q
port 2 nsew signal output
rlabel locali s 1220 70 1327 168 6 Q
port 2 nsew signal output
rlabel locali s 1087 270 1153 356 6 RESET_B
port 3 nsew signal input
rlabel locali s 186 290 257 356 6 GATE
port 4 nsew clock input
rlabel metal1 s 0 -49 1344 49 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1344 715 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1344 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2934316
string GDS_START 2924030
<< end >>
