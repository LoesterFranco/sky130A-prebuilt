magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 386 1766 704
rect -38 341 641 386
rect -38 332 443 341
rect 895 332 1766 386
<< pwell >>
rect 0 0 1728 49
<< scnmos >>
rect 84 74 114 222
rect 256 80 286 208
rect 334 80 364 208
rect 461 124 491 208
rect 581 189 611 273
rect 724 125 754 273
rect 931 74 961 222
rect 1017 74 1047 222
rect 1095 74 1125 222
rect 1342 74 1372 222
rect 1428 74 1458 222
rect 1528 74 1558 222
rect 1614 74 1644 222
<< pmoshvt >>
rect 105 368 135 592
rect 253 392 283 592
rect 337 392 367 592
rect 494 508 524 592
rect 578 508 608 592
rect 702 424 732 592
rect 904 422 934 590
rect 1014 368 1044 592
rect 1111 368 1141 592
rect 1332 368 1362 592
rect 1425 368 1455 592
rect 1522 368 1552 592
rect 1612 368 1642 592
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 208 164 222
rect 769 306 827 318
rect 769 273 781 306
rect 511 208 581 273
rect 114 120 256 208
rect 114 86 130 120
rect 164 86 256 120
rect 114 80 256 86
rect 286 80 334 208
rect 364 180 461 208
rect 364 146 395 180
rect 429 146 461 180
rect 364 124 461 146
rect 491 189 581 208
rect 611 189 724 273
rect 491 124 541 189
rect 364 80 414 124
rect 667 170 724 189
rect 667 136 679 170
rect 713 136 724 170
rect 667 125 724 136
rect 754 272 781 273
rect 815 272 827 306
rect 754 243 827 272
rect 754 125 804 243
rect 881 166 931 222
rect 860 154 931 166
rect 114 74 181 80
rect 860 120 872 154
rect 906 120 931 154
rect 860 74 931 120
rect 961 154 1017 222
rect 961 120 972 154
rect 1006 120 1017 154
rect 961 74 1017 120
rect 1047 74 1095 222
rect 1125 210 1182 222
rect 1125 176 1136 210
rect 1170 176 1182 210
rect 1125 120 1182 176
rect 1125 86 1136 120
rect 1170 86 1182 120
rect 1292 96 1342 222
rect 1125 74 1182 86
rect 1236 84 1342 96
rect 1236 50 1264 84
rect 1298 74 1342 84
rect 1372 210 1428 222
rect 1372 176 1383 210
rect 1417 176 1428 210
rect 1372 120 1428 176
rect 1372 86 1383 120
rect 1417 86 1428 120
rect 1372 74 1428 86
rect 1458 192 1528 222
rect 1458 158 1483 192
rect 1517 158 1528 192
rect 1458 120 1528 158
rect 1458 86 1483 120
rect 1517 86 1528 120
rect 1458 74 1528 86
rect 1558 210 1614 222
rect 1558 176 1569 210
rect 1603 176 1614 210
rect 1558 120 1614 176
rect 1558 86 1569 120
rect 1603 86 1614 120
rect 1558 74 1614 86
rect 1644 192 1701 222
rect 1644 158 1655 192
rect 1689 158 1701 192
rect 1644 120 1701 158
rect 1644 86 1655 120
rect 1689 86 1701 120
rect 1644 74 1701 86
rect 1298 50 1327 74
rect 1236 38 1327 50
<< pdiff >>
rect 626 622 684 634
rect 626 592 638 622
rect 46 580 105 592
rect 46 546 58 580
rect 92 546 105 580
rect 46 497 105 546
rect 46 463 58 497
rect 92 463 105 497
rect 46 414 105 463
rect 46 380 58 414
rect 92 380 105 414
rect 46 368 105 380
rect 135 580 253 592
rect 135 546 176 580
rect 210 546 253 580
rect 135 499 253 546
rect 135 465 176 499
rect 210 465 253 499
rect 135 392 253 465
rect 283 392 337 592
rect 367 554 494 592
rect 367 520 413 554
rect 447 520 494 554
rect 367 508 494 520
rect 524 508 578 592
rect 608 588 638 592
rect 672 592 684 622
rect 672 588 702 592
rect 608 508 702 588
rect 367 392 420 508
rect 135 368 188 392
rect 649 424 702 508
rect 732 470 791 592
rect 952 590 1014 592
rect 732 436 745 470
rect 779 436 791 470
rect 732 424 791 436
rect 845 578 904 590
rect 845 544 857 578
rect 891 544 904 578
rect 845 468 904 544
rect 845 434 857 468
rect 891 434 904 468
rect 845 422 904 434
rect 934 580 1014 590
rect 934 546 964 580
rect 998 546 1014 580
rect 934 468 1014 546
rect 934 434 964 468
rect 998 434 1014 468
rect 934 422 1014 434
rect 952 368 1014 422
rect 1044 580 1111 592
rect 1044 546 1064 580
rect 1098 546 1111 580
rect 1044 497 1111 546
rect 1044 463 1064 497
rect 1098 463 1111 497
rect 1044 414 1111 463
rect 1044 380 1064 414
rect 1098 380 1111 414
rect 1044 368 1111 380
rect 1141 580 1332 592
rect 1141 546 1164 580
rect 1198 546 1275 580
rect 1309 546 1332 580
rect 1141 469 1332 546
rect 1141 435 1164 469
rect 1198 435 1275 469
rect 1309 435 1332 469
rect 1141 368 1332 435
rect 1362 580 1425 592
rect 1362 546 1375 580
rect 1409 546 1425 580
rect 1362 497 1425 546
rect 1362 463 1375 497
rect 1409 463 1425 497
rect 1362 414 1425 463
rect 1362 380 1375 414
rect 1409 380 1425 414
rect 1362 368 1425 380
rect 1455 580 1522 592
rect 1455 546 1475 580
rect 1509 546 1522 580
rect 1455 504 1522 546
rect 1455 470 1475 504
rect 1509 470 1522 504
rect 1455 428 1522 470
rect 1455 394 1475 428
rect 1509 394 1522 428
rect 1455 368 1522 394
rect 1552 580 1612 592
rect 1552 546 1565 580
rect 1599 546 1612 580
rect 1552 497 1612 546
rect 1552 463 1565 497
rect 1599 463 1612 497
rect 1552 414 1612 463
rect 1552 380 1565 414
rect 1599 380 1612 414
rect 1552 368 1612 380
rect 1642 580 1701 592
rect 1642 546 1655 580
rect 1689 546 1701 580
rect 1642 502 1701 546
rect 1642 468 1655 502
rect 1689 468 1701 502
rect 1642 424 1701 468
rect 1642 390 1655 424
rect 1689 390 1701 424
rect 1642 368 1701 390
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 130 86 164 120
rect 395 146 429 180
rect 679 136 713 170
rect 781 272 815 306
rect 872 120 906 154
rect 972 120 1006 154
rect 1136 176 1170 210
rect 1136 86 1170 120
rect 1264 50 1298 84
rect 1383 176 1417 210
rect 1383 86 1417 120
rect 1483 158 1517 192
rect 1483 86 1517 120
rect 1569 176 1603 210
rect 1569 86 1603 120
rect 1655 158 1689 192
rect 1655 86 1689 120
<< pdiffc >>
rect 58 546 92 580
rect 58 463 92 497
rect 58 380 92 414
rect 176 546 210 580
rect 176 465 210 499
rect 413 520 447 554
rect 638 588 672 622
rect 745 436 779 470
rect 857 544 891 578
rect 857 434 891 468
rect 964 546 998 580
rect 964 434 998 468
rect 1064 546 1098 580
rect 1064 463 1098 497
rect 1064 380 1098 414
rect 1164 546 1198 580
rect 1275 546 1309 580
rect 1164 435 1198 469
rect 1275 435 1309 469
rect 1375 546 1409 580
rect 1375 463 1409 497
rect 1375 380 1409 414
rect 1475 546 1509 580
rect 1475 470 1509 504
rect 1475 394 1509 428
rect 1565 546 1599 580
rect 1565 463 1599 497
rect 1565 380 1599 414
rect 1655 546 1689 580
rect 1655 468 1689 502
rect 1655 390 1689 424
<< poly >>
rect 105 592 135 618
rect 253 592 283 618
rect 337 592 367 618
rect 494 592 524 618
rect 578 592 608 618
rect 702 592 732 618
rect 494 493 524 508
rect 578 493 608 508
rect 491 476 527 493
rect 461 460 527 476
rect 461 426 477 460
rect 511 426 527 460
rect 461 410 527 426
rect 253 377 283 392
rect 337 377 367 392
rect 105 353 135 368
rect 250 360 286 377
rect 102 310 138 353
rect 220 344 286 360
rect 220 310 236 344
rect 270 310 286 344
rect 334 368 370 377
rect 334 345 527 368
rect 334 338 477 345
rect 84 294 172 310
rect 220 294 286 310
rect 461 311 477 338
rect 511 311 527 345
rect 84 260 122 294
rect 156 260 172 294
rect 84 244 172 260
rect 84 222 114 244
rect 256 208 286 294
rect 334 280 413 296
rect 334 246 363 280
rect 397 246 413 280
rect 334 230 413 246
rect 461 295 527 311
rect 334 208 364 230
rect 461 208 491 295
rect 575 288 611 493
rect 904 590 934 616
rect 1014 592 1044 618
rect 1111 592 1141 618
rect 1332 592 1362 618
rect 1425 592 1455 618
rect 1522 592 1552 618
rect 1612 592 1642 618
rect 702 409 732 424
rect 699 392 735 409
rect 904 407 934 422
rect 665 376 754 392
rect 665 342 681 376
rect 715 342 754 376
rect 665 326 754 342
rect 901 336 937 407
rect 1014 353 1044 368
rect 1111 353 1141 368
rect 1332 353 1362 368
rect 1425 353 1455 368
rect 1522 353 1552 368
rect 1612 353 1642 368
rect 1011 336 1047 353
rect 581 273 611 288
rect 724 273 754 326
rect 880 320 1047 336
rect 1108 326 1144 353
rect 1329 336 1365 353
rect 1422 336 1458 353
rect 1519 336 1555 353
rect 1609 336 1645 353
rect 461 98 491 124
rect 581 109 611 189
rect 880 286 896 320
rect 930 286 964 320
rect 998 286 1047 320
rect 880 270 1047 286
rect 931 222 961 270
rect 1017 222 1047 270
rect 1095 310 1161 326
rect 1095 276 1111 310
rect 1145 276 1161 310
rect 1095 260 1161 276
rect 1204 320 1645 336
rect 1204 286 1220 320
rect 1254 306 1645 320
rect 1254 286 1644 306
rect 1204 280 1644 286
rect 1095 222 1125 260
rect 1204 252 1270 280
rect 563 93 629 109
rect 84 48 114 74
rect 256 54 286 80
rect 334 54 364 80
rect 563 59 579 93
rect 613 59 629 93
rect 563 43 629 59
rect 724 103 754 125
rect 724 87 829 103
rect 724 53 779 87
rect 813 53 829 87
rect 1204 218 1220 252
rect 1254 218 1270 252
rect 1342 222 1372 280
rect 1428 222 1458 280
rect 1528 222 1558 280
rect 1614 222 1644 280
rect 1204 184 1270 218
rect 1204 150 1220 184
rect 1254 150 1270 184
rect 1204 134 1270 150
rect 724 37 829 53
rect 931 48 961 74
rect 1017 48 1047 74
rect 1095 48 1125 74
rect 1342 48 1372 74
rect 1428 48 1458 74
rect 1528 48 1558 74
rect 1614 48 1644 74
<< polycont >>
rect 477 426 511 460
rect 236 310 270 344
rect 477 311 511 345
rect 122 260 156 294
rect 363 246 397 280
rect 681 342 715 376
rect 896 286 930 320
rect 964 286 998 320
rect 1111 276 1145 310
rect 1220 286 1254 320
rect 579 59 613 93
rect 779 53 813 87
rect 1220 218 1254 252
rect 1220 150 1254 184
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 23 580 108 596
rect 23 546 58 580
rect 92 546 108 580
rect 23 497 108 546
rect 23 463 58 497
rect 92 463 108 497
rect 23 414 108 463
rect 157 580 232 649
rect 157 546 176 580
rect 210 546 232 580
rect 622 622 688 649
rect 622 588 638 622
rect 672 588 688 622
rect 622 572 688 588
rect 841 578 907 594
rect 157 499 232 546
rect 157 465 176 499
rect 210 465 232 499
rect 157 462 232 465
rect 287 554 497 570
rect 287 520 413 554
rect 447 520 497 554
rect 841 544 857 578
rect 891 544 907 578
rect 841 538 907 544
rect 287 504 497 520
rect 661 504 907 538
rect 287 428 321 504
rect 661 470 695 504
rect 23 380 58 414
rect 92 380 108 414
rect 23 364 108 380
rect 142 394 321 428
rect 355 460 695 470
rect 355 426 477 460
rect 511 426 695 460
rect 729 436 745 470
rect 779 436 799 470
rect 355 410 695 426
rect 23 210 73 364
rect 142 310 176 394
rect 107 294 176 310
rect 217 344 286 360
rect 217 310 236 344
rect 270 310 286 344
rect 217 306 286 310
rect 107 260 122 294
rect 156 272 176 294
rect 355 280 413 410
rect 661 392 695 410
rect 661 376 731 392
rect 156 260 321 272
rect 107 238 321 260
rect 23 176 39 210
rect 73 176 253 204
rect 23 170 253 176
rect 23 120 73 170
rect 23 86 39 120
rect 23 70 73 86
rect 110 120 185 136
rect 110 86 130 120
rect 164 86 185 120
rect 110 17 185 86
rect 219 85 253 170
rect 287 196 321 238
rect 355 246 363 280
rect 397 246 413 280
rect 461 345 527 361
rect 461 311 477 345
rect 511 311 527 345
rect 661 342 681 376
rect 715 342 731 376
rect 661 340 731 342
rect 461 306 527 311
rect 765 322 799 436
rect 841 468 907 504
rect 841 434 857 468
rect 891 434 907 468
rect 841 418 907 434
rect 948 580 1014 649
rect 948 546 964 580
rect 998 546 1014 580
rect 948 468 1014 546
rect 948 434 964 468
rect 998 434 1014 468
rect 948 418 1014 434
rect 1048 580 1114 596
rect 1048 546 1064 580
rect 1098 546 1114 580
rect 1048 497 1114 546
rect 1048 463 1064 497
rect 1098 463 1114 497
rect 1048 414 1114 463
rect 1148 580 1325 649
rect 1148 546 1164 580
rect 1198 546 1275 580
rect 1309 546 1325 580
rect 1148 469 1325 546
rect 1148 435 1164 469
rect 1198 435 1275 469
rect 1309 435 1325 469
rect 1148 432 1325 435
rect 1359 580 1425 596
rect 1359 546 1375 580
rect 1409 546 1425 580
rect 1359 497 1425 546
rect 1359 463 1375 497
rect 1409 463 1425 497
rect 1048 380 1064 414
rect 1098 398 1114 414
rect 1359 414 1425 463
rect 1098 380 1270 398
rect 1048 364 1270 380
rect 765 306 831 322
rect 461 272 781 306
rect 815 272 831 306
rect 880 320 1014 356
rect 880 286 896 320
rect 930 286 964 320
rect 998 286 1014 320
rect 880 272 1014 286
rect 1052 310 1161 326
rect 1052 276 1111 310
rect 1145 276 1161 310
rect 355 230 413 246
rect 1052 260 1161 276
rect 1195 320 1270 364
rect 1195 286 1220 320
rect 1254 286 1270 320
rect 1359 380 1375 414
rect 1409 380 1425 414
rect 1359 344 1425 380
rect 1459 580 1509 649
rect 1459 546 1475 580
rect 1459 504 1509 546
rect 1459 470 1475 504
rect 1459 428 1509 470
rect 1459 394 1475 428
rect 1459 378 1509 394
rect 1549 580 1599 596
rect 1549 546 1565 580
rect 1549 497 1599 546
rect 1549 463 1565 497
rect 1549 414 1599 463
rect 1549 380 1565 414
rect 1639 580 1705 649
rect 1639 546 1655 580
rect 1689 546 1705 580
rect 1639 502 1705 546
rect 1639 468 1655 502
rect 1689 468 1705 502
rect 1639 424 1705 468
rect 1639 390 1655 424
rect 1689 390 1705 424
rect 1549 356 1599 380
rect 1549 344 1703 356
rect 1359 310 1703 344
rect 1052 238 1086 260
rect 563 204 1086 238
rect 1195 252 1270 286
rect 1561 276 1603 310
rect 1195 226 1220 252
rect 1120 218 1220 226
rect 1254 218 1270 252
rect 1120 210 1270 218
rect 287 180 466 196
rect 287 146 395 180
rect 429 146 466 180
rect 287 130 466 146
rect 563 93 629 204
rect 1120 176 1136 210
rect 1170 184 1270 210
rect 1170 176 1220 184
rect 563 85 579 93
rect 219 59 579 85
rect 613 59 629 93
rect 219 51 629 59
rect 663 136 679 170
rect 713 136 729 170
rect 663 17 729 136
rect 856 154 922 170
rect 856 120 872 154
rect 906 120 922 154
rect 856 103 922 120
rect 763 87 922 103
rect 763 53 779 87
rect 813 53 922 87
rect 763 51 922 53
rect 956 154 1022 170
rect 956 120 972 154
rect 1006 120 1022 154
rect 956 17 1022 120
rect 1120 150 1220 176
rect 1254 150 1270 184
rect 1120 134 1270 150
rect 1367 242 1603 276
rect 1367 210 1433 242
rect 1367 176 1383 210
rect 1417 176 1433 210
rect 1553 210 1603 242
rect 1120 120 1195 134
rect 1120 86 1136 120
rect 1170 86 1195 120
rect 1367 120 1433 176
rect 1120 70 1195 86
rect 1232 84 1331 100
rect 1232 50 1264 84
rect 1298 50 1331 84
rect 1367 86 1383 120
rect 1417 86 1433 120
rect 1367 70 1433 86
rect 1467 192 1517 208
rect 1467 158 1483 192
rect 1467 120 1517 158
rect 1467 86 1483 120
rect 1232 17 1331 50
rect 1467 17 1517 86
rect 1553 176 1569 210
rect 1553 120 1603 176
rect 1553 86 1569 120
rect 1553 70 1603 86
rect 1639 192 1705 208
rect 1639 158 1655 192
rect 1689 158 1705 192
rect 1639 120 1705 158
rect 1639 86 1655 120
rect 1689 86 1705 120
rect 1639 17 1705 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
<< metal1 >>
rect 0 683 1728 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 0 617 1728 649
rect 0 17 1728 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
rect 0 -49 1728 -17
<< labels >>
flabel comment s 738 315 738 315 0 FreeSans 200 0 0 0 no_jumper_check
rlabel comment s 0 0 0 0 4 dlclkp_4
flabel pwell s 0 0 1728 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nwell s 0 617 1728 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 0 617 1728 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 1728 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 GATE
port 2 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 1567 316 1601 350 0 FreeSans 340 0 0 0 GCLK
port 7 nsew
flabel corelocali s 1663 316 1697 350 0 FreeSans 340 0 0 0 GCLK
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 1728 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2896904
string GDS_START 2883982
<< end >>
