magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 25 260 91 356
rect 193 210 263 344
rect 593 270 659 578
rect 848 364 943 596
rect 697 270 767 356
rect 909 226 943 364
rect 869 70 943 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 23 496 89 596
rect 123 530 189 649
rect 223 581 551 615
rect 223 496 257 581
rect 23 462 257 496
rect 23 420 159 462
rect 125 226 159 420
rect 230 378 331 428
rect 28 192 159 226
rect 297 340 331 378
rect 369 374 449 547
rect 297 206 381 340
rect 28 70 94 192
rect 297 176 331 206
rect 128 17 194 158
rect 228 70 331 176
rect 415 204 449 374
rect 485 238 551 581
rect 748 390 814 649
rect 801 260 875 326
rect 801 236 835 260
rect 662 204 835 236
rect 415 202 835 204
rect 415 170 728 202
rect 365 17 415 136
rect 449 70 515 170
rect 549 17 628 136
rect 662 70 728 170
rect 762 17 828 168
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
rlabel locali s 697 270 767 356 6 A
port 1 nsew signal input
rlabel locali s 593 270 659 578 6 B
port 2 nsew signal input
rlabel locali s 25 260 91 356 6 C_N
port 3 nsew signal input
rlabel locali s 193 210 263 344 6 D_N
port 4 nsew signal input
rlabel locali s 909 226 943 364 6 X
port 5 nsew signal output
rlabel locali s 869 70 943 226 6 X
port 5 nsew signal output
rlabel locali s 848 364 943 596 6 X
port 5 nsew signal output
rlabel metal1 s 0 -49 960 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 960 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 919306
string GDS_START 910970
<< end >>
