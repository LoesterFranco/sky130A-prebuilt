magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 902 704
<< pwell >>
rect 0 0 864 49
<< scnmos >>
rect 86 74 116 222
rect 223 94 253 222
rect 301 94 331 222
rect 558 74 588 202
rect 644 74 674 202
rect 750 74 780 202
<< pmoshvt >>
rect 86 368 116 592
rect 203 384 233 552
rect 304 384 334 552
rect 561 384 591 552
rect 663 384 693 584
rect 747 384 777 584
<< ndiff >>
rect 29 210 86 222
rect 29 176 41 210
rect 75 176 86 210
rect 29 120 86 176
rect 29 86 41 120
rect 75 86 86 120
rect 29 74 86 86
rect 116 182 223 222
rect 116 148 174 182
rect 208 148 223 182
rect 116 116 223 148
rect 116 82 127 116
rect 161 94 223 116
rect 253 94 301 222
rect 331 189 388 222
rect 331 155 342 189
rect 376 155 388 189
rect 331 94 388 155
rect 501 184 558 202
rect 501 150 513 184
rect 547 150 558 184
rect 501 116 558 150
rect 161 82 187 94
rect 116 74 187 82
rect 501 82 513 116
rect 547 82 558 116
rect 501 74 558 82
rect 588 186 644 202
rect 588 152 599 186
rect 633 152 644 186
rect 588 118 644 152
rect 588 84 599 118
rect 633 84 644 118
rect 588 74 644 84
rect 674 127 750 202
rect 674 93 699 127
rect 733 93 750 127
rect 674 74 750 93
rect 780 186 837 202
rect 780 152 791 186
rect 825 152 837 186
rect 780 118 837 152
rect 780 84 791 118
rect 825 84 837 118
rect 780 74 837 84
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 497 86 546
rect 27 463 39 497
rect 73 463 86 497
rect 27 414 86 463
rect 27 380 39 414
rect 73 380 86 414
rect 27 368 86 380
rect 116 580 185 592
rect 116 546 139 580
rect 173 552 185 580
rect 610 552 663 584
rect 173 546 203 552
rect 116 500 203 546
rect 116 466 139 500
rect 173 466 203 500
rect 116 426 203 466
rect 116 392 139 426
rect 173 392 203 426
rect 116 384 203 392
rect 233 440 304 552
rect 233 406 246 440
rect 280 406 304 440
rect 233 384 304 406
rect 334 533 561 552
rect 334 499 347 533
rect 381 499 430 533
rect 464 499 514 533
rect 548 499 561 533
rect 334 384 561 499
rect 591 540 663 552
rect 591 506 614 540
rect 648 506 663 540
rect 591 430 663 506
rect 591 396 614 430
rect 648 396 663 430
rect 591 384 663 396
rect 693 384 747 584
rect 777 572 836 584
rect 777 538 790 572
rect 824 538 836 572
rect 777 501 836 538
rect 777 467 790 501
rect 824 467 836 501
rect 777 430 836 467
rect 777 396 790 430
rect 824 396 836 430
rect 777 384 836 396
rect 116 368 169 384
<< ndiffc >>
rect 41 176 75 210
rect 41 86 75 120
rect 174 148 208 182
rect 127 82 161 116
rect 342 155 376 189
rect 513 150 547 184
rect 513 82 547 116
rect 599 152 633 186
rect 599 84 633 118
rect 699 93 733 127
rect 791 152 825 186
rect 791 84 825 118
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 139 546 173 580
rect 139 466 173 500
rect 139 392 173 426
rect 246 406 280 440
rect 347 499 381 533
rect 430 499 464 533
rect 514 499 548 533
rect 614 506 648 540
rect 614 396 648 430
rect 790 538 824 572
rect 790 467 824 501
rect 790 396 824 430
<< poly >>
rect 86 592 116 618
rect 663 584 693 610
rect 747 584 777 610
rect 203 552 233 578
rect 304 552 334 578
rect 561 552 591 578
rect 203 369 233 384
rect 304 369 334 384
rect 561 369 591 384
rect 663 369 693 384
rect 747 369 777 384
rect 86 353 116 368
rect 83 326 119 353
rect 200 342 236 369
rect 301 352 337 369
rect 193 326 259 342
rect 83 310 151 326
rect 83 276 101 310
rect 135 276 151 310
rect 83 260 151 276
rect 193 292 209 326
rect 243 292 259 326
rect 193 270 259 292
rect 301 336 367 352
rect 301 302 317 336
rect 351 302 367 336
rect 301 286 367 302
rect 410 336 476 352
rect 410 302 426 336
rect 460 302 476 336
rect 86 222 116 260
rect 223 222 253 270
rect 301 222 331 286
rect 410 268 476 302
rect 410 234 426 268
rect 460 248 476 268
rect 558 350 591 369
rect 558 248 588 350
rect 660 302 696 369
rect 747 350 780 369
rect 750 302 780 350
rect 460 234 588 248
rect 636 286 702 302
rect 636 252 652 286
rect 686 252 702 286
rect 636 236 702 252
rect 750 286 843 302
rect 750 252 793 286
rect 827 252 843 286
rect 750 236 843 252
rect 410 218 588 234
rect 558 202 588 218
rect 644 202 674 236
rect 750 202 780 236
rect 86 48 116 74
rect 223 68 253 94
rect 301 68 331 94
rect 558 48 588 74
rect 644 48 674 74
rect 750 48 780 74
<< polycont >>
rect 101 276 135 310
rect 209 292 243 326
rect 317 302 351 336
rect 426 302 460 336
rect 426 234 460 268
rect 652 252 686 286
rect 793 252 827 286
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 17 580 89 596
rect 17 546 39 580
rect 73 546 89 580
rect 17 497 89 546
rect 17 463 39 497
rect 73 463 89 497
rect 17 414 89 463
rect 17 380 39 414
rect 73 380 89 414
rect 123 580 189 649
rect 123 546 139 580
rect 173 546 189 580
rect 123 500 189 546
rect 123 466 139 500
rect 173 466 189 500
rect 331 533 564 649
rect 774 572 840 649
rect 331 499 347 533
rect 381 499 430 533
rect 464 499 514 533
rect 548 499 564 533
rect 331 490 564 499
rect 598 540 664 556
rect 598 506 614 540
rect 648 506 664 540
rect 123 426 189 466
rect 123 392 139 426
rect 173 392 189 426
rect 123 390 189 392
rect 230 440 476 456
rect 230 406 246 440
rect 280 406 476 440
rect 598 430 664 506
rect 598 414 614 430
rect 230 390 476 406
rect 17 364 89 380
rect 17 226 51 364
rect 217 342 263 356
rect 193 326 263 342
rect 85 310 159 326
rect 85 276 101 310
rect 135 276 159 310
rect 193 292 209 326
rect 243 292 263 326
rect 193 284 263 292
rect 301 336 367 356
rect 301 302 317 336
rect 351 302 367 336
rect 301 286 367 302
rect 410 336 476 390
rect 410 302 426 336
rect 460 302 476 336
rect 85 260 159 276
rect 125 250 159 260
rect 410 268 476 302
rect 410 252 426 268
rect 17 210 91 226
rect 125 216 292 250
rect 17 176 41 210
rect 75 176 91 210
rect 17 120 91 176
rect 17 86 41 120
rect 75 86 91 120
rect 17 70 91 86
rect 125 148 174 182
rect 208 148 224 182
rect 125 116 224 148
rect 125 82 127 116
rect 161 82 224 116
rect 125 17 224 82
rect 258 85 292 216
rect 326 234 426 252
rect 460 234 476 268
rect 326 218 476 234
rect 529 396 614 414
rect 648 396 664 430
rect 529 380 664 396
rect 774 538 790 572
rect 824 538 840 572
rect 774 501 840 538
rect 774 467 790 501
rect 824 467 840 501
rect 774 430 840 467
rect 774 396 790 430
rect 824 396 840 430
rect 774 380 840 396
rect 326 189 376 218
rect 326 155 342 189
rect 529 184 563 380
rect 601 286 743 302
rect 601 252 652 286
rect 686 252 743 286
rect 601 236 743 252
rect 777 286 843 302
rect 777 252 793 286
rect 827 252 843 286
rect 777 236 843 252
rect 326 119 376 155
rect 497 150 513 184
rect 547 150 563 184
rect 497 116 563 150
rect 497 85 513 116
rect 258 82 513 85
rect 547 82 563 116
rect 258 51 563 82
rect 599 186 841 202
rect 633 168 791 186
rect 633 152 649 168
rect 599 118 649 152
rect 825 152 841 186
rect 633 84 649 118
rect 599 68 649 84
rect 683 127 749 134
rect 683 93 699 127
rect 733 93 749 127
rect 683 17 749 93
rect 791 118 841 152
rect 825 84 841 118
rect 791 68 841 84
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o2bb2a_1
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 607 242 641 276 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 703 242 737 276 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A2_N
port 2 nsew
flabel corelocali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 799 242 833 276 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A1_N
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 864 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1550420
string GDS_START 1542546
<< end >>
