magic
tech sky130A
magscale 1 2
timestamp 1599588232
<< locali >>
rect 21 192 74 430
rect 291 236 353 330
rect 2121 364 2191 596
rect 2157 230 2191 364
rect 2118 88 2191 230
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 22 504 88 649
rect 128 470 174 596
rect 208 504 274 649
rect 414 504 480 649
rect 634 470 684 547
rect 108 436 684 470
rect 724 436 815 547
rect 892 462 958 649
rect 108 158 142 436
rect 303 364 433 402
rect 176 350 257 356
rect 176 316 223 350
rect 176 249 257 316
rect 387 202 433 364
rect 29 70 142 158
rect 209 17 259 162
rect 295 133 433 202
rect 467 145 501 436
rect 775 428 815 436
rect 994 428 1060 547
rect 1098 472 1164 649
rect 1198 428 1340 596
rect 1374 541 1520 573
rect 1374 507 1580 541
rect 535 249 741 402
rect 535 165 588 249
rect 467 141 507 145
rect 467 137 510 141
rect 295 70 361 133
rect 467 131 515 137
rect 623 131 673 215
rect 467 125 673 131
rect 471 121 673 125
rect 474 119 673 121
rect 479 113 673 119
rect 482 109 673 113
rect 483 105 673 109
rect 488 97 673 105
rect 707 93 741 249
rect 775 394 1139 428
rect 775 127 815 394
rect 855 260 931 355
rect 971 350 1031 360
rect 971 316 991 350
rect 1025 316 1031 350
rect 971 294 1031 316
rect 1067 294 1139 394
rect 1173 394 1340 428
rect 1173 260 1207 394
rect 1462 360 1512 473
rect 1241 326 1512 360
rect 1241 294 1302 326
rect 855 226 1239 260
rect 1350 259 1484 291
rect 937 158 1139 192
rect 937 93 971 158
rect 404 17 451 93
rect 707 51 971 93
rect 1005 17 1071 124
rect 1105 85 1139 158
rect 1173 119 1239 226
rect 1273 225 1484 259
rect 1546 259 1580 507
rect 1628 504 1694 649
rect 1736 467 1802 596
rect 1842 504 1892 649
rect 1614 427 1810 467
rect 1930 461 1996 596
rect 1614 393 1912 427
rect 1657 350 1742 359
rect 1657 316 1663 350
rect 1697 316 1742 350
rect 1657 293 1742 316
rect 1784 259 1844 359
rect 1546 225 1844 259
rect 1273 85 1307 225
rect 1546 191 1580 225
rect 1878 191 1912 393
rect 1341 125 1580 191
rect 1105 51 1307 85
rect 1623 17 1711 181
rect 1809 115 1912 191
rect 1946 330 1996 461
rect 2030 420 2080 649
rect 1946 264 2123 330
rect 1946 106 1996 264
rect 2032 17 2082 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 223 316 257 350
rect 991 316 1025 350
rect 1663 316 1697 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
<< metal1 >>
rect 0 683 2208 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 0 617 2208 649
rect 0 616 50 617
rect 211 350 269 356
rect 211 316 223 350
rect 257 347 269 350
rect 979 350 1037 356
rect 979 347 991 350
rect 257 319 991 347
rect 257 316 269 319
rect 211 310 269 316
rect 979 316 991 319
rect 1025 347 1037 350
rect 1651 350 1709 356
rect 1651 347 1663 350
rect 1025 319 1663 347
rect 1025 316 1037 319
rect 979 310 1037 316
rect 1651 316 1663 319
rect 1697 316 1709 350
rect 1651 310 1709 316
rect 0 49 50 50
rect 0 17 2208 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
rect 0 -49 2208 -17
<< labels >>
rlabel locali s 21 192 74 430 6 D
port 1 nsew signal input
rlabel locali s 2157 230 2191 364 6 Q
port 2 nsew signal output
rlabel locali s 2121 364 2191 596 6 Q
port 2 nsew signal output
rlabel locali s 2118 88 2191 230 6 Q
port 2 nsew signal output
rlabel metal1 s 1651 347 1709 356 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 1651 310 1709 319 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 979 347 1037 356 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 979 310 1037 319 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 211 347 269 356 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 211 319 1709 347 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 211 310 269 319 6 RESET_B
port 3 nsew signal input
rlabel locali s 291 236 353 330 6 CLK_N
port 4 nsew clock input
rlabel metal1 s 0 -49 2208 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 6 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 617 2208 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2208 666
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 2976988
string GDS_START 2960264
<< end >>
