magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 1694 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 79 47 109 177
rect 173 47 203 177
rect 267 47 297 177
rect 371 47 401 177
rect 455 47 485 177
rect 549 47 579 177
rect 757 47 787 177
rect 851 47 881 177
rect 935 47 965 177
rect 1029 47 1059 177
rect 1256 47 1286 177
rect 1350 47 1380 177
rect 1443 47 1473 177
rect 1537 47 1567 177
<< pmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 457 297 493 497
rect 551 297 587 497
rect 749 297 785 497
rect 843 297 879 497
rect 937 297 973 497
rect 1031 297 1067 497
rect 1257 297 1293 497
rect 1351 297 1387 497
rect 1445 297 1481 497
rect 1539 297 1575 497
<< ndiff >>
rect 27 93 79 177
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 101 173 177
rect 109 67 129 101
rect 163 67 173 101
rect 109 47 173 67
rect 203 93 267 177
rect 203 59 223 93
rect 257 59 267 93
rect 203 47 267 59
rect 297 101 371 177
rect 297 67 317 101
rect 351 67 371 101
rect 297 47 371 67
rect 401 93 455 177
rect 401 59 411 93
rect 445 59 455 93
rect 401 47 455 59
rect 485 101 549 177
rect 485 67 505 101
rect 539 67 549 101
rect 485 47 549 67
rect 579 93 641 177
rect 579 59 599 93
rect 633 59 641 93
rect 579 47 641 59
rect 695 93 757 177
rect 695 59 703 93
rect 737 59 757 93
rect 695 47 757 59
rect 787 165 851 177
rect 787 131 797 165
rect 831 131 851 165
rect 787 47 851 131
rect 881 93 935 177
rect 881 59 891 93
rect 925 59 935 93
rect 881 47 935 59
rect 965 161 1029 177
rect 965 127 985 161
rect 1019 127 1029 161
rect 965 47 1029 127
rect 1059 93 1121 177
rect 1059 59 1079 93
rect 1113 59 1121 93
rect 1059 47 1121 59
rect 1194 93 1256 177
rect 1194 59 1202 93
rect 1236 59 1256 93
rect 1194 47 1256 59
rect 1286 161 1350 177
rect 1286 127 1296 161
rect 1330 127 1350 161
rect 1286 47 1350 127
rect 1380 101 1443 177
rect 1380 67 1399 101
rect 1433 67 1443 101
rect 1380 47 1443 67
rect 1473 93 1537 177
rect 1473 59 1493 93
rect 1527 59 1537 93
rect 1473 47 1537 59
rect 1567 101 1629 177
rect 1567 67 1587 101
rect 1621 67 1629 101
rect 1567 47 1629 67
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 297 81 383
rect 117 477 175 497
rect 117 443 129 477
rect 163 443 175 477
rect 117 409 175 443
rect 117 375 129 409
rect 163 375 175 409
rect 117 297 175 375
rect 211 485 269 497
rect 211 451 223 485
rect 257 451 269 485
rect 211 417 269 451
rect 211 383 223 417
rect 257 383 269 417
rect 211 297 269 383
rect 305 477 363 497
rect 305 443 317 477
rect 351 443 363 477
rect 305 409 363 443
rect 305 375 317 409
rect 351 375 363 409
rect 305 297 363 375
rect 399 485 457 497
rect 399 451 411 485
rect 445 451 457 485
rect 399 417 457 451
rect 399 383 411 417
rect 445 383 457 417
rect 399 297 457 383
rect 493 477 551 497
rect 493 443 505 477
rect 539 443 551 477
rect 493 297 551 443
rect 587 485 641 497
rect 587 451 599 485
rect 633 451 641 485
rect 587 297 641 451
rect 695 477 749 497
rect 695 443 703 477
rect 737 443 749 477
rect 695 297 749 443
rect 785 485 843 497
rect 785 451 797 485
rect 831 451 843 485
rect 785 297 843 451
rect 879 477 937 497
rect 879 443 891 477
rect 925 443 937 477
rect 879 297 937 443
rect 973 485 1031 497
rect 973 451 985 485
rect 1019 451 1031 485
rect 973 297 1031 451
rect 1067 485 1257 497
rect 1067 451 1211 485
rect 1245 451 1257 485
rect 1067 297 1257 451
rect 1293 417 1351 497
rect 1293 383 1305 417
rect 1339 383 1351 417
rect 1293 297 1351 383
rect 1387 485 1445 497
rect 1387 451 1399 485
rect 1433 451 1445 485
rect 1387 297 1445 451
rect 1481 417 1539 497
rect 1481 383 1493 417
rect 1527 383 1539 417
rect 1481 297 1539 383
rect 1575 485 1629 497
rect 1575 451 1587 485
rect 1621 451 1629 485
rect 1575 401 1629 451
rect 1575 367 1587 401
rect 1621 367 1629 401
rect 1575 297 1629 367
<< ndiffc >>
rect 35 59 69 93
rect 129 67 163 101
rect 223 59 257 93
rect 317 67 351 101
rect 411 59 445 93
rect 505 67 539 101
rect 599 59 633 93
rect 703 59 737 93
rect 797 131 831 165
rect 891 59 925 93
rect 985 127 1019 161
rect 1079 59 1113 93
rect 1202 59 1236 93
rect 1296 127 1330 161
rect 1399 67 1433 101
rect 1493 59 1527 93
rect 1587 67 1621 101
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 129 443 163 477
rect 129 375 163 409
rect 223 451 257 485
rect 223 383 257 417
rect 317 443 351 477
rect 317 375 351 409
rect 411 451 445 485
rect 411 383 445 417
rect 505 443 539 477
rect 599 451 633 485
rect 703 443 737 477
rect 797 451 831 485
rect 891 443 925 477
rect 985 451 1019 485
rect 1211 451 1245 485
rect 1305 383 1339 417
rect 1399 451 1433 485
rect 1493 383 1527 417
rect 1587 451 1621 485
rect 1587 367 1621 401
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 457 497 493 523
rect 551 497 587 523
rect 749 497 785 523
rect 843 497 879 523
rect 937 497 973 523
rect 1031 497 1067 523
rect 1257 497 1293 523
rect 1351 497 1387 523
rect 1445 497 1481 523
rect 1539 497 1575 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 457 282 493 297
rect 551 282 587 297
rect 749 282 785 297
rect 843 282 879 297
rect 937 282 973 297
rect 1031 282 1067 297
rect 1257 282 1293 297
rect 1351 282 1387 297
rect 1445 282 1481 297
rect 1539 282 1575 297
rect 79 265 119 282
rect 173 265 213 282
rect 267 265 307 282
rect 361 265 401 282
rect 79 249 401 265
rect 79 215 124 249
rect 158 215 198 249
rect 232 215 282 249
rect 316 215 401 249
rect 79 199 401 215
rect 79 177 109 199
rect 173 177 203 199
rect 267 177 297 199
rect 371 177 401 199
rect 455 265 495 282
rect 549 265 589 282
rect 747 269 787 282
rect 841 269 881 282
rect 455 261 602 265
rect 455 249 636 261
rect 747 259 881 269
rect 455 215 508 249
rect 542 215 576 249
rect 610 215 636 249
rect 455 203 636 215
rect 727 249 881 259
rect 727 215 743 249
rect 777 215 821 249
rect 855 215 881 249
rect 727 205 881 215
rect 455 199 612 203
rect 757 199 881 205
rect 455 177 485 199
rect 549 177 579 199
rect 757 177 787 199
rect 851 177 881 199
rect 935 269 975 282
rect 1029 269 1069 282
rect 935 261 1069 269
rect 1255 265 1295 282
rect 1349 265 1389 282
rect 935 249 1115 261
rect 1255 259 1389 265
rect 935 215 987 249
rect 1021 215 1055 249
rect 1089 215 1115 249
rect 935 205 1115 215
rect 1235 249 1389 259
rect 1235 215 1251 249
rect 1285 215 1329 249
rect 1363 215 1389 249
rect 1235 205 1389 215
rect 1443 265 1483 282
rect 1537 265 1577 282
rect 1443 261 1577 265
rect 1443 249 1634 261
rect 1443 215 1506 249
rect 1540 215 1584 249
rect 1618 215 1634 249
rect 1443 205 1634 215
rect 935 177 965 205
rect 1029 203 1115 205
rect 1029 177 1059 203
rect 1256 177 1286 205
rect 1350 177 1380 205
rect 1443 177 1473 205
rect 1537 177 1567 205
rect 79 21 109 47
rect 173 21 203 47
rect 267 21 297 47
rect 371 21 401 47
rect 455 21 485 47
rect 549 21 579 47
rect 757 21 787 47
rect 851 21 881 47
rect 935 21 965 47
rect 1029 21 1059 47
rect 1256 21 1286 47
rect 1350 21 1380 47
rect 1443 21 1473 47
rect 1537 21 1567 47
<< polycont >>
rect 124 215 158 249
rect 198 215 232 249
rect 282 215 316 249
rect 508 215 542 249
rect 576 215 610 249
rect 743 215 777 249
rect 821 215 855 249
rect 987 215 1021 249
rect 1055 215 1089 249
rect 1251 215 1285 249
rect 1329 215 1363 249
rect 1506 215 1540 249
rect 1584 215 1618 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 19 485 85 527
rect 19 451 35 485
rect 69 451 85 485
rect 19 417 85 451
rect 19 383 35 417
rect 69 383 85 417
rect 129 477 163 493
rect 129 409 163 443
rect 197 485 273 527
rect 197 451 223 485
rect 257 451 273 485
rect 197 417 273 451
rect 197 383 223 417
rect 257 383 273 417
rect 317 477 351 493
rect 317 409 351 443
rect 129 333 163 375
rect 385 485 461 527
rect 385 451 411 485
rect 445 451 461 485
rect 385 417 461 451
rect 385 383 411 417
rect 445 383 461 417
rect 505 477 539 493
rect 573 485 649 527
rect 573 451 599 485
rect 633 451 649 485
rect 703 477 737 493
rect 505 417 539 443
rect 771 485 847 527
rect 771 451 797 485
rect 831 451 847 485
rect 891 477 925 493
rect 703 417 737 443
rect 959 485 1035 527
rect 959 451 985 485
rect 1019 451 1035 485
rect 1079 451 1211 485
rect 1245 451 1399 485
rect 1433 451 1587 485
rect 1621 451 1637 485
rect 891 417 925 443
rect 1079 417 1113 451
rect 505 383 1113 417
rect 1289 415 1305 417
rect 1156 383 1305 415
rect 1339 383 1493 417
rect 1527 383 1543 417
rect 1587 401 1637 451
rect 317 333 351 375
rect 1156 381 1302 383
rect 1156 333 1190 381
rect 1621 367 1637 401
rect 1587 351 1637 367
rect 24 299 351 333
rect 390 299 1190 333
rect 24 161 68 299
rect 390 265 434 299
rect 124 249 434 265
rect 158 215 198 249
rect 232 215 282 249
rect 316 215 434 249
rect 482 249 681 259
rect 482 215 508 249
rect 542 215 576 249
rect 610 215 681 249
rect 727 249 886 265
rect 727 215 743 249
rect 777 215 821 249
rect 855 215 886 249
rect 936 249 1115 265
rect 936 215 987 249
rect 1021 215 1055 249
rect 1089 215 1115 249
rect 124 199 434 215
rect 24 127 351 161
rect 129 101 163 127
rect 19 59 35 93
rect 69 59 85 93
rect 19 17 85 59
rect 317 101 351 127
rect 129 51 163 67
rect 197 59 223 93
rect 257 59 273 93
rect 197 17 273 59
rect 505 131 797 165
rect 831 131 847 165
rect 1156 161 1190 299
rect 1224 249 1428 325
rect 1224 215 1251 249
rect 1285 215 1329 249
rect 1363 215 1428 249
rect 1488 259 1527 327
rect 1488 249 1634 259
rect 1488 215 1506 249
rect 1540 215 1584 249
rect 1618 215 1634 249
rect 505 101 539 131
rect 959 127 985 161
rect 1019 127 1296 161
rect 1330 127 1347 161
rect 1399 129 1621 163
rect 317 51 351 67
rect 385 59 411 93
rect 445 59 461 93
rect 385 17 461 59
rect 1399 101 1433 129
rect 505 51 539 67
rect 573 59 599 93
rect 633 59 649 93
rect 687 59 703 93
rect 737 59 891 93
rect 925 59 1079 93
rect 1113 59 1129 93
rect 1186 59 1202 93
rect 1236 67 1399 93
rect 1587 101 1621 129
rect 1236 59 1433 67
rect 573 17 649 59
rect 1399 51 1433 59
rect 1467 59 1493 93
rect 1527 59 1543 93
rect 1467 17 1543 59
rect 1587 51 1621 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
<< metal1 >>
rect 0 561 1656 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 0 496 1656 527
rect 0 17 1656 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
rect 0 -48 1656 -17
<< labels >>
flabel corelocali s 491 221 525 255 0 FreeSans 200 0 0 0 A3
port 3 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 200 0 0 0 X
port 10 nsew
flabel corelocali s 30 289 64 323 0 FreeSans 200 0 0 0 X
port 10 nsew
flabel corelocali s 30 153 64 187 0 FreeSans 200 0 0 0 X
port 10 nsew
flabel corelocali s 1393 289 1427 323 0 FreeSans 200 0 0 0 B1
port 4 nsew
flabel corelocali s 1393 221 1427 255 0 FreeSans 200 0 0 0 B1
port 4 nsew
flabel corelocali s 1490 221 1524 255 0 FreeSans 200 0 0 0 B2
port 5 nsew
flabel corelocali s 1307 306 1307 306 0 FreeSans 200 0 0 0 B1
port 4 nsew
flabel corelocali s 1044 221 1078 255 0 FreeSans 200 0 0 0 A1
port 1 nsew
flabel corelocali s 1307 238 1307 238 0 FreeSans 200 0 0 0 B1
port 4 nsew
flabel corelocali s 1490 289 1524 323 0 FreeSans 200 0 0 0 B2
port 5 nsew
flabel corelocali s 1583 238 1583 238 0 FreeSans 200 0 0 0 B2
port 5 nsew
flabel corelocali s 807 221 841 255 0 FreeSans 200 0 0 0 A2
port 2 nsew
flabel corelocali s 583 221 617 255 0 FreeSans 200 0 0 0 A3
port 3 nsew
flabel corelocali s 950 221 984 255 0 FreeSans 200 0 0 0 A1
port 1 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 1656 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1444274
string GDS_START 1432108
<< end >>
