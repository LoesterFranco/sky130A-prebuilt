magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 614 704
<< pwell >>
rect 0 0 576 49
<< scnmos >>
rect 84 74 114 222
rect 170 74 200 222
rect 362 74 392 222
rect 452 74 482 222
<< pmoshvt >>
rect 89 368 119 592
rect 173 368 203 592
rect 287 368 317 592
rect 455 368 485 592
<< ndiff >>
rect 27 202 84 222
rect 27 168 39 202
rect 73 168 84 202
rect 27 120 84 168
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 210 170 222
rect 114 176 125 210
rect 159 176 170 210
rect 114 120 170 176
rect 114 86 125 120
rect 159 86 170 120
rect 114 74 170 86
rect 200 90 362 222
rect 200 74 227 90
rect 215 56 227 74
rect 261 56 301 90
rect 335 74 362 90
rect 392 131 452 222
rect 392 97 403 131
rect 437 97 452 131
rect 392 74 452 97
rect 482 210 549 222
rect 482 176 503 210
rect 537 176 549 210
rect 482 120 549 176
rect 482 86 503 120
rect 537 86 549 120
rect 482 74 549 86
rect 335 56 347 74
rect 215 44 347 56
<< pdiff >>
rect 30 580 89 592
rect 30 546 42 580
rect 76 546 89 580
rect 30 497 89 546
rect 30 463 42 497
rect 76 463 89 497
rect 30 414 89 463
rect 30 380 42 414
rect 76 380 89 414
rect 30 368 89 380
rect 119 368 173 592
rect 203 368 287 592
rect 317 580 455 592
rect 317 546 330 580
rect 364 546 408 580
rect 442 546 455 580
rect 317 510 455 546
rect 317 476 330 510
rect 364 476 408 510
rect 442 476 455 510
rect 317 440 455 476
rect 317 406 330 440
rect 364 406 408 440
rect 442 406 455 440
rect 317 368 455 406
rect 485 580 544 592
rect 485 546 498 580
rect 532 546 544 580
rect 485 510 544 546
rect 485 476 498 510
rect 532 476 544 510
rect 485 440 544 476
rect 485 406 498 440
rect 532 406 544 440
rect 485 368 544 406
<< ndiffc >>
rect 39 168 73 202
rect 39 86 73 120
rect 125 176 159 210
rect 125 86 159 120
rect 227 56 261 90
rect 301 56 335 90
rect 403 97 437 131
rect 503 176 537 210
rect 503 86 537 120
<< pdiffc >>
rect 42 546 76 580
rect 42 463 76 497
rect 42 380 76 414
rect 330 546 364 580
rect 408 546 442 580
rect 330 476 364 510
rect 408 476 442 510
rect 330 406 364 440
rect 408 406 442 440
rect 498 546 532 580
rect 498 476 532 510
rect 498 406 532 440
<< poly >>
rect 89 592 119 618
rect 173 592 203 618
rect 287 592 317 618
rect 455 592 485 618
rect 89 353 119 368
rect 173 353 203 368
rect 287 353 317 368
rect 455 353 485 368
rect 86 310 122 353
rect 21 294 122 310
rect 21 260 37 294
rect 71 280 122 294
rect 170 326 206 353
rect 284 336 320 353
rect 170 310 236 326
rect 71 260 114 280
rect 21 244 114 260
rect 84 222 114 244
rect 170 276 186 310
rect 220 276 236 310
rect 284 320 404 336
rect 284 306 354 320
rect 170 260 236 276
rect 338 286 354 306
rect 388 286 404 320
rect 338 270 404 286
rect 452 326 488 353
rect 452 310 555 326
rect 452 276 505 310
rect 539 276 555 310
rect 170 222 200 260
rect 362 222 392 270
rect 452 260 555 276
rect 452 222 482 260
rect 84 48 114 74
rect 170 48 200 74
rect 362 48 392 74
rect 452 48 482 74
<< polycont >>
rect 37 260 71 294
rect 186 276 220 310
rect 354 286 388 320
rect 505 276 539 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 26 580 76 649
rect 26 546 42 580
rect 270 580 446 596
rect 26 497 76 546
rect 26 463 42 497
rect 26 414 76 463
rect 26 380 42 414
rect 26 364 76 380
rect 121 310 236 578
rect 21 294 87 310
rect 21 260 37 294
rect 71 260 87 294
rect 121 276 186 310
rect 220 276 236 310
rect 121 260 236 276
rect 270 546 330 580
rect 364 546 408 580
rect 442 546 446 580
rect 270 510 446 546
rect 270 476 330 510
rect 364 476 408 510
rect 442 476 446 510
rect 270 440 446 476
rect 270 406 330 440
rect 364 406 408 440
rect 442 406 446 440
rect 270 390 446 406
rect 482 580 548 649
rect 482 546 498 580
rect 532 546 548 580
rect 482 510 548 546
rect 482 476 498 510
rect 532 476 548 510
rect 482 440 548 476
rect 482 406 498 440
rect 532 406 548 440
rect 482 390 548 406
rect 21 236 87 260
rect 270 226 304 390
rect 338 320 455 356
rect 338 286 354 320
rect 388 286 455 320
rect 338 270 455 286
rect 489 310 555 356
rect 489 276 505 310
rect 539 276 555 310
rect 489 260 555 276
rect 125 210 175 226
rect 23 168 39 202
rect 73 168 89 202
rect 23 120 89 168
rect 23 86 39 120
rect 73 86 89 120
rect 23 17 89 86
rect 159 176 175 210
rect 270 210 553 226
rect 270 192 503 210
rect 125 158 175 176
rect 487 176 503 192
rect 537 176 553 210
rect 125 131 453 158
rect 125 124 403 131
rect 125 120 175 124
rect 159 86 175 120
rect 387 97 403 124
rect 437 97 453 131
rect 125 70 175 86
rect 211 56 227 90
rect 261 56 301 90
rect 335 56 351 90
rect 387 70 453 97
rect 487 120 553 176
rect 487 86 503 120
rect 537 86 553 120
rect 487 70 553 86
rect 211 17 351 56
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o31ai_1
flabel pwell s 0 0 576 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nwell s 0 617 576 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 576 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 576 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 127 390 161 424 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 127 464 161 498 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 127 538 161 572 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 B1
port 4 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 319 464 353 498 0 FreeSans 340 0 0 0 Y
port 9 nsew
flabel corelocali s 319 538 353 572 0 FreeSans 340 0 0 0 Y
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 576 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 814634
string GDS_START 808462
<< end >>
