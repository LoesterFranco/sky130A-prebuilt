magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1104 561
rect 103 427 169 527
rect 17 197 66 325
rect 103 17 169 93
rect 391 367 449 527
rect 755 435 819 527
rect 287 191 353 265
rect 944 314 1001 527
rect 1035 334 1087 491
rect 1053 149 1087 334
rect 375 17 441 89
rect 755 17 809 109
rect 951 17 996 143
rect 1035 83 1087 149
rect 0 -17 1104 17
<< obsli1 >>
rect 35 393 69 493
rect 35 359 156 393
rect 122 323 156 359
rect 122 280 156 289
rect 203 391 248 493
rect 203 357 214 391
rect 203 337 248 357
rect 122 214 168 280
rect 122 161 156 214
rect 35 127 156 161
rect 35 69 69 127
rect 203 69 237 337
rect 286 333 357 483
rect 549 451 721 485
rect 659 421 721 451
rect 659 418 724 421
rect 678 417 724 418
rect 678 413 726 417
rect 678 409 729 413
rect 681 407 729 409
rect 686 402 729 407
rect 489 391 556 401
rect 523 357 556 391
rect 286 299 423 333
rect 389 247 423 299
rect 489 271 556 357
rect 590 323 657 382
rect 624 312 657 323
rect 624 289 653 312
rect 691 290 729 402
rect 859 373 908 487
rect 763 307 908 373
rect 389 157 464 247
rect 590 208 653 289
rect 302 153 464 157
rect 302 123 423 153
rect 512 147 653 208
rect 687 265 729 290
rect 874 265 908 307
rect 687 199 840 265
rect 874 199 1019 265
rect 302 69 341 123
rect 687 107 721 199
rect 874 144 908 199
rect 553 73 721 107
rect 859 52 908 144
<< obsli1c >>
rect 122 289 156 323
rect 214 357 248 391
rect 489 357 523 391
rect 590 289 624 323
<< metal1 >>
rect 0 496 1104 592
rect 0 -48 1104 48
<< obsm1 >>
rect 202 391 260 397
rect 202 357 214 391
rect 248 388 260 391
rect 477 391 535 397
rect 477 388 489 391
rect 248 360 489 388
rect 248 357 260 360
rect 202 351 260 357
rect 477 357 489 360
rect 523 357 535 391
rect 477 351 535 357
rect 110 323 168 329
rect 110 289 122 323
rect 156 320 168 323
rect 578 323 636 329
rect 578 320 590 323
rect 156 292 590 320
rect 156 289 168 292
rect 110 283 168 289
rect 578 289 590 292
rect 624 289 636 323
rect 578 283 636 289
<< labels >>
rlabel locali s 287 191 353 265 6 D
port 1 nsew signal input
rlabel locali s 1053 149 1087 334 6 Q
port 2 nsew signal output
rlabel locali s 1035 334 1087 491 6 Q
port 2 nsew signal output
rlabel locali s 1035 83 1087 149 6 Q
port 2 nsew signal output
rlabel locali s 17 197 66 325 6 GATE_N
port 3 nsew clock input
rlabel locali s 951 17 996 143 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 755 17 809 109 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 375 17 441 89 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 103 17 169 93 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 1104 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1104 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 944 314 1001 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 755 435 819 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 391 367 449 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 103 427 169 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 1104 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 1104 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1104 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2774062
string GDS_START 2763460
<< end >>
