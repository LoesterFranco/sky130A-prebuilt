magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 22 289 419 323
rect 22 215 128 289
rect 171 215 289 255
rect 343 215 419 289
rect 489 181 555 425
rect 695 215 894 255
rect 944 215 1087 255
rect 197 145 555 181
rect 197 129 273 145
rect 479 51 555 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 27 391 77 493
rect 121 427 171 527
rect 215 391 265 493
rect 309 427 359 527
rect 403 459 641 493
rect 403 391 453 459
rect 27 357 453 391
rect 591 359 641 459
rect 695 393 745 493
rect 789 427 839 527
rect 883 459 1121 493
rect 883 393 933 459
rect 695 357 933 393
rect 977 323 1027 425
rect 623 289 1027 323
rect 1071 291 1121 459
rect 623 265 657 289
rect 599 199 657 265
rect 35 17 69 179
rect 103 95 163 179
rect 623 181 657 199
rect 623 145 1035 181
rect 103 51 367 95
rect 411 17 445 111
rect 599 17 737 111
rect 771 51 847 145
rect 891 17 925 111
rect 959 51 1035 145
rect 1079 17 1113 181
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
rlabel locali s 695 215 894 255 6 A1_N
port 1 nsew signal input
rlabel locali s 944 215 1087 255 6 A2_N
port 2 nsew signal input
rlabel locali s 343 215 419 289 6 B1
port 3 nsew signal input
rlabel locali s 22 289 419 323 6 B1
port 3 nsew signal input
rlabel locali s 22 215 128 289 6 B1
port 3 nsew signal input
rlabel locali s 171 215 289 255 6 B2
port 4 nsew signal input
rlabel locali s 489 181 555 425 6 Y
port 5 nsew signal output
rlabel locali s 479 51 555 145 6 Y
port 5 nsew signal output
rlabel locali s 197 145 555 181 6 Y
port 5 nsew signal output
rlabel locali s 197 129 273 145 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -48 1196 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 1196 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1348520
string GDS_START 1339322
<< end >>
