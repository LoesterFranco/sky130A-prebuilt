magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 1970 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 81 47 111 177
rect 181 47 211 177
rect 305 93 335 177
rect 548 49 578 177
rect 667 49 697 177
rect 939 47 969 177
rect 1145 49 1175 177
rect 1307 49 1337 133
rect 1466 49 1496 177
rect 1606 47 1636 167
rect 1716 47 1746 175
rect 1810 47 1840 175
<< pmoshvt >>
rect 83 297 119 497
rect 177 297 213 497
rect 307 297 343 425
rect 531 325 567 493
rect 647 325 683 493
rect 898 297 934 497
rect 1137 297 1173 465
rect 1299 297 1335 425
rect 1484 329 1520 457
rect 1597 329 1633 497
rect 1708 297 1744 497
rect 1802 297 1838 497
<< ndiff >>
rect 27 93 81 177
rect 27 59 37 93
rect 71 59 81 93
rect 27 47 81 59
rect 111 129 181 177
rect 111 95 136 129
rect 170 95 181 129
rect 111 47 181 95
rect 211 93 305 177
rect 335 169 429 177
rect 335 135 383 169
rect 417 135 429 169
rect 335 93 429 135
rect 483 165 548 177
rect 483 131 493 165
rect 527 131 548 165
rect 211 89 290 93
rect 211 55 237 89
rect 271 55 290 89
rect 211 47 290 55
rect 483 49 548 131
rect 578 91 667 177
rect 578 57 588 91
rect 622 57 667 91
rect 578 49 667 57
rect 697 169 796 177
rect 697 135 749 169
rect 783 135 796 169
rect 697 49 796 135
rect 869 157 939 177
rect 869 123 885 157
rect 919 123 939 157
rect 869 89 939 123
rect 869 55 885 89
rect 919 55 939 89
rect 869 47 939 55
rect 969 161 1031 177
rect 969 127 989 161
rect 1023 127 1031 161
rect 969 121 1031 127
rect 969 47 1029 121
rect 1085 105 1145 177
rect 1083 97 1145 105
rect 1083 63 1091 97
rect 1125 63 1145 97
rect 1083 49 1145 63
rect 1175 133 1276 177
rect 1362 169 1466 177
rect 1362 135 1408 169
rect 1442 135 1466 169
rect 1362 133 1466 135
rect 1175 126 1307 133
rect 1175 92 1185 126
rect 1219 92 1307 126
rect 1175 49 1307 92
rect 1337 49 1466 133
rect 1496 167 1556 177
rect 1656 167 1716 175
rect 1496 93 1606 167
rect 1496 59 1518 93
rect 1552 59 1606 93
rect 1496 49 1606 59
rect 1523 47 1606 49
rect 1636 142 1716 167
rect 1636 108 1662 142
rect 1696 108 1716 142
rect 1636 47 1716 108
rect 1746 97 1810 175
rect 1746 63 1756 97
rect 1790 63 1810 97
rect 1746 47 1810 63
rect 1840 101 1892 175
rect 1840 67 1850 101
rect 1884 67 1892 101
rect 1840 47 1892 67
<< pdiff >>
rect 29 477 83 497
rect 29 443 37 477
rect 71 443 83 477
rect 29 297 83 443
rect 119 477 177 497
rect 119 443 131 477
rect 165 443 177 477
rect 119 409 177 443
rect 119 375 131 409
rect 165 375 177 409
rect 119 341 177 375
rect 119 307 131 341
rect 165 307 177 341
rect 119 297 177 307
rect 213 477 290 497
rect 213 443 242 477
rect 276 443 290 477
rect 213 425 290 443
rect 213 297 307 425
rect 343 341 401 425
rect 343 307 355 341
rect 389 307 401 341
rect 465 413 531 493
rect 465 379 485 413
rect 519 379 531 413
rect 465 325 531 379
rect 567 481 647 493
rect 567 447 588 481
rect 622 447 647 481
rect 567 325 647 447
rect 683 481 790 493
rect 683 447 745 481
rect 779 447 790 481
rect 683 325 790 447
rect 844 481 898 497
rect 844 447 852 481
rect 886 447 898 481
rect 343 297 401 307
rect 844 297 898 447
rect 934 349 996 497
rect 1537 489 1597 497
rect 1050 405 1137 465
rect 1050 371 1058 405
rect 1092 371 1137 405
rect 1050 365 1137 371
rect 934 343 998 349
rect 934 309 946 343
rect 980 309 998 343
rect 934 297 998 309
rect 1052 297 1137 365
rect 1173 425 1275 465
rect 1537 457 1549 489
rect 1397 425 1484 457
rect 1173 409 1299 425
rect 1173 375 1226 409
rect 1260 375 1299 409
rect 1173 341 1299 375
rect 1173 307 1226 341
rect 1260 307 1299 341
rect 1173 297 1299 307
rect 1335 421 1484 425
rect 1335 387 1438 421
rect 1472 387 1484 421
rect 1335 329 1484 387
rect 1520 455 1549 457
rect 1583 455 1597 489
rect 1520 329 1597 455
rect 1633 341 1708 497
rect 1633 329 1662 341
rect 1335 297 1432 329
rect 1650 307 1662 329
rect 1696 307 1708 341
rect 1650 297 1708 307
rect 1744 489 1802 497
rect 1744 455 1756 489
rect 1790 455 1802 489
rect 1744 297 1802 455
rect 1838 477 1893 497
rect 1838 443 1851 477
rect 1885 443 1893 477
rect 1838 409 1893 443
rect 1838 375 1851 409
rect 1885 375 1893 409
rect 1838 297 1893 375
<< ndiffc >>
rect 37 59 71 93
rect 136 95 170 129
rect 383 135 417 169
rect 493 131 527 165
rect 237 55 271 89
rect 588 57 622 91
rect 749 135 783 169
rect 885 123 919 157
rect 885 55 919 89
rect 989 127 1023 161
rect 1091 63 1125 97
rect 1408 135 1442 169
rect 1185 92 1219 126
rect 1518 59 1552 93
rect 1662 108 1696 142
rect 1756 63 1790 97
rect 1850 67 1884 101
<< pdiffc >>
rect 37 443 71 477
rect 131 443 165 477
rect 131 375 165 409
rect 131 307 165 341
rect 242 443 276 477
rect 355 307 389 341
rect 485 379 519 413
rect 588 447 622 481
rect 745 447 779 481
rect 852 447 886 481
rect 1058 371 1092 405
rect 946 309 980 343
rect 1226 375 1260 409
rect 1226 307 1260 341
rect 1438 387 1472 421
rect 1549 455 1583 489
rect 1662 307 1696 341
rect 1756 455 1790 489
rect 1851 443 1885 477
rect 1851 375 1885 409
<< poly >>
rect 83 497 119 523
rect 177 497 213 523
rect 531 493 567 519
rect 647 493 683 519
rect 898 497 934 523
rect 305 451 345 483
rect 307 425 343 451
rect 531 310 567 325
rect 647 310 683 325
rect 83 282 119 297
rect 177 282 213 297
rect 307 282 343 297
rect 81 265 121 282
rect 175 265 215 282
rect 305 265 345 282
rect 529 271 569 310
rect 529 265 578 271
rect 645 265 685 310
rect 1135 493 1522 523
rect 1597 497 1633 523
rect 1708 497 1744 523
rect 1802 497 1838 523
rect 1135 491 1175 493
rect 1137 465 1173 491
rect 1482 483 1522 493
rect 1484 457 1520 483
rect 1299 425 1335 451
rect 1484 314 1520 329
rect 1597 314 1633 329
rect 898 282 934 297
rect 1137 282 1173 297
rect 1299 282 1335 297
rect 81 249 263 265
rect 81 215 219 249
rect 253 215 263 249
rect 81 199 263 215
rect 305 249 578 265
rect 305 215 456 249
rect 490 215 524 249
rect 558 215 578 249
rect 305 199 578 215
rect 633 249 697 265
rect 633 215 643 249
rect 677 215 697 249
rect 896 247 936 282
rect 1135 247 1175 282
rect 1297 265 1337 282
rect 1482 265 1522 314
rect 896 217 1175 247
rect 633 199 697 215
rect 81 177 111 199
rect 181 177 211 199
rect 305 177 335 199
rect 548 177 578 199
rect 667 177 697 199
rect 939 177 969 217
rect 1145 177 1175 217
rect 1217 249 1337 265
rect 1217 215 1227 249
rect 1261 215 1337 249
rect 1217 199 1337 215
rect 305 67 335 93
rect 81 21 111 47
rect 181 21 211 47
rect 548 21 578 49
rect 667 21 697 49
rect 1307 133 1337 199
rect 1466 249 1522 265
rect 1595 256 1635 314
rect 1708 282 1744 297
rect 1802 282 1838 297
rect 1706 265 1746 282
rect 1800 265 1840 282
rect 1595 255 1636 256
rect 1466 215 1476 249
rect 1510 215 1522 249
rect 1466 199 1522 215
rect 1574 239 1636 255
rect 1574 205 1584 239
rect 1618 205 1636 239
rect 1466 177 1496 199
rect 1574 189 1636 205
rect 1678 249 1746 265
rect 1678 215 1688 249
rect 1722 215 1746 249
rect 1678 199 1746 215
rect 1788 249 1852 265
rect 1788 215 1798 249
rect 1832 215 1852 249
rect 1788 199 1852 215
rect 1606 167 1636 189
rect 1716 175 1746 199
rect 1810 175 1840 199
rect 939 21 969 47
rect 1145 21 1175 49
rect 1307 23 1337 49
rect 1466 21 1496 49
rect 1606 21 1636 47
rect 1716 21 1746 47
rect 1810 21 1840 47
<< polycont >>
rect 219 215 253 249
rect 456 215 490 249
rect 524 215 558 249
rect 643 215 677 249
rect 1227 215 1261 249
rect 1476 215 1510 249
rect 1584 205 1618 239
rect 1688 215 1722 249
rect 1798 215 1832 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 21 477 87 527
rect 21 443 37 477
rect 71 443 87 477
rect 131 477 181 493
rect 165 443 181 477
rect 225 477 292 527
rect 836 481 902 527
rect 1730 489 1807 527
rect 225 443 242 477
rect 276 443 292 477
rect 329 447 588 481
rect 622 447 668 481
rect 721 447 745 481
rect 779 447 802 481
rect 836 447 852 481
rect 886 447 902 481
rect 989 455 1549 489
rect 1583 455 1648 489
rect 1730 455 1756 489
rect 1790 455 1807 489
rect 1851 477 1910 493
rect 131 409 181 443
rect 329 409 373 447
rect 768 413 802 447
rect 989 413 1023 455
rect 66 375 131 409
rect 165 375 181 409
rect 66 341 181 375
rect 66 307 131 341
rect 165 307 181 341
rect 66 288 181 307
rect 225 375 373 409
rect 453 379 485 413
rect 519 379 734 413
rect 768 379 1023 413
rect 1058 405 1092 421
rect 66 185 139 288
rect 225 265 259 375
rect 306 307 355 341
rect 389 307 656 341
rect 219 249 259 265
rect 253 215 259 249
rect 219 199 259 215
rect 66 132 186 185
rect 225 173 259 199
rect 225 139 349 173
rect 136 129 186 132
rect 170 95 186 129
rect 21 59 37 93
rect 71 59 87 93
rect 136 70 186 95
rect 221 89 271 105
rect 21 17 87 59
rect 221 55 237 89
rect 221 17 271 55
rect 305 85 349 139
rect 383 169 417 307
rect 622 265 656 307
rect 700 339 734 379
rect 700 323 806 339
rect 700 305 772 323
rect 749 289 772 305
rect 749 275 806 289
rect 451 249 588 265
rect 451 215 456 249
rect 490 215 524 249
rect 558 215 588 249
rect 451 199 588 215
rect 622 249 687 265
rect 622 215 643 249
rect 677 215 687 249
rect 622 199 687 215
rect 749 169 783 275
rect 840 241 874 379
rect 920 309 946 343
rect 980 309 1023 343
rect 920 289 1023 309
rect 383 119 417 135
rect 473 131 493 165
rect 527 131 715 165
rect 557 85 588 91
rect 305 57 588 85
rect 622 57 638 91
rect 305 51 638 57
rect 672 85 715 131
rect 749 119 783 135
rect 817 207 874 241
rect 817 85 851 207
rect 965 187 1023 289
rect 672 51 851 85
rect 885 157 919 173
rect 885 89 919 123
rect 965 153 966 187
rect 1000 161 1023 187
rect 965 127 989 153
rect 965 83 1023 127
rect 1058 119 1092 371
rect 1126 178 1160 455
rect 1885 443 1910 477
rect 1851 421 1910 443
rect 1208 375 1226 409
rect 1260 375 1291 409
rect 1208 341 1291 375
rect 1208 307 1226 341
rect 1260 323 1291 341
rect 1408 387 1438 421
rect 1472 409 1910 421
rect 1472 387 1851 409
rect 1260 307 1262 323
rect 1208 289 1262 307
rect 1296 289 1374 323
rect 1211 249 1296 254
rect 1211 215 1227 249
rect 1261 215 1296 249
rect 1211 199 1296 215
rect 1253 187 1296 199
rect 1126 165 1180 178
rect 1126 144 1219 165
rect 1136 131 1219 144
rect 1185 126 1219 131
rect 1253 153 1262 187
rect 1253 126 1296 153
rect 1058 85 1068 119
rect 885 17 919 55
rect 1058 63 1091 85
rect 1125 63 1141 97
rect 1185 64 1219 92
rect 1340 85 1374 289
rect 1408 169 1442 387
rect 1803 375 1851 387
rect 1885 375 1910 409
rect 1476 289 1602 333
rect 1646 307 1662 341
rect 1696 307 1820 341
rect 1646 299 1820 307
rect 1476 249 1520 289
rect 1786 265 1820 299
rect 1510 215 1520 249
rect 1476 199 1520 215
rect 1554 239 1618 255
rect 1554 205 1584 239
rect 1660 249 1752 265
rect 1660 215 1688 249
rect 1722 215 1752 249
rect 1786 249 1842 265
rect 1786 215 1798 249
rect 1832 215 1842 249
rect 1554 189 1618 205
rect 1786 199 1842 215
rect 1554 187 1595 189
rect 1554 153 1558 187
rect 1592 153 1595 187
rect 1786 181 1820 199
rect 1554 146 1595 153
rect 1662 150 1820 181
rect 1654 147 1820 150
rect 1408 119 1442 135
rect 1654 142 1712 147
rect 1654 119 1662 142
rect 1476 85 1518 93
rect 1058 53 1141 63
rect 1340 59 1518 85
rect 1552 59 1579 93
rect 1654 85 1660 119
rect 1696 108 1712 142
rect 1876 117 1910 375
rect 1694 85 1712 108
rect 1654 59 1712 85
rect 1756 97 1790 113
rect 1340 51 1579 59
rect 1756 17 1790 63
rect 1850 101 1910 117
rect 1884 67 1910 101
rect 1850 51 1910 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 772 289 806 323
rect 966 161 1000 187
rect 966 153 989 161
rect 989 153 1000 161
rect 1262 289 1296 323
rect 1262 153 1296 187
rect 1068 97 1102 119
rect 1068 85 1091 97
rect 1091 85 1102 97
rect 1558 153 1592 187
rect 1660 108 1662 119
rect 1662 108 1694 119
rect 1660 85 1694 108
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
rect 760 323 818 329
rect 760 289 772 323
rect 806 320 818 323
rect 1250 323 1308 329
rect 1250 320 1262 323
rect 806 292 1262 320
rect 806 289 818 292
rect 760 283 818 289
rect 1250 289 1262 292
rect 1296 289 1308 323
rect 1250 283 1308 289
rect 954 187 1012 193
rect 954 153 966 187
rect 1000 184 1012 187
rect 1250 187 1308 193
rect 1250 184 1262 187
rect 1000 156 1262 184
rect 1000 153 1012 156
rect 954 147 1012 153
rect 1250 153 1262 156
rect 1296 184 1308 187
rect 1546 187 1604 193
rect 1546 184 1558 187
rect 1296 156 1558 184
rect 1296 153 1308 156
rect 1250 147 1308 153
rect 1546 153 1558 156
rect 1592 153 1604 187
rect 1546 147 1604 153
rect 1056 119 1114 125
rect 1056 85 1068 119
rect 1102 116 1114 119
rect 1648 119 1706 125
rect 1648 116 1660 119
rect 1102 88 1660 116
rect 1102 85 1114 88
rect 1056 79 1114 85
rect 1648 85 1660 88
rect 1694 85 1706 119
rect 1648 79 1706 85
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< labels >>
flabel corelocali s 121 357 155 391 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 490 221 524 255 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 1502 289 1536 323 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 1679 238 1679 238 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
rlabel comment s 0 0 0 0 4 xor3_2
<< properties >>
string FIXED_BBOX 0 0 1932 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 805980
string GDS_START 793160
<< end >>
