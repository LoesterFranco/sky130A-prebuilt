magic
tech sky130A
magscale 1 2
timestamp 1604502741
<< locali >>
rect 191 236 257 350
rect 984 236 1050 310
rect 1375 236 1425 337
rect 1741 74 1807 596
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 17 452 119 591
rect 153 452 219 649
rect 262 581 779 615
rect 17 255 51 452
rect 262 418 328 581
rect 745 551 779 581
rect 85 415 328 418
rect 370 513 711 547
rect 370 415 436 513
rect 85 384 325 415
rect 85 289 149 384
rect 17 166 89 255
rect 291 200 325 384
rect 470 313 536 479
rect 577 375 643 479
rect 359 279 536 313
rect 359 166 393 279
rect 502 245 536 279
rect 17 132 393 166
rect 17 130 89 132
rect 427 119 461 245
rect 502 153 575 245
rect 609 119 643 375
rect 125 17 239 98
rect 427 85 643 119
rect 677 85 711 513
rect 745 381 879 551
rect 745 287 811 347
rect 745 153 779 287
rect 845 253 879 381
rect 813 187 879 253
rect 916 202 950 596
rect 990 364 1040 649
rect 1081 384 1168 596
rect 1202 581 1490 615
rect 1102 237 1136 384
rect 1202 337 1236 581
rect 1170 271 1236 337
rect 1270 305 1320 540
rect 1357 405 1410 538
rect 1456 500 1490 581
rect 1456 439 1561 500
rect 1357 371 1493 405
rect 1270 271 1341 305
rect 1102 203 1273 237
rect 916 153 961 202
rect 745 119 961 153
rect 995 135 1205 169
rect 995 85 1029 135
rect 677 51 1029 85
rect 1063 17 1113 101
rect 1155 85 1205 135
rect 1239 153 1273 203
rect 1307 187 1341 271
rect 1459 253 1493 371
rect 1527 321 1561 439
rect 1595 464 1706 649
rect 1595 364 1629 464
rect 1663 330 1705 430
rect 1527 287 1605 321
rect 1459 219 1521 253
rect 1377 153 1453 185
rect 1239 119 1453 153
rect 1487 85 1521 219
rect 1155 51 1521 85
rect 1555 74 1605 287
rect 1639 264 1705 330
rect 1641 17 1707 230
rect 1847 364 1897 649
rect 1843 17 1893 230
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
<< metal1 >>
rect 0 683 1920 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 0 617 1920 649
rect 0 17 1920 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
rect 0 -49 1920 -17
<< obsm1 >>
rect 595 421 653 430
rect 1075 421 1133 430
rect 595 393 1133 421
rect 595 384 653 393
rect 1075 384 1133 393
rect 1267 421 1325 430
rect 1651 421 1709 430
rect 1267 393 1709 421
rect 1267 384 1325 393
rect 1651 384 1709 393
<< labels >>
rlabel locali s 191 236 257 350 6 A
port 1 nsew signal input
rlabel locali s 984 236 1050 310 6 B
port 2 nsew signal input
rlabel locali s 1375 236 1425 337 6 C
port 3 nsew signal input
rlabel locali s 1741 74 1807 596 6 X
port 4 nsew signal output
rlabel metal1 s 0 -49 1920 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 617 1920 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1920 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 586836
string GDS_START 572620
<< end >>
