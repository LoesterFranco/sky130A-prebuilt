magic
tech sky130A
magscale 1 2
timestamp 1604502705
<< nwell >>
rect -38 332 518 704
<< pwell >>
rect 0 0 480 49
<< scnmos >>
rect 88 74 118 222
rect 166 74 196 222
rect 268 74 298 222
rect 354 74 384 222
<< pmoshvt >>
rect 85 392 115 592
rect 175 392 205 592
rect 276 368 306 592
rect 366 368 396 592
<< ndiff >>
rect 31 210 88 222
rect 31 176 43 210
rect 77 176 88 210
rect 31 120 88 176
rect 31 86 43 120
rect 77 86 88 120
rect 31 74 88 86
rect 118 74 166 222
rect 196 131 268 222
rect 196 97 207 131
rect 241 97 268 131
rect 196 74 268 97
rect 298 131 354 222
rect 298 97 309 131
rect 343 97 354 131
rect 298 74 354 97
rect 384 120 453 222
rect 384 86 401 120
rect 435 86 453 120
rect 384 74 453 86
<< pdiff >>
rect 27 580 85 592
rect 27 546 38 580
rect 72 546 85 580
rect 27 510 85 546
rect 27 476 38 510
rect 72 476 85 510
rect 27 440 85 476
rect 27 406 38 440
rect 72 406 85 440
rect 27 392 85 406
rect 115 580 175 592
rect 115 546 128 580
rect 162 546 175 580
rect 115 510 175 546
rect 115 476 128 510
rect 162 476 175 510
rect 115 440 175 476
rect 115 406 128 440
rect 162 406 175 440
rect 115 392 175 406
rect 205 580 276 592
rect 205 546 228 580
rect 262 546 276 580
rect 205 508 276 546
rect 205 474 228 508
rect 262 474 276 508
rect 205 392 276 474
rect 223 368 276 392
rect 306 580 366 592
rect 306 546 319 580
rect 353 546 366 580
rect 306 497 366 546
rect 306 463 319 497
rect 353 463 366 497
rect 306 414 366 463
rect 306 380 319 414
rect 353 380 366 414
rect 306 368 366 380
rect 396 580 453 592
rect 396 546 409 580
rect 443 546 453 580
rect 396 462 453 546
rect 396 428 409 462
rect 443 428 453 462
rect 396 368 453 428
<< ndiffc >>
rect 43 176 77 210
rect 43 86 77 120
rect 207 97 241 131
rect 309 97 343 131
rect 401 86 435 120
<< pdiffc >>
rect 38 546 72 580
rect 38 476 72 510
rect 38 406 72 440
rect 128 546 162 580
rect 128 476 162 510
rect 128 406 162 440
rect 228 546 262 580
rect 228 474 262 508
rect 319 546 353 580
rect 319 463 353 497
rect 319 380 353 414
rect 409 546 443 580
rect 409 428 443 462
<< poly >>
rect 85 592 115 618
rect 175 592 205 618
rect 276 592 306 618
rect 366 592 396 618
rect 85 377 115 392
rect 175 377 205 392
rect 82 326 118 377
rect 172 326 208 377
rect 276 353 306 368
rect 366 353 396 368
rect 21 310 118 326
rect 21 276 37 310
rect 71 276 118 310
rect 21 260 118 276
rect 160 310 226 326
rect 273 310 309 353
rect 363 310 399 353
rect 160 276 176 310
rect 210 276 226 310
rect 160 260 226 276
rect 268 294 399 310
rect 268 260 284 294
rect 318 260 399 294
rect 88 222 118 260
rect 166 222 196 260
rect 268 244 399 260
rect 268 222 298 244
rect 354 222 384 244
rect 88 48 118 74
rect 166 48 196 74
rect 268 48 298 74
rect 354 48 384 74
<< polycont >>
rect 37 276 71 310
rect 176 276 210 310
rect 284 260 318 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 22 580 88 649
rect 22 546 38 580
rect 72 546 88 580
rect 22 510 88 546
rect 22 476 38 510
rect 72 476 88 510
rect 22 440 88 476
rect 22 406 38 440
rect 72 406 88 440
rect 22 390 88 406
rect 128 580 178 596
rect 162 546 178 580
rect 128 510 178 546
rect 162 476 178 510
rect 128 440 178 476
rect 212 580 278 649
rect 212 546 228 580
rect 262 546 278 580
rect 212 508 278 546
rect 212 474 228 508
rect 262 474 278 508
rect 212 458 278 474
rect 319 580 369 596
rect 353 546 369 580
rect 319 497 369 546
rect 353 463 369 497
rect 162 424 178 440
rect 162 406 285 424
rect 128 390 285 406
rect 21 310 87 356
rect 21 276 37 310
rect 71 276 87 310
rect 21 260 87 276
rect 121 310 217 356
rect 121 276 176 310
rect 210 276 217 310
rect 121 260 217 276
rect 251 310 285 390
rect 319 414 369 463
rect 353 380 369 414
rect 409 580 459 649
rect 443 546 459 580
rect 409 462 459 546
rect 443 428 459 462
rect 409 412 459 428
rect 319 378 369 380
rect 319 344 402 378
rect 251 294 334 310
rect 251 260 284 294
rect 318 260 334 294
rect 251 244 334 260
rect 251 226 285 244
rect 27 210 285 226
rect 27 176 43 210
rect 77 192 285 210
rect 368 204 402 344
rect 77 176 93 192
rect 27 120 93 176
rect 325 170 402 204
rect 325 158 359 170
rect 27 86 43 120
rect 77 86 93 120
rect 27 70 93 86
rect 191 131 257 158
rect 191 97 207 131
rect 241 97 257 131
rect 191 17 257 97
rect 293 131 359 158
rect 293 97 309 131
rect 343 97 359 131
rect 293 70 359 97
rect 395 120 457 136
rect 395 86 401 120
rect 435 86 457 120
rect 395 17 457 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< metal1 >>
rect 0 683 480 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 0 617 480 649
rect 0 17 480 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
rect 0 -49 480 -17
<< labels >>
rlabel comment s 0 0 0 0 4 and2_2
flabel pwell s 0 0 480 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 0 617 480 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 0 617 480 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 480 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 319 390 353 424 0 FreeSans 340 0 0 0 X
port 7 nsew
flabel corelocali s 319 464 353 498 0 FreeSans 340 0 0 0 X
port 7 nsew
flabel corelocali s 319 538 353 572 0 FreeSans 340 0 0 0 X
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 480 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3808312
string GDS_START 3803110
<< end >>
