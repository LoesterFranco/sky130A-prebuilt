magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 828 561
rect 147 359 197 527
rect 17 199 83 257
rect 299 265 363 341
rect 185 215 251 257
rect 287 215 363 265
rect 401 257 476 341
rect 578 359 644 527
rect 678 375 811 493
rect 401 215 498 257
rect 536 215 626 257
rect 761 181 811 375
rect 438 17 472 111
rect 606 17 640 181
rect 674 53 811 181
rect 0 -17 828 17
<< obsli1 >>
rect 48 325 108 493
rect 315 409 476 493
rect 231 375 544 409
rect 231 325 265 375
rect 48 291 265 325
rect 117 165 151 291
rect 510 325 544 375
rect 510 291 694 325
rect 660 257 694 291
rect 660 215 727 257
rect 49 129 151 165
rect 232 147 572 181
rect 232 129 309 147
rect 49 51 115 129
rect 149 61 386 95
rect 506 54 572 147
<< metal1 >>
rect 0 496 828 592
rect 0 -48 828 48
<< labels >>
rlabel locali s 536 215 626 257 6 A1
port 1 nsew signal input
rlabel locali s 401 257 476 341 6 A2
port 2 nsew signal input
rlabel locali s 401 215 498 257 6 A2
port 2 nsew signal input
rlabel locali s 185 215 251 257 6 B1
port 3 nsew signal input
rlabel locali s 299 265 363 341 6 B2
port 4 nsew signal input
rlabel locali s 287 215 363 265 6 B2
port 4 nsew signal input
rlabel locali s 17 199 83 257 6 C1
port 5 nsew signal input
rlabel locali s 761 181 811 375 6 X
port 6 nsew signal output
rlabel locali s 678 375 811 493 6 X
port 6 nsew signal output
rlabel locali s 674 53 811 181 6 X
port 6 nsew signal output
rlabel locali s 606 17 640 181 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 438 17 472 111 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 828 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 828 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 578 359 644 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 147 359 197 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 828 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 828 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1419676
string GDS_START 1412446
<< end >>
