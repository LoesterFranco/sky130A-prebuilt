magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 1263 436 1318 596
rect 1459 436 1509 596
rect 25 290 110 356
rect 217 290 359 356
rect 597 290 663 356
rect 697 290 1031 356
rect 1065 290 1131 356
rect 1263 370 1509 436
rect 1459 330 1509 370
rect 1459 296 1607 330
rect 1561 236 1607 296
rect 1237 202 1607 236
rect 1237 70 1303 202
rect 1437 70 1503 202
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 23 424 89 564
rect 123 463 189 649
rect 223 424 289 564
rect 323 463 389 649
rect 430 424 496 564
rect 537 463 603 649
rect 644 581 910 615
rect 644 424 710 581
rect 744 492 810 547
rect 844 526 910 581
rect 956 526 1022 649
rect 1056 492 1122 596
rect 744 458 1122 492
rect 1163 458 1229 649
rect 1353 470 1419 649
rect 23 390 1229 424
rect 144 226 178 390
rect 430 388 496 390
rect 1195 336 1229 390
rect 1195 270 1425 336
rect 1543 364 1609 649
rect 473 256 555 260
rect 23 120 76 223
rect 110 154 178 226
rect 212 120 246 226
rect 23 85 246 120
rect 282 176 348 226
rect 473 222 1101 256
rect 473 210 711 222
rect 282 142 625 176
rect 282 119 348 142
rect 384 85 450 108
rect 575 104 625 142
rect 661 104 711 210
rect 23 51 450 85
rect 747 17 813 188
rect 847 104 913 222
rect 965 17 1031 188
rect 1067 70 1101 222
rect 1137 17 1203 226
rect 1337 17 1403 163
rect 1537 17 1603 163
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
rlabel locali s 1065 290 1131 356 6 A1
port 1 nsew signal input
rlabel locali s 697 290 1031 356 6 A2
port 2 nsew signal input
rlabel locali s 597 290 663 356 6 B1
port 3 nsew signal input
rlabel locali s 217 290 359 356 6 C1
port 4 nsew signal input
rlabel locali s 25 290 110 356 6 D1
port 5 nsew signal input
rlabel locali s 1561 236 1607 296 6 X
port 6 nsew signal output
rlabel locali s 1459 436 1509 596 6 X
port 6 nsew signal output
rlabel locali s 1459 330 1509 370 6 X
port 6 nsew signal output
rlabel locali s 1459 296 1607 330 6 X
port 6 nsew signal output
rlabel locali s 1437 70 1503 202 6 X
port 6 nsew signal output
rlabel locali s 1263 436 1318 596 6 X
port 6 nsew signal output
rlabel locali s 1263 370 1509 436 6 X
port 6 nsew signal output
rlabel locali s 1237 202 1607 236 6 X
port 6 nsew signal output
rlabel locali s 1237 70 1303 202 6 X
port 6 nsew signal output
rlabel metal1 s 0 -49 1632 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 617 1632 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1733404
string GDS_START 1720482
<< end >>
