magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 17 370 98 596
rect 17 236 51 370
rect 217 286 337 356
rect 457 352 551 356
rect 457 286 715 352
rect 17 96 89 236
rect 697 114 743 134
rect 529 51 743 114
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 132 390 198 649
rect 313 424 379 588
rect 487 458 568 649
rect 679 424 745 588
rect 313 390 745 424
rect 85 270 157 336
rect 123 252 157 270
rect 379 252 413 390
rect 679 386 745 390
rect 123 218 740 252
rect 123 17 198 182
rect 296 116 362 218
rect 461 148 570 182
rect 674 168 740 218
rect 461 17 495 148
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel locali s 697 114 743 134 6 A
port 1 nsew signal input
rlabel locali s 529 51 743 114 6 A
port 1 nsew signal input
rlabel locali s 217 286 337 356 6 B
port 2 nsew signal input
rlabel locali s 457 352 551 356 6 C
port 3 nsew signal input
rlabel locali s 457 286 715 352 6 C
port 3 nsew signal input
rlabel locali s 17 370 98 596 6 X
port 4 nsew signal output
rlabel locali s 17 236 51 370 6 X
port 4 nsew signal output
rlabel locali s 17 96 89 236 6 X
port 4 nsew signal output
rlabel metal1 s 0 -49 768 49 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 617 768 715 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2420170
string GDS_START 2413322
<< end >>
