magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 92 47 122 177
rect 176 47 206 177
rect 366 47 396 177
rect 464 47 494 177
rect 548 47 578 177
<< pmoshvt >>
rect 84 297 120 497
rect 178 297 214 497
rect 358 297 394 497
rect 456 297 492 497
rect 550 297 586 497
<< ndiff >>
rect 27 163 92 177
rect 27 129 35 163
rect 69 129 92 163
rect 27 95 92 129
rect 27 61 35 95
rect 69 61 92 95
rect 27 47 92 61
rect 122 47 176 177
rect 206 163 258 177
rect 206 129 216 163
rect 250 129 258 163
rect 206 95 258 129
rect 206 61 216 95
rect 250 61 258 95
rect 206 47 258 61
rect 312 138 366 177
rect 312 104 322 138
rect 356 104 366 138
rect 312 47 366 104
rect 396 138 464 177
rect 396 104 420 138
rect 454 104 464 138
rect 396 47 464 104
rect 494 95 548 177
rect 494 61 504 95
rect 538 61 548 95
rect 494 47 548 61
rect 578 163 640 177
rect 578 129 598 163
rect 632 129 640 163
rect 578 95 640 129
rect 578 61 598 95
rect 632 61 640 95
rect 578 47 640 61
<< pdiff >>
rect 27 479 84 497
rect 27 445 38 479
rect 72 445 84 479
rect 27 411 84 445
rect 27 377 38 411
rect 72 377 84 411
rect 27 343 84 377
rect 27 309 38 343
rect 72 309 84 343
rect 27 297 84 309
rect 120 477 178 497
rect 120 443 132 477
rect 166 443 178 477
rect 120 409 178 443
rect 120 375 132 409
rect 166 375 178 409
rect 120 297 178 375
rect 214 477 358 497
rect 214 443 234 477
rect 268 443 304 477
rect 338 443 358 477
rect 214 409 358 443
rect 214 375 234 409
rect 268 375 304 409
rect 338 375 358 409
rect 214 297 358 375
rect 394 477 456 497
rect 394 443 406 477
rect 440 443 456 477
rect 394 409 456 443
rect 394 375 406 409
rect 440 375 456 409
rect 394 341 456 375
rect 394 307 406 341
rect 440 307 456 341
rect 394 297 456 307
rect 492 297 550 497
rect 586 479 640 497
rect 586 445 598 479
rect 632 445 640 479
rect 586 411 640 445
rect 586 377 598 411
rect 632 377 640 411
rect 586 343 640 377
rect 586 309 598 343
rect 632 309 640 343
rect 586 297 640 309
<< ndiffc >>
rect 35 129 69 163
rect 35 61 69 95
rect 216 129 250 163
rect 216 61 250 95
rect 322 104 356 138
rect 420 104 454 138
rect 504 61 538 95
rect 598 129 632 163
rect 598 61 632 95
<< pdiffc >>
rect 38 445 72 479
rect 38 377 72 411
rect 38 309 72 343
rect 132 443 166 477
rect 132 375 166 409
rect 234 443 268 477
rect 304 443 338 477
rect 234 375 268 409
rect 304 375 338 409
rect 406 443 440 477
rect 406 375 440 409
rect 406 307 440 341
rect 598 445 632 479
rect 598 377 632 411
rect 598 309 632 343
<< poly >>
rect 84 497 120 523
rect 178 497 214 523
rect 358 497 394 523
rect 456 497 492 523
rect 550 497 586 523
rect 84 282 120 297
rect 178 282 214 297
rect 358 282 394 297
rect 456 282 492 297
rect 550 282 586 297
rect 82 265 122 282
rect 21 249 122 265
rect 21 215 37 249
rect 71 215 122 249
rect 21 199 122 215
rect 92 177 122 199
rect 176 265 216 282
rect 356 265 396 282
rect 454 265 494 282
rect 176 249 230 265
rect 176 215 186 249
rect 220 215 230 249
rect 176 199 230 215
rect 272 249 396 265
rect 272 215 282 249
rect 316 215 396 249
rect 272 199 396 215
rect 440 249 494 265
rect 440 215 450 249
rect 484 215 494 249
rect 440 199 494 215
rect 176 177 206 199
rect 366 177 396 199
rect 464 177 494 199
rect 548 265 588 282
rect 548 249 649 265
rect 548 215 599 249
rect 633 215 649 249
rect 548 199 649 215
rect 548 177 578 199
rect 92 21 122 47
rect 176 21 206 47
rect 366 21 396 47
rect 464 21 494 47
rect 548 21 578 47
<< polycont >>
rect 37 215 71 249
rect 186 215 220 249
rect 282 215 316 249
rect 450 215 484 249
rect 599 215 633 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 30 479 80 527
rect 30 445 38 479
rect 72 445 80 479
rect 30 411 80 445
rect 30 377 38 411
rect 72 377 80 411
rect 30 343 80 377
rect 30 309 38 343
rect 72 309 80 343
rect 30 291 80 309
rect 124 477 174 493
rect 124 443 132 477
rect 166 443 174 477
rect 124 409 174 443
rect 124 375 132 409
rect 166 375 174 409
rect 124 333 174 375
rect 218 477 356 527
rect 218 443 234 477
rect 268 443 304 477
rect 338 443 356 477
rect 218 409 356 443
rect 218 375 234 409
rect 268 375 304 409
rect 338 375 356 409
rect 218 367 356 375
rect 390 477 455 493
rect 390 443 406 477
rect 440 443 455 477
rect 390 409 455 443
rect 390 375 406 409
rect 440 375 455 409
rect 390 341 455 375
rect 390 333 406 341
rect 124 299 288 333
rect 254 265 288 299
rect 352 307 406 333
rect 440 307 455 341
rect 352 289 455 307
rect 17 249 87 257
rect 17 215 37 249
rect 71 215 87 249
rect 17 197 87 215
rect 121 249 220 265
rect 121 215 186 249
rect 121 199 220 215
rect 254 249 316 265
rect 254 215 282 249
rect 254 199 316 215
rect 18 129 35 163
rect 69 129 85 163
rect 18 95 85 129
rect 18 61 35 95
rect 69 61 85 95
rect 18 17 85 61
rect 121 56 165 199
rect 254 165 288 199
rect 200 163 288 165
rect 200 129 216 163
rect 250 129 288 163
rect 352 158 386 289
rect 489 255 523 485
rect 590 479 640 527
rect 590 445 598 479
rect 632 445 640 479
rect 590 411 640 445
rect 590 377 598 411
rect 632 377 640 411
rect 590 343 640 377
rect 590 309 598 343
rect 632 309 640 343
rect 590 291 640 309
rect 430 249 523 255
rect 430 215 450 249
rect 484 215 523 249
rect 573 249 649 257
rect 573 215 599 249
rect 633 215 649 249
rect 200 95 288 129
rect 200 61 216 95
rect 250 61 288 95
rect 322 138 386 158
rect 356 104 386 138
rect 322 86 386 104
rect 420 163 648 181
rect 420 145 598 163
rect 420 138 470 145
rect 454 104 470 138
rect 572 129 598 145
rect 632 129 648 163
rect 420 85 470 104
rect 504 95 538 111
rect 200 56 288 61
rect 504 17 538 61
rect 572 95 648 129
rect 572 61 598 95
rect 632 61 648 95
rect 572 55 648 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel corelocali s 397 357 431 391 0 FreeSans 400 0 0 0 Y
port 9 nsew
flabel corelocali s 29 221 63 255 0 FreeSans 200 0 0 0 A1_N
port 1 nsew
flabel corelocali s 121 221 155 255 0 FreeSans 400 0 0 0 A2_N
port 2 nsew
flabel corelocali s 489 289 523 323 0 FreeSans 400 0 0 0 B2
port 4 nsew
flabel corelocali s 581 221 615 255 0 FreeSans 400 0 0 0 B1
port 3 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
rlabel comment s 0 0 0 0 4 o2bb2ai_1
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 912454
string GDS_START 906012
<< end >>
