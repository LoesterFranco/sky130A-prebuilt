magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 590 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 79 47 109 177
rect 183 47 213 177
rect 267 47 297 177
rect 371 47 401 177
<< pmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
<< ndiff >>
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 93 183 177
rect 109 59 129 93
rect 163 59 183 93
rect 109 47 183 59
rect 213 161 267 177
rect 213 127 223 161
rect 257 127 267 161
rect 213 93 267 127
rect 213 59 223 93
rect 257 59 267 93
rect 213 47 267 59
rect 297 165 371 177
rect 297 131 317 165
rect 351 131 371 165
rect 297 47 371 131
rect 401 93 453 177
rect 401 59 411 93
rect 445 59 453 93
rect 401 47 453 59
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 485 175 497
rect 117 451 129 485
rect 163 451 175 485
rect 117 417 175 451
rect 117 383 129 417
rect 163 383 175 417
rect 117 349 175 383
rect 117 315 129 349
rect 163 315 175 349
rect 117 297 175 315
rect 211 485 269 497
rect 211 451 223 485
rect 257 451 269 485
rect 211 417 269 451
rect 211 383 223 417
rect 257 383 269 417
rect 211 297 269 383
rect 305 485 363 497
rect 305 451 317 485
rect 351 451 363 485
rect 305 417 363 451
rect 305 383 317 417
rect 351 383 363 417
rect 305 349 363 383
rect 305 315 317 349
rect 351 315 363 349
rect 305 297 363 315
rect 399 485 453 497
rect 399 451 411 485
rect 445 451 453 485
rect 399 417 453 451
rect 399 383 411 417
rect 445 383 453 417
rect 399 297 453 383
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 129 59 163 93
rect 223 127 257 161
rect 223 59 257 93
rect 317 131 351 165
rect 411 59 445 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 451 163 485
rect 129 383 163 417
rect 129 315 163 349
rect 223 451 257 485
rect 223 383 257 417
rect 317 451 351 485
rect 317 383 351 417
rect 317 315 351 349
rect 411 451 445 485
rect 411 383 445 417
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 79 265 119 282
rect 173 265 213 282
rect 79 249 213 265
rect 79 215 129 249
rect 163 215 213 249
rect 79 199 213 215
rect 79 177 109 199
rect 183 177 213 199
rect 267 265 307 282
rect 361 265 401 282
rect 267 249 401 265
rect 267 215 290 249
rect 324 215 401 249
rect 267 199 401 215
rect 267 177 297 199
rect 371 177 401 199
rect 79 21 109 47
rect 183 21 213 47
rect 267 21 297 47
rect 371 21 401 47
<< polycont >>
rect 129 215 163 249
rect 290 215 324 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 17 485 69 527
rect 17 451 35 485
rect 17 417 69 451
rect 17 383 35 417
rect 17 349 69 383
rect 17 315 35 349
rect 17 299 69 315
rect 103 485 179 493
rect 103 451 129 485
rect 163 451 179 485
rect 103 417 179 451
rect 103 383 129 417
rect 163 383 179 417
rect 103 349 179 383
rect 223 485 257 527
rect 223 417 257 451
rect 223 367 257 383
rect 291 485 367 493
rect 291 451 317 485
rect 351 451 367 485
rect 291 417 367 451
rect 291 383 317 417
rect 351 383 367 417
rect 103 315 129 349
rect 163 333 179 349
rect 291 349 367 383
rect 411 485 462 527
rect 445 451 462 485
rect 411 417 462 451
rect 445 383 462 417
rect 411 367 462 383
rect 291 333 317 349
rect 163 315 317 333
rect 351 333 367 349
rect 351 315 446 333
rect 103 299 446 315
rect 17 249 179 265
rect 17 215 129 249
rect 163 215 179 249
rect 213 249 356 265
rect 213 215 290 249
rect 324 215 356 249
rect 390 181 446 299
rect 17 161 257 177
rect 17 127 35 161
rect 69 143 223 161
rect 69 127 85 143
rect 17 93 85 127
rect 197 127 223 143
rect 291 165 446 181
rect 291 131 317 165
rect 351 131 446 165
rect 17 59 35 93
rect 69 59 85 93
rect 17 51 85 59
rect 129 93 163 109
rect 129 17 163 59
rect 197 97 257 127
rect 197 93 461 97
rect 197 59 223 93
rect 257 59 411 93
rect 445 59 461 93
rect 197 51 461 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
flabel corelocali s 401 153 435 187 0 FreeSans 250 0 0 0 Y
port 7 nsew
flabel corelocali s 401 221 435 255 0 FreeSans 250 0 0 0 Y
port 7 nsew
flabel corelocali s 401 289 435 323 0 FreeSans 250 0 0 0 Y
port 7 nsew
flabel corelocali s 309 221 343 255 0 FreeSans 250 0 0 0 A
port 1 nsew
flabel corelocali s 132 221 166 255 0 FreeSans 250 0 0 0 B
port 2 nsew
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew
rlabel comment s 0 0 0 0 4 nand2_2
<< properties >>
string FIXED_BBOX 0 0 552 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2196566
string GDS_START 2191314
<< end >>
