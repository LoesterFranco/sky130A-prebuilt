magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 1418 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 80 47 110 177
rect 174 47 204 177
rect 268 47 298 177
rect 362 47 392 177
rect 577 47 607 177
rect 649 47 679 177
rect 788 47 818 177
rect 865 47 895 177
rect 960 47 990 177
rect 1068 47 1098 177
rect 1164 47 1194 177
rect 1260 47 1290 177
<< pmoshvt >>
rect 170 297 206 497
rect 266 297 302 497
rect 362 297 398 497
rect 458 297 494 497
rect 553 297 589 497
rect 684 297 720 497
rect 780 297 816 497
rect 879 297 915 497
rect 974 297 1010 497
rect 1070 297 1106 497
rect 1166 297 1202 497
rect 1262 297 1298 497
<< ndiff >>
rect 27 93 80 177
rect 27 59 35 93
rect 69 59 80 93
rect 27 47 80 59
rect 110 101 174 177
rect 110 67 129 101
rect 163 67 174 101
rect 110 47 174 67
rect 204 89 268 177
rect 204 55 223 89
rect 257 55 268 89
rect 204 47 268 55
rect 298 101 362 177
rect 298 67 317 101
rect 351 67 362 101
rect 298 47 362 67
rect 392 93 460 177
rect 392 59 411 93
rect 445 59 460 93
rect 392 47 460 59
rect 524 93 577 177
rect 524 59 532 93
rect 566 59 577 93
rect 524 47 577 59
rect 607 47 649 177
rect 679 163 788 177
rect 679 129 704 163
rect 738 129 788 163
rect 679 47 788 129
rect 818 47 865 177
rect 895 169 960 177
rect 895 135 911 169
rect 945 135 960 169
rect 895 101 960 135
rect 895 67 911 101
rect 945 67 960 101
rect 895 47 960 67
rect 990 89 1068 177
rect 990 55 1009 89
rect 1043 55 1068 89
rect 990 47 1068 55
rect 1098 157 1164 177
rect 1098 123 1119 157
rect 1153 123 1164 157
rect 1098 89 1164 123
rect 1098 55 1119 89
rect 1153 55 1164 89
rect 1098 47 1164 55
rect 1194 89 1260 177
rect 1194 55 1215 89
rect 1249 55 1260 89
rect 1194 47 1260 55
rect 1290 161 1353 177
rect 1290 127 1311 161
rect 1345 127 1353 161
rect 1290 93 1353 127
rect 1290 59 1311 93
rect 1345 59 1353 93
rect 1290 47 1353 59
<< pdiff >>
rect 104 485 170 497
rect 104 451 122 485
rect 156 451 170 485
rect 104 408 170 451
rect 104 374 122 408
rect 156 374 170 408
rect 104 297 170 374
rect 206 477 266 497
rect 206 443 218 477
rect 252 443 266 477
rect 206 386 266 443
rect 206 352 218 386
rect 252 352 266 386
rect 206 297 266 352
rect 302 485 362 497
rect 302 451 314 485
rect 348 451 362 485
rect 302 408 362 451
rect 302 374 314 408
rect 348 374 362 408
rect 302 297 362 374
rect 398 477 458 497
rect 398 443 410 477
rect 444 443 458 477
rect 398 386 458 443
rect 398 352 410 386
rect 444 352 458 386
rect 398 297 458 352
rect 494 481 553 497
rect 494 447 506 481
rect 540 447 553 481
rect 494 297 553 447
rect 589 477 684 497
rect 589 443 622 477
rect 656 443 684 477
rect 589 297 684 443
rect 720 489 780 497
rect 720 455 733 489
rect 767 455 780 489
rect 720 297 780 455
rect 816 477 879 497
rect 816 443 833 477
rect 867 443 879 477
rect 816 297 879 443
rect 915 489 974 497
rect 915 455 928 489
rect 962 455 974 489
rect 915 297 974 455
rect 1010 297 1070 497
rect 1106 489 1166 497
rect 1106 455 1119 489
rect 1153 455 1166 489
rect 1106 421 1166 455
rect 1106 387 1119 421
rect 1153 387 1166 421
rect 1106 297 1166 387
rect 1202 297 1262 497
rect 1298 485 1353 497
rect 1298 451 1311 485
rect 1345 451 1353 485
rect 1298 417 1353 451
rect 1298 383 1311 417
rect 1345 383 1353 417
rect 1298 297 1353 383
<< ndiffc >>
rect 35 59 69 93
rect 129 67 163 101
rect 223 55 257 89
rect 317 67 351 101
rect 411 59 445 93
rect 532 59 566 93
rect 704 129 738 163
rect 911 135 945 169
rect 911 67 945 101
rect 1009 55 1043 89
rect 1119 123 1153 157
rect 1119 55 1153 89
rect 1215 55 1249 89
rect 1311 127 1345 161
rect 1311 59 1345 93
<< pdiffc >>
rect 122 451 156 485
rect 122 374 156 408
rect 218 443 252 477
rect 218 352 252 386
rect 314 451 348 485
rect 314 374 348 408
rect 410 443 444 477
rect 410 352 444 386
rect 506 447 540 481
rect 622 443 656 477
rect 733 455 767 489
rect 833 443 867 477
rect 928 455 962 489
rect 1119 455 1153 489
rect 1119 387 1153 421
rect 1311 451 1345 485
rect 1311 383 1345 417
<< poly >>
rect 170 497 206 523
rect 266 497 302 523
rect 362 497 398 523
rect 458 497 494 523
rect 553 497 589 523
rect 684 497 720 523
rect 780 497 816 523
rect 879 497 915 523
rect 974 497 1010 523
rect 1070 497 1106 523
rect 1166 497 1202 523
rect 1262 497 1298 523
rect 170 282 206 297
rect 266 282 302 297
rect 362 282 398 297
rect 458 282 494 297
rect 553 282 589 297
rect 684 282 720 297
rect 780 282 816 297
rect 879 282 915 297
rect 974 282 1010 297
rect 1070 282 1106 297
rect 1166 282 1202 297
rect 1262 282 1298 297
rect 168 265 208 282
rect 264 265 304 282
rect 360 265 400 282
rect 456 265 496 282
rect 551 265 591 282
rect 682 265 722 282
rect 778 265 818 282
rect 877 265 917 282
rect 972 265 1012 282
rect 1068 265 1108 282
rect 1164 265 1204 282
rect 1260 265 1300 282
rect 80 249 496 265
rect 80 215 133 249
rect 167 215 211 249
rect 245 215 279 249
rect 313 215 357 249
rect 391 215 435 249
rect 469 215 496 249
rect 80 199 496 215
rect 548 249 607 265
rect 548 215 558 249
rect 592 215 607 249
rect 548 199 607 215
rect 80 177 110 199
rect 174 177 204 199
rect 268 177 298 199
rect 362 177 392 199
rect 577 177 607 199
rect 649 249 818 265
rect 649 215 680 249
rect 714 215 758 249
rect 792 215 818 249
rect 649 199 818 215
rect 860 249 917 265
rect 860 215 870 249
rect 904 215 917 249
rect 860 199 917 215
rect 960 249 1026 265
rect 960 215 981 249
rect 1015 215 1026 249
rect 960 199 1026 215
rect 1068 249 1218 265
rect 1068 215 1084 249
rect 1118 215 1162 249
rect 1196 215 1218 249
rect 1068 199 1218 215
rect 1260 249 1350 265
rect 1260 215 1282 249
rect 1316 215 1350 249
rect 1260 199 1350 215
rect 649 177 679 199
rect 788 177 818 199
rect 865 177 895 199
rect 960 177 990 199
rect 1068 177 1098 199
rect 1164 177 1194 199
rect 1260 177 1290 199
rect 80 21 110 47
rect 174 21 204 47
rect 268 21 298 47
rect 362 21 392 47
rect 577 21 607 47
rect 649 21 679 47
rect 788 21 818 47
rect 865 21 895 47
rect 960 21 990 47
rect 1068 21 1098 47
rect 1164 21 1194 47
rect 1260 21 1290 47
<< polycont >>
rect 133 215 167 249
rect 211 215 245 249
rect 279 215 313 249
rect 357 215 391 249
rect 435 215 469 249
rect 558 215 592 249
rect 680 215 714 249
rect 758 215 792 249
rect 870 215 904 249
rect 981 215 1015 249
rect 1084 215 1118 249
rect 1162 215 1196 249
rect 1282 215 1316 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 96 485 172 527
rect 96 451 122 485
rect 156 451 172 485
rect 96 408 172 451
rect 96 374 122 408
rect 156 374 172 408
rect 216 477 252 493
rect 216 443 218 477
rect 216 386 252 443
rect 216 352 218 386
rect 288 485 364 527
rect 288 451 314 485
rect 348 451 364 485
rect 288 408 364 451
rect 288 374 314 408
rect 348 374 364 408
rect 408 477 446 493
rect 408 443 410 477
rect 444 443 446 477
rect 408 386 446 443
rect 480 481 556 527
rect 480 447 506 481
rect 540 447 556 481
rect 480 440 556 447
rect 600 477 672 493
rect 600 443 622 477
rect 656 443 672 477
rect 600 405 672 443
rect 707 489 783 527
rect 707 455 733 489
rect 767 455 783 489
rect 707 439 783 455
rect 817 477 883 493
rect 817 443 833 477
rect 867 443 883 477
rect 817 405 883 443
rect 919 489 972 527
rect 919 455 928 489
rect 962 455 972 489
rect 919 439 972 455
rect 1093 489 1169 493
rect 1093 455 1119 489
rect 1153 455 1169 489
rect 1093 421 1169 455
rect 1093 405 1119 421
rect 216 340 252 352
rect 408 352 410 386
rect 444 352 446 386
rect 408 340 446 352
rect 17 287 446 340
rect 480 387 1119 405
rect 1153 387 1169 421
rect 480 371 1169 387
rect 1285 485 1361 527
rect 1285 451 1311 485
rect 1345 451 1361 485
rect 1285 417 1361 451
rect 1285 383 1311 417
rect 1345 383 1361 417
rect 17 161 73 287
rect 480 253 524 371
rect 107 249 524 253
rect 107 215 133 249
rect 167 215 211 249
rect 245 215 279 249
rect 313 215 357 249
rect 391 215 435 249
rect 469 215 524 249
rect 107 213 524 215
rect 480 163 524 213
rect 558 289 920 337
rect 558 249 617 289
rect 592 215 617 249
rect 558 199 617 215
rect 651 249 818 255
rect 651 215 680 249
rect 714 215 758 249
rect 792 215 818 249
rect 651 207 818 215
rect 854 249 920 289
rect 854 215 870 249
rect 904 215 920 249
rect 854 207 920 215
rect 965 299 1363 337
rect 965 249 1031 299
rect 965 215 981 249
rect 1015 215 1031 249
rect 965 207 1031 215
rect 1068 249 1223 265
rect 1068 215 1084 249
rect 1118 215 1162 249
rect 1196 215 1223 249
rect 1068 207 1223 215
rect 1260 249 1363 299
rect 1260 215 1282 249
rect 1316 215 1363 249
rect 1260 207 1363 215
rect 895 169 1361 173
rect 17 127 351 161
rect 480 129 704 163
rect 738 129 764 163
rect 480 127 764 129
rect 895 135 911 169
rect 945 161 1361 169
rect 945 157 1311 161
rect 945 139 1119 157
rect 945 135 961 139
rect 129 123 351 127
rect 129 101 163 123
rect 19 59 35 93
rect 69 59 85 93
rect 19 17 85 59
rect 317 101 351 123
rect 129 51 163 67
rect 207 55 223 89
rect 257 55 273 89
rect 207 17 273 55
rect 895 101 961 135
rect 1093 123 1119 139
rect 1153 139 1311 157
rect 1153 123 1169 139
rect 895 93 911 101
rect 317 51 351 67
rect 385 59 411 93
rect 445 59 468 93
rect 385 17 468 59
rect 516 59 532 93
rect 566 67 911 93
rect 945 67 961 101
rect 566 59 961 67
rect 516 51 961 59
rect 996 89 1059 105
rect 996 55 1009 89
rect 1043 55 1059 89
rect 996 17 1059 55
rect 1093 89 1169 123
rect 1285 127 1311 139
rect 1345 127 1361 161
rect 1093 55 1119 89
rect 1153 55 1169 89
rect 1093 51 1169 55
rect 1213 89 1251 105
rect 1213 55 1215 89
rect 1249 55 1251 89
rect 1213 17 1251 55
rect 1285 93 1361 127
rect 1285 59 1311 93
rect 1345 59 1361 93
rect 1285 51 1361 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
<< metal1 >>
rect 0 561 1380 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 0 496 1380 527
rect 0 17 1380 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
rect 0 -48 1380 -17
<< labels >>
flabel corelocali s 1316 289 1350 323 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 29 153 63 187 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 671 221 705 255 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 1129 221 1163 255 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 854 289 888 323 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
rlabel comment s 0 0 0 0 4 o211a_4
<< properties >>
string FIXED_BBOX 0 0 1380 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2584542
string GDS_START 2575002
<< end >>
