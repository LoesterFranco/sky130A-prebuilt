magic
tech sky130A
magscale 1 2
timestamp 1599588238
<< locali >>
rect 121 310 199 412
rect 146 150 199 310
rect 301 252 359 356
rect 393 290 459 356
rect 501 290 567 356
rect 601 252 743 356
rect 777 288 843 356
rect 146 70 212 150
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 43 514 109 649
rect 223 514 289 649
rect 327 514 393 596
rect 427 548 533 649
rect 567 514 633 596
rect 21 446 267 480
rect 327 458 633 514
rect 21 270 87 446
rect 233 424 267 446
rect 741 424 807 596
rect 60 17 110 226
rect 233 390 807 424
rect 233 218 267 390
rect 233 184 808 218
rect 246 17 326 150
rect 526 70 600 184
rect 634 17 708 150
rect 742 70 808 184
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel locali s 501 290 567 356 6 A1
port 1 nsew signal input
rlabel locali s 393 290 459 356 6 A2
port 2 nsew signal input
rlabel locali s 301 252 359 356 6 A3
port 3 nsew signal input
rlabel locali s 601 252 743 356 6 B1
port 4 nsew signal input
rlabel locali s 777 288 843 356 6 C1
port 5 nsew signal input
rlabel locali s 146 150 199 310 6 X
port 6 nsew signal output
rlabel locali s 146 70 212 150 6 X
port 6 nsew signal output
rlabel locali s 121 310 199 412 6 X
port 6 nsew signal output
rlabel metal1 s 0 -49 864 49 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 617 864 715 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3601780
string GDS_START 3594564
<< end >>
