magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 111 299 179 493
rect 306 459 775 493
rect 111 51 161 299
rect 306 265 346 459
rect 291 199 346 265
rect 448 323 707 357
rect 448 162 482 323
rect 550 51 615 283
rect 649 51 707 323
rect 741 326 775 459
rect 741 288 891 326
rect 853 211 891 288
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 27 299 76 527
rect 215 299 265 527
rect 27 17 77 131
rect 195 165 229 265
rect 380 391 669 425
rect 380 165 414 391
rect 195 131 414 165
rect 379 124 414 131
rect 195 17 271 97
rect 379 51 516 124
rect 809 367 855 527
rect 889 367 969 493
rect 757 173 791 237
rect 935 173 969 367
rect 757 139 969 173
rect 742 17 845 105
rect 899 51 948 139
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
rlabel locali s 550 51 615 283 6 A0
port 1 nsew signal input
rlabel locali s 649 51 707 323 6 A1
port 2 nsew signal input
rlabel locali s 448 323 707 357 6 A1
port 2 nsew signal input
rlabel locali s 448 162 482 323 6 A1
port 2 nsew signal input
rlabel locali s 853 211 891 288 6 S
port 3 nsew signal input
rlabel locali s 741 326 775 459 6 S
port 3 nsew signal input
rlabel locali s 741 288 891 326 6 S
port 3 nsew signal input
rlabel locali s 306 459 775 493 6 S
port 3 nsew signal input
rlabel locali s 306 265 346 459 6 S
port 3 nsew signal input
rlabel locali s 291 199 346 265 6 S
port 3 nsew signal input
rlabel locali s 111 299 179 493 6 X
port 4 nsew signal output
rlabel locali s 111 51 161 299 6 X
port 4 nsew signal output
rlabel metal1 s 0 -48 1012 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 1012 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1012 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3284060
string GDS_START 3276300
<< end >>
