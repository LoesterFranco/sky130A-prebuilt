magic
tech sky130A
magscale 1 2
timestamp 1604502705
<< nwell >>
rect -38 332 1958 704
rect 136 305 852 332
<< pwell >>
rect 0 0 1920 49
<< scnmos >>
rect 84 74 114 202
rect 234 74 264 202
rect 312 74 342 202
rect 420 74 450 202
rect 600 74 630 202
rect 738 74 768 202
rect 816 74 846 202
rect 949 74 979 202
rect 1027 74 1057 202
rect 1308 125 1338 253
rect 1396 125 1426 253
rect 1677 104 1707 232
rect 1791 84 1821 232
<< pmoshvt >>
rect 108 368 138 568
rect 225 341 255 541
rect 417 341 447 541
rect 507 341 537 541
rect 609 341 639 541
rect 733 341 763 541
rect 834 387 864 587
rect 1035 387 1065 587
rect 1119 387 1149 587
rect 1321 392 1351 592
rect 1421 392 1451 592
rect 1643 387 1673 587
rect 1801 368 1831 592
<< ndiff >>
rect 27 190 84 202
rect 27 156 39 190
rect 73 156 84 190
rect 27 120 84 156
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 127 234 202
rect 114 93 162 127
rect 196 93 234 127
rect 114 74 234 93
rect 264 74 312 202
rect 342 179 420 202
rect 342 145 375 179
rect 409 145 420 179
rect 342 74 420 145
rect 450 74 600 202
rect 630 120 738 202
rect 630 86 667 120
rect 701 86 738 120
rect 630 74 738 86
rect 768 74 816 202
rect 846 125 949 202
rect 846 91 880 125
rect 914 91 949 125
rect 846 74 949 91
rect 979 74 1027 202
rect 1057 184 1114 202
rect 1258 194 1308 253
rect 1057 150 1068 184
rect 1102 150 1114 184
rect 1057 116 1114 150
rect 1057 82 1068 116
rect 1102 82 1114 116
rect 1057 74 1114 82
rect 1199 181 1308 194
rect 1199 147 1213 181
rect 1247 147 1308 181
rect 1199 125 1308 147
rect 1338 241 1396 253
rect 1338 207 1350 241
rect 1384 207 1396 241
rect 1338 125 1396 207
rect 1426 171 1483 253
rect 1426 137 1437 171
rect 1471 137 1483 171
rect 1426 125 1483 137
rect 1620 220 1677 232
rect 1620 186 1632 220
rect 1666 186 1677 220
rect 1620 150 1677 186
rect 1199 89 1293 125
rect 1199 55 1213 89
rect 1247 55 1293 89
rect 1199 43 1293 55
rect 1620 116 1632 150
rect 1666 116 1677 150
rect 1620 104 1677 116
rect 1707 220 1791 232
rect 1707 186 1732 220
rect 1766 186 1791 220
rect 1707 150 1791 186
rect 1707 116 1732 150
rect 1766 116 1791 150
rect 1707 104 1791 116
rect 1741 84 1791 104
rect 1821 220 1878 232
rect 1821 186 1832 220
rect 1866 186 1878 220
rect 1821 130 1878 186
rect 1821 96 1832 130
rect 1866 96 1878 130
rect 1821 84 1878 96
<< pdiff >>
rect 49 560 108 568
rect 49 526 61 560
rect 95 526 108 560
rect 49 492 108 526
rect 49 458 61 492
rect 95 458 108 492
rect 49 424 108 458
rect 49 390 61 424
rect 95 390 108 424
rect 49 368 108 390
rect 138 560 207 568
rect 138 526 161 560
rect 195 541 207 560
rect 657 585 715 597
rect 657 551 669 585
rect 703 551 715 585
rect 657 541 715 551
rect 781 541 834 587
rect 195 526 225 541
rect 138 492 225 526
rect 138 458 161 492
rect 195 458 225 492
rect 138 424 225 458
rect 138 390 161 424
rect 195 390 225 424
rect 138 368 225 390
rect 172 341 225 368
rect 255 341 417 541
rect 447 529 507 541
rect 447 495 460 529
rect 494 495 507 529
rect 447 458 507 495
rect 447 424 460 458
rect 494 424 507 458
rect 447 387 507 424
rect 447 353 460 387
rect 494 353 507 387
rect 447 341 507 353
rect 537 341 609 541
rect 639 341 733 541
rect 763 387 834 541
rect 864 531 1035 587
rect 864 497 877 531
rect 911 497 988 531
rect 1022 497 1035 531
rect 864 433 1035 497
rect 864 399 877 433
rect 911 399 988 433
rect 1022 399 1035 433
rect 864 387 1035 399
rect 1065 387 1119 587
rect 1149 572 1208 587
rect 1149 538 1162 572
rect 1196 538 1208 572
rect 1149 387 1208 538
rect 1262 580 1321 592
rect 1262 546 1274 580
rect 1308 546 1321 580
rect 1262 510 1321 546
rect 1262 476 1274 510
rect 1308 476 1321 510
rect 1262 440 1321 476
rect 1262 406 1274 440
rect 1308 406 1321 440
rect 1262 392 1321 406
rect 1351 580 1421 592
rect 1351 546 1374 580
rect 1408 546 1421 580
rect 1351 509 1421 546
rect 1351 475 1374 509
rect 1408 475 1421 509
rect 1351 438 1421 475
rect 1351 404 1374 438
rect 1408 404 1421 438
rect 1351 392 1421 404
rect 1451 531 1520 592
rect 1742 587 1801 592
rect 1451 497 1474 531
rect 1508 497 1520 531
rect 1451 439 1520 497
rect 1451 405 1474 439
rect 1508 405 1520 439
rect 1451 392 1520 405
rect 1574 531 1643 587
rect 1574 497 1586 531
rect 1620 497 1643 531
rect 1574 440 1643 497
rect 1574 406 1586 440
rect 1620 406 1643 440
rect 763 341 816 387
rect 1574 387 1643 406
rect 1673 580 1801 587
rect 1673 546 1754 580
rect 1788 546 1801 580
rect 1673 508 1801 546
rect 1673 474 1754 508
rect 1788 474 1801 508
rect 1673 387 1801 474
rect 1748 368 1801 387
rect 1831 562 1893 592
rect 1831 528 1845 562
rect 1879 528 1893 562
rect 1831 368 1893 528
<< ndiffc >>
rect 39 156 73 190
rect 39 86 73 120
rect 162 93 196 127
rect 375 145 409 179
rect 667 86 701 120
rect 880 91 914 125
rect 1068 150 1102 184
rect 1068 82 1102 116
rect 1213 147 1247 181
rect 1350 207 1384 241
rect 1437 137 1471 171
rect 1632 186 1666 220
rect 1213 55 1247 89
rect 1632 116 1666 150
rect 1732 186 1766 220
rect 1732 116 1766 150
rect 1832 186 1866 220
rect 1832 96 1866 130
<< pdiffc >>
rect 61 526 95 560
rect 61 458 95 492
rect 61 390 95 424
rect 161 526 195 560
rect 669 551 703 585
rect 161 458 195 492
rect 161 390 195 424
rect 460 495 494 529
rect 460 424 494 458
rect 460 353 494 387
rect 877 497 911 531
rect 988 497 1022 531
rect 877 399 911 433
rect 988 399 1022 433
rect 1162 538 1196 572
rect 1274 546 1308 580
rect 1274 476 1308 510
rect 1274 406 1308 440
rect 1374 546 1408 580
rect 1374 475 1408 509
rect 1374 404 1408 438
rect 1474 497 1508 531
rect 1474 405 1508 439
rect 1586 497 1620 531
rect 1586 406 1620 440
rect 1754 546 1788 580
rect 1754 474 1788 508
rect 1845 528 1879 562
<< poly >>
rect 105 615 867 645
rect 105 583 141 615
rect 108 568 138 583
rect 225 541 255 567
rect 414 556 450 615
rect 831 602 867 615
rect 834 587 864 602
rect 1035 587 1065 613
rect 1119 587 1149 613
rect 1321 592 1351 618
rect 1421 592 1451 618
rect 417 541 447 556
rect 507 541 537 567
rect 609 541 639 567
rect 733 541 763 567
rect 108 353 138 368
rect 105 309 141 353
rect 1643 587 1673 613
rect 1801 592 1831 618
rect 834 372 864 387
rect 1035 372 1065 387
rect 1119 372 1149 387
rect 1321 377 1351 392
rect 1421 377 1451 392
rect 831 368 867 372
rect 225 326 255 341
rect 417 326 447 341
rect 507 326 537 341
rect 609 326 639 341
rect 733 326 763 341
rect 831 338 960 368
rect 1032 355 1068 372
rect 1119 355 1152 372
rect 222 309 258 326
rect 84 293 156 309
rect 84 259 106 293
rect 140 259 156 293
rect 84 243 156 259
rect 198 293 264 309
rect 198 259 214 293
rect 248 259 264 293
rect 198 243 264 259
rect 84 202 114 243
rect 234 202 264 243
rect 306 290 372 306
rect 306 256 322 290
rect 356 256 372 290
rect 306 240 372 256
rect 312 202 342 240
rect 414 217 450 326
rect 504 290 540 326
rect 606 309 642 326
rect 730 309 766 326
rect 600 293 666 309
rect 492 274 558 290
rect 492 240 508 274
rect 542 240 558 274
rect 492 224 558 240
rect 600 259 616 293
rect 650 259 666 293
rect 600 243 666 259
rect 708 293 774 309
rect 708 259 724 293
rect 758 259 774 293
rect 708 243 774 259
rect 816 274 882 290
rect 420 202 450 217
rect 600 202 630 243
rect 738 202 768 243
rect 816 240 832 274
rect 866 240 882 274
rect 816 224 882 240
rect 930 247 960 338
rect 1002 339 1068 355
rect 1002 305 1018 339
rect 1052 305 1068 339
rect 1002 289 1068 305
rect 1122 339 1236 355
rect 1122 305 1186 339
rect 1220 305 1236 339
rect 1122 247 1236 305
rect 1318 298 1354 377
rect 1418 318 1454 377
rect 1643 372 1673 387
rect 1526 339 1592 355
rect 1526 318 1542 339
rect 1308 268 1354 298
rect 1396 305 1542 318
rect 1576 305 1592 339
rect 1640 336 1676 372
rect 1801 353 1831 368
rect 1798 336 1834 353
rect 1396 288 1592 305
rect 1641 320 1707 336
rect 1308 253 1338 268
rect 1396 253 1426 288
rect 1641 286 1657 320
rect 1691 286 1707 320
rect 1641 270 1707 286
rect 1749 320 1834 336
rect 1749 286 1765 320
rect 1799 286 1834 320
rect 1749 270 1834 286
rect 816 202 846 224
rect 930 217 979 247
rect 949 202 979 217
rect 1027 217 1236 247
rect 1027 202 1057 217
rect 1677 232 1707 270
rect 1791 232 1821 270
rect 84 48 114 74
rect 234 48 264 74
rect 312 48 342 74
rect 420 48 450 74
rect 600 48 630 74
rect 738 48 768 74
rect 816 48 846 74
rect 949 48 979 74
rect 1027 48 1057 74
rect 1308 51 1338 125
rect 1396 99 1426 125
rect 1677 51 1707 104
rect 1791 58 1821 84
rect 1308 21 1707 51
<< polycont >>
rect 106 259 140 293
rect 214 259 248 293
rect 322 256 356 290
rect 508 240 542 274
rect 616 259 650 293
rect 724 259 758 293
rect 832 240 866 274
rect 1018 305 1052 339
rect 1186 305 1220 339
rect 1542 305 1576 339
rect 1657 286 1691 320
rect 1765 286 1799 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 22 560 111 576
rect 22 526 61 560
rect 95 526 111 560
rect 22 492 111 526
rect 22 458 61 492
rect 95 458 111 492
rect 22 424 111 458
rect 22 390 61 424
rect 95 390 111 424
rect 145 560 211 649
rect 145 526 161 560
rect 195 526 211 560
rect 653 585 719 649
rect 653 551 669 585
rect 703 551 719 585
rect 145 492 211 526
rect 145 458 161 492
rect 195 458 211 492
rect 145 424 211 458
rect 145 390 161 424
rect 195 390 211 424
rect 406 529 510 545
rect 653 535 719 551
rect 759 581 1110 615
rect 406 495 460 529
rect 494 501 510 529
rect 759 501 804 581
rect 494 495 804 501
rect 406 467 804 495
rect 861 531 1033 547
rect 861 497 877 531
rect 911 497 988 531
rect 1022 497 1033 531
rect 406 458 510 467
rect 406 424 460 458
rect 494 424 510 458
rect 861 433 1033 497
rect 1070 501 1110 581
rect 1146 572 1212 649
rect 1146 538 1162 572
rect 1196 538 1212 572
rect 1146 535 1212 538
rect 1258 580 1324 596
rect 1258 546 1274 580
rect 1308 546 1324 580
rect 1258 510 1324 546
rect 1258 501 1274 510
rect 1070 476 1274 501
rect 1308 476 1324 510
rect 1070 467 1324 476
rect 1258 440 1324 467
rect 22 206 56 390
rect 406 387 510 424
rect 90 293 164 356
rect 90 259 106 293
rect 140 259 164 293
rect 90 243 164 259
rect 198 293 264 356
rect 406 353 460 387
rect 494 353 510 387
rect 406 337 510 353
rect 198 259 214 293
rect 248 259 264 293
rect 198 243 264 259
rect 306 290 372 306
rect 306 256 322 290
rect 356 256 372 290
rect 306 240 372 256
rect 306 206 340 240
rect 406 206 440 337
rect 600 293 666 430
rect 22 190 340 206
rect 22 156 39 190
rect 73 172 340 190
rect 73 156 89 172
rect 22 120 89 156
rect 22 86 39 120
rect 73 86 89 120
rect 22 70 89 86
rect 140 127 218 136
rect 140 93 162 127
rect 196 93 218 127
rect 140 17 218 93
rect 306 85 340 172
rect 375 179 440 206
rect 409 145 440 179
rect 375 119 440 145
rect 492 274 558 290
rect 492 240 508 274
rect 542 240 558 274
rect 600 259 616 293
rect 650 259 666 293
rect 600 243 666 259
rect 700 293 774 430
rect 861 399 877 433
rect 911 399 988 433
rect 1022 399 1136 433
rect 700 259 724 293
rect 758 259 774 293
rect 916 339 1068 355
rect 916 305 1018 339
rect 1052 305 1068 339
rect 700 243 774 259
rect 816 274 882 290
rect 492 209 558 240
rect 816 240 832 274
rect 866 240 882 274
rect 816 209 882 240
rect 916 289 1068 305
rect 916 209 950 289
rect 1102 255 1136 399
rect 1258 406 1274 440
rect 1308 406 1324 440
rect 1258 390 1324 406
rect 1358 581 1704 615
rect 1358 580 1424 581
rect 1358 546 1374 580
rect 1408 546 1424 580
rect 1358 509 1424 546
rect 1358 475 1374 509
rect 1408 475 1424 509
rect 1358 438 1424 475
rect 1358 404 1374 438
rect 1408 404 1424 438
rect 1170 339 1236 356
rect 1170 305 1186 339
rect 1220 305 1236 339
rect 1170 289 1236 305
rect 492 175 950 209
rect 984 221 1247 255
rect 492 85 526 175
rect 984 141 1018 221
rect 306 51 526 85
rect 625 120 743 136
rect 625 86 667 120
rect 701 86 743 120
rect 625 17 743 86
rect 842 125 1018 141
rect 842 91 880 125
rect 914 91 1018 125
rect 842 75 1018 91
rect 1052 184 1118 187
rect 1052 150 1068 184
rect 1102 150 1118 184
rect 1052 116 1118 150
rect 1052 82 1068 116
rect 1102 82 1118 116
rect 1052 17 1118 82
rect 1197 181 1247 221
rect 1197 147 1213 181
rect 1197 89 1247 147
rect 1281 157 1315 390
rect 1358 257 1424 404
rect 1349 241 1424 257
rect 1349 207 1350 241
rect 1384 223 1424 241
rect 1458 531 1524 547
rect 1458 497 1474 531
rect 1508 497 1524 531
rect 1458 439 1524 497
rect 1458 405 1474 439
rect 1508 405 1524 439
rect 1458 389 1524 405
rect 1570 531 1636 547
rect 1570 497 1586 531
rect 1620 497 1636 531
rect 1570 440 1636 497
rect 1570 406 1586 440
rect 1620 406 1636 440
rect 1570 390 1636 406
rect 1670 424 1704 581
rect 1738 580 1804 649
rect 1738 546 1754 580
rect 1788 546 1804 580
rect 1738 508 1804 546
rect 1844 562 1897 578
rect 1844 528 1845 562
rect 1879 528 1897 562
rect 1844 512 1897 528
rect 1738 474 1754 508
rect 1788 474 1804 508
rect 1738 458 1804 474
rect 1670 390 1783 424
rect 1458 255 1492 389
rect 1570 355 1607 390
rect 1526 339 1607 355
rect 1526 305 1542 339
rect 1576 305 1607 339
rect 1526 289 1607 305
rect 1384 207 1385 223
rect 1458 221 1539 255
rect 1349 191 1385 207
rect 1421 171 1471 187
rect 1421 157 1437 171
rect 1281 137 1437 157
rect 1281 123 1471 137
rect 1421 121 1471 123
rect 1197 55 1213 89
rect 1247 87 1297 89
rect 1505 87 1539 221
rect 1573 236 1607 289
rect 1641 320 1707 356
rect 1641 286 1657 320
rect 1691 286 1707 320
rect 1641 270 1707 286
rect 1749 336 1783 390
rect 1749 320 1815 336
rect 1749 286 1765 320
rect 1799 286 1815 320
rect 1749 270 1815 286
rect 1849 236 1897 512
rect 1573 220 1682 236
rect 1573 186 1632 220
rect 1666 186 1682 220
rect 1573 150 1682 186
rect 1573 116 1632 150
rect 1666 116 1682 150
rect 1573 100 1682 116
rect 1716 220 1782 236
rect 1716 186 1732 220
rect 1766 186 1782 220
rect 1716 150 1782 186
rect 1716 116 1732 150
rect 1766 116 1782 150
rect 1247 55 1539 87
rect 1197 53 1539 55
rect 1716 17 1782 116
rect 1816 220 1897 236
rect 1816 186 1832 220
rect 1866 186 1897 220
rect 1816 130 1897 186
rect 1816 96 1832 130
rect 1866 96 1897 130
rect 1816 80 1897 96
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
<< metal1 >>
rect 0 683 1920 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 0 617 1920 649
rect 0 17 1920 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
rect 0 -49 1920 -17
<< labels >>
rlabel comment s 0 0 0 0 4 mux4_1
flabel pwell s 0 0 1920 49 0 FreeSans 200 0 0 0 VNB
port 8 nsew
flabel nbase s 0 617 1920 666 0 FreeSans 200 0 0 0 VPB
port 9 nsew
flabel metal1 s 0 617 1920 666 0 FreeSans 340 0 0 0 VPWR
port 10 nsew
flabel metal1 s 0 0 1920 49 0 FreeSans 340 0 0 0 VGND
port 7 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 S0
port 5 nsew
flabel corelocali s 1183 316 1217 350 0 FreeSans 340 0 0 0 A3
port 4 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 A2
port 3 nsew
flabel corelocali s 703 390 737 424 0 FreeSans 340 0 0 0 A2
port 3 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 A1
port 2 nsew
flabel corelocali s 607 390 641 424 0 FreeSans 340 0 0 0 A1
port 2 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A0
port 1 nsew
flabel corelocali s 1663 316 1697 350 0 FreeSans 340 0 0 0 S1
port 6 nsew
flabel corelocali s 1855 94 1889 128 0 FreeSans 340 0 0 0 X
port 11 nsew
flabel corelocali s 1855 168 1889 202 0 FreeSans 340 0 0 0 X
port 11 nsew
flabel corelocali s 1855 242 1889 276 0 FreeSans 340 0 0 0 X
port 11 nsew
flabel corelocali s 1855 316 1889 350 0 FreeSans 340 0 0 0 X
port 11 nsew
flabel corelocali s 1855 390 1889 424 0 FreeSans 340 0 0 0 X
port 11 nsew
flabel corelocali s 1855 464 1889 498 0 FreeSans 340 0 0 0 X
port 11 nsew
flabel corelocali s 1855 538 1889 572 0 FreeSans 340 0 0 0 X
port 11 nsew
<< properties >>
string FIXED_BBOX 0 0 1920 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1685028
string GDS_START 1670566
<< end >>
