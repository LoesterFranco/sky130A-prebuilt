magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 2246 704
rect 188 314 1286 332
rect 1078 305 1286 314
<< pwell >>
rect 0 0 2208 49
<< scnmos >>
rect 84 74 114 158
rect 282 74 312 222
rect 368 74 398 222
rect 574 74 604 158
rect 710 74 740 158
rect 788 74 818 158
rect 997 118 1027 202
rect 1069 118 1099 202
rect 1185 74 1215 202
rect 1290 74 1320 202
rect 1392 74 1422 158
rect 1470 74 1500 158
rect 1548 74 1578 158
rect 1761 74 1791 158
rect 1959 74 1989 184
rect 2075 74 2105 222
<< pmoshvt >>
rect 84 508 114 592
rect 281 350 311 574
rect 371 350 401 574
rect 579 463 609 547
rect 679 463 709 547
rect 763 463 793 547
rect 928 463 958 547
rect 1018 463 1048 547
rect 1167 341 1197 541
rect 1268 392 1298 592
rect 1427 508 1457 592
rect 1511 508 1541 592
rect 1601 508 1631 592
rect 1796 508 1826 592
rect 1990 403 2020 571
rect 2094 368 2124 592
<< ndiff >>
rect 225 196 282 222
rect 225 162 237 196
rect 271 162 282 196
rect 27 133 84 158
rect 27 99 39 133
rect 73 99 84 133
rect 27 74 84 99
rect 114 133 171 158
rect 114 99 125 133
rect 159 99 171 133
rect 114 74 171 99
rect 225 120 282 162
rect 225 86 237 120
rect 271 86 282 120
rect 225 74 282 86
rect 312 186 368 222
rect 312 152 323 186
rect 357 152 368 186
rect 312 116 368 152
rect 312 82 323 116
rect 357 82 368 116
rect 312 74 368 82
rect 398 202 451 222
rect 398 168 409 202
rect 443 168 451 202
rect 398 120 451 168
rect 398 86 409 120
rect 443 86 451 120
rect 398 74 451 86
rect 505 169 559 181
rect 505 135 513 169
rect 547 158 559 169
rect 941 177 997 202
rect 547 135 574 158
rect 505 74 574 135
rect 604 133 710 158
rect 604 99 665 133
rect 699 99 710 133
rect 604 74 710 99
rect 740 74 788 158
rect 818 120 887 158
rect 818 86 835 120
rect 869 86 887 120
rect 941 143 952 177
rect 986 143 997 177
rect 941 118 997 143
rect 1027 118 1069 202
rect 1099 190 1185 202
rect 1099 156 1140 190
rect 1174 156 1185 190
rect 1099 120 1185 156
rect 1099 118 1140 120
rect 818 74 887 86
rect 1128 86 1140 118
rect 1174 86 1185 120
rect 1128 74 1185 86
rect 1215 74 1290 202
rect 1320 169 1377 202
rect 1320 135 1331 169
rect 1365 158 1377 169
rect 2004 203 2075 222
rect 2004 184 2016 203
rect 1365 135 1392 158
rect 1320 74 1392 135
rect 1422 74 1470 158
rect 1500 74 1548 158
rect 1578 120 1761 158
rect 1578 86 1590 120
rect 1624 86 1702 120
rect 1736 86 1761 120
rect 1578 74 1761 86
rect 1791 133 1848 158
rect 1791 99 1802 133
rect 1836 99 1848 133
rect 1791 74 1848 99
rect 1902 138 1959 184
rect 1902 104 1914 138
rect 1948 104 1959 138
rect 1902 74 1959 104
rect 1989 169 2016 184
rect 2050 169 2075 203
rect 1989 116 2075 169
rect 1989 82 2016 116
rect 2050 82 2075 116
rect 1989 74 2075 82
rect 2105 194 2162 222
rect 2105 160 2116 194
rect 2150 160 2162 194
rect 2105 120 2162 160
rect 2105 86 2116 120
rect 2150 86 2162 120
rect 2105 74 2162 86
<< pdiff >>
rect 27 567 84 592
rect 27 533 37 567
rect 71 533 84 567
rect 27 508 84 533
rect 114 572 170 592
rect 114 538 127 572
rect 161 538 170 572
rect 114 508 170 538
rect 224 396 281 574
rect 224 362 234 396
rect 268 362 281 396
rect 224 350 281 362
rect 311 555 371 574
rect 311 521 324 555
rect 358 521 371 555
rect 311 350 371 521
rect 401 546 460 574
rect 401 512 414 546
rect 448 512 460 546
rect 401 350 460 512
rect 1095 582 1149 594
rect 1095 548 1107 582
rect 1141 548 1149 582
rect 1095 547 1149 548
rect 520 520 579 547
rect 520 486 532 520
rect 566 486 579 520
rect 520 463 579 486
rect 609 520 679 547
rect 609 486 632 520
rect 666 486 679 520
rect 609 463 679 486
rect 709 463 763 547
rect 793 535 928 547
rect 793 501 809 535
rect 843 501 928 535
rect 793 463 928 501
rect 958 522 1018 547
rect 958 488 971 522
rect 1005 488 1018 522
rect 958 463 1018 488
rect 1048 541 1149 547
rect 1215 541 1268 592
rect 1048 463 1167 541
rect 1114 341 1167 463
rect 1197 392 1268 541
rect 1298 584 1427 592
rect 1298 550 1311 584
rect 1345 550 1380 584
rect 1414 550 1427 584
rect 1298 516 1427 550
rect 1298 482 1311 516
rect 1345 508 1427 516
rect 1457 508 1511 592
rect 1541 580 1601 592
rect 1541 546 1554 580
rect 1588 546 1601 580
rect 1541 508 1601 546
rect 1631 570 1686 592
rect 1631 536 1644 570
rect 1678 536 1686 570
rect 1631 508 1686 536
rect 1740 580 1796 592
rect 1740 546 1749 580
rect 1783 546 1796 580
rect 1740 508 1796 546
rect 1826 580 1881 592
rect 1826 546 1839 580
rect 1873 546 1881 580
rect 2038 580 2094 592
rect 2038 571 2047 580
rect 1826 508 1881 546
rect 1935 559 1990 571
rect 1935 525 1943 559
rect 1977 525 1990 559
rect 1345 482 1354 508
rect 1298 448 1354 482
rect 1298 414 1312 448
rect 1346 414 1354 448
rect 1298 392 1354 414
rect 1197 341 1250 392
rect 1935 449 1990 525
rect 1935 415 1943 449
rect 1977 415 1990 449
rect 1935 403 1990 415
rect 2020 546 2047 571
rect 2081 546 2094 580
rect 2020 497 2094 546
rect 2020 463 2047 497
rect 2081 463 2094 497
rect 2020 414 2094 463
rect 2020 403 2047 414
rect 2038 380 2047 403
rect 2081 380 2094 414
rect 2038 368 2094 380
rect 2124 580 2181 592
rect 2124 546 2137 580
rect 2171 546 2181 580
rect 2124 497 2181 546
rect 2124 463 2137 497
rect 2171 463 2181 497
rect 2124 414 2181 463
rect 2124 380 2137 414
rect 2171 380 2181 414
rect 2124 368 2181 380
<< ndiffc >>
rect 237 162 271 196
rect 39 99 73 133
rect 125 99 159 133
rect 237 86 271 120
rect 323 152 357 186
rect 323 82 357 116
rect 409 168 443 202
rect 409 86 443 120
rect 513 135 547 169
rect 665 99 699 133
rect 835 86 869 120
rect 952 143 986 177
rect 1140 156 1174 190
rect 1140 86 1174 120
rect 1331 135 1365 169
rect 1590 86 1624 120
rect 1702 86 1736 120
rect 1802 99 1836 133
rect 1914 104 1948 138
rect 2016 169 2050 203
rect 2016 82 2050 116
rect 2116 160 2150 194
rect 2116 86 2150 120
<< pdiffc >>
rect 37 533 71 567
rect 127 538 161 572
rect 234 362 268 396
rect 324 521 358 555
rect 414 512 448 546
rect 1107 548 1141 582
rect 532 486 566 520
rect 632 486 666 520
rect 809 501 843 535
rect 971 488 1005 522
rect 1311 550 1345 584
rect 1380 550 1414 584
rect 1311 482 1345 516
rect 1554 546 1588 580
rect 1644 536 1678 570
rect 1749 546 1783 580
rect 1839 546 1873 580
rect 1943 525 1977 559
rect 1312 414 1346 448
rect 1943 415 1977 449
rect 2047 546 2081 580
rect 2047 463 2081 497
rect 2047 380 2081 414
rect 2137 546 2171 580
rect 2137 463 2171 497
rect 2137 380 2171 414
<< poly >>
rect 84 592 114 618
rect 475 615 1301 645
rect 281 574 311 600
rect 371 574 401 600
rect 84 493 114 508
rect 81 398 117 493
rect 81 382 161 398
rect 81 348 111 382
rect 145 348 161 382
rect 81 314 161 348
rect 281 335 311 350
rect 371 335 401 350
rect 81 280 111 314
rect 145 280 161 314
rect 278 310 314 335
rect 368 318 404 335
rect 475 318 505 615
rect 579 547 609 573
rect 676 562 712 615
rect 1265 607 1301 615
rect 1268 592 1298 607
rect 1427 592 1457 618
rect 1511 592 1541 618
rect 1601 592 1631 618
rect 1796 592 1826 618
rect 679 547 709 562
rect 763 547 793 573
rect 928 547 958 573
rect 1018 547 1048 573
rect 1167 541 1197 567
rect 579 448 609 463
rect 576 421 612 448
rect 679 437 709 463
rect 763 448 793 463
rect 928 448 958 463
rect 1018 448 1048 463
rect 760 425 796 448
rect 81 246 161 280
rect 81 212 111 246
rect 145 212 161 246
rect 260 294 326 310
rect 260 260 276 294
rect 310 260 326 294
rect 260 244 326 260
rect 368 302 505 318
rect 368 268 413 302
rect 447 268 505 302
rect 557 405 623 421
rect 557 371 573 405
rect 607 371 623 405
rect 760 395 841 425
rect 557 337 623 371
rect 811 393 841 395
rect 811 377 877 393
rect 557 303 573 337
rect 607 317 623 337
rect 701 337 767 353
rect 701 317 717 337
rect 607 303 717 317
rect 751 303 767 337
rect 811 343 827 377
rect 861 343 877 377
rect 811 318 877 343
rect 925 318 961 448
rect 1015 430 1051 448
rect 1015 414 1099 430
rect 1015 380 1032 414
rect 1066 380 1099 414
rect 1015 364 1099 380
rect 557 287 767 303
rect 368 252 505 268
rect 282 222 312 244
rect 368 222 398 252
rect 475 239 505 252
rect 81 196 161 212
rect 84 158 114 196
rect 475 209 604 239
rect 574 158 604 209
rect 710 158 740 287
rect 847 246 877 318
rect 931 293 1027 318
rect 931 288 977 293
rect 961 259 977 288
rect 1011 259 1027 293
rect 847 230 919 246
rect 961 243 1027 259
rect 847 210 869 230
rect 788 196 869 210
rect 903 196 919 230
rect 997 202 1027 243
rect 1069 202 1099 364
rect 1990 571 2020 597
rect 2094 592 2124 618
rect 1427 493 1457 508
rect 1511 493 1541 508
rect 1601 493 1631 508
rect 1796 493 1826 508
rect 1424 470 1460 493
rect 1386 454 1460 470
rect 1386 420 1402 454
rect 1436 420 1460 454
rect 1386 404 1460 420
rect 1268 377 1298 392
rect 1265 362 1301 377
rect 1167 326 1197 341
rect 1265 332 1422 362
rect 1164 309 1200 326
rect 1147 293 1215 309
rect 1147 259 1163 293
rect 1197 259 1215 293
rect 1147 243 1215 259
rect 1185 202 1215 243
rect 1263 274 1329 290
rect 1263 240 1279 274
rect 1313 240 1329 274
rect 1263 224 1329 240
rect 1290 202 1320 224
rect 788 180 919 196
rect 788 158 818 180
rect 997 92 1027 118
rect 1069 92 1099 118
rect 1392 158 1422 332
rect 1508 311 1544 493
rect 1598 428 1634 493
rect 1793 476 1829 493
rect 1755 460 1829 476
rect 1604 412 1703 428
rect 1604 378 1653 412
rect 1687 378 1703 412
rect 1604 344 1703 378
rect 1470 295 1556 311
rect 1470 261 1506 295
rect 1540 261 1556 295
rect 1470 245 1556 261
rect 1604 310 1653 344
rect 1687 310 1703 344
rect 1604 276 1703 310
rect 1470 158 1500 245
rect 1604 242 1653 276
rect 1687 242 1703 276
rect 1755 426 1771 460
rect 1805 446 1829 460
rect 1805 426 1823 446
rect 1755 392 1823 426
rect 1755 358 1771 392
rect 1805 388 1823 392
rect 1990 388 2020 403
rect 1805 358 2023 388
rect 1755 324 1823 358
rect 1755 290 1771 324
rect 1805 290 1823 324
rect 1755 274 1823 290
rect 1604 226 1703 242
rect 1604 203 1634 226
rect 1548 173 1634 203
rect 1548 158 1578 173
rect 1761 158 1791 274
rect 1959 184 1989 358
rect 2094 353 2124 368
rect 2091 310 2127 353
rect 2037 294 2127 310
rect 2037 260 2053 294
rect 2087 260 2127 294
rect 2037 244 2127 260
rect 2075 222 2105 244
rect 84 48 114 74
rect 282 48 312 74
rect 368 48 398 74
rect 574 48 604 74
rect 710 48 740 74
rect 788 48 818 74
rect 1185 48 1215 74
rect 1290 48 1320 74
rect 1392 48 1422 74
rect 1470 48 1500 74
rect 1548 48 1578 74
rect 1761 48 1791 74
rect 1959 48 1989 74
rect 2075 48 2105 74
<< polycont >>
rect 111 348 145 382
rect 111 280 145 314
rect 111 212 145 246
rect 276 260 310 294
rect 413 268 447 302
rect 573 371 607 405
rect 573 303 607 337
rect 717 303 751 337
rect 827 343 861 377
rect 1032 380 1066 414
rect 977 259 1011 293
rect 869 196 903 230
rect 1402 420 1436 454
rect 1163 259 1197 293
rect 1279 240 1313 274
rect 1653 378 1687 412
rect 1506 261 1540 295
rect 1653 310 1687 344
rect 1653 242 1687 276
rect 1771 426 1805 460
rect 1771 358 1805 392
rect 1771 290 1805 324
rect 2053 260 2087 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 21 567 71 596
rect 21 533 37 567
rect 21 480 71 533
rect 111 572 177 649
rect 111 538 127 572
rect 161 538 177 572
rect 111 514 177 538
rect 308 555 374 649
rect 308 521 324 555
rect 358 521 374 555
rect 308 514 374 521
rect 414 581 751 615
rect 414 546 464 581
rect 448 512 464 546
rect 414 480 464 512
rect 498 520 582 547
rect 498 486 532 520
rect 566 486 582 520
rect 21 446 352 480
rect 498 459 582 486
rect 616 520 683 547
rect 616 486 632 520
rect 666 486 683 520
rect 616 459 683 486
rect 498 446 532 459
rect 21 162 55 446
rect 318 412 532 446
rect 95 382 161 398
rect 95 348 111 382
rect 145 348 161 382
rect 95 314 161 348
rect 95 280 111 314
rect 145 280 161 314
rect 95 246 161 280
rect 95 212 111 246
rect 145 212 161 246
rect 95 196 161 212
rect 195 396 284 412
rect 195 362 234 396
rect 268 378 284 396
rect 268 362 463 378
rect 195 344 463 362
rect 195 202 229 344
rect 263 294 359 310
rect 263 260 276 294
rect 310 260 359 294
rect 263 236 359 260
rect 397 302 463 344
rect 397 268 413 302
rect 447 268 463 302
rect 397 252 463 268
rect 393 202 459 218
rect 195 196 287 202
rect 195 162 237 196
rect 271 162 287 196
rect 21 133 73 162
rect 21 99 39 133
rect 21 70 73 99
rect 109 133 159 162
rect 109 99 125 133
rect 109 17 159 99
rect 195 120 287 162
rect 195 86 237 120
rect 271 86 287 120
rect 195 70 287 86
rect 323 186 357 202
rect 323 116 357 152
rect 323 17 357 82
rect 393 168 409 202
rect 443 168 459 202
rect 393 120 459 168
rect 393 86 409 120
rect 443 86 459 120
rect 497 185 532 412
rect 566 405 615 421
rect 566 371 573 405
rect 607 371 615 405
rect 566 337 615 371
rect 566 303 573 337
rect 607 303 615 337
rect 566 287 615 303
rect 497 169 547 185
rect 497 135 513 169
rect 497 119 547 135
rect 393 85 459 86
rect 581 85 615 287
rect 393 51 615 85
rect 649 204 683 459
rect 717 451 751 581
rect 790 535 846 649
rect 790 501 809 535
rect 843 501 846 535
rect 790 485 846 501
rect 880 581 1073 615
rect 880 451 914 581
rect 717 417 914 451
rect 948 522 1005 547
rect 948 488 971 522
rect 948 464 1005 488
rect 1039 498 1073 581
rect 1107 582 1157 649
rect 1141 548 1157 582
rect 1107 532 1157 548
rect 1295 584 1520 596
rect 1295 550 1311 584
rect 1345 550 1380 584
rect 1414 550 1520 584
rect 1295 525 1520 550
rect 1554 580 1588 649
rect 1554 530 1588 546
rect 1628 570 1694 586
rect 1628 536 1644 570
rect 1678 536 1694 570
rect 1295 516 1362 525
rect 1039 464 1195 498
rect 717 337 751 417
rect 948 383 982 464
rect 811 377 982 383
rect 811 343 827 377
rect 861 349 982 377
rect 1016 424 1127 430
rect 1016 414 1087 424
rect 1016 380 1032 414
rect 1066 390 1087 414
rect 1121 390 1127 424
rect 1066 380 1127 390
rect 1016 364 1127 380
rect 1161 377 1195 464
rect 1295 482 1311 516
rect 1345 482 1362 516
rect 1295 448 1362 482
rect 1486 496 1520 525
rect 1628 496 1694 536
rect 1733 580 1783 649
rect 1733 546 1749 580
rect 1733 530 1783 546
rect 1823 580 1889 596
rect 1823 546 1839 580
rect 1873 546 1889 580
rect 2031 580 2097 649
rect 1823 530 1889 546
rect 1295 414 1312 448
rect 1346 414 1362 448
rect 1295 410 1362 414
rect 861 343 877 349
rect 1161 343 1281 377
rect 811 337 877 343
rect 961 303 1213 309
rect 717 287 751 303
rect 785 293 1213 303
rect 785 269 977 293
rect 785 204 819 269
rect 961 259 977 269
rect 1011 259 1163 293
rect 1197 259 1213 293
rect 961 243 1213 259
rect 1247 290 1281 343
rect 1315 360 1362 410
rect 1396 454 1452 471
rect 1486 462 1821 496
rect 1396 420 1402 454
rect 1436 428 1452 454
rect 1755 460 1821 462
rect 1436 420 1465 428
rect 1396 394 1465 420
rect 1315 326 1397 360
rect 1247 274 1329 290
rect 1247 240 1279 274
rect 1313 240 1329 274
rect 649 170 819 204
rect 853 230 925 235
rect 853 196 869 230
rect 903 206 925 230
rect 1247 224 1329 240
rect 903 196 1002 206
rect 853 177 1002 196
rect 853 172 952 177
rect 649 133 715 170
rect 925 143 952 172
rect 986 143 1002 177
rect 649 99 665 133
rect 699 99 715 133
rect 649 83 715 99
rect 813 120 891 136
rect 813 86 835 120
rect 869 86 891 120
rect 925 114 1002 143
rect 1124 190 1190 206
rect 1124 156 1140 190
rect 1174 156 1190 190
rect 1124 120 1190 156
rect 813 17 891 86
rect 1124 86 1140 120
rect 1174 86 1190 120
rect 1124 17 1190 86
rect 1247 85 1281 224
rect 1363 185 1397 326
rect 1315 169 1397 185
rect 1315 135 1331 169
rect 1365 135 1397 169
rect 1315 119 1397 135
rect 1431 85 1465 394
rect 1637 424 1703 428
rect 1637 412 1663 424
rect 1637 378 1653 412
rect 1697 390 1703 424
rect 1687 378 1703 390
rect 1637 344 1703 378
rect 1499 295 1546 311
rect 1499 261 1506 295
rect 1540 261 1546 295
rect 1499 192 1546 261
rect 1637 310 1653 344
rect 1687 310 1703 344
rect 1637 276 1703 310
rect 1637 242 1653 276
rect 1687 242 1703 276
rect 1755 426 1771 460
rect 1805 426 1821 460
rect 1755 392 1821 426
rect 1755 358 1771 392
rect 1805 358 1821 392
rect 1755 324 1821 358
rect 1755 290 1771 324
rect 1805 290 1821 324
rect 1755 274 1821 290
rect 1637 226 1703 242
rect 1855 240 1889 530
rect 1818 206 1889 240
rect 1927 559 1993 575
rect 1927 525 1943 559
rect 1977 525 1993 559
rect 1927 449 1993 525
rect 1927 415 1943 449
rect 1977 415 1993 449
rect 1927 310 1993 415
rect 2031 546 2047 580
rect 2081 546 2097 580
rect 2031 497 2097 546
rect 2031 463 2047 497
rect 2081 463 2097 497
rect 2031 414 2097 463
rect 2031 380 2047 414
rect 2081 380 2097 414
rect 2031 364 2097 380
rect 2137 580 2187 596
rect 2171 546 2187 580
rect 2137 497 2187 546
rect 2171 463 2187 497
rect 2137 414 2187 463
rect 2171 380 2187 414
rect 1927 294 2103 310
rect 1927 260 2053 294
rect 2087 260 2103 294
rect 1927 244 2103 260
rect 1818 192 1852 206
rect 1499 158 1852 192
rect 1927 172 1964 244
rect 2137 210 2187 380
rect 1786 133 1852 158
rect 1247 51 1465 85
rect 1574 86 1590 120
rect 1624 86 1702 120
rect 1736 86 1752 120
rect 1574 17 1752 86
rect 1786 99 1802 133
rect 1836 99 1852 133
rect 1786 70 1852 99
rect 1898 138 1964 172
rect 1898 104 1914 138
rect 1948 104 1964 138
rect 1898 70 1964 104
rect 2000 203 2066 206
rect 2000 169 2016 203
rect 2050 169 2066 203
rect 2000 116 2066 169
rect 2000 82 2016 116
rect 2050 82 2066 116
rect 2000 17 2066 82
rect 2100 194 2187 210
rect 2100 160 2116 194
rect 2150 160 2187 194
rect 2100 120 2187 160
rect 2100 86 2116 120
rect 2150 86 2187 120
rect 2100 70 2187 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 1087 390 1121 424
rect 1663 412 1697 424
rect 1663 390 1687 412
rect 1687 390 1697 412
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
<< metal1 >>
rect 0 683 2208 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 0 617 2208 649
rect 1075 424 1133 430
rect 1075 390 1087 424
rect 1121 421 1133 424
rect 1651 424 1709 430
rect 1651 421 1663 424
rect 1121 393 1663 421
rect 1121 390 1133 393
rect 1075 384 1133 390
rect 1651 390 1663 393
rect 1697 390 1709 424
rect 1651 384 1709 390
rect 0 17 2208 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
rect 0 -49 2208 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dfstp_1
flabel comment s 866 259 866 259 0 FreeSans 200 0 0 0 no_jumper_check
flabel comment s 693 302 693 302 0 FreeSans 200 0 0 0 no_jumper_check
flabel pwell s 0 0 2208 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 0 617 2208 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 1663 390 1697 424 0 FreeSans 340 0 0 0 SET_B
port 3 nsew
flabel metal1 s 0 617 2208 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 2208 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 2143 94 2177 128 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 2143 168 2177 202 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 2143 242 2177 276 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 2143 316 2177 350 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 2143 390 2177 424 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 2143 464 2177 498 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 2143 538 2177 572 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 127 242 161 276 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 319 242 353 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 2208 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2749860
string GDS_START 2732446
<< end >>
