magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1656 561
rect 103 427 169 527
rect 17 197 66 325
rect 103 17 169 93
rect 391 367 454 527
rect 292 191 358 265
rect 764 427 918 527
rect 1020 371 1070 527
rect 1130 332 1183 493
rect 1217 366 1271 527
rect 1130 299 1195 332
rect 1158 265 1195 299
rect 1407 367 1466 527
rect 1500 289 1551 493
rect 1585 299 1639 527
rect 1509 265 1551 289
rect 878 199 1028 265
rect 1158 177 1271 265
rect 1509 211 1639 265
rect 1158 172 1195 177
rect 1148 165 1195 172
rect 375 17 441 89
rect 748 17 814 165
rect 1130 137 1195 165
rect 1130 131 1190 137
rect 1020 17 1096 97
rect 1130 83 1182 131
rect 1217 17 1271 109
rect 1509 165 1551 211
rect 1405 17 1466 109
rect 1500 51 1551 165
rect 1585 17 1639 177
rect 0 -17 1656 17
<< obsli1 >>
rect 17 393 69 493
rect 17 359 156 393
rect 121 323 156 359
rect 121 289 122 323
rect 121 280 156 289
rect 203 391 248 493
rect 203 357 214 391
rect 203 337 248 357
rect 121 214 168 280
rect 121 161 156 214
rect 17 127 156 161
rect 17 69 69 127
rect 203 69 237 337
rect 291 333 357 483
rect 580 451 730 485
rect 494 391 551 401
rect 528 357 551 391
rect 291 299 428 333
rect 394 219 428 299
rect 494 271 551 357
rect 585 323 653 399
rect 585 289 586 323
rect 620 289 653 323
rect 585 283 653 289
rect 394 157 468 219
rect 585 207 619 283
rect 696 265 730 451
rect 952 373 986 487
rect 768 333 986 373
rect 768 299 1096 333
rect 1062 265 1096 299
rect 1305 265 1371 493
rect 696 233 840 265
rect 307 153 468 157
rect 307 123 428 153
rect 543 141 619 207
rect 666 199 840 233
rect 1062 199 1124 265
rect 307 69 341 123
rect 666 107 700 199
rect 1062 165 1096 199
rect 1305 199 1475 265
rect 568 73 700 107
rect 868 131 1096 165
rect 868 83 912 131
rect 1305 51 1371 199
<< obsli1c >>
rect 122 289 156 323
rect 214 357 248 391
rect 494 357 528 391
rect 586 289 620 323
<< metal1 >>
rect 0 496 1656 592
rect 0 -48 1656 48
<< obsm1 >>
rect 202 391 260 397
rect 202 357 214 391
rect 248 388 260 391
rect 482 391 540 397
rect 482 388 494 391
rect 248 360 494 388
rect 248 357 260 360
rect 202 351 260 357
rect 482 357 494 360
rect 528 357 540 391
rect 482 351 540 357
rect 110 323 168 329
rect 110 289 122 323
rect 156 320 168 323
rect 574 323 632 329
rect 574 320 586 323
rect 156 292 586 320
rect 156 289 168 292
rect 110 283 168 289
rect 574 289 586 292
rect 620 289 632 323
rect 574 283 632 289
<< labels >>
rlabel locali s 292 191 358 265 6 D
port 1 nsew signal input
rlabel locali s 1158 265 1195 299 6 Q
port 2 nsew signal output
rlabel locali s 1158 177 1271 265 6 Q
port 2 nsew signal output
rlabel locali s 1158 172 1195 177 6 Q
port 2 nsew signal output
rlabel locali s 1148 165 1195 172 6 Q
port 2 nsew signal output
rlabel locali s 1130 332 1183 493 6 Q
port 2 nsew signal output
rlabel locali s 1130 299 1195 332 6 Q
port 2 nsew signal output
rlabel locali s 1130 137 1195 165 6 Q
port 2 nsew signal output
rlabel locali s 1130 131 1190 137 6 Q
port 2 nsew signal output
rlabel locali s 1130 83 1182 131 6 Q
port 2 nsew signal output
rlabel locali s 1509 265 1551 289 6 Q_N
port 3 nsew signal output
rlabel locali s 1509 211 1639 265 6 Q_N
port 3 nsew signal output
rlabel locali s 1509 165 1551 211 6 Q_N
port 3 nsew signal output
rlabel locali s 1500 289 1551 493 6 Q_N
port 3 nsew signal output
rlabel locali s 1500 51 1551 165 6 Q_N
port 3 nsew signal output
rlabel locali s 878 199 1028 265 6 RESET_B
port 4 nsew signal input
rlabel locali s 17 197 66 325 6 GATE_N
port 5 nsew clock input
rlabel locali s 1585 17 1639 177 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1405 17 1466 109 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1217 17 1271 109 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1020 17 1096 97 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 748 17 814 165 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 375 17 441 89 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 103 17 169 93 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 1656 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1656 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1585 299 1639 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1407 367 1466 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1217 366 1271 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1020 371 1070 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 764 427 918 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 391 367 454 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 103 427 169 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 1656 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 1656 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1656 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2697216
string GDS_START 2683874
<< end >>
