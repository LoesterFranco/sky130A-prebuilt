magic
tech sky130A
magscale 1 2
timestamp 1599588209
<< nwell >>
rect -38 332 422 704
<< pwell >>
rect 0 0 384 49
<< scpmos >>
rect 84 368 114 592
rect 174 368 204 592
rect 264 368 294 592
<< nmoslvt >>
rect 84 74 114 158
rect 170 74 200 158
rect 270 74 300 158
<< ndiff >>
rect 27 131 84 158
rect 27 97 39 131
rect 73 97 84 131
rect 27 74 84 97
rect 114 131 170 158
rect 114 97 125 131
rect 159 97 170 131
rect 114 74 170 97
rect 200 133 270 158
rect 200 99 211 133
rect 245 99 270 133
rect 200 74 270 99
rect 300 133 357 158
rect 300 99 311 133
rect 345 99 357 133
rect 300 74 357 99
<< pdiff >>
rect 27 573 84 592
rect 27 539 37 573
rect 71 539 84 573
rect 27 368 84 539
rect 114 414 174 592
rect 114 380 127 414
rect 161 380 174 414
rect 114 368 174 380
rect 204 573 264 592
rect 204 539 217 573
rect 251 539 264 573
rect 204 368 264 539
rect 294 580 357 592
rect 294 546 309 580
rect 343 546 357 580
rect 294 498 357 546
rect 294 464 309 498
rect 343 464 357 498
rect 294 368 357 464
<< ndiffc >>
rect 39 97 73 131
rect 125 97 159 131
rect 211 99 245 133
rect 311 99 345 133
<< pdiffc >>
rect 37 539 71 573
rect 127 380 161 414
rect 217 539 251 573
rect 309 546 343 580
rect 309 464 343 498
<< poly >>
rect 84 592 114 618
rect 174 592 204 618
rect 264 592 294 618
rect 84 353 114 368
rect 174 353 204 368
rect 264 353 294 368
rect 81 326 117 353
rect 171 326 207 353
rect 261 336 297 353
rect 43 310 207 326
rect 43 276 59 310
rect 93 276 207 310
rect 43 242 207 276
rect 43 208 59 242
rect 93 208 207 242
rect 43 192 207 208
rect 249 320 315 336
rect 249 286 265 320
rect 299 286 315 320
rect 249 252 315 286
rect 249 218 265 252
rect 299 218 315 252
rect 249 202 315 218
rect 84 158 114 192
rect 170 158 200 192
rect 270 158 300 202
rect 84 48 114 74
rect 170 48 200 74
rect 270 48 300 74
<< polycont >>
rect 59 276 93 310
rect 59 208 93 242
rect 265 286 299 320
rect 265 218 299 252
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 384 683
rect 21 573 87 649
rect 21 539 37 573
rect 71 539 87 573
rect 21 532 87 539
rect 201 573 267 649
rect 201 539 217 573
rect 251 539 267 573
rect 201 532 267 539
rect 307 580 367 596
rect 307 546 309 580
rect 343 546 367 580
rect 307 498 367 546
rect 43 464 309 498
rect 343 464 367 498
rect 43 326 77 464
rect 111 414 177 430
rect 111 380 127 414
rect 161 380 177 414
rect 111 364 177 380
rect 43 310 109 326
rect 43 276 59 310
rect 93 276 109 310
rect 43 242 109 276
rect 43 208 59 242
rect 93 208 109 242
rect 43 192 109 208
rect 143 158 177 364
rect 217 320 299 430
rect 217 286 265 320
rect 217 252 299 286
rect 217 218 265 252
rect 217 202 299 218
rect 333 162 367 464
rect 23 131 73 158
rect 23 97 39 131
rect 23 17 73 97
rect 109 131 177 158
rect 109 97 125 131
rect 159 97 177 131
rect 109 70 177 97
rect 211 133 261 162
rect 245 99 261 133
rect 211 17 261 99
rect 295 133 367 162
rect 295 99 311 133
rect 345 99 367 133
rect 295 70 367 99
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 384 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
<< metal1 >>
rect 0 683 384 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 384 683
rect 0 617 384 649
rect 0 17 384 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 384 17
rect 0 -49 384 -17
<< labels >>
rlabel comment s 0 0 0 0 4 clkbuf_2
flabel pwell s 0 0 384 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew
flabel nwell s 0 617 384 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew
flabel metal1 s 0 617 384 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew
flabel metal1 s 0 0 384 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew
flabel corelocali s 127 94 161 128 0 FreeSans 340 0 0 0 X
port 6 nsew
flabel corelocali s 223 242 257 276 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 223 390 257 424 0 FreeSans 340 0 0 0 A
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 384 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3428484
string GDS_START 3424318
<< end >>
