magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 88 153 168 327
rect 206 309 472 343
rect 206 164 272 309
rect 574 199 624 265
rect 206 130 456 164
rect 666 151 728 265
rect 762 147 838 265
rect 206 51 268 130
rect 422 51 456 130
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 17 417 69 493
rect 103 451 179 527
rect 302 451 378 527
rect 490 451 566 527
rect 702 451 778 527
rect 914 451 990 527
rect 17 383 977 417
rect 17 117 52 383
rect 506 309 906 343
rect 506 265 540 309
rect 306 199 540 265
rect 872 162 906 309
rect 943 199 977 383
rect 17 51 69 117
rect 113 17 163 109
rect 302 17 378 94
rect 872 128 980 162
rect 507 17 573 89
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
rlabel locali s 88 153 168 327 6 A_N
port 1 nsew signal input
rlabel locali s 762 147 838 265 6 B
port 2 nsew signal input
rlabel locali s 666 151 728 265 6 C
port 3 nsew signal input
rlabel locali s 574 199 624 265 6 D
port 4 nsew signal input
rlabel locali s 422 51 456 130 6 X
port 5 nsew signal output
rlabel locali s 206 309 472 343 6 X
port 5 nsew signal output
rlabel locali s 206 164 272 309 6 X
port 5 nsew signal output
rlabel locali s 206 130 456 164 6 X
port 5 nsew signal output
rlabel locali s 206 51 268 130 6 X
port 5 nsew signal output
rlabel metal1 s 0 -48 1012 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 1012 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1012 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1597714
string GDS_START 1589860
<< end >>
