magic
tech sky130A
magscale 1 2
timestamp 1604502693
<< nwell >>
rect -38 261 1510 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 415 47 445 177
rect 499 47 529 177
rect 687 47 717 177
rect 771 47 801 177
rect 855 47 885 177
rect 939 47 969 177
rect 1023 47 1053 177
rect 1107 47 1137 177
rect 1191 47 1221 177
rect 1275 47 1305 177
<< pmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 415 297 445 497
rect 499 297 529 497
rect 687 297 717 497
rect 771 297 801 497
rect 855 297 885 497
rect 939 297 969 497
rect 1023 297 1053 497
rect 1107 297 1137 497
rect 1191 297 1221 497
rect 1275 297 1305 497
<< ndiff >>
rect 27 163 79 177
rect 27 129 35 163
rect 69 129 79 163
rect 27 95 79 129
rect 27 61 35 95
rect 69 61 79 95
rect 27 47 79 61
rect 109 163 163 177
rect 109 129 119 163
rect 153 129 163 163
rect 109 95 163 129
rect 109 61 119 95
rect 153 61 163 95
rect 109 47 163 61
rect 193 163 247 177
rect 193 129 203 163
rect 237 129 247 163
rect 193 47 247 129
rect 277 95 331 177
rect 277 61 287 95
rect 321 61 331 95
rect 277 47 331 61
rect 361 95 415 177
rect 361 61 371 95
rect 405 61 415 95
rect 361 47 415 61
rect 445 163 499 177
rect 445 129 455 163
rect 489 129 499 163
rect 445 95 499 129
rect 445 61 455 95
rect 489 61 499 95
rect 445 47 499 61
rect 529 95 687 177
rect 529 61 539 95
rect 573 61 643 95
rect 677 61 687 95
rect 529 47 687 61
rect 717 163 771 177
rect 717 129 727 163
rect 761 129 771 163
rect 717 95 771 129
rect 717 61 727 95
rect 761 61 771 95
rect 717 47 771 61
rect 801 95 855 177
rect 801 61 811 95
rect 845 61 855 95
rect 801 47 855 61
rect 885 163 939 177
rect 885 129 895 163
rect 929 129 939 163
rect 885 95 939 129
rect 885 61 895 95
rect 929 61 939 95
rect 885 47 939 61
rect 969 163 1023 177
rect 969 129 979 163
rect 1013 129 1023 163
rect 969 95 1023 129
rect 969 61 979 95
rect 1013 61 1023 95
rect 969 47 1023 61
rect 1053 163 1107 177
rect 1053 129 1063 163
rect 1097 129 1107 163
rect 1053 95 1107 129
rect 1053 61 1063 95
rect 1097 61 1107 95
rect 1053 47 1107 61
rect 1137 95 1191 177
rect 1137 61 1147 95
rect 1181 61 1191 95
rect 1137 47 1191 61
rect 1221 163 1275 177
rect 1221 129 1231 163
rect 1265 129 1275 163
rect 1221 95 1275 129
rect 1221 61 1231 95
rect 1265 61 1275 95
rect 1221 47 1275 61
rect 1305 95 1357 177
rect 1305 61 1315 95
rect 1349 61 1357 95
rect 1305 47 1357 61
<< pdiff >>
rect 27 477 79 497
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 297 79 375
rect 109 477 163 497
rect 109 443 119 477
rect 153 443 163 477
rect 109 297 163 443
rect 193 477 247 497
rect 193 443 203 477
rect 237 443 247 477
rect 193 409 247 443
rect 193 375 203 409
rect 237 375 247 409
rect 193 297 247 375
rect 277 477 331 497
rect 277 443 287 477
rect 321 443 331 477
rect 277 297 331 443
rect 361 477 415 497
rect 361 443 371 477
rect 405 443 415 477
rect 361 409 415 443
rect 361 375 371 409
rect 405 375 415 409
rect 361 341 415 375
rect 361 307 371 341
rect 405 307 415 341
rect 361 297 415 307
rect 445 409 499 497
rect 445 375 455 409
rect 489 375 499 409
rect 445 341 499 375
rect 445 307 455 341
rect 489 307 499 341
rect 445 297 499 307
rect 529 477 581 497
rect 529 443 539 477
rect 573 443 581 477
rect 529 297 581 443
rect 635 485 687 497
rect 635 451 643 485
rect 677 451 687 485
rect 635 297 687 451
rect 717 477 771 497
rect 717 443 727 477
rect 761 443 771 477
rect 717 297 771 443
rect 801 409 855 497
rect 801 375 811 409
rect 845 375 855 409
rect 801 297 855 375
rect 885 477 939 497
rect 885 443 895 477
rect 929 443 939 477
rect 885 409 939 443
rect 885 375 895 409
rect 929 375 939 409
rect 885 297 939 375
rect 969 477 1023 497
rect 969 443 979 477
rect 1013 443 1023 477
rect 969 409 1023 443
rect 969 375 979 409
rect 1013 375 1023 409
rect 969 297 1023 375
rect 1053 477 1107 497
rect 1053 443 1063 477
rect 1097 443 1107 477
rect 1053 409 1107 443
rect 1053 375 1063 409
rect 1097 375 1107 409
rect 1053 297 1107 375
rect 1137 483 1191 497
rect 1137 449 1147 483
rect 1181 449 1191 483
rect 1137 297 1191 449
rect 1221 477 1275 497
rect 1221 443 1231 477
rect 1265 443 1275 477
rect 1221 409 1275 443
rect 1221 375 1231 409
rect 1265 375 1275 409
rect 1221 341 1275 375
rect 1221 307 1231 341
rect 1265 307 1275 341
rect 1221 297 1275 307
rect 1305 483 1357 497
rect 1305 449 1315 483
rect 1349 449 1357 483
rect 1305 415 1357 449
rect 1305 381 1315 415
rect 1349 381 1357 415
rect 1305 297 1357 381
<< ndiffc >>
rect 35 129 69 163
rect 35 61 69 95
rect 119 129 153 163
rect 119 61 153 95
rect 203 129 237 163
rect 287 61 321 95
rect 371 61 405 95
rect 455 129 489 163
rect 455 61 489 95
rect 539 61 573 95
rect 643 61 677 95
rect 727 129 761 163
rect 727 61 761 95
rect 811 61 845 95
rect 895 129 929 163
rect 895 61 929 95
rect 979 129 1013 163
rect 979 61 1013 95
rect 1063 129 1097 163
rect 1063 61 1097 95
rect 1147 61 1181 95
rect 1231 129 1265 163
rect 1231 61 1265 95
rect 1315 61 1349 95
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 443 153 477
rect 203 443 237 477
rect 203 375 237 409
rect 287 443 321 477
rect 371 443 405 477
rect 371 375 405 409
rect 371 307 405 341
rect 455 375 489 409
rect 455 307 489 341
rect 539 443 573 477
rect 643 451 677 485
rect 727 443 761 477
rect 811 375 845 409
rect 895 443 929 477
rect 895 375 929 409
rect 979 443 1013 477
rect 979 375 1013 409
rect 1063 443 1097 477
rect 1063 375 1097 409
rect 1147 449 1181 483
rect 1231 443 1265 477
rect 1231 375 1265 409
rect 1231 307 1265 341
rect 1315 449 1349 483
rect 1315 381 1349 415
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 415 497 445 523
rect 499 497 529 523
rect 687 497 717 523
rect 771 497 801 523
rect 855 497 885 523
rect 939 497 969 523
rect 1023 497 1053 523
rect 1107 497 1137 523
rect 1191 497 1221 523
rect 1275 497 1305 523
rect 79 265 109 297
rect 55 249 109 265
rect 55 215 65 249
rect 99 215 109 249
rect 55 199 109 215
rect 79 177 109 199
rect 163 265 193 297
rect 247 265 277 297
rect 331 265 361 297
rect 415 265 445 297
rect 499 265 529 297
rect 687 265 717 297
rect 771 265 801 297
rect 855 265 885 297
rect 939 265 969 297
rect 1023 265 1053 297
rect 1107 265 1137 297
rect 1191 265 1221 297
rect 1275 265 1305 297
rect 163 249 277 265
rect 163 215 203 249
rect 237 215 277 249
rect 163 199 277 215
rect 319 249 373 265
rect 319 215 329 249
rect 363 215 373 249
rect 319 199 373 215
rect 415 249 589 265
rect 415 215 539 249
rect 573 215 589 249
rect 415 199 589 215
rect 663 249 729 265
rect 663 215 679 249
rect 713 215 729 249
rect 663 199 729 215
rect 771 249 885 265
rect 771 215 812 249
rect 846 215 885 249
rect 771 199 885 215
rect 927 249 981 265
rect 927 215 937 249
rect 971 215 981 249
rect 927 199 981 215
rect 1023 249 1305 265
rect 1023 215 1089 249
rect 1123 215 1157 249
rect 1191 215 1225 249
rect 1259 215 1305 249
rect 1023 199 1305 215
rect 163 177 193 199
rect 247 177 277 199
rect 331 177 361 199
rect 415 177 445 199
rect 499 177 529 199
rect 687 177 717 199
rect 771 177 801 199
rect 855 177 885 199
rect 939 177 969 199
rect 1023 177 1053 199
rect 1107 177 1137 199
rect 1191 177 1221 199
rect 1275 177 1305 199
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 415 21 445 47
rect 499 21 529 47
rect 687 21 717 47
rect 771 21 801 47
rect 855 21 885 47
rect 939 21 969 47
rect 1023 21 1053 47
rect 1107 21 1137 47
rect 1191 21 1221 47
rect 1275 21 1305 47
<< polycont >>
rect 65 215 99 249
rect 203 215 237 249
rect 329 215 363 249
rect 539 215 573 249
rect 679 215 713 249
rect 812 215 846 249
rect 937 215 971 249
rect 1089 215 1123 249
rect 1157 215 1191 249
rect 1225 215 1259 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 27 477 77 493
rect 27 443 35 477
rect 69 443 77 477
rect 27 409 77 443
rect 111 477 161 527
rect 111 443 119 477
rect 153 443 161 477
rect 111 425 161 443
rect 195 477 245 493
rect 195 443 203 477
rect 237 443 245 477
rect 27 375 35 409
rect 69 391 77 409
rect 195 409 245 443
rect 279 477 329 527
rect 279 443 287 477
rect 321 443 329 477
rect 279 425 329 443
rect 363 477 581 493
rect 363 443 371 477
rect 405 459 539 477
rect 405 443 413 459
rect 195 391 203 409
rect 69 375 203 391
rect 237 391 245 409
rect 363 409 413 443
rect 531 443 539 459
rect 573 443 581 477
rect 531 427 581 443
rect 635 485 685 527
rect 635 451 643 485
rect 677 451 685 485
rect 635 427 685 451
rect 719 477 937 493
rect 719 443 727 477
rect 761 459 895 477
rect 761 443 769 459
rect 719 427 769 443
rect 887 443 895 459
rect 929 443 937 477
rect 363 391 371 409
rect 237 375 371 391
rect 405 375 413 409
rect 27 357 413 375
rect 371 341 413 357
rect 17 289 337 323
rect 405 307 413 341
rect 371 291 413 307
rect 447 409 497 425
rect 447 375 455 409
rect 489 393 497 409
rect 803 409 853 425
rect 803 393 811 409
rect 489 375 524 393
rect 447 341 524 375
rect 447 307 455 341
rect 489 323 524 341
rect 627 375 811 393
rect 845 375 853 409
rect 627 357 853 375
rect 887 409 937 443
rect 887 375 895 409
rect 929 375 937 409
rect 887 357 937 375
rect 971 477 1021 527
rect 971 443 979 477
rect 1013 443 1021 477
rect 971 409 1021 443
rect 971 375 979 409
rect 1013 375 1021 409
rect 971 359 1021 375
rect 1055 477 1105 493
rect 1055 443 1063 477
rect 1097 443 1105 477
rect 1055 409 1105 443
rect 1139 483 1189 527
rect 1139 449 1147 483
rect 1181 449 1189 483
rect 1139 433 1189 449
rect 1223 477 1273 493
rect 1223 443 1231 477
rect 1265 443 1273 477
rect 1055 375 1063 409
rect 1097 391 1105 409
rect 1223 409 1273 443
rect 1223 391 1231 409
rect 1097 375 1231 391
rect 1265 375 1273 409
rect 1055 357 1273 375
rect 1307 483 1357 527
rect 1307 449 1315 483
rect 1349 449 1357 483
rect 1307 415 1357 449
rect 1307 381 1315 415
rect 1349 381 1357 415
rect 1307 365 1357 381
rect 627 333 661 357
rect 489 307 490 323
rect 17 249 115 289
rect 17 215 65 249
rect 99 215 115 249
rect 161 249 269 255
rect 161 215 203 249
rect 237 215 269 249
rect 303 249 337 289
rect 447 289 490 307
rect 447 283 524 289
rect 591 299 661 333
rect 1223 341 1273 357
rect 303 215 329 249
rect 363 215 379 249
rect 447 181 489 283
rect 591 249 629 299
rect 695 289 993 323
rect 695 265 729 289
rect 523 215 539 249
rect 573 215 629 249
rect 663 249 729 265
rect 663 215 679 249
rect 713 215 729 249
rect 763 249 887 255
rect 763 215 812 249
rect 846 215 887 249
rect 921 249 993 289
rect 921 215 937 249
rect 971 215 993 249
rect 1027 289 1046 323
rect 1080 289 1092 323
rect 1027 249 1092 289
rect 1223 307 1231 341
rect 1265 331 1273 341
rect 1265 307 1384 331
rect 1223 283 1384 307
rect 1027 215 1089 249
rect 1123 215 1157 249
rect 1191 215 1225 249
rect 1259 215 1288 249
rect 591 181 629 215
rect 1322 181 1384 283
rect 35 163 69 179
rect 35 95 69 129
rect 35 17 69 61
rect 103 163 153 181
rect 103 129 119 163
rect 187 163 505 181
rect 187 129 203 163
rect 237 147 455 163
rect 237 129 254 147
rect 439 129 455 147
rect 489 129 505 163
rect 591 163 945 181
rect 591 145 727 163
rect 103 95 153 129
rect 371 95 405 111
rect 103 61 119 95
rect 153 61 287 95
rect 321 61 337 95
rect 103 51 337 61
rect 371 17 405 61
rect 439 95 505 129
rect 711 129 727 145
rect 761 145 895 163
rect 761 129 777 145
rect 439 61 455 95
rect 489 61 505 95
rect 439 51 505 61
rect 539 95 677 111
rect 573 61 643 95
rect 539 17 677 61
rect 711 95 777 129
rect 879 129 895 145
rect 929 129 945 163
rect 711 61 727 95
rect 761 61 777 95
rect 711 51 777 61
rect 811 95 845 111
rect 811 17 845 61
rect 879 95 945 129
rect 879 61 895 95
rect 929 61 945 95
rect 879 51 945 61
rect 979 163 1013 179
rect 979 95 1013 129
rect 979 17 1013 61
rect 1047 163 1384 181
rect 1047 129 1063 163
rect 1097 145 1231 163
rect 1097 129 1113 145
rect 1047 95 1113 129
rect 1215 129 1231 145
rect 1265 145 1384 163
rect 1265 129 1281 145
rect 1047 61 1063 95
rect 1097 61 1113 95
rect 1047 55 1113 61
rect 1147 95 1181 111
rect 1147 17 1181 61
rect 1215 95 1281 129
rect 1215 61 1231 95
rect 1265 61 1281 95
rect 1215 55 1281 61
rect 1315 95 1349 111
rect 1315 17 1349 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 490 289 524 323
rect 1046 289 1080 323
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 478 323 536 329
rect 478 289 490 323
rect 524 320 536 323
rect 1034 323 1092 329
rect 1034 320 1046 323
rect 524 292 1046 320
rect 524 289 536 292
rect 478 283 536 289
rect 1034 289 1046 292
rect 1080 289 1092 323
rect 1034 283 1092 289
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< labels >>
flabel corelocali s 30 221 64 255 0 FreeSans 400 0 0 0 B1
port 3 nsew
flabel corelocali s 214 221 248 255 0 FreeSans 400 0 0 0 B2
port 4 nsew
flabel corelocali s 1322 289 1356 323 0 FreeSans 400 180 0 0 X
port 9 nsew
flabel corelocali s 954 221 988 255 0 FreeSans 400 180 0 0 A1_N
port 1 nsew
flabel corelocali s 770 221 804 255 0 FreeSans 400 180 0 0 A2_N
port 2 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
rlabel comment s 0 0 0 0 4 a2bb2o_4
<< properties >>
string FIXED_BBOX 0 0 1472 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3475012
string GDS_START 3463608
string path 0.000 0.000 36.800 0.000 
<< end >>
