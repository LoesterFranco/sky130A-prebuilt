magic
tech sky130A
magscale 1 2
timestamp 1599588232
<< locali >>
rect 25 290 114 356
rect 377 209 455 356
rect 491 236 557 356
rect 599 270 665 356
rect 767 364 847 596
rect 813 226 847 364
rect 767 70 847 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 24 424 90 596
rect 124 458 190 649
rect 263 424 329 572
rect 667 458 733 649
rect 24 390 196 424
rect 162 382 196 390
rect 263 390 733 424
rect 162 316 228 382
rect 162 256 196 316
rect 23 222 196 256
rect 23 70 89 222
rect 123 17 189 188
rect 263 175 329 390
rect 699 326 733 390
rect 699 260 779 326
rect 699 236 733 260
rect 591 202 733 236
rect 591 188 625 202
rect 223 109 418 175
rect 452 17 518 175
rect 552 70 625 188
rect 659 17 725 168
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel locali s 599 270 665 356 6 A
port 1 nsew signal input
rlabel locali s 491 236 557 356 6 B
port 2 nsew signal input
rlabel locali s 377 209 455 356 6 C
port 3 nsew signal input
rlabel locali s 25 290 114 356 6 D_N
port 4 nsew signal input
rlabel locali s 813 226 847 364 6 X
port 5 nsew signal output
rlabel locali s 767 364 847 596 6 X
port 5 nsew signal output
rlabel locali s 767 70 847 226 6 X
port 5 nsew signal output
rlabel metal1 s 0 -49 864 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 7 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 617 864 715 6 VPWR
port 9 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 858036
string GDS_START 850552
<< end >>
