magic
tech sky130A
magscale 1 2
timestamp 1604502741
<< locali >>
rect 493 378 559 596
rect 493 344 659 378
rect 21 236 167 310
rect 211 236 277 310
rect 313 236 391 310
rect 593 70 659 344
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 67 364 133 649
rect 265 378 331 572
rect 393 412 459 649
rect 593 412 659 649
rect 265 344 459 378
rect 425 310 459 344
rect 425 244 529 310
rect 425 202 459 244
rect 50 168 347 202
rect 50 68 116 168
rect 150 17 247 120
rect 281 68 347 168
rect 381 68 459 202
rect 493 17 559 210
rect 695 17 745 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel locali s 21 236 167 310 6 A1
port 1 nsew signal input
rlabel locali s 211 236 277 310 6 A2
port 2 nsew signal input
rlabel locali s 313 236 391 310 6 B1
port 3 nsew signal input
rlabel locali s 593 70 659 344 6 X
port 4 nsew signal output
rlabel locali s 493 378 559 596 6 X
port 4 nsew signal output
rlabel locali s 493 344 659 378 6 X
port 4 nsew signal output
rlabel metal1 s 0 -49 768 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 617 768 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1034154
string GDS_START 1027326
<< end >>
