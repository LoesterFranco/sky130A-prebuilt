magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 89 53 119 137
rect 287 53 317 137
rect 381 53 411 137
rect 453 53 483 137
rect 593 47 623 177
rect 687 47 717 177
<< pmoshvt >>
rect 81 311 117 395
rect 279 311 315 395
rect 373 311 409 395
rect 478 297 514 381
rect 585 297 621 497
rect 679 297 715 497
<< ndiff >>
rect 524 137 593 177
rect 27 99 89 137
rect 27 65 35 99
rect 69 65 89 99
rect 27 53 89 65
rect 119 111 175 137
rect 119 77 133 111
rect 167 77 175 111
rect 119 53 175 77
rect 229 111 287 137
rect 229 77 237 111
rect 271 77 287 111
rect 229 53 287 77
rect 317 53 381 137
rect 411 53 453 137
rect 483 116 593 137
rect 483 82 538 116
rect 572 82 593 116
rect 483 53 593 82
rect 527 47 593 53
rect 623 123 687 177
rect 623 89 633 123
rect 667 89 687 123
rect 623 47 687 89
rect 717 120 795 177
rect 717 86 753 120
rect 787 86 795 120
rect 717 47 795 86
<< pdiff >>
rect 531 477 585 497
rect 531 443 539 477
rect 573 443 585 477
rect 531 408 585 443
rect 27 365 81 395
rect 27 331 35 365
rect 69 331 81 365
rect 27 311 81 331
rect 117 365 171 395
rect 117 331 129 365
rect 163 331 171 365
rect 117 311 171 331
rect 225 369 279 395
rect 225 335 233 369
rect 267 335 279 369
rect 225 311 279 335
rect 315 387 373 395
rect 315 353 327 387
rect 361 353 373 387
rect 315 311 373 353
rect 409 381 461 395
rect 531 381 539 408
rect 409 362 478 381
rect 409 328 432 362
rect 466 328 478 362
rect 409 311 478 328
rect 426 297 478 311
rect 514 374 539 381
rect 573 374 585 408
rect 514 297 585 374
rect 621 477 679 497
rect 621 443 633 477
rect 667 443 679 477
rect 621 409 679 443
rect 621 375 633 409
rect 667 375 679 409
rect 621 297 679 375
rect 715 477 795 497
rect 715 443 753 477
rect 787 443 795 477
rect 715 409 795 443
rect 715 375 753 409
rect 787 375 795 409
rect 715 297 795 375
<< ndiffc >>
rect 35 65 69 99
rect 133 77 167 111
rect 237 77 271 111
rect 538 82 572 116
rect 633 89 667 123
rect 753 86 787 120
<< pdiffc >>
rect 539 443 573 477
rect 35 331 69 365
rect 129 331 163 365
rect 233 335 267 369
rect 327 353 361 387
rect 432 328 466 362
rect 539 374 573 408
rect 633 443 667 477
rect 633 375 667 409
rect 753 443 787 477
rect 753 375 787 409
<< poly >>
rect 371 477 437 500
rect 585 497 621 523
rect 679 497 715 523
rect 371 443 383 477
rect 417 443 437 477
rect 371 427 437 443
rect 81 395 117 425
rect 279 395 315 425
rect 371 421 411 427
rect 373 395 409 421
rect 478 381 514 407
rect 81 296 117 311
rect 279 296 315 311
rect 373 296 409 311
rect 79 265 119 296
rect 277 265 317 296
rect 28 259 119 265
rect 21 249 119 259
rect 21 215 37 249
rect 71 215 119 249
rect 21 205 119 215
rect 28 199 119 205
rect 227 249 317 265
rect 227 215 237 249
rect 271 215 317 249
rect 371 240 411 296
rect 478 282 514 297
rect 585 282 621 297
rect 679 282 715 297
rect 476 265 516 282
rect 583 265 623 282
rect 677 265 717 282
rect 227 199 317 215
rect 89 137 119 199
rect 287 137 317 199
rect 381 137 411 240
rect 453 249 516 265
rect 453 215 463 249
rect 497 215 516 249
rect 453 199 516 215
rect 560 249 717 265
rect 560 215 570 249
rect 604 215 717 249
rect 560 199 717 215
rect 453 137 483 199
rect 593 177 623 199
rect 687 177 717 199
rect 89 27 119 53
rect 287 27 317 53
rect 381 27 411 53
rect 453 27 483 53
rect 593 21 623 47
rect 687 21 717 47
<< polycont >>
rect 383 443 417 477
rect 37 215 71 249
rect 237 215 271 249
rect 463 215 497 249
rect 570 215 604 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 17 365 80 527
rect 216 426 349 527
rect 17 331 35 365
rect 69 331 80 365
rect 17 315 80 331
rect 126 365 181 381
rect 126 331 129 365
rect 163 331 181 365
rect 29 249 82 265
rect 29 215 37 249
rect 71 215 82 249
rect 29 149 82 215
rect 126 249 181 331
rect 220 369 267 392
rect 220 335 233 369
rect 301 391 349 426
rect 383 477 498 493
rect 417 443 498 477
rect 383 425 498 443
rect 532 477 575 527
rect 532 443 539 477
rect 573 443 575 477
rect 532 408 575 443
rect 301 387 377 391
rect 301 353 327 387
rect 361 353 377 387
rect 432 362 470 378
rect 220 319 267 335
rect 466 328 470 362
rect 532 374 539 408
rect 573 374 575 408
rect 532 358 575 374
rect 625 477 718 493
rect 625 443 633 477
rect 667 443 718 477
rect 625 409 718 443
rect 625 375 633 409
rect 667 375 718 409
rect 625 359 718 375
rect 432 319 470 328
rect 220 285 604 319
rect 126 215 237 249
rect 271 215 293 249
rect 126 203 293 215
rect 17 99 71 115
rect 17 65 35 99
rect 69 65 71 99
rect 17 17 71 65
rect 126 111 181 203
rect 329 114 363 285
rect 558 249 604 285
rect 126 77 133 111
rect 167 77 181 111
rect 126 61 181 77
rect 221 111 363 114
rect 221 77 237 111
rect 271 77 363 111
rect 221 61 363 77
rect 397 215 463 249
rect 497 215 524 249
rect 397 153 524 215
rect 558 215 570 249
rect 558 199 604 215
rect 648 289 718 359
rect 752 477 805 527
rect 752 443 753 477
rect 787 443 805 477
rect 752 409 805 443
rect 752 375 753 409
rect 787 375 805 409
rect 752 325 805 375
rect 648 185 808 289
rect 397 61 474 153
rect 648 143 714 185
rect 633 123 714 143
rect 522 82 538 116
rect 572 82 588 116
rect 522 17 588 82
rect 667 89 714 123
rect 633 51 714 89
rect 752 120 805 149
rect 752 86 753 120
rect 787 86 805 120
rect 752 17 805 86
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
flabel corelocali s 401 425 435 459 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel corelocali s 672 85 706 119 0 FreeSans 200 0 0 0 X
port 8 nsew
flabel corelocali s 675 425 709 459 0 FreeSans 200 0 0 0 X
port 8 nsew
flabel corelocali s 29 221 63 255 0 FreeSans 400 0 0 0 A_N
port 1 nsew
flabel corelocali s 403 153 437 187 0 FreeSans 400 0 0 0 C
port 3 nsew
flabel corelocali s 747 238 747 238 0 FreeSans 200 0 0 0 X
port 8 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
rlabel comment s 0 0 0 0 4 and3b_2
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1544568
string GDS_START 1537716
<< end >>
