magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1472 561
rect 18 299 69 527
rect 103 333 169 493
rect 203 367 237 527
rect 271 333 337 493
rect 371 367 405 527
rect 439 333 505 493
rect 539 367 573 527
rect 607 333 673 493
rect 707 367 741 527
rect 775 333 841 493
rect 875 367 909 527
rect 943 333 1009 493
rect 1043 367 1077 527
rect 1111 333 1177 493
rect 1211 367 1245 527
rect 1279 333 1345 493
rect 103 293 1345 333
rect 1383 299 1454 527
rect 102 215 673 259
rect 728 215 824 293
rect 858 215 1261 255
rect 775 181 824 215
rect 1295 181 1345 293
rect 119 17 153 113
rect 287 17 321 113
rect 455 17 489 113
rect 623 17 657 113
rect 775 131 1345 181
rect 0 -17 1472 17
<< obsli1 >>
rect 18 147 741 181
rect 18 51 85 147
rect 187 51 253 147
rect 355 51 421 147
rect 523 51 589 147
rect 691 97 741 147
rect 1379 97 1454 181
rect 691 51 1454 97
<< metal1 >>
rect 0 496 1472 592
rect 0 -48 1472 48
<< labels >>
rlabel locali s 858 215 1261 255 6 A
port 1 nsew signal input
rlabel locali s 102 215 673 259 6 B
port 2 nsew signal input
rlabel locali s 1295 181 1345 293 6 Y
port 3 nsew signal output
rlabel locali s 1279 333 1345 493 6 Y
port 3 nsew signal output
rlabel locali s 1111 333 1177 493 6 Y
port 3 nsew signal output
rlabel locali s 943 333 1009 493 6 Y
port 3 nsew signal output
rlabel locali s 775 333 841 493 6 Y
port 3 nsew signal output
rlabel locali s 775 181 824 215 6 Y
port 3 nsew signal output
rlabel locali s 775 131 1345 181 6 Y
port 3 nsew signal output
rlabel locali s 728 215 824 293 6 Y
port 3 nsew signal output
rlabel locali s 607 333 673 493 6 Y
port 3 nsew signal output
rlabel locali s 439 333 505 493 6 Y
port 3 nsew signal output
rlabel locali s 271 333 337 493 6 Y
port 3 nsew signal output
rlabel locali s 103 333 169 493 6 Y
port 3 nsew signal output
rlabel locali s 103 293 1345 333 6 Y
port 3 nsew signal output
rlabel locali s 623 17 657 113 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 455 17 489 113 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 287 17 321 113 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 119 17 153 113 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 1472 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1472 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 1383 299 1454 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 1211 367 1245 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 1043 367 1077 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 875 367 909 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 707 367 741 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 539 367 573 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 371 367 405 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 203 367 237 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 18 299 69 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 1472 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 1472 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1472 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1710792
string GDS_START 1698500
<< end >>
