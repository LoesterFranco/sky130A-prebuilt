magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 301 333 377 493
rect 489 333 565 493
rect 677 333 753 493
rect 865 333 941 493
rect 1157 333 1233 493
rect 1345 333 1421 493
rect 1533 333 1609 493
rect 1721 333 1797 493
rect 301 289 1797 333
rect 22 215 88 255
rect 482 181 568 289
rect 636 215 1008 255
rect 1048 215 1422 255
rect 1533 215 1901 255
rect 301 127 568 181
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 18 333 85 493
rect 129 367 267 527
rect 18 299 171 333
rect 209 299 267 367
rect 421 367 455 527
rect 609 367 643 527
rect 797 367 831 527
rect 985 367 1123 527
rect 1277 367 1311 527
rect 1465 367 1499 527
rect 1653 367 1687 527
rect 132 255 171 299
rect 1841 289 1892 527
rect 132 215 395 255
rect 132 181 171 215
rect 18 147 171 181
rect 18 51 85 147
rect 129 17 179 109
rect 217 93 267 181
rect 677 127 1421 181
rect 1465 147 1892 181
rect 1465 93 1515 147
rect 217 51 1035 93
rect 1073 51 1515 93
rect 1559 17 1593 109
rect 1627 51 1703 147
rect 1747 17 1781 109
rect 1815 51 1892 147
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< labels >>
rlabel locali s 22 215 88 255 6 A_N
port 1 nsew signal input
rlabel locali s 636 215 1008 255 6 B
port 2 nsew signal input
rlabel locali s 1048 215 1422 255 6 C
port 3 nsew signal input
rlabel locali s 1533 215 1901 255 6 D
port 4 nsew signal input
rlabel locali s 1721 333 1797 493 6 Y
port 5 nsew signal output
rlabel locali s 1533 333 1609 493 6 Y
port 5 nsew signal output
rlabel locali s 1345 333 1421 493 6 Y
port 5 nsew signal output
rlabel locali s 1157 333 1233 493 6 Y
port 5 nsew signal output
rlabel locali s 865 333 941 493 6 Y
port 5 nsew signal output
rlabel locali s 677 333 753 493 6 Y
port 5 nsew signal output
rlabel locali s 489 333 565 493 6 Y
port 5 nsew signal output
rlabel locali s 482 181 568 289 6 Y
port 5 nsew signal output
rlabel locali s 301 333 377 493 6 Y
port 5 nsew signal output
rlabel locali s 301 289 1797 333 6 Y
port 5 nsew signal output
rlabel locali s 301 127 568 181 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -48 1932 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 1932 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1932 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2347334
string GDS_START 2331984
<< end >>
