magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 552 561
rect 55 208 395 346
rect 57 17 123 174
rect 429 108 495 527
rect 0 -17 552 17
<< metal1 >>
rect 0 496 552 592
rect 0 -48 552 48
<< labels >>
rlabel locali s 55 208 395 346 6 SHORT
port 1 nsew signal input
rlabel locali s 57 17 123 174 6 VGND
port 2 nsew ground bidirectional abutment
rlabel locali s 0 -17 552 17 8 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 552 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel locali s 429 108 495 527 6 VPWR
port 3 nsew power bidirectional abutment
rlabel locali s 0 527 552 561 6 VPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 0 496 552 592 6 VPWR
port 3 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 552 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2216638
string GDS_START 2213646
<< end >>
