magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 828 561
rect 37 289 71 527
rect 105 305 156 493
rect 190 447 256 527
rect 37 17 71 186
rect 105 162 139 305
rect 269 199 335 323
rect 369 199 427 275
rect 105 51 156 162
rect 675 435 725 527
rect 610 271 706 331
rect 654 153 706 271
rect 746 153 798 331
rect 190 17 276 106
rect 391 17 538 97
rect 721 17 801 119
rect 0 -17 828 17
<< obsli1 >>
rect 500 474 534 493
rect 308 440 534 474
rect 575 451 641 485
rect 308 395 342 440
rect 190 361 342 395
rect 488 413 534 440
rect 190 265 224 361
rect 395 343 429 381
rect 488 379 570 413
rect 173 199 224 265
rect 395 309 502 343
rect 468 165 502 309
rect 323 131 502 165
rect 536 174 570 379
rect 607 401 641 451
rect 759 401 793 493
rect 607 367 793 401
rect 536 140 606 174
rect 323 51 357 131
rect 572 51 606 140
<< metal1 >>
rect 0 496 828 592
rect 0 -48 828 48
<< labels >>
rlabel locali s 269 199 335 323 6 A1_N
port 1 nsew signal input
rlabel locali s 369 199 427 275 6 A2_N
port 2 nsew signal input
rlabel locali s 746 153 798 331 6 B1
port 3 nsew signal input
rlabel locali s 654 153 706 271 6 B2
port 4 nsew signal input
rlabel locali s 610 271 706 331 6 B2
port 4 nsew signal input
rlabel locali s 105 305 156 493 6 X
port 5 nsew signal output
rlabel locali s 105 162 139 305 6 X
port 5 nsew signal output
rlabel locali s 105 51 156 162 6 X
port 5 nsew signal output
rlabel locali s 721 17 801 119 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 391 17 538 97 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 190 17 276 106 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 37 17 71 186 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 828 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 828 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 675 435 725 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 190 447 256 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 37 289 71 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 828 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 828 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3463550
string GDS_START 3455822
<< end >>
