magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 1670 704
<< pwell >>
rect 0 0 1632 49
<< scnmos >>
rect 85 74 115 222
rect 171 74 201 222
rect 257 74 287 222
rect 343 74 373 222
rect 550 108 580 256
rect 636 108 666 256
rect 722 108 752 256
rect 820 108 850 256
rect 1026 74 1056 222
rect 1112 74 1142 222
rect 1212 74 1242 222
rect 1298 74 1328 222
rect 1412 74 1442 222
rect 1498 74 1528 222
<< pmoshvt >>
rect 86 392 116 560
rect 196 392 226 560
rect 286 392 316 560
rect 386 392 416 560
rect 510 392 540 560
rect 600 392 630 560
rect 717 392 747 592
rect 817 392 847 592
rect 1029 392 1059 592
rect 1119 392 1149 592
rect 1226 368 1256 592
rect 1326 368 1356 592
rect 1416 368 1446 592
rect 1506 368 1536 592
<< ndiff >>
rect 477 244 550 256
rect 27 207 85 222
rect 27 173 39 207
rect 73 173 85 207
rect 27 120 85 173
rect 27 86 39 120
rect 73 86 85 120
rect 27 74 85 86
rect 115 207 171 222
rect 115 173 126 207
rect 160 173 171 207
rect 115 74 171 173
rect 201 210 257 222
rect 201 176 212 210
rect 246 176 257 210
rect 201 120 257 176
rect 201 86 212 120
rect 246 86 257 120
rect 201 74 257 86
rect 287 189 343 222
rect 287 155 298 189
rect 332 155 343 189
rect 287 74 343 155
rect 373 104 423 222
rect 477 210 497 244
rect 531 210 550 244
rect 477 198 550 210
rect 500 108 550 198
rect 580 157 636 256
rect 580 123 591 157
rect 625 123 636 157
rect 580 108 636 123
rect 666 240 722 256
rect 666 206 677 240
rect 711 206 722 240
rect 666 154 722 206
rect 666 120 677 154
rect 711 120 722 154
rect 666 108 722 120
rect 752 163 820 256
rect 752 129 763 163
rect 797 129 820 163
rect 752 108 820 129
rect 850 240 909 256
rect 850 206 863 240
rect 897 206 909 240
rect 850 154 909 206
rect 850 120 863 154
rect 897 120 909 154
rect 850 108 909 120
rect 969 188 1026 222
rect 969 154 981 188
rect 1015 154 1026 188
rect 969 120 1026 154
rect 373 92 446 104
rect 373 74 400 92
rect 388 58 400 74
rect 434 58 446 92
rect 969 86 981 120
rect 1015 86 1026 120
rect 969 74 1026 86
rect 1056 210 1112 222
rect 1056 176 1067 210
rect 1101 176 1112 210
rect 1056 120 1112 176
rect 1056 86 1067 120
rect 1101 86 1112 120
rect 1056 74 1112 86
rect 1142 210 1212 222
rect 1142 176 1153 210
rect 1187 176 1212 210
rect 1142 120 1212 176
rect 1142 86 1153 120
rect 1187 86 1212 120
rect 1142 74 1212 86
rect 1242 210 1298 222
rect 1242 176 1253 210
rect 1287 176 1298 210
rect 1242 120 1298 176
rect 1242 86 1253 120
rect 1287 86 1298 120
rect 1242 74 1298 86
rect 1328 147 1412 222
rect 1328 113 1353 147
rect 1387 113 1412 147
rect 1328 74 1412 113
rect 1442 210 1498 222
rect 1442 176 1453 210
rect 1487 176 1498 210
rect 1442 120 1498 176
rect 1442 86 1453 120
rect 1487 86 1498 120
rect 1442 74 1498 86
rect 1528 147 1599 222
rect 1528 113 1553 147
rect 1587 113 1599 147
rect 1528 74 1599 113
rect 388 46 446 58
<< pdiff >>
rect 648 580 717 592
rect 648 560 660 580
rect 27 548 86 560
rect 27 514 39 548
rect 73 514 86 548
rect 27 440 86 514
rect 27 406 39 440
rect 73 406 86 440
rect 27 392 86 406
rect 116 513 196 560
rect 116 479 139 513
rect 173 479 196 513
rect 116 392 196 479
rect 226 548 286 560
rect 226 514 239 548
rect 273 514 286 548
rect 226 440 286 514
rect 226 406 239 440
rect 273 406 286 440
rect 226 392 286 406
rect 316 513 386 560
rect 316 479 339 513
rect 373 479 386 513
rect 316 392 386 479
rect 416 548 510 560
rect 416 514 446 548
rect 480 514 510 548
rect 416 438 510 514
rect 416 404 446 438
rect 480 404 510 438
rect 416 392 510 404
rect 540 513 600 560
rect 540 479 553 513
rect 587 479 600 513
rect 540 392 600 479
rect 630 546 660 560
rect 694 546 717 580
rect 630 512 717 546
rect 630 478 660 512
rect 694 478 717 512
rect 630 440 717 478
rect 630 406 660 440
rect 694 406 717 440
rect 630 392 717 406
rect 747 519 817 592
rect 747 485 760 519
rect 794 485 817 519
rect 747 392 817 485
rect 847 578 906 592
rect 847 544 860 578
rect 894 544 906 578
rect 847 392 906 544
rect 960 578 1029 592
rect 960 544 972 578
rect 1006 544 1029 578
rect 960 392 1029 544
rect 1059 580 1119 592
rect 1059 546 1072 580
rect 1106 546 1119 580
rect 1059 508 1119 546
rect 1059 474 1072 508
rect 1106 474 1119 508
rect 1059 392 1119 474
rect 1149 580 1226 592
rect 1149 546 1179 580
rect 1213 546 1226 580
rect 1149 508 1226 546
rect 1149 474 1179 508
rect 1213 474 1226 508
rect 1149 392 1226 474
rect 1173 368 1226 392
rect 1256 580 1326 592
rect 1256 546 1279 580
rect 1313 546 1326 580
rect 1256 497 1326 546
rect 1256 463 1279 497
rect 1313 463 1326 497
rect 1256 420 1326 463
rect 1256 386 1279 420
rect 1313 386 1326 420
rect 1256 368 1326 386
rect 1356 580 1416 592
rect 1356 546 1369 580
rect 1403 546 1416 580
rect 1356 504 1416 546
rect 1356 470 1369 504
rect 1403 470 1416 504
rect 1356 368 1416 470
rect 1446 580 1506 592
rect 1446 546 1459 580
rect 1493 546 1506 580
rect 1446 497 1506 546
rect 1446 463 1459 497
rect 1493 463 1506 497
rect 1446 414 1506 463
rect 1446 380 1459 414
rect 1493 380 1506 414
rect 1446 368 1506 380
rect 1536 580 1605 592
rect 1536 546 1559 580
rect 1593 546 1605 580
rect 1536 497 1605 546
rect 1536 463 1559 497
rect 1593 463 1605 497
rect 1536 414 1605 463
rect 1536 380 1559 414
rect 1593 380 1605 414
rect 1536 368 1605 380
<< ndiffc >>
rect 39 173 73 207
rect 39 86 73 120
rect 126 173 160 207
rect 212 176 246 210
rect 212 86 246 120
rect 298 155 332 189
rect 497 210 531 244
rect 591 123 625 157
rect 677 206 711 240
rect 677 120 711 154
rect 763 129 797 163
rect 863 206 897 240
rect 863 120 897 154
rect 981 154 1015 188
rect 400 58 434 92
rect 981 86 1015 120
rect 1067 176 1101 210
rect 1067 86 1101 120
rect 1153 176 1187 210
rect 1153 86 1187 120
rect 1253 176 1287 210
rect 1253 86 1287 120
rect 1353 113 1387 147
rect 1453 176 1487 210
rect 1453 86 1487 120
rect 1553 113 1587 147
<< pdiffc >>
rect 39 514 73 548
rect 39 406 73 440
rect 139 479 173 513
rect 239 514 273 548
rect 239 406 273 440
rect 339 479 373 513
rect 446 514 480 548
rect 446 404 480 438
rect 553 479 587 513
rect 660 546 694 580
rect 660 478 694 512
rect 660 406 694 440
rect 760 485 794 519
rect 860 544 894 578
rect 972 544 1006 578
rect 1072 546 1106 580
rect 1072 474 1106 508
rect 1179 546 1213 580
rect 1179 474 1213 508
rect 1279 546 1313 580
rect 1279 463 1313 497
rect 1279 386 1313 420
rect 1369 546 1403 580
rect 1369 470 1403 504
rect 1459 546 1493 580
rect 1459 463 1493 497
rect 1459 380 1493 414
rect 1559 546 1593 580
rect 1559 463 1593 497
rect 1559 380 1593 414
<< poly >>
rect 717 592 747 618
rect 817 592 847 618
rect 1029 592 1059 618
rect 1119 592 1149 618
rect 1226 592 1256 618
rect 1326 592 1356 618
rect 1416 592 1446 618
rect 1506 592 1536 618
rect 86 560 116 586
rect 196 560 226 586
rect 286 560 316 586
rect 386 560 416 586
rect 510 560 540 586
rect 600 560 630 586
rect 86 377 116 392
rect 196 377 226 392
rect 286 377 316 392
rect 386 377 416 392
rect 510 377 540 392
rect 600 377 630 392
rect 717 377 747 392
rect 817 377 847 392
rect 1029 377 1059 392
rect 1119 377 1149 392
rect 83 356 119 377
rect 193 356 229 377
rect 44 340 229 356
rect 44 306 60 340
rect 94 326 229 340
rect 283 356 319 377
rect 383 356 419 377
rect 283 340 419 356
rect 94 306 119 326
rect 44 290 119 306
rect 85 222 115 290
rect 171 222 201 326
rect 283 306 299 340
rect 333 306 419 340
rect 507 356 543 377
rect 597 356 633 377
rect 714 356 750 377
rect 814 356 850 377
rect 507 340 666 356
rect 507 326 613 340
rect 283 290 419 306
rect 550 306 613 326
rect 647 306 666 340
rect 550 290 666 306
rect 714 340 850 356
rect 714 306 730 340
rect 764 306 798 340
rect 832 306 850 340
rect 714 290 850 306
rect 283 267 373 290
rect 257 237 373 267
rect 550 256 580 290
rect 636 256 666 290
rect 722 256 752 290
rect 820 256 850 290
rect 1026 356 1062 377
rect 1116 356 1149 377
rect 1026 340 1146 356
rect 1226 353 1256 368
rect 1326 353 1356 368
rect 1416 353 1446 368
rect 1506 353 1536 368
rect 1026 306 1081 340
rect 1115 306 1146 340
rect 1026 290 1146 306
rect 1223 336 1259 353
rect 1323 336 1359 353
rect 1413 336 1449 353
rect 1223 320 1449 336
rect 1223 300 1239 320
rect 257 222 287 237
rect 343 222 373 237
rect 1026 222 1056 290
rect 1112 222 1142 290
rect 1212 286 1239 300
rect 1273 286 1307 320
rect 1341 286 1375 320
rect 1409 300 1449 320
rect 1503 300 1539 353
rect 1409 286 1539 300
rect 1212 270 1539 286
rect 1212 222 1242 270
rect 1298 222 1328 270
rect 1412 222 1442 270
rect 1498 222 1528 270
rect 85 48 115 74
rect 171 48 201 74
rect 257 48 287 74
rect 343 48 373 74
rect 550 82 580 108
rect 636 82 666 108
rect 722 82 752 108
rect 820 82 850 108
rect 1026 48 1056 74
rect 1112 48 1142 74
rect 1212 48 1242 74
rect 1298 48 1328 74
rect 1412 48 1442 74
rect 1498 48 1528 74
<< polycont >>
rect 60 306 94 340
rect 299 306 333 340
rect 613 306 647 340
rect 730 306 764 340
rect 798 306 832 340
rect 1081 306 1115 340
rect 1239 286 1273 320
rect 1307 286 1341 320
rect 1375 286 1409 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 23 548 89 564
rect 23 514 39 548
rect 73 514 89 548
rect 23 440 89 514
rect 123 513 189 649
rect 123 479 139 513
rect 173 479 189 513
rect 123 463 189 479
rect 223 548 289 564
rect 223 514 239 548
rect 273 514 289 548
rect 23 406 39 440
rect 73 424 89 440
rect 223 440 289 514
rect 323 513 389 649
rect 323 479 339 513
rect 373 479 389 513
rect 323 463 389 479
rect 430 548 496 564
rect 430 514 446 548
rect 480 514 496 548
rect 223 424 239 440
rect 73 406 239 424
rect 273 424 289 440
rect 430 438 496 514
rect 537 513 603 649
rect 537 479 553 513
rect 587 479 603 513
rect 537 463 603 479
rect 644 581 910 615
rect 644 580 710 581
rect 644 546 660 580
rect 694 546 710 580
rect 844 578 910 581
rect 644 512 710 546
rect 644 478 660 512
rect 694 478 710 512
rect 430 424 446 438
rect 273 406 446 424
rect 23 404 446 406
rect 480 424 496 438
rect 644 440 710 478
rect 744 519 810 547
rect 844 544 860 578
rect 894 544 910 578
rect 844 526 910 544
rect 956 578 1022 649
rect 956 544 972 578
rect 1006 544 1022 578
rect 956 526 1022 544
rect 1056 580 1122 596
rect 1056 546 1072 580
rect 1106 546 1122 580
rect 744 485 760 519
rect 794 492 810 519
rect 1056 508 1122 546
rect 1056 492 1072 508
rect 794 485 1072 492
rect 744 474 1072 485
rect 1106 474 1122 508
rect 744 458 1122 474
rect 1163 580 1229 649
rect 1163 546 1179 580
rect 1213 546 1229 580
rect 1163 508 1229 546
rect 1163 474 1179 508
rect 1213 474 1229 508
rect 1163 458 1229 474
rect 1263 580 1318 596
rect 1263 546 1279 580
rect 1313 546 1318 580
rect 1263 497 1318 546
rect 1263 463 1279 497
rect 1313 463 1318 497
rect 1353 580 1419 649
rect 1353 546 1369 580
rect 1403 546 1419 580
rect 1353 504 1419 546
rect 1353 470 1369 504
rect 1403 470 1419 504
rect 1459 580 1509 596
rect 1493 546 1509 580
rect 1459 497 1509 546
rect 644 424 660 440
rect 480 406 660 424
rect 694 424 710 440
rect 1263 436 1318 463
rect 1493 463 1509 497
rect 1459 436 1509 463
rect 694 406 1229 424
rect 480 404 1229 406
rect 23 390 1229 404
rect 25 340 110 356
rect 25 306 60 340
rect 94 306 110 340
rect 25 290 110 306
rect 144 226 178 390
rect 430 388 496 390
rect 217 340 359 356
rect 217 306 299 340
rect 333 306 359 340
rect 217 290 359 306
rect 597 340 663 356
rect 597 306 613 340
rect 647 306 663 340
rect 597 290 663 306
rect 697 340 1031 356
rect 697 306 730 340
rect 764 306 798 340
rect 832 306 1031 340
rect 697 290 1031 306
rect 1065 340 1131 356
rect 1065 306 1081 340
rect 1115 306 1131 340
rect 1065 290 1131 306
rect 1195 336 1229 390
rect 1263 420 1509 436
rect 1263 386 1279 420
rect 1313 414 1509 420
rect 1313 386 1459 414
rect 1263 380 1459 386
rect 1493 380 1509 414
rect 1263 370 1509 380
rect 1195 320 1425 336
rect 1195 286 1239 320
rect 1273 286 1307 320
rect 1341 286 1375 320
rect 1409 286 1425 320
rect 1459 330 1509 370
rect 1543 580 1609 649
rect 1543 546 1559 580
rect 1593 546 1609 580
rect 1543 497 1609 546
rect 1543 463 1559 497
rect 1593 463 1609 497
rect 1543 414 1609 463
rect 1543 380 1559 414
rect 1593 380 1609 414
rect 1543 364 1609 380
rect 1459 296 1607 330
rect 1195 270 1425 286
rect 473 256 555 260
rect 473 244 1101 256
rect 23 207 76 223
rect 23 173 39 207
rect 73 173 76 207
rect 23 120 76 173
rect 110 207 178 226
rect 110 173 126 207
rect 160 173 178 207
rect 110 154 178 173
rect 212 210 246 226
rect 212 120 246 176
rect 23 86 39 120
rect 73 86 212 120
rect 282 189 348 226
rect 473 210 497 244
rect 531 240 1101 244
rect 531 210 677 240
rect 282 155 298 189
rect 332 176 348 189
rect 661 206 677 210
rect 711 222 863 240
rect 332 157 625 176
rect 332 155 591 157
rect 282 142 591 155
rect 282 119 348 142
rect 575 123 591 142
rect 23 85 246 86
rect 384 92 450 108
rect 575 104 625 123
rect 661 154 711 206
rect 847 206 863 222
rect 897 222 1101 240
rect 1561 236 1607 296
rect 897 206 913 222
rect 661 120 677 154
rect 661 104 711 120
rect 747 163 813 188
rect 747 129 763 163
rect 797 129 813 163
rect 384 85 400 92
rect 23 58 400 85
rect 434 58 450 92
rect 23 51 450 58
rect 747 17 813 129
rect 847 154 913 206
rect 1067 210 1101 222
rect 847 120 863 154
rect 897 120 913 154
rect 847 104 913 120
rect 965 154 981 188
rect 1015 154 1031 188
rect 965 120 1031 154
rect 965 86 981 120
rect 1015 86 1031 120
rect 965 17 1031 86
rect 1067 120 1101 176
rect 1067 70 1101 86
rect 1137 210 1203 226
rect 1137 176 1153 210
rect 1187 176 1203 210
rect 1137 120 1203 176
rect 1137 86 1153 120
rect 1187 86 1203 120
rect 1137 17 1203 86
rect 1237 210 1607 236
rect 1237 176 1253 210
rect 1287 202 1453 210
rect 1287 176 1303 202
rect 1237 120 1303 176
rect 1437 176 1453 202
rect 1487 202 1607 210
rect 1487 176 1503 202
rect 1237 86 1253 120
rect 1287 86 1303 120
rect 1237 70 1303 86
rect 1337 147 1403 163
rect 1337 113 1353 147
rect 1387 113 1403 147
rect 1337 17 1403 113
rect 1437 120 1503 176
rect 1437 86 1453 120
rect 1487 86 1503 120
rect 1437 70 1503 86
rect 1537 147 1603 163
rect 1537 113 1553 147
rect 1587 113 1603 147
rect 1537 17 1603 113
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o2111a_4
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nwell s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 D1
port 5 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 1567 242 1601 276 0 FreeSans 340 0 0 0 X
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 1632 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1240600
string GDS_START 1227710
<< end >>
